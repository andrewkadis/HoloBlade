// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Fri Aug 28 16:25:58 2020
//
// Verilog Description of module top
//

module top (ICE_SYSCLK, DCD, DSR, DTR, CTS, RST, UART_RX, UART_TX, 
            SEN, SCK, SOUT, SDAT, UPDATE, RESET, SLM_CLK, INVERT, 
            SYNC, VALID, DATA31, DATA0, DATA30, DATA29, DATA1, 
            DATA28, DATA27, DATA2, DATA26, DATA25, DATA3, DATA24, 
            DATA23, DATA4, DATA22, DATA21, DATA5, DATA20, DATA19, 
            DATA6, DATA18, DATA17, DATA7, DATA16, DATA15, DATA8, 
            DATA14, DATA13, DATA12, DATA11, DATA9, DATA10, FT_OE, 
            FT_RD, FT_WR, FT_SIWU, FR_RXF, FT_TXE, FIFO_BE3, FIFO_BE2, 
            FIFO_BE1, FIFO_BE0, FIFO_D31, FIFO_D30, FIFO_D29, FIFO_D28, 
            FIFO_D27, FIFO_CLK, FIFO_D26, FIFO_D25, FIFO_D24, FIFO_D23, 
            FIFO_D22, FIFO_D21, FIFO_D20, FIFO_D19, FIFO_D18, FIFO_D17, 
            FIFO_D16, FIFO_D15, FIFO_D14, FIFO_D13, FIFO_D12, FIFO_D11, 
            FIFO_D10, FIFO_D9, FIFO_D8, FIFO_D7, FIFO_D6, FIFO_D5, 
            FIFO_D4, FIFO_D3, FIFO_D2, FIFO_D1, FIFO_D0, DEBUG_0, 
            DEBUG_1, DEBUG_2, DEBUG_3, DEBUG_5, DEBUG_6, DEBUG_8, 
            DEBUG_9, ICE_CLK, ICE_CDONE, ICE_CREST) /* synthesis syn_module_defined=1 */ ;   // src/top.v(5[8:11])
    input ICE_SYSCLK;   // src/top.v(8[11:21])
    output DCD;   // src/top.v(11[12:15])
    output DSR;   // src/top.v(12[12:15])
    output DTR;   // src/top.v(13[12:15])
    output CTS;   // src/top.v(14[12:15])
    output RST;   // src/top.v(15[12:15])
    input UART_RX;   // src/top.v(16[12:19])
    output UART_TX;   // src/top.v(17[12:19])
    output SEN;   // src/top.v(20[12:15])
    output SCK;   // src/top.v(21[12:15])
    input SOUT;   // src/top.v(22[12:16])
    output SDAT;   // src/top.v(23[12:16])
    output UPDATE;   // src/top.v(27[12:18])
    output RESET;   // src/top.v(28[12:17])
    output SLM_CLK;   // src/top.v(29[12:19])
    output INVERT;   // src/top.v(30[12:18])
    output SYNC;   // src/top.v(31[12:16])
    output VALID;   // src/top.v(32[12:17])
    output DATA31;   // src/top.v(34[12:18])
    output DATA0;   // src/top.v(35[12:17])
    output DATA30;   // src/top.v(36[12:18])
    output DATA29;   // src/top.v(37[12:18])
    output DATA1;   // src/top.v(38[12:17])
    output DATA28;   // src/top.v(39[12:18])
    output DATA27;   // src/top.v(40[12:18])
    output DATA2;   // src/top.v(41[12:17])
    output DATA26;   // src/top.v(42[12:18])
    output DATA25;   // src/top.v(43[12:18])
    output DATA3;   // src/top.v(44[12:17])
    output DATA24;   // src/top.v(45[12:18])
    output DATA23;   // src/top.v(46[12:18])
    output DATA4;   // src/top.v(47[12:17])
    output DATA22;   // src/top.v(48[12:18])
    output DATA21;   // src/top.v(49[12:18])
    output DATA5;   // src/top.v(50[12:17])
    output DATA20;   // src/top.v(51[12:18])
    output DATA19;   // src/top.v(52[12:18])
    output DATA6;   // src/top.v(53[12:17])
    output DATA18;   // src/top.v(54[12:18])
    output DATA17;   // src/top.v(55[12:18])
    output DATA7;   // src/top.v(56[12:17])
    output DATA16;   // src/top.v(57[12:18])
    output DATA15;   // src/top.v(58[12:18])
    output DATA8;   // src/top.v(59[12:17])
    output DATA14;   // src/top.v(60[12:18])
    output DATA13;   // src/top.v(61[12:18])
    output DATA12;   // src/top.v(62[12:18])
    output DATA11;   // src/top.v(63[12:18])
    output DATA9;   // src/top.v(64[12:17])
    output DATA10;   // src/top.v(65[12:18])
    output FT_OE;   // src/top.v(69[12:17])
    output FT_RD;   // src/top.v(70[12:17])
    output FT_WR;   // src/top.v(71[12:17])
    output FT_SIWU;   // src/top.v(72[12:19])
    input FR_RXF;   // src/top.v(73[12:18])
    input FT_TXE;   // src/top.v(74[12:18])
    input FIFO_BE3;   // src/top.v(75[12:20])
    input FIFO_BE2;   // src/top.v(76[12:20])
    input FIFO_BE1;   // src/top.v(77[12:20])
    input FIFO_BE0;   // src/top.v(78[12:20])
    input FIFO_D31;   // src/top.v(79[12:20])
    input FIFO_D30;   // src/top.v(80[12:20])
    input FIFO_D29;   // src/top.v(81[12:20])
    input FIFO_D28;   // src/top.v(82[12:20])
    input FIFO_D27;   // src/top.v(83[12:20])
    input FIFO_CLK;   // src/top.v(84[12:20])
    input FIFO_D26;   // src/top.v(85[12:20])
    input FIFO_D25;   // src/top.v(86[12:20])
    input FIFO_D24;   // src/top.v(87[12:20])
    input FIFO_D23;   // src/top.v(88[12:20])
    input FIFO_D22;   // src/top.v(89[12:20])
    input FIFO_D21;   // src/top.v(90[12:20])
    input FIFO_D20;   // src/top.v(91[12:20])
    input FIFO_D19;   // src/top.v(92[12:20])
    input FIFO_D18;   // src/top.v(93[12:20])
    input FIFO_D17;   // src/top.v(94[12:20])
    input FIFO_D16;   // src/top.v(95[12:20])
    input FIFO_D15;   // src/top.v(97[11:19])
    input FIFO_D14;   // src/top.v(98[11:19])
    input FIFO_D13;   // src/top.v(99[11:19])
    input FIFO_D12;   // src/top.v(100[11:19])
    input FIFO_D11;   // src/top.v(101[11:19])
    input FIFO_D10;   // src/top.v(102[11:19])
    input FIFO_D9;   // src/top.v(103[11:18])
    input FIFO_D8;   // src/top.v(104[11:18])
    input FIFO_D7;   // src/top.v(105[11:18])
    input FIFO_D6;   // src/top.v(106[11:18])
    input FIFO_D5;   // src/top.v(107[11:18])
    input FIFO_D4;   // src/top.v(108[11:18])
    input FIFO_D3;   // src/top.v(109[11:18])
    input FIFO_D2;   // src/top.v(110[11:18])
    input FIFO_D1;   // src/top.v(111[11:18])
    input FIFO_D0;   // src/top.v(112[11:18])
    output DEBUG_0;   // src/top.v(115[12:19])
    output DEBUG_1;   // src/top.v(116[12:19])
    output DEBUG_2;   // src/top.v(117[12:19])
    output DEBUG_3;   // src/top.v(118[12:19])
    output DEBUG_5;   // src/top.v(119[12:19])
    output DEBUG_6;   // src/top.v(120[12:19])
    output DEBUG_8;   // src/top.v(121[12:19])
    output DEBUG_9;   // src/top.v(122[12:19])
    output ICE_CLK;   // src/top.v(125[12:19])
    output ICE_CDONE;   // src/top.v(126[12:21])
    output ICE_CREST;   // src/top.v(127[12:21])
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    
    wire GND_net, VCC_net, ICE_SYSCLK_c, UART_RX_c, UART_TX_c, SEN_c_1, 
        SCK_c_0, SOUT_c, SDAT_c_15, UPDATE_c_2, RESET_c, INVERT_c_3, 
        SYNC_c, DEBUG_9_c, DEBUG_6_c, DATA1_c_1, DATA2_c_2, DATA3_c_3, 
        DATA4_c_4, DATA5_c_5, DATA6_c_6, DATA7_c_7, DATA15_c_15, DATA8_c_8, 
        DATA14_c_14, DATA13_c_13, DATA12_c_12, DATA11_c_11, DATA9_c_9, 
        DATA10_c_10, FT_OE_c, DEBUG_2_c, DEBUG_1_c_c, FIFO_D15_c_15, 
        FIFO_D14_c_14, FIFO_D13_c_13, FIFO_D12_c_12, FIFO_D11_c_11, 
        FIFO_D10_c_10, FIFO_D9_c_9, FIFO_D8_c_8, FIFO_D7_c_7, FIFO_D6_c_6, 
        FIFO_D5_c_5, FIFO_D4_c_4, FIFO_D3_c_3, FIFO_D2_c_2, FIFO_D1_c_1, 
        DEBUG_8_c_0_c, DEBUG_0_c_24, DEBUG_3_c, DEBUG_5_c, debug_led3, 
        reset_all_w;
    wire [3:0]reset_clk_counter;   // src/top.v(242[10:27])
    
    wire reset_per_frame, buffer_switch_done, dc32_fifo_almost_full, \REG.mem_13_13 , 
        \REG.mem_13_12 , \REG.mem_13_11 , \REG.mem_13_10 , \REG.mem_13_9 , 
        \REG.mem_13_8 , \REG.mem_13_7 , \REG.mem_13_6 , \REG.mem_11_15 , 
        \REG.mem_11_14 , \REG.mem_11_13 , \REG.mem_11_12 , \REG.mem_11_11 , 
        \REG.mem_11_10 , \REG.mem_11_9 ;
    wire [31:0]dc32_fifo_data_in;   // src/top.v(510[13:30])
    
    wire dc32_fifo_almost_empty, get_next_word, \REG.mem_9_14 , \REG.mem_9_13 , 
        \REG.mem_9_12 , \REG.mem_9_11 , \REG.mem_9_10 , \REG.mem_9_9 , 
        \REG.mem_9_8 , \REG.mem_9_7 , \REG.mem_9_6 , \REG.mem_9_5 , 
        \REG.mem_9_4 , \REG.mem_9_3 , \REG.mem_9_2 , \REG.mem_9_1 , 
        \REG.mem_9_0 ;
    wire [31:0]fifo_data_out;   // src/top.v(545[12:25])
    wire [7:0]pc_data_rx;   // src/top.v(685[11:21])
    
    wire \REG.mem_15_15 , tx_uart_active_flag, spi_start_transfer_r, multi_byte_spi_trans_flag_r;
    wire [7:0]tx_addr_byte;   // src/top.v(807[11:23])
    wire [7:0]tx_data_byte;   // src/top.v(809[11:23])
    wire [7:0]rx_buf_byte;   // src/top.v(816[11:22])
    
    wire is_tx_fifo_full_flag, fifo_write_cmd, spi_rx_byte_ready, fifo_read_cmd, 
        is_fifo_empty_flag;
    wire [31:0]fifo_temp_output;   // src/top.v(906[12:28])
    
    wire even_byte_flag, uart_rx_complete_rising_edge, uart_rx_complete_prev, 
        reset_all_w_N_61, \REG.mem_11_8 , \REG.mem_11_7 , start_tx_N_64, 
        pll_clk_unbuf, n7258;
    wire [3:0]state;   // src/timing_controller.v(48[11:16])
    
    wire n771, multi_byte_spi_trans_flag_r_N_72, \REG.mem_8_15 , \REG.mem_18_15 , 
        \REG.mem_18_14 , \REG.mem_18_13 , \REG.mem_18_12 , \REG.mem_18_11 , 
        \REG.mem_18_10 , \REG.mem_18_9 , \REG.mem_18_8 , \REG.mem_18_7 , 
        \REG.mem_18_6 , \REG.mem_18_5 , \REG.mem_18_4 , \REG.mem_18_3 , 
        \REG.mem_18_2 , \REG.mem_18_1 , \REG.mem_18_0 , n4253, \REG.mem_16_15 , 
        \REG.mem_16_14 , \REG.mem_16_13 , \REG.mem_16_12 , \REG.mem_16_11 , 
        \REG.mem_16_10 , \REG.mem_16_9 , \REG.mem_16_8 , \REG.mem_16_7 , 
        \REG.mem_16_6 , \REG.mem_16_5 , \REG.mem_16_4 , \REG.mem_16_3 , 
        \REG.mem_16_2 , \REG.mem_8_14 , \REG.mem_8_13 , \REG.mem_8_12 , 
        \REG.mem_8_11 , \REG.mem_8_10 , \REG.mem_8_9 , \REG.mem_8_8 , 
        \REG.mem_8_7 , \REG.mem_8_6 , \REG.mem_8_5 , \REG.mem_8_4 , 
        \REG.mem_8_3 , \REG.mem_8_2 , \REG.mem_8_1 , \REG.mem_8_0 , 
        \REG.mem_7_15 , \REG.mem_15_14 , reset_per_frame_latched, \REG.mem_11_6 , 
        n32, buffer_switch_done_latched, \REG.mem_11_5 , \REG.mem_11_4 , 
        \REG.mem_11_3 , \REG.mem_11_2 , \REG.mem_11_1 , \REG.mem_11_0 , 
        n2352, n4, \REG.mem_16_1 , \REG.mem_16_0 , n2034, n4945, 
        n2086, \REG.mem_22_15 , n4942, n4941, \REG.mem_22_14 , \REG.mem_12_2 , 
        \REG.mem_12_3 , write_to_dc32_fifo_latched_N_425, FT_OE_N_420, 
        \REG.mem_22_13 , \REG.mem_10_15 , \REG.mem_10_14 , \REG.mem_10_13 , 
        \REG.mem_22_12 , n4938, \REG.mem_10_12 , \REG.mem_22_11 , \REG.mem_22_10 , 
        \REG.mem_10_11 , \REG.mem_10_10 , \REG.mem_10_9 , \REG.mem_10_8 , 
        \REG.mem_10_7 , \REG.mem_10_6 , \REG.mem_14_11 , \REG.mem_14_12 , 
        \REG.mem_14_13 , \REG.mem_14_14 , \REG.mem_14_15 , \REG.mem_10_5 , 
        \REG.mem_10_4 , \REG.mem_10_3 , \REG.mem_10_2 , \REG.mem_10_1 , 
        \REG.mem_10_0 , \REG.mem_15_13 , \REG.mem_15_12 , \REG.mem_15_11 , 
        \REG.mem_15_10 , n4923, n4922, n4919, \REG.mem_9_15 , \REG.mem_3_0 , 
        \REG.mem_7_14 , \REG.mem_7_13 , \REG.mem_7_12 , \REG.mem_7_11 , 
        \REG.mem_13_5 , \REG.mem_15_9 , n4662, \REG.mem_15_8 , \REG.mem_15_7 , 
        \REG.mem_15_6 , \REG.mem_13_0 , n4916, \REG.mem_22_9 , n4911, 
        n4910, \REG.mem_22_8 , \REG.mem_22_7 , n4909, \REG.mem_22_6 , 
        \REG.mem_22_5 , \REG.mem_15_5 , \REG.mem_22_4 , \REG.mem_22_3 , 
        \REG.mem_22_2 , \REG.mem_22_1 , \REG.mem_22_0 , n4907, n4658, 
        n10700, n4904, n4903, n4901, n4899, n4898, n4897, n4896, 
        \REG.mem_7_10 , \REG.mem_7_9 , \REG.mem_7_8 , \REG.mem_7_7 , 
        \REG.mem_7_6 , \REG.mem_7_5 , \REG.mem_7_4 , \REG.mem_7_3 , 
        bluejay_data_out_31__N_736, bluejay_data_out_31__N_737, n575, 
        r_Rx_Data, n1879, n4893, \REG.mem_12_1 , \REG.mem_12_0 , \REG.mem_15_4 , 
        n4666, \REG.mem_14_10 , \REG.mem_14_8 , \REG.mem_14_7 , \REG.mem_15_3 , 
        n10662, n10681, n4661;
    wire [2:0]r_SM_Main_adj_1261;   // src/uart_tx.v(31[16:25])
    wire [7:0]r_Tx_Data;   // src/uart_tx.v(34[16:25])
    
    wire n10149;
    wire [2:0]r_SM_Main_2__N_844;
    wire [2:0]r_SM_Main_2__N_841;
    
    wire \REG.mem_15_2 , \REG.mem_14_6 , \REG.mem_14_5 , \REG.mem_15_1 , 
        n4667, \REG.mem_14_9 ;
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    wire [15:0]rx_shift_reg;   // src/spi.v(72[12:24])
    
    wire \REG.mem_15_0 , n4660, n4668, n4245, n4890, n4669, n4889, 
        n571, n24, n4888, n4887, n4883, n4882, \REG.mem_7_2 , 
        \REG.mem_7_1 , \REG.mem_7_0 , \REG.mem_14_2 , \REG.mem_14_1 , 
        \REG.mem_14_3 , \REG.mem_14_4 , \REG.mem_6_15 , \REG.mem_6_14 , 
        \REG.mem_6_13 , \REG.mem_6_12 , \REG.mem_6_11 , \REG.mem_6_10 , 
        \REG.mem_6_9 , \REG.mem_6_8 , \REG.mem_6_7 , \REG.mem_6_6 , 
        \REG.mem_6_5 , \REG.mem_6_4 , \REG.mem_6_3 , \REG.mem_6_2 , 
        \REG.mem_6_1 , \REG.mem_6_0 , \REG.mem_13_1 , \REG.mem_13_15 , 
        \REG.mem_13_2 , \REG.mem_13_3 ;
    wire [6:0]wr_addr_nxt_c;   // src/fifo_dc_32_lut_gen.v(198[29:42])
    wire [6:0]rp_sync1_r;   // src/fifo_dc_32_lut_gen.v(201[37:47])
    wire [6:0]wr_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(204[37:51])
    wire [6:0]rd_addr_r;   // src/fifo_dc_32_lut_gen.v(217[29:38])
    
    wire \REG.mem_14_0 ;
    wire [6:0]rd_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(221[30:42])
    wire [6:0]wp_sync1_r;   // src/fifo_dc_32_lut_gen.v(222[37:47])
    wire [6:0]rd_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(225[37:51])
    wire [6:0]rd_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(233[30:44])
    
    wire rd_fifo_en_w, \aempty_flag_impl.ae_flag_nxt_w , t_rd_fifo_en_w;
    wire [31:0]\REG.out_raw ;   // src/fifo_dc_32_lut_gen.v(879[47:54])
    wire [6:0]rd_addr_nxt_c_6__N_498;
    
    wire n4_adj_1220, \REG.mem_5_15 , \REG.mem_5_14 , \REG.mem_5_13 , 
        \REG.mem_5_12 , \REG.mem_5_11 , \REG.mem_5_10 , \REG.mem_5_9 , 
        \REG.mem_5_8 , \REG.mem_5_7 , \REG.mem_5_6 , \REG.mem_5_5 , 
        \REG.mem_5_4 , \REG.mem_5_3 , \REG.mem_5_2 , \REG.mem_5_1 , 
        \REG.mem_5_0 , n8, n4878, n4877, \REG.mem_4_15 , \REG.mem_4_14 , 
        \REG.mem_4_13 , \REG.mem_4_12 , \REG.mem_4_11 , \REG.mem_4_10 , 
        \REG.mem_4_9 , \REG.mem_4_8 , \REG.mem_4_7 , \REG.mem_4_6 , 
        \REG.mem_4_5 , \REG.mem_4_4 , \REG.mem_4_3 , \REG.mem_4_2 , 
        \REG.mem_4_1 , \REG.mem_4_0 , \REG.mem_13_14 , \REG.mem_13_4 , 
        wr_fifo_en_w, rd_fifo_en_w_adj_1221, rd_fifo_en_prev_r;
    wire [2:0]wr_addr_r_adj_1284;   // src/fifo_quad_word_mod.v(65[31:40])
    wire [2:0]wr_addr_p1_w_adj_1286;   // src/fifo_quad_word_mod.v(67[32:44])
    wire [2:0]rd_addr_r_adj_1287;   // src/fifo_quad_word_mod.v(69[31:40])
    wire [2:0]rd_addr_p1_w_adj_1289;   // src/fifo_quad_word_mod.v(71[32:44])
    
    wire n7462, n7440;
    wire [31:0]\mem_LUT.data_raw_r ;   // src/fifo_quad_word_mod.v(449[42:52])
    
    wire empty_o_N_1149, n15, n2944, \REG.mem_3_15 , \REG.mem_3_14 , 
        \REG.mem_3_13 , \REG.mem_3_12 , \REG.mem_3_11 , \REG.mem_3_10 , 
        \REG.mem_3_9 , \REG.mem_3_8 , \REG.mem_3_7 , \REG.mem_3_6 , 
        \REG.mem_3_5 , \REG.mem_3_4 , \REG.mem_3_3 , \REG.mem_3_2 , 
        \REG.mem_3_1 , n3022, n4875, n7347, n4872, n4869, n4864, 
        n4860, n4859, \REG.mem_12_9 , \REG.mem_12_8 , \REG.mem_12_7 , 
        n843, \REG.mem_12_6 , n6112, n10632, n4459, \REG.mem_12_15 , 
        \REG.mem_12_14 , \REG.mem_12_13 , \REG.mem_12_12 , n10098, \REG.mem_12_11 , 
        \REG.mem_12_10 , \REG.mem_12_4 , \REG.mem_12_5 , n6106, n1774, 
        n6103, \REG.mem_23_0 , \REG.mem_23_1 , \REG.mem_23_2 , \REG.mem_23_3 , 
        \REG.mem_23_4 , \REG.mem_23_5 , \REG.mem_23_6 , \REG.mem_23_7 , 
        \REG.mem_23_8 , \REG.mem_23_9 , \REG.mem_23_10 , \REG.mem_23_11 , 
        \REG.mem_23_12 , \REG.mem_23_13 , \REG.mem_23_14 , \REG.mem_23_15 , 
        n4192, \REG.mem_25_0 , \REG.mem_25_1 , \REG.mem_25_2 , \REG.mem_25_3 , 
        \REG.mem_25_4 , \REG.mem_25_5 , \REG.mem_25_6 , \REG.mem_25_7 , 
        \REG.mem_25_8 , \REG.mem_25_9 , \REG.mem_25_10 , \REG.mem_25_11 , 
        \REG.mem_25_12 , \REG.mem_25_13 , \REG.mem_25_14 , \REG.mem_25_15 , 
        n4659, \REG.mem_30_0 , \REG.mem_30_1 , \REG.mem_30_2 , \REG.mem_30_3 , 
        \REG.mem_30_4 , \REG.mem_30_5 , \REG.mem_30_6 , \REG.mem_30_7 , 
        \REG.mem_30_8 , \REG.mem_30_9 , \REG.mem_30_10 , \REG.mem_30_11 , 
        \REG.mem_30_12 , \REG.mem_30_13 , \REG.mem_30_14 , \REG.mem_30_15 , 
        n6098, n4664, \REG.mem_31_0 , \REG.mem_31_1 , \REG.mem_31_2 , 
        \REG.mem_31_3 , \REG.mem_31_4 , \REG.mem_31_5 , \REG.mem_31_6 , 
        \REG.mem_31_7 , \REG.mem_31_8 , \REG.mem_31_9 , \REG.mem_31_10 , 
        \REG.mem_31_11 , \REG.mem_31_12 , \REG.mem_31_13 , \REG.mem_31_14 , 
        \REG.mem_31_15 , n4665, n10384, n4676, \REG.mem_35_0 , \REG.mem_35_1 , 
        \REG.mem_35_2 , \REG.mem_35_3 , \REG.mem_35_4 , \REG.mem_35_5 , 
        \REG.mem_35_6 , \REG.mem_35_7 , \REG.mem_35_8 , \REG.mem_35_9 , 
        \REG.mem_35_10 , \REG.mem_35_11 , \REG.mem_35_12 , \REG.mem_35_13 , 
        \REG.mem_35_14 , \REG.mem_35_15 , n10300, \REG.mem_36_0 , \REG.mem_36_1 , 
        \REG.mem_36_2 , \REG.mem_36_3 , \REG.mem_36_4 , \REG.mem_36_5 , 
        \REG.mem_36_6 , \REG.mem_36_7 , \REG.mem_36_8 , \REG.mem_36_9 , 
        \REG.mem_36_10 , \REG.mem_36_11 , \REG.mem_36_12 , \REG.mem_36_13 , 
        \REG.mem_36_14 , \REG.mem_36_15 , \REG.mem_37_0 , \REG.mem_37_1 , 
        \REG.mem_37_2 , \REG.mem_37_3 , \REG.mem_37_4 , \REG.mem_37_5 , 
        \REG.mem_37_6 , \REG.mem_37_7 , \REG.mem_37_8 , \REG.mem_37_9 , 
        \REG.mem_37_10 , \REG.mem_37_11 , \REG.mem_37_12 , \REG.mem_37_13 , 
        \REG.mem_37_14 , \REG.mem_37_15 , n11939, \REG.mem_38_0 , \REG.mem_38_1 , 
        \REG.mem_38_2 , \REG.mem_38_3 , \REG.mem_38_4 , \REG.mem_38_5 , 
        \REG.mem_38_6 , \REG.mem_38_7 , \REG.mem_38_8 , \REG.mem_38_9 , 
        \REG.mem_38_10 , \REG.mem_38_11 , \REG.mem_38_12 , \REG.mem_38_13 , 
        \REG.mem_38_14 , \REG.mem_38_15 , \REG.mem_39_0 , \REG.mem_39_1 , 
        \REG.mem_39_2 , \REG.mem_39_3 , \REG.mem_39_4 , \REG.mem_39_5 , 
        \REG.mem_39_6 , \REG.mem_39_7 , \REG.mem_39_8 , \REG.mem_39_9 , 
        \REG.mem_39_10 , \REG.mem_39_11 , \REG.mem_39_12 , \REG.mem_39_13 , 
        \REG.mem_39_14 , \REG.mem_39_15 , n13895, \REG.mem_40_0 , \REG.mem_40_1 , 
        \REG.mem_40_2 , \REG.mem_40_3 , \REG.mem_40_4 , \REG.mem_40_5 , 
        \REG.mem_40_6 , \REG.mem_40_7 , \REG.mem_40_8 , \REG.mem_40_9 , 
        \REG.mem_40_10 , \REG.mem_40_11 , \REG.mem_40_12 , \REG.mem_40_13 , 
        \REG.mem_40_14 , \REG.mem_40_15 , \REG.mem_41_0 , \REG.mem_41_1 , 
        \REG.mem_41_2 , \REG.mem_41_3 , \REG.mem_41_4 , \REG.mem_41_5 , 
        \REG.mem_41_6 , \REG.mem_41_7 , \REG.mem_41_8 , \REG.mem_41_9 , 
        \REG.mem_41_10 , \REG.mem_41_11 , \REG.mem_41_12 , \REG.mem_41_13 , 
        \REG.mem_41_14 , \REG.mem_41_15 , n10302, \REG.mem_42_0 , \REG.mem_42_1 , 
        \REG.mem_42_2 , \REG.mem_42_3 , \REG.mem_42_4 , \REG.mem_42_5 , 
        \REG.mem_42_6 , \REG.mem_42_7 , \REG.mem_42_8 , \REG.mem_42_9 , 
        \REG.mem_42_10 , \REG.mem_42_11 , \REG.mem_42_12 , \REG.mem_42_13 , 
        \REG.mem_42_14 , \REG.mem_42_15 , \REG.mem_43_0 , \REG.mem_43_1 , 
        \REG.mem_43_2 , \REG.mem_43_3 , \REG.mem_43_4 , \REG.mem_43_5 , 
        \REG.mem_43_6 , \REG.mem_43_7 , \REG.mem_43_8 , \REG.mem_43_9 , 
        \REG.mem_43_10 , \REG.mem_43_11 , \REG.mem_43_12 , \REG.mem_43_13 , 
        \REG.mem_43_14 , \REG.mem_43_15 , \REG.mem_44_0 , \REG.mem_44_1 , 
        \REG.mem_44_2 , \REG.mem_44_3 , \REG.mem_44_4 , \REG.mem_44_5 , 
        \REG.mem_44_6 , \REG.mem_44_7 , \REG.mem_44_8 , \REG.mem_44_9 , 
        \REG.mem_44_10 , \REG.mem_44_11 , \REG.mem_44_12 , \REG.mem_44_13 , 
        \REG.mem_44_14 , \REG.mem_44_15 , n6087, \REG.mem_45_0 , \REG.mem_45_1 , 
        \REG.mem_45_2 , \REG.mem_45_3 , \REG.mem_45_4 , \REG.mem_45_5 , 
        \REG.mem_45_6 , \REG.mem_45_7 , \REG.mem_45_8 , \REG.mem_45_9 , 
        \REG.mem_45_10 , \REG.mem_45_11 , \REG.mem_45_12 , \REG.mem_45_13 , 
        \REG.mem_45_14 , \REG.mem_45_15 , n10748, \REG.mem_46_0 , \REG.mem_46_1 , 
        \REG.mem_46_2 , \REG.mem_46_3 , \REG.mem_46_4 , \REG.mem_46_5 , 
        \REG.mem_46_6 , \REG.mem_46_7 , \REG.mem_46_8 , \REG.mem_46_9 , 
        \REG.mem_46_10 , \REG.mem_46_11 , \REG.mem_46_12 , \REG.mem_46_13 , 
        \REG.mem_46_14 , \REG.mem_46_15 , \REG.mem_47_0 , \REG.mem_47_1 , 
        \REG.mem_47_2 , \REG.mem_47_3 , \REG.mem_47_4 , \REG.mem_47_5 , 
        \REG.mem_47_6 , \REG.mem_47_7 , \REG.mem_47_8 , \REG.mem_47_9 , 
        \REG.mem_47_10 , \REG.mem_47_11 , \REG.mem_47_12 , \REG.mem_47_13 , 
        \REG.mem_47_14 , \REG.mem_47_15 , n3495, \REG.mem_48_0 , \REG.mem_48_1 , 
        \REG.mem_48_2 , \REG.mem_48_3 , \REG.mem_48_4 , \REG.mem_48_5 , 
        \REG.mem_48_6 , \REG.mem_48_7 , \REG.mem_48_8 , \REG.mem_48_9 , 
        \REG.mem_48_10 , \REG.mem_48_11 , \REG.mem_48_12 , \REG.mem_48_13 , 
        \REG.mem_48_14 , \REG.mem_48_15 , n6083, n4663, n4672, \REG.mem_50_0 , 
        \REG.mem_50_1 , \REG.mem_50_2 , \REG.mem_50_3 , \REG.mem_50_4 , 
        \REG.mem_50_5 , \REG.mem_50_6 , \REG.mem_50_7 , \REG.mem_50_8 , 
        \REG.mem_50_9 , \REG.mem_50_10 , \REG.mem_50_11 , \REG.mem_50_12 , 
        \REG.mem_50_13 , \REG.mem_50_14 , \REG.mem_50_15 , \REG.mem_54_0 , 
        \REG.mem_54_1 , \REG.mem_54_2 , \REG.mem_54_3 , \REG.mem_54_4 , 
        \REG.mem_54_5 , \REG.mem_54_6 , \REG.mem_54_7 , \REG.mem_54_8 , 
        \REG.mem_54_9 , \REG.mem_54_10 , \REG.mem_54_11 , \REG.mem_54_12 , 
        \REG.mem_54_13 , \REG.mem_54_14 , \REG.mem_54_15 , \REG.mem_55_0 , 
        \REG.mem_55_1 , \REG.mem_55_2 , \REG.mem_55_3 , \REG.mem_55_4 , 
        \REG.mem_55_5 , \REG.mem_55_6 , \REG.mem_55_7 , \REG.mem_55_8 , 
        \REG.mem_55_9 , \REG.mem_55_10 , \REG.mem_55_11 , \REG.mem_55_12 , 
        \REG.mem_55_13 , \REG.mem_55_14 , \REG.mem_55_15 , n10834, \REG.mem_57_0 , 
        \REG.mem_57_1 , \REG.mem_57_2 , \REG.mem_57_3 , \REG.mem_57_4 , 
        \REG.mem_57_5 , \REG.mem_57_6 , \REG.mem_57_7 , \REG.mem_57_8 , 
        \REG.mem_57_9 , \REG.mem_57_10 , \REG.mem_57_11 , \REG.mem_57_12 , 
        \REG.mem_57_13 , \REG.mem_57_14 , \REG.mem_57_15 , \REG.mem_62_0 , 
        \REG.mem_62_1 , \REG.mem_62_2 , \REG.mem_62_3 , \REG.mem_62_4 , 
        \REG.mem_62_5 , \REG.mem_62_6 , \REG.mem_62_7 , \REG.mem_62_8 , 
        \REG.mem_62_9 , \REG.mem_62_10 , \REG.mem_62_11 , \REG.mem_62_12 , 
        \REG.mem_62_13 , \REG.mem_62_14 , \REG.mem_62_15 , \REG.mem_63_0 , 
        \REG.mem_63_1 , \REG.mem_63_2 , \REG.mem_63_3 , \REG.mem_63_4 , 
        \REG.mem_63_5 , \REG.mem_63_6 , \REG.mem_63_7 , \REG.mem_63_8 , 
        \REG.mem_63_9 , \REG.mem_63_10 , \REG.mem_63_11 , \REG.mem_63_12 , 
        \REG.mem_63_13 , \REG.mem_63_14 , \REG.mem_63_15 , n2, n3, 
        n8_adj_1223, n10, n11, n15_adj_1224, n17, n18, n19, n20, 
        n21, n22, n23, n24_adj_1225, n25, n26, n27, n28, n29, 
        n30, n34, n35, n40, n42, n43, n47, n49, n50, n51, 
        n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, 
        n62, n6073, n6070, n6067, n6066, n6064, n6063, n6062, 
        n63, n6060, n6049, n6048, n6047, n6046, n6045, n6044, 
        n6043, n6034, n6032, n6030, n10790, n6013, n6012, n6011, 
        n6010, n6009, n6008, n4858, n6007, n6006, n6005, n6004, 
        n6003, n6002, n6001, n6000, n5999, n5998, n5997, n5996, 
        n5995, n5994, n5993, n5992, n5991, n5990, n5989, n5988, 
        n5987, n5986, n5985, n5984, n5983, n5982, n5981, n5963, 
        n5946, n5945, n5944, n5943, n5942, n5941, n5940, n5939, 
        n5938, n5921, n5920, n5919, n5917, n5916, n5914, n5894, 
        n5893, n5892, n5891, n5890, n5889, n5888, n5887, n5886, 
        n5885, n5884, n5883, n5882, n5881, n5880, n5879, n5861, 
        n5860, n5859, n5858, n5857, n5856, n5855, n5854, n5853, 
        n5852, n5851, n5850, n5849, n5848, n5847, n5846, n5845, 
        n5844, n5843, n5842, n5841, n5840, n5839, n5838, n5836, 
        n5835, n5834, n5833, n5832, n5831, n5830, n5829, n5828, 
        n5827, n5826, n5825, n5824, n5823, n5822, n5821, n5820, 
        n5819, n5818, n5817, n5768, n5767, n5766, n5765, n5764, 
        n5763, n5762, n5761, n5760, n5759, n5758, n5757, n5756, 
        n5755, n5754, n5750, n10211, n3794, n5733, n5732, n5731, 
        n5730, n5729, n5728, n5727, n5726, n5725, n5724, n5723, 
        n5722, n5721, n5720, n5719, n5718, n5717, n5716, n5715, 
        n5714, n5713, n5712, n5711, n5710, n5709, n5708, n5707, 
        n5706, n5705, n5704, n5703, n5702, n5701, n5700, n5699, 
        n5698, n5697, n5696, n5695, n5694, n5693, n5692, n5691, 
        n5690, n5689, n5688, n5687, n4671, n5686, n5685, n5684, 
        n5683, n5682, n5681, n5680, n5679, n5678, n5677, n5676, 
        n5675, n5674, n5673, n5672, n5671, n5670, n5668, n5667, 
        n10754, n5665, n5664, n5663, n5661, n5660, n5659, n5658, 
        n5657, n5656, n5655, n5654, n5653, n5652, n5651, n5650, 
        n5649, n5648, n5647, n5646, n5645, n5644, n5643, n5642, 
        n5641, n5640, n5639, n5638, n5637, n5636, n5635, n5634, 
        n5633, n5632, n5631, n5630, n5629, n5628, n5627, n5626, 
        n5625, n5624, n5623, n5622, n5621, n5620, n5619, n5618, 
        n5617, n5616, n5615, n5614, n5613, n5612, n5611, n5610, 
        n5609, n5608, n5607, n5606, n5605, n5604, n5603, n5602, 
        n5601, n5600, n5599, n5598, n5597, n5596, n5595, n5594, 
        n5593, n5592, n5591, n5590, n5589, n5588, n5587, n5586, 
        n5585, n5584, n5583, n5582, n5581, n5580, n5579, n5578, 
        n5577, n5576, n5575, n5574, n5573, n5572, n5570, n5569, 
        n5568, n5567, n5566, n5565, n5564, n5563, n5562, n5561, 
        n5560, n5559, n5558, n5557, n5556, n5555, n5554, n5553, 
        n5552, n5551, n5550, n5549, n5548, n5547, n5546, n5545, 
        n5544, n5543, n5542, n5541, n5540, n5539, n5538, n5537, 
        n5534, n5531, n5530, n5529, n5528, n5527, n4248, n10067, 
        n5526, n5525, n5524, n5523, n5522, n5521, n5520, n5519, 
        n5518, n5517, n5516, n5515, n5514, n5513, n5512, n5511, 
        n10066, n5510, n5509, n5508, n5505, n5504, n5503, n5502, 
        n5501, n5500, n5499, n5498, n5497, n5496, n5495, n10065, 
        n10064, n5494, n5493, n5492, n5491, n5490, n10063, n10062, 
        n10061, n10060, n10059, n10058, n10057, n130, n129, n128, 
        n127, n126, n125, n124, n123, n122, n121, n120, n5440, 
        n5439, n5438, n5437, n5436, n5435, n5434, n5433, n5432, 
        n5431, n119, n118, n117, n116, n115, n114, n113, n112, 
        n111, n110, n109, n108, n107, n106, n5430, n5429, n5428, 
        n5427, n5426, n5425, n5424, n5423, n5422, n5421, n5420, 
        n5419, n5418, n5417, n5416, n5415, n10056, n10055, n5414, 
        n5413, n5412, n5411, n5410, n5409, n10054, n10053, n10052, 
        n10051, n10050, n10049, n25_adj_1226, n24_adj_1227, n23_adj_1228, 
        n22_adj_1229, n21_adj_1230, n5344, n5343, n5342, n5341, 
        n5340, n5339, n5338, n5337, n5336, n5335, n20_adj_1231, 
        n19_adj_1232, n18_adj_1233, n17_adj_1234, n16, n15_adj_1235, 
        n14, n13, n12, n11_adj_1236, n10_adj_1237, n9, n8_adj_1238, 
        n7, n6, n5, n5334, n5333, n5332, n5331, n5330, n5329, 
        n4_adj_1239, n3_adj_1240, n2_adj_1241, n10048, n10047, n10046, 
        n25_adj_1242, n10045, n5313, n5310, n5306, n5305, n5304, 
        n5303, n10044, n5302, n5301, n5300, n5299, n5298, n5297, 
        n5296, n5295, n5294, n5293, n5292, n5291, n5290, n5289, 
        n5288, n5287, n5286, n5285, n5284, n5283, n5282, n5281, 
        n5280, n5279, n5278, n5277, n4855, n4854, n4851, n4848, 
        n5276, n5275, n9936, n5226, n5225, n5224, n5223, n5222, 
        n5221, n5220, n5219, n5218, n5217, n5216, n5215, n5214, 
        n5213, n5212, n5211, n4845, n4844, n4841, n4838, n5194, 
        n5193, n5192, n5191, n5190, n5189, n5188, n5187, n5186, 
        n5185, n5184, n5183, n5182, n5181, n5180, n5179, n5178, 
        n5177, n5176, n5175, n5174, n5173, n5172, n5171, n5170, 
        n5169, n5168, n5167, n5166, n5165, n5164, n5163, n5162, 
        n5161, n5160, n5159, n5158, n5157, n5156, n5155, n5154, 
        n4824, n5153, n5152, n5151, n5150, n5149, n5148, n5147, 
        n5146, n5145, n5144, n5143, n5142, n5141, n5140, n5139, 
        n5138, n5137, n5136, n5135, n5134, n5133, n5132, n5131, 
        n5130, n5129, n5128, n4836, n4834, n4830, n4827, n5127, 
        n5126, n5125, n5124, n5123, n5122, n5121, n5120, n5119, 
        n5118, n5117, n5116, n5115, n5114, n5113, n5112, n5111, 
        n5110, n5109, n5108, n5107, n5106, n5105, n5104, n5103, 
        n5102, n5101, n5100, n5099, n5098, n5097, n5096, n5095, 
        n5094, n5093, n5092, n5091, n5090, n5089, n5088, n5087, 
        n5086, n5085, n5084, n5083, n5082, n5081, n5080, n5079, 
        n5078, n5077, n5076, n5075, n5074, n5073, n5072, n5071, 
        n5070, n5069, n5068, n5067, n5066, n5065, n5064, n5063, 
        n5062, n5061, n5060, n5059, n5058, n5057, n5056, n5055, 
        n5054, n5053, n5052, n5051, n5050, n5049, n5048, n5047, 
        n5046, n5045, n5044, n5043, n5042, n5041, n5040, n5039, 
        n5038, n5037, n5036, n5035, n5034, n5033, n5032, n5031, 
        n5030, n5029, n5028, n5027, n5026, n5025, n5024, n5023, 
        n5022, n5021, n5020, n5019, n5018, n5017, n5016, n5015, 
        n10712, n5014, n5013, n5012, n5011, n5010, n5009, n5008, 
        n5007, n5006, n5005, n10653, n5004, n5003, n5002, n5001, 
        n5000, n4999, n4998, n4997, n4996, n4995, n4994, n4993, 
        n4992, n4991, n4990, n4989, n4988, n4987, n4986, n4985, 
        n4984, n4983, n4982, n4981, n4980, n4979, n4978, n4977, 
        n4976, n4319, n4975, n4670, n4974, n10706, n4973, n4972, 
        n4312, n4_adj_1243, n4971, n4970, n4_adj_1244, n4969, n4968, 
        n4967, n4966, n4965, n4964, n10167, n1, n13737, n10165, 
        n10163;
    
    VCC i2 (.Y(VCC_net));
    timing_controller timing_controller_inst (.state({state}), .SLM_CLK_c(SLM_CLK_c), 
            .n1879(n1879), .GND_net(GND_net), .n10384(n10384), .VCC_net(VCC_net), 
            .n10662(n10662), .reset_per_frame(reset_per_frame), .n1774(n1774), 
            .n7258(n7258), .INVERT_c_3(INVERT_c_3), .buffer_switch_done(buffer_switch_done), 
            .n4245(n4245), .n7440(n7440), .n7462(n7462), .n4192(n4192), 
            .n63(n63), .n10681(n10681), .UPDATE_c_2(UPDATE_c_2)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(452[19] 464[2])
    SB_LUT4 i4607_3_lut (.I0(\REG.mem_62_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n3), .I3(GND_net), .O(n5990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4270_3_lut (.I0(\REG.mem_44_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n21), .I3(GND_net), .O(n5653));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4207_3_lut (.I0(\REG.mem_40_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n25), .I3(GND_net), .O(n5590));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4271_3_lut (.I0(\REG.mem_44_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n21), .I3(GND_net), .O(n5654));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4608_3_lut (.I0(\REG.mem_62_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n3), .I3(GND_net), .O(n5991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4208_3_lut (.I0(\REG.mem_40_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n25), .I3(GND_net), .O(n5591));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4272_3_lut (.I0(\REG.mem_44_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n21), .I3(GND_net), .O(n5655));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4232_3_lut (.I0(\REG.mem_41_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4209_3_lut (.I0(\REG.mem_40_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n25), .I3(GND_net), .O(n5592));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4209_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF uart_rx_complete_prev_83 (.Q(uart_rx_complete_prev), .C(SLM_CLK_c), 
           .D(debug_led3));   // src/top.v(1065[8] 1071[4])
    bluejay_data bluejay_data_inst (.dc32_fifo_almost_full(dc32_fifo_almost_full), 
            .n843(n843), .GND_net(GND_net), .DEBUG_9_c(DEBUG_9_c), .SLM_CLK_c(SLM_CLK_c), 
            .n771(n771), .buffer_switch_done_latched(buffer_switch_done_latched), 
            .dc32_fifo_almost_empty(dc32_fifo_almost_empty), .bluejay_data_out_31__N_736(bluejay_data_out_31__N_736), 
            .buffer_switch_done(buffer_switch_done), .bluejay_data_out_31__N_737(bluejay_data_out_31__N_737), 
            .n6087(n6087), .DEBUG_6_c(DEBUG_6_c), .VCC_net(VCC_net), .SYNC_c(SYNC_c), 
            .n10149(n10149), .\rd_sig_diff0_w[1] (rd_sig_diff0_w[1]), .get_next_word(get_next_word), 
            .\rd_sig_diff0_w[0] (rd_sig_diff0_w[0]), .\rd_sig_diff0_w[2] (rd_sig_diff0_w[2]), 
            .n10700(n10700), .n10748(n10748), .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .DATA10_c_10(DATA10_c_10), .n4672(n4672), .DATA9_c_9(DATA9_c_9), 
            .n4671(n4671), .DATA11_c_11(DATA11_c_11), .n4670(n4670), .DATA12_c_12(DATA12_c_12), 
            .n4669(n4669), .DATA13_c_13(DATA13_c_13), .n4668(n4668), .DATA14_c_14(DATA14_c_14), 
            .n4667(n4667), .DATA8_c_8(DATA8_c_8), .n4666(n4666), .DATA15_c_15(DATA15_c_15), 
            .n4665(n4665), .DATA7_c_7(DATA7_c_7), .n4664(n4664), .DATA6_c_6(DATA6_c_6), 
            .n4663(n4663), .DATA5_c_5(DATA5_c_5), .n4662(n4662), .DATA4_c_4(DATA4_c_4), 
            .n4661(n4661), .DATA3_c_3(DATA3_c_3), .n4660(n4660), .DATA2_c_2(DATA2_c_2), 
            .n4659(n4659), .DATA1_c_1(DATA1_c_1), .n4658(n4658)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(626[14] 639[2])
    SB_LUT4 i4210_3_lut (.I0(\REG.mem_40_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n25), .I3(GND_net), .O(n5593));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4210_3_lut.LUT_INIT = 16'hcaca;
    SB_GB clk_gb (.GLOBAL_BUFFER_OUTPUT(SLM_CLK_c), .USER_SIGNAL_TO_GLOBAL_BUFFER(pll_clk_unbuf)) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/clock.v(82[7:96])
    SB_LUT4 i4211_3_lut (.I0(\REG.mem_40_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n25), .I3(GND_net), .O(n5594));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4212_3_lut (.I0(\REG.mem_40_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n25), .I3(GND_net), .O(n5595));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4213_3_lut (.I0(\REG.mem_40_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n25), .I3(GND_net), .O(n5596));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4233_3_lut (.I0(\REG.mem_41_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5616));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4233_3_lut.LUT_INIT = 16'hcaca;
    SB_IO RST_pad (.PACKAGE_PIN(RST), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RST_pad.PIN_TYPE = 6'b011001;
    defparam RST_pad.PULLUP = 1'b0;
    defparam RST_pad.NEG_TRIGGER = 1'b0;
    defparam RST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4234_3_lut (.I0(\REG.mem_41_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5617));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3458_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [5]), .I3(fifo_data_out[5]), .O(n4841));
    defparam i3458_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4273_3_lut (.I0(\REG.mem_44_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n21), .I3(GND_net), .O(n5656));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4609_3_lut (.I0(\REG.mem_62_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n3), .I3(GND_net), .O(n5992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3516_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4899));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i3516_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3520_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4903));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i3520_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4610_3_lut (.I0(\REG.mem_62_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n3), .I3(GND_net), .O(n5993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3521_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4904));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i3521_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3461_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [6]), .I3(fifo_data_out[6]), .O(n4844));
    defparam i3461_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4274_3_lut (.I0(\REG.mem_44_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n21), .I3(GND_net), .O(n5657));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4275_3_lut (.I0(\REG.mem_44_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n21), .I3(GND_net), .O(n5658));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4276_3_lut (.I0(\REG.mem_44_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n21), .I3(GND_net), .O(n5659));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4277_3_lut (.I0(\REG.mem_44_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n21), .I3(GND_net), .O(n5660));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3524_2_lut (.I0(n2352), .I1(DEBUG_8_c_0_c), .I2(GND_net), 
            .I3(GND_net), .O(n4907));   // src/usb3_if.v(88[8] 191[4])
    defparam i3524_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3526_2_lut (.I0(uart_rx_complete_prev), .I1(debug_led3), .I2(GND_net), 
            .I3(GND_net), .O(n4909));   // src/top.v(1065[8] 1071[4])
    defparam i3526_2_lut.LUT_INIT = 16'h4444;
    SB_DFF reset_all_r_77 (.Q(reset_all_w), .C(SLM_CLK_c), .D(reset_all_w_N_61));   // src/top.v(246[8] 264[4])
    SB_LUT4 i3527_2_lut (.I0(reset_per_frame_latched), .I1(n571), .I2(GND_net), 
            .I3(GND_net), .O(n4910));   // src/usb3_if.v(98[9] 189[16])
    defparam i3527_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3465_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [7]), .I3(fifo_data_out[7]), .O(n4848));
    defparam i3465_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3468_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [8]), .I3(fifo_data_out[8]), .O(n4851));
    defparam i3468_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4214_3_lut (.I0(\REG.mem_40_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n25), .I3(GND_net), .O(n5597));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4215_3_lut (.I0(\REG.mem_40_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n25), .I3(GND_net), .O(n5598));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4216_3_lut (.I0(\REG.mem_40_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n25), .I3(GND_net), .O(n5599));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4217_3_lut (.I0(\REG.mem_40_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n25), .I3(GND_net), .O(n5600));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4218_3_lut (.I0(\REG.mem_40_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n25), .I3(GND_net), .O(n5601));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4611_3_lut (.I0(\REG.mem_62_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n3), .I3(GND_net), .O(n5994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4219_3_lut (.I0(\REG.mem_40_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n25), .I3(GND_net), .O(n5602));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4220_3_lut (.I0(\REG.mem_41_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5603));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4221_3_lut (.I0(\REG.mem_41_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5604));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4222_3_lut (.I0(\REG.mem_41_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5605));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4223_3_lut (.I0(\REG.mem_41_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5606));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4235_3_lut (.I0(\REG.mem_41_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5618));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4224_3_lut (.I0(\REG.mem_41_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5607));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4225_3_lut (.I0(\REG.mem_41_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5608));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4226_3_lut (.I0(\REG.mem_41_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5609));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3471_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [9]), .I3(fifo_data_out[9]), .O(n4854));
    defparam i3471_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4227_3_lut (.I0(\REG.mem_41_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4236_3_lut (.I0(\REG.mem_42_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n23), .I3(GND_net), .O(n5619));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4237_3_lut (.I0(\REG.mem_42_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n23), .I3(GND_net), .O(n5620));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4612_3_lut (.I0(\REG.mem_62_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n3), .I3(GND_net), .O(n5995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4228_3_lut (.I0(\REG.mem_41_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5611));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3528_2_lut (.I0(reset_per_frame_latched), .I1(n575), .I2(GND_net), 
            .I3(GND_net), .O(n4911));   // src/usb3_if.v(98[9] 189[16])
    defparam i3528_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4238_3_lut (.I0(\REG.mem_42_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n23), .I3(GND_net), .O(n5621));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4229_3_lut (.I0(\REG.mem_41_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5612));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4230_3_lut (.I0(\REG.mem_41_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5613));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4239_3_lut (.I0(\REG.mem_42_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n23), .I3(GND_net), .O(n5622));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4240_3_lut (.I0(\REG.mem_42_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n23), .I3(GND_net), .O(n5623));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4231_3_lut (.I0(\REG.mem_41_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n24_adj_1225), .I3(GND_net), .O(n5614));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3475_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [10]), .I3(fifo_data_out[10]), .O(n4858));
    defparam i3475_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4241_3_lut (.I0(\REG.mem_42_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n23), .I3(GND_net), .O(n5624));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4242_3_lut (.I0(\REG.mem_42_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n23), .I3(GND_net), .O(n5625));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4613_3_lut (.I0(\REG.mem_62_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n3), .I3(GND_net), .O(n5996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4614_3_lut (.I0(\REG.mem_63_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n2), .I3(GND_net), .O(n5997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4243_3_lut (.I0(\REG.mem_42_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n23), .I3(GND_net), .O(n5626));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4244_3_lut (.I0(\REG.mem_42_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n23), .I3(GND_net), .O(n5627));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4615_3_lut (.I0(\REG.mem_63_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n2), .I3(GND_net), .O(n5998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4245_3_lut (.I0(\REG.mem_42_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n23), .I3(GND_net), .O(n5628));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4616_3_lut (.I0(\REG.mem_63_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n2), .I3(GND_net), .O(n5999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4617_3_lut (.I0(\REG.mem_63_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n2), .I3(GND_net), .O(n6000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(rd_addr_r_adj_1287[1]), .I1(rd_addr_r_adj_1287[0]), 
            .I2(wr_addr_r_adj_1284[1]), .I3(wr_addr_r_adj_1284[0]), .O(n32));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 i3481_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [11]), .I3(fifo_data_out[11]), .O(n4864));
    defparam i3481_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4618_3_lut (.I0(\REG.mem_63_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n2), .I3(GND_net), .O(n6001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4687_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [0]), .I3(fifo_data_out[0]), .O(n6070));
    defparam i4687_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3489_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [12]), .I3(fifo_data_out[12]), .O(n4872));
    defparam i3489_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i1_3_lut (.I0(is_fifo_empty_flag), .I1(fifo_write_cmd), .I2(n32), 
            .I3(GND_net), .O(n24));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i8857_4_lut (.I0(rd_addr_p1_w_adj_1289[2]), .I1(n13895), .I2(wr_addr_r_adj_1284[2]), 
            .I3(wr_addr_r_adj_1284[1]), .O(n10706));
    defparam i8857_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_73 (.I0(reset_all_w), .I1(n10706), .I2(n24), 
            .I3(n4), .O(n10632));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_73.LUT_INIT = 16'hfbfa;
    SB_LUT4 i4619_3_lut (.I0(\REG.mem_63_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n2), .I3(GND_net), .O(n6002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3492_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [13]), .I3(fifo_data_out[13]), .O(n4875));
    defparam i3492_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3510_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [14]), .I3(fifo_data_out[14]), .O(n4893));
    defparam i3510_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4620_3_lut (.I0(\REG.mem_63_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n2), .I3(GND_net), .O(n6003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4620_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_data_byte_r_i0_i7 (.Q(tx_data_byte[7]), .C(SLM_CLK_c), .D(n4945));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i4621_3_lut (.I0(\REG.mem_63_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n2), .I3(GND_net), .O(n6004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4622_3_lut (.I0(\REG.mem_63_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n2), .I3(GND_net), .O(n6005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4623_3_lut (.I0(\REG.mem_63_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n2), .I3(GND_net), .O(n6006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4278_3_lut (.I0(\REG.mem_44_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n21), .I3(GND_net), .O(n5661));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3513_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [15]), .I3(fifo_data_out[15]), .O(n4896));
    defparam i3513_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4280_3_lut (.I0(\REG.mem_44_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n21), .I3(GND_net), .O(n5663));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4624_3_lut (.I0(\REG.mem_63_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n2), .I3(GND_net), .O(n6007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4281_3_lut (.I0(\REG.mem_44_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n21), .I3(GND_net), .O(n5664));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4246_3_lut (.I0(\REG.mem_42_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n23), .I3(GND_net), .O(n5629));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4247_3_lut (.I0(\REG.mem_42_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n23), .I3(GND_net), .O(n5630));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4282_3_lut (.I0(\REG.mem_44_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n21), .I3(GND_net), .O(n5665));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4248_3_lut (.I0(\REG.mem_42_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n23), .I3(GND_net), .O(n5631));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4249_3_lut (.I0(\REG.mem_42_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n23), .I3(GND_net), .O(n5632));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3539_4_lut (.I0(RESET_c), .I1(rd_addr_r_adj_1287[2]), .I2(rd_addr_p1_w_adj_1289[2]), 
            .I3(empty_o_N_1149), .O(n4922));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i3539_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i4107_3_lut (.I0(\REG.mem_35_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n30), .I3(GND_net), .O(n5490));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4625_3_lut (.I0(\REG.mem_63_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n2), .I3(GND_net), .O(n6008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4284_3_lut (.I0(\REG.mem_44_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n21), .I3(GND_net), .O(n5667));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4250_3_lut (.I0(\REG.mem_42_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n23), .I3(GND_net), .O(n5633));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4108_3_lut (.I0(\REG.mem_35_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n30), .I3(GND_net), .O(n5491));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4626_3_lut (.I0(\REG.mem_63_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n2), .I3(GND_net), .O(n6009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4285_3_lut (.I0(\REG.mem_44_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n21), .I3(GND_net), .O(n5668));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4285_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF fifo_write_cmd_79 (.Q(fifo_write_cmd), .C(SLM_CLK_c), .D(n4942));   // src/top.v(889[8] 898[4])
    SB_LUT4 i4627_3_lut (.I0(\REG.mem_63_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n2), .I3(GND_net), .O(n6010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4628_3_lut (.I0(\REG.mem_63_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n2), .I3(GND_net), .O(n6011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4287_3_lut (.I0(\REG.mem_45_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n20), .I3(GND_net), .O(n5670));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4288_3_lut (.I0(\REG.mem_45_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n20), .I3(GND_net), .O(n5671));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4289_3_lut (.I0(\REG.mem_45_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n20), .I3(GND_net), .O(n5672));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4251_3_lut (.I0(\REG.mem_42_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n23), .I3(GND_net), .O(n5634));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4290_3_lut (.I0(\REG.mem_45_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n20), .I3(GND_net), .O(n5673));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4291_3_lut (.I0(\REG.mem_45_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n20), .I3(GND_net), .O(n5674));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4252_3_lut (.I0(\REG.mem_43_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n22), .I3(GND_net), .O(n5635));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4292_3_lut (.I0(\REG.mem_45_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n20), .I3(GND_net), .O(n5675));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4109_3_lut (.I0(\REG.mem_35_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n30), .I3(GND_net), .O(n5492));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4293_3_lut (.I0(\REG.mem_45_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n20), .I3(GND_net), .O(n5676));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4253_3_lut (.I0(\REG.mem_43_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n22), .I3(GND_net), .O(n5636));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4254_3_lut (.I0(\REG.mem_43_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n22), .I3(GND_net), .O(n5637));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4294_3_lut (.I0(\REG.mem_45_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n20), .I3(GND_net), .O(n5677));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4110_3_lut (.I0(\REG.mem_35_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n30), .I3(GND_net), .O(n5493));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4295_3_lut (.I0(\REG.mem_45_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n20), .I3(GND_net), .O(n5678));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4111_3_lut (.I0(\REG.mem_35_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n30), .I3(GND_net), .O(n5494));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4629_3_lut (.I0(\REG.mem_63_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n2), .I3(GND_net), .O(n6012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4255_3_lut (.I0(\REG.mem_43_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n22), .I3(GND_net), .O(n5638));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4112_3_lut (.I0(\REG.mem_35_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n30), .I3(GND_net), .O(n5495));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4113_3_lut (.I0(\REG.mem_35_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n30), .I3(GND_net), .O(n5496));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4256_3_lut (.I0(\REG.mem_43_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n22), .I3(GND_net), .O(n5639));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4296_3_lut (.I0(\REG.mem_45_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n20), .I3(GND_net), .O(n5679));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4296_3_lut.LUT_INIT = 16'hcaca;
    SB_IO CTS_pad (.PACKAGE_PIN(CTS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CTS_pad.PIN_TYPE = 6'b011001;
    defparam CTS_pad.PULLUP = 1'b0;
    defparam CTS_pad.NEG_TRIGGER = 1'b0;
    defparam CTS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4257_3_lut (.I0(\REG.mem_43_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n22), .I3(GND_net), .O(n5640));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4297_3_lut (.I0(\REG.mem_45_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n20), .I3(GND_net), .O(n5680));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4297_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DTR_pad (.PACKAGE_PIN(DTR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DTR_pad.PIN_TYPE = 6'b011001;
    defparam DTR_pad.PULLUP = 1'b0;
    defparam DTR_pad.NEG_TRIGGER = 1'b0;
    defparam DTR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4114_3_lut (.I0(\REG.mem_35_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n30), .I3(GND_net), .O(n5497));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4114_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DSR_pad (.PACKAGE_PIN(DSR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DSR_pad.PIN_TYPE = 6'b011001;
    defparam DSR_pad.PULLUP = 1'b0;
    defparam DSR_pad.NEG_TRIGGER = 1'b0;
    defparam DSR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4115_3_lut (.I0(\REG.mem_35_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n30), .I3(GND_net), .O(n5498));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4115_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DCD_pad (.PACKAGE_PIN(DCD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DCD_pad.PIN_TYPE = 6'b011001;
    defparam DCD_pad.PULLUP = 1'b0;
    defparam DCD_pad.NEG_TRIGGER = 1'b0;
    defparam DCD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4258_3_lut (.I0(\REG.mem_43_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n22), .I3(GND_net), .O(n5641));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4116_3_lut (.I0(\REG.mem_35_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n30), .I3(GND_net), .O(n5499));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4116_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DEBUG_8_c_0_pad (.PACKAGE_PIN(FIFO_D0), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(DEBUG_8_c_0_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_8_c_0_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_8_c_0_pad.PULLUP = 1'b0;
    defparam DEBUG_8_c_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_8_c_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4259_3_lut (.I0(\REG.mem_43_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n22), .I3(GND_net), .O(n5642));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4260_3_lut (.I0(\REG.mem_43_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n22), .I3(GND_net), .O(n5643));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4298_3_lut (.I0(\REG.mem_45_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n20), .I3(GND_net), .O(n5681));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4299_3_lut (.I0(\REG.mem_45_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n20), .I3(GND_net), .O(n5682));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4117_3_lut (.I0(\REG.mem_35_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n30), .I3(GND_net), .O(n5500));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4300_3_lut (.I0(\REG.mem_45_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n20), .I3(GND_net), .O(n5683));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4301_3_lut (.I0(\REG.mem_45_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n20), .I3(GND_net), .O(n5684));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4630_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[5]), .I2(GND_net), 
            .I3(GND_net), .O(n6013));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4630_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4261_3_lut (.I0(\REG.mem_43_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n22), .I3(GND_net), .O(n5644));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4118_3_lut (.I0(\REG.mem_35_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n30), .I3(GND_net), .O(n5501));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4302_3_lut (.I0(\REG.mem_45_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n20), .I3(GND_net), .O(n5685));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_74 (.I0(buffer_switch_done_latched), .I1(n843), 
            .I2(n771), .I3(GND_net), .O(n10149));
    defparam i1_3_lut_adj_74.LUT_INIT = 16'heaea;
    SB_LUT4 i4262_3_lut (.I0(\REG.mem_43_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n22), .I3(GND_net), .O(n5645));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4303_3_lut (.I0(\REG.mem_46_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n19), .I3(GND_net), .O(n5686));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4263_3_lut (.I0(\REG.mem_43_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n22), .I3(GND_net), .O(n5646));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4304_3_lut (.I0(\REG.mem_46_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n19), .I3(GND_net), .O(n5687));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4305_3_lut (.I0(\REG.mem_46_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n19), .I3(GND_net), .O(n5688));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4306_3_lut (.I0(\REG.mem_46_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n19), .I3(GND_net), .O(n5689));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4264_3_lut (.I0(\REG.mem_43_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n22), .I3(GND_net), .O(n5647));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4119_3_lut (.I0(\REG.mem_35_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n30), .I3(GND_net), .O(n5502));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4265_3_lut (.I0(\REG.mem_43_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n22), .I3(GND_net), .O(n5648));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4120_3_lut (.I0(\REG.mem_35_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n30), .I3(GND_net), .O(n5503));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4307_3_lut (.I0(\REG.mem_46_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n19), .I3(GND_net), .O(n5690));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4121_3_lut (.I0(\REG.mem_35_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n30), .I3(GND_net), .O(n5504));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4308_3_lut (.I0(\REG.mem_46_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n19), .I3(GND_net), .O(n5691));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4309_3_lut (.I0(\REG.mem_46_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n19), .I3(GND_net), .O(n5692));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4266_3_lut (.I0(\REG.mem_43_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n22), .I3(GND_net), .O(n5649));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4310_3_lut (.I0(\REG.mem_46_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n19), .I3(GND_net), .O(n5693));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4267_3_lut (.I0(\REG.mem_43_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n22), .I3(GND_net), .O(n5650));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4267_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i0 (.Q(n25_adj_1226), .C(SLM_CLK_c), .D(n130));   // src/top.v(203[20:35])
    SB_LUT4 i4311_3_lut (.I0(\REG.mem_46_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n19), .I3(GND_net), .O(n5694));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4268_3_lut (.I0(\REG.mem_44_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n21), .I3(GND_net), .O(n5651));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4312_3_lut (.I0(\REG.mem_46_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n19), .I3(GND_net), .O(n5695));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4122_3_lut (.I0(\REG.mem_35_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n30), .I3(GND_net), .O(n5505));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4313_3_lut (.I0(\REG.mem_46_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n19), .I3(GND_net), .O(n5696));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4314_3_lut (.I0(\REG.mem_46_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n19), .I3(GND_net), .O(n5697));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4125_3_lut (.I0(tx_data_byte[6]), .I1(pc_data_rx[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5508));   // src/top.v(1074[8] 1141[4])
    defparam i4125_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_1187__i3 (.Q(reset_clk_counter[3]), .C(SLM_CLK_c), 
           .D(n10165));   // src/top.v(259[27:51])
    SB_LUT4 i4126_3_lut (.I0(\REG.mem_36_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n29), .I3(GND_net), .O(n5509));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4315_3_lut (.I0(\REG.mem_46_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n19), .I3(GND_net), .O(n5698));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4316_3_lut (.I0(\REG.mem_46_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n19), .I3(GND_net), .O(n5699));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4317_3_lut (.I0(\REG.mem_46_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n19), .I3(GND_net), .O(n5700));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4127_3_lut (.I0(\REG.mem_36_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n29), .I3(GND_net), .O(n5510));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4128_3_lut (.I0(\REG.mem_36_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n29), .I3(GND_net), .O(n5511));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4129_3_lut (.I0(\REG.mem_36_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n29), .I3(GND_net), .O(n5512));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4130_3_lut (.I0(\REG.mem_36_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n29), .I3(GND_net), .O(n5513));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4318_3_lut (.I0(\REG.mem_46_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n19), .I3(GND_net), .O(n5701));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4319_3_lut (.I0(\REG.mem_47_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n18), .I3(GND_net), .O(n5702));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3540_3_lut (.I0(tx_addr_byte[0]), .I1(tx_data_byte[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4923));   // src/top.v(1074[8] 1141[4])
    defparam i3540_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_1187__i2 (.Q(reset_clk_counter[2]), .C(SLM_CLK_c), 
           .D(n10167));   // src/top.v(259[27:51])
    SB_DFF reset_clk_counter_i3_1187__i1 (.Q(reset_clk_counter[1]), .C(SLM_CLK_c), 
           .D(n10163));   // src/top.v(259[27:51])
    SB_DFF led_counter_1186_1260__i24 (.Q(DEBUG_0_c_24), .C(SLM_CLK_c), 
           .D(n106));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i23 (.Q(n2_adj_1241), .C(SLM_CLK_c), .D(n107));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i22 (.Q(n3_adj_1240), .C(SLM_CLK_c), .D(n108));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i21 (.Q(n4_adj_1239), .C(SLM_CLK_c), .D(n109));   // src/top.v(203[20:35])
    SB_LUT4 i4131_3_lut (.I0(\REG.mem_36_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n29), .I3(GND_net), .O(n5514));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4131_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i20 (.Q(n5), .C(SLM_CLK_c), .D(n110));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i19 (.Q(n6), .C(SLM_CLK_c), .D(n111));   // src/top.v(203[20:35])
    SB_LUT4 i4320_3_lut (.I0(\REG.mem_47_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n18), .I3(GND_net), .O(n5703));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4321_3_lut (.I0(\REG.mem_47_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n18), .I3(GND_net), .O(n5704));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4322_3_lut (.I0(\REG.mem_47_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n18), .I3(GND_net), .O(n5705));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4323_3_lut (.I0(\REG.mem_47_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n18), .I3(GND_net), .O(n5706));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4132_3_lut (.I0(\REG.mem_36_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n29), .I3(GND_net), .O(n5515));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4132_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i18 (.Q(n7), .C(SLM_CLK_c), .D(n112));   // src/top.v(203[20:35])
    SB_LUT4 i4324_3_lut (.I0(\REG.mem_47_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n18), .I3(GND_net), .O(n5707));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4324_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i17 (.Q(n8_adj_1238), .C(SLM_CLK_c), .D(n113));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i16 (.Q(n9), .C(SLM_CLK_c), .D(n114));   // src/top.v(203[20:35])
    SB_LUT4 i4325_3_lut (.I0(\REG.mem_47_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n18), .I3(GND_net), .O(n5708));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4325_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i15 (.Q(n10_adj_1237), .C(SLM_CLK_c), 
           .D(n115));   // src/top.v(203[20:35])
    SB_LUT4 i4133_3_lut (.I0(\REG.mem_36_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n29), .I3(GND_net), .O(n5516));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4133_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i14 (.Q(n11_adj_1236), .C(SLM_CLK_c), 
           .D(n116));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i13 (.Q(n12), .C(SLM_CLK_c), .D(n117));   // src/top.v(203[20:35])
    SB_LUT4 i4134_3_lut (.I0(\REG.mem_36_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n29), .I3(GND_net), .O(n5517));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4134_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i12 (.Q(n13), .C(SLM_CLK_c), .D(n118));   // src/top.v(203[20:35])
    SB_LUT4 i4135_3_lut (.I0(\REG.mem_36_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n29), .I3(GND_net), .O(n5518));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4135_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i11 (.Q(n14), .C(SLM_CLK_c), .D(n119));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i10 (.Q(n15_adj_1235), .C(SLM_CLK_c), 
           .D(n120));   // src/top.v(203[20:35])
    SB_LUT4 i4136_3_lut (.I0(\REG.mem_36_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n29), .I3(GND_net), .O(n5519));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4136_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i9 (.Q(n16), .C(SLM_CLK_c), .D(n121));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i8 (.Q(n17_adj_1234), .C(SLM_CLK_c), .D(n122));   // src/top.v(203[20:35])
    SB_LUT4 i4326_3_lut (.I0(\REG.mem_47_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n18), .I3(GND_net), .O(n5709));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4326_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i7 (.Q(n18_adj_1233), .C(SLM_CLK_c), .D(n123));   // src/top.v(203[20:35])
    SB_LUT4 i4137_3_lut (.I0(\REG.mem_36_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n29), .I3(GND_net), .O(n5520));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4137_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i6 (.Q(n19_adj_1232), .C(SLM_CLK_c), .D(n124));   // src/top.v(203[20:35])
    SB_LUT4 i4138_3_lut (.I0(\REG.mem_36_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n29), .I3(GND_net), .O(n5521));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4138_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i5 (.Q(n20_adj_1231), .C(SLM_CLK_c), .D(n125));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i4 (.Q(n21_adj_1230), .C(SLM_CLK_c), .D(n126));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i3 (.Q(n22_adj_1229), .C(SLM_CLK_c), .D(n127));   // src/top.v(203[20:35])
    SB_LUT4 i4327_3_lut (.I0(\REG.mem_47_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n18), .I3(GND_net), .O(n5710));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4328_3_lut (.I0(\REG.mem_47_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n18), .I3(GND_net), .O(n5711));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4328_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1186_1260_add_4_6 (.CI(n10047), .I0(GND_net), .I1(n21_adj_1230), 
            .CO(n10048));
    SB_LUT4 i4329_3_lut (.I0(\REG.mem_47_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n18), .I3(GND_net), .O(n5712));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4330_3_lut (.I0(\REG.mem_47_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n18), .I3(GND_net), .O(n5713));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4331_3_lut (.I0(\REG.mem_47_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n18), .I3(GND_net), .O(n5714));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4139_3_lut (.I0(\REG.mem_36_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n29), .I3(GND_net), .O(n5522));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4139_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1186_1260__i2 (.Q(n23_adj_1228), .C(SLM_CLK_c), .D(n128));   // src/top.v(203[20:35])
    SB_DFF led_counter_1186_1260__i1 (.Q(n24_adj_1227), .C(SLM_CLK_c), .D(n129));   // src/top.v(203[20:35])
    SB_LUT4 i4140_3_lut (.I0(\REG.mem_36_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n29), .I3(GND_net), .O(n5523));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4332_3_lut (.I0(\REG.mem_47_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n18), .I3(GND_net), .O(n5715));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4333_3_lut (.I0(\REG.mem_47_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n18), .I3(GND_net), .O(n5716));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4334_3_lut (.I0(\REG.mem_47_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n18), .I3(GND_net), .O(n5717));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4335_3_lut (.I0(\REG.mem_48_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n17), .I3(GND_net), .O(n5718));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4647_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[1]), .I2(n4_adj_1243), 
            .I3(n4253), .O(n6030));   // src/uart_rx.v(49[10] 144[8])
    defparam i4647_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4336_3_lut (.I0(\REG.mem_48_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n17), .I3(GND_net), .O(n5719));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4337_3_lut (.I0(\REG.mem_48_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n17), .I3(GND_net), .O(n5720));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4141_3_lut (.I0(\REG.mem_36_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n29), .I3(GND_net), .O(n5524));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4338_3_lut (.I0(\REG.mem_48_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n17), .I3(GND_net), .O(n5721));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4142_3_lut (.I0(tx_addr_byte[7]), .I1(tx_data_byte[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5525));   // src/top.v(1074[8] 1141[4])
    defparam i4142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4143_3_lut (.I0(tx_addr_byte[6]), .I1(tx_data_byte[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5526));   // src/top.v(1074[8] 1141[4])
    defparam i4143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4339_3_lut (.I0(\REG.mem_48_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n17), .I3(GND_net), .O(n5722));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4649_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[3]), .I2(GND_net), 
            .I3(GND_net), .O(n6032));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4649_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4340_3_lut (.I0(\REG.mem_48_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n17), .I3(GND_net), .O(n5723));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4341_3_lut (.I0(\REG.mem_48_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n17), .I3(GND_net), .O(n5724));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4342_3_lut (.I0(\REG.mem_48_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n17), .I3(GND_net), .O(n5725));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4343_3_lut (.I0(\REG.mem_48_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n17), .I3(GND_net), .O(n5726));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4344_3_lut (.I0(\REG.mem_48_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n17), .I3(GND_net), .O(n5727));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4345_3_lut (.I0(\REG.mem_48_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n17), .I3(GND_net), .O(n5728));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4346_3_lut (.I0(\REG.mem_48_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n17), .I3(GND_net), .O(n5729));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4144_3_lut (.I0(tx_addr_byte[5]), .I1(tx_data_byte[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5527));   // src/top.v(1074[8] 1141[4])
    defparam i4144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4347_3_lut (.I0(\REG.mem_48_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n17), .I3(GND_net), .O(n5730));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4145_3_lut (.I0(tx_addr_byte[4]), .I1(tx_data_byte[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5528));   // src/top.v(1074[8] 1141[4])
    defparam i4145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4146_3_lut (.I0(tx_addr_byte[3]), .I1(tx_data_byte[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5529));   // src/top.v(1074[8] 1141[4])
    defparam i4146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4147_3_lut (.I0(tx_addr_byte[2]), .I1(tx_data_byte[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5530));   // src/top.v(1074[8] 1141[4])
    defparam i4147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4651_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[1]), .I2(GND_net), 
            .I3(GND_net), .O(n6034));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4651_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4148_3_lut (.I0(tx_addr_byte[1]), .I1(tx_data_byte[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5531));   // src/top.v(1074[8] 1141[4])
    defparam i4148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4348_3_lut (.I0(\REG.mem_48_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n17), .I3(GND_net), .O(n5731));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4349_3_lut (.I0(\REG.mem_48_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n17), .I3(GND_net), .O(n5732));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4350_3_lut (.I0(\REG.mem_48_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n17), .I3(GND_net), .O(n5733));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4660_3_lut (.I0(rx_buf_byte[7]), .I1(rx_shift_reg[7]), .I2(n3495), 
            .I3(GND_net), .O(n6043));   // src/spi.v(76[8] 221[4])
    defparam i4660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4661_3_lut (.I0(rx_buf_byte[6]), .I1(rx_shift_reg[6]), .I2(n3495), 
            .I3(GND_net), .O(n6044));   // src/spi.v(76[8] 221[4])
    defparam i4661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 reset_all_w_I_0_1_lut (.I0(reset_all_w), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(RESET_c));   // src/top.v(295[16:28])
    defparam reset_all_w_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4662_3_lut (.I0(rx_buf_byte[5]), .I1(rx_shift_reg[5]), .I2(n3495), 
            .I3(GND_net), .O(n6045));   // src/spi.v(76[8] 221[4])
    defparam i4662_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4663_3_lut (.I0(rx_buf_byte[4]), .I1(rx_shift_reg[4]), .I2(n3495), 
            .I3(GND_net), .O(n6046));   // src/spi.v(76[8] 221[4])
    defparam i4663_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4155_3_lut (.I0(\REG.mem_37_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n28), .I3(GND_net), .O(n5538));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4664_3_lut (.I0(rx_buf_byte[3]), .I1(rx_shift_reg[3]), .I2(n3495), 
            .I3(GND_net), .O(n6047));   // src/spi.v(76[8] 221[4])
    defparam i4664_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4156_3_lut (.I0(\REG.mem_37_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n28), .I3(GND_net), .O(n5539));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4157_3_lut (.I0(\REG.mem_37_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n28), .I3(GND_net), .O(n5540));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4158_3_lut (.I0(\REG.mem_37_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n28), .I3(GND_net), .O(n5541));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4159_3_lut (.I0(\REG.mem_37_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n28), .I3(GND_net), .O(n5542));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4160_3_lut (.I0(\REG.mem_37_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n28), .I3(GND_net), .O(n5543));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4665_3_lut (.I0(rx_buf_byte[2]), .I1(rx_shift_reg[2]), .I2(n3495), 
            .I3(GND_net), .O(n6048));   // src/spi.v(76[8] 221[4])
    defparam i4665_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4161_3_lut (.I0(\REG.mem_37_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n28), .I3(GND_net), .O(n5544));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4162_3_lut (.I0(\REG.mem_37_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n28), .I3(GND_net), .O(n5545));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1186_1260_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_1229), .I3(n10046), .O(n127)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4163_3_lut (.I0(\REG.mem_37_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n28), .I3(GND_net), .O(n5546));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4666_3_lut (.I0(rx_buf_byte[1]), .I1(rx_shift_reg[1]), .I2(n3495), 
            .I3(GND_net), .O(n6049));   // src/spi.v(76[8] 221[4])
    defparam i4666_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4164_3_lut (.I0(\REG.mem_37_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n28), .I3(GND_net), .O(n5547));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4165_3_lut (.I0(\REG.mem_37_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n28), .I3(GND_net), .O(n5548));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4367_3_lut (.I0(\REG.mem_50_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5750));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3504_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[3]), .I2(\mem_LUT.data_raw_r [3]), 
            .I3(n4459), .O(n4887));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3504_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4677_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[2]), .I2(n4_adj_1220), 
            .I3(n4248), .O(n6060));   // src/uart_rx.v(49[10] 144[8])
    defparam i4677_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4371_3_lut (.I0(\REG.mem_50_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5754));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1655_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n3022));   // src/top.v(1074[8] 1141[4])
    defparam i1655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4372_3_lut (.I0(\REG.mem_50_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5755));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4679_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[3]), .I2(n4_adj_1220), 
            .I3(n4253), .O(n6062));   // src/uart_rx.v(49[10] 144[8])
    defparam i4679_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4680_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[4]), .I2(n4_adj_1244), 
            .I3(n4248), .O(n6063));   // src/uart_rx.v(49[10] 144[8])
    defparam i4680_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4681_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[5]), .I2(n4_adj_1244), 
            .I3(n4253), .O(n6064));   // src/uart_rx.v(49[10] 144[8])
    defparam i4681_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4373_3_lut (.I0(\REG.mem_50_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5756));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4373_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1186_1260_add_4_5 (.CI(n10046), .I0(GND_net), .I1(n22_adj_1229), 
            .CO(n10047));
    SB_LUT4 i4683_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[6]), .I2(n7347), 
            .I3(n4248), .O(n6066));   // src/uart_rx.v(49[10] 144[8])
    defparam i4683_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i4684_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[7]), .I2(n7347), 
            .I3(n4253), .O(n6067));   // src/uart_rx.v(49[10] 144[8])
    defparam i4684_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i4374_3_lut (.I0(\REG.mem_50_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5757));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4374_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF start_tx_81 (.Q(r_SM_Main_2__N_844[0]), .C(SLM_CLK_c), .D(n6098));   // src/top.v(910[8] 928[4])
    SB_LUT4 i4375_3_lut (.I0(\REG.mem_50_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5758));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4376_3_lut (.I0(\REG.mem_50_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5759));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4377_3_lut (.I0(\REG.mem_50_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5760));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4378_3_lut (.I0(\REG.mem_50_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5761));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4379_3_lut (.I0(\REG.mem_50_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4380_3_lut (.I0(\REG.mem_50_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5763));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4381_3_lut (.I0(\REG.mem_50_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5764));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4382_3_lut (.I0(\REG.mem_50_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5765));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4383_3_lut (.I0(\REG.mem_50_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4690_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[0]), .I2(\mem_LUT.data_raw_r [0]), 
            .I3(n4459), .O(n6073));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4690_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4384_3_lut (.I0(\REG.mem_50_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5767));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4384_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF spi_start_transfer_r_84 (.Q(spi_start_transfer_r), .C(SLM_CLK_c), 
           .D(n3022));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i4385_3_lut (.I0(\REG.mem_50_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n15_adj_1224), .I3(GND_net), .O(n5768));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4700_3_lut (.I0(pc_data_rx[0]), .I1(r_Rx_Data), .I2(n10211), 
            .I3(GND_net), .O(n6083));   // src/uart_rx.v(49[10] 144[8])
    defparam i4700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8863_4_lut (.I0(n1), .I1(fifo_read_cmd), .I2(wr_addr_r_adj_1284[1]), 
            .I3(rd_addr_r_adj_1287[1]), .O(n10712));
    defparam i8863_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i1_4_lut_adj_75 (.I0(reset_all_w), .I1(n15), .I2(wr_fifo_en_w), 
            .I3(n10098), .O(n10302));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_75.LUT_INIT = 16'h5444;
    SB_LUT4 i4166_3_lut (.I0(\REG.mem_37_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n28), .I3(GND_net), .O(n5549));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4167_3_lut (.I0(\REG.mem_37_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n28), .I3(GND_net), .O(n5550));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut (.I0(tx_shift_reg[0]), .I1(n2086), .I2(n4319), .I3(tx_data_byte[0]), 
            .O(n10300));   // src/spi.v(76[8] 221[4])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    GND i1 (.Y(GND_net));
    SB_LUT4 i4168_3_lut (.I0(\REG.mem_37_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n28), .I3(GND_net), .O(n5551));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4169_3_lut (.I0(\REG.mem_37_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n28), .I3(GND_net), .O(n5552));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10188_2_lut (.I0(is_fifo_empty_flag), .I1(tx_uart_active_flag), 
            .I2(GND_net), .I3(GND_net), .O(start_tx_N_64));
    defparam i10188_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 led_counter_1186_1260_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_1228), .I3(n10045), .O(n128)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8941_2_lut (.I0(n63), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n10790));
    defparam i8941_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19_4_lut (.I0(n4245), .I1(n11939), .I2(state[3]), .I3(n10790), 
            .O(n10384));   // src/timing_controller.v(53[8] 129[4])
    defparam i19_4_lut.LUT_INIT = 16'hfcac;
    SB_CARRY led_counter_1186_1260_add_4_4 (.CI(n10045), .I0(GND_net), .I1(n23_adj_1228), 
            .CO(n10046));
    SB_LUT4 i4729_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[1]), .I2(\mem_LUT.data_raw_r [1]), 
            .I3(n4459), .O(n6112));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4729_4_lut.LUT_INIT = 16'h5044;
    SB_DFF tx_data_byte_r_i0_i5 (.Q(tx_data_byte[5]), .C(SLM_CLK_c), .D(n5963));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 led_counter_1186_1260_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_1227), .I3(n10044), .O(n129)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_3 (.CI(n10044), .I0(GND_net), .I1(n24_adj_1227), 
            .CO(n10045));
    SB_LUT4 led_counter_1186_1260_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_1226), .I3(VCC_net), .O(n130)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 led_counter_1186_1260_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(DEBUG_0_c_24), .I3(n10067), .O(n106)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(n25_adj_1226), .CO(n10044));
    SB_LUT4 led_counter_1186_1260_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n2_adj_1241), .I3(n10066), .O(n107)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_25 (.CI(n10066), .I0(GND_net), 
            .I1(n2_adj_1241), .CO(n10067));
    SB_LUT4 led_counter_1186_1260_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_1240), .I3(n10065), .O(n108)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_24 (.CI(n10065), .I0(GND_net), 
            .I1(n3_adj_1240), .CO(n10066));
    SB_LUT4 led_counter_1186_1260_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_1239), .I3(n10064), .O(n109)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_23 (.CI(n10064), .I0(GND_net), 
            .I1(n4_adj_1239), .CO(n10065));
    SB_LUT4 led_counter_1186_1260_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5), .I3(n10063), .O(n110)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4170_3_lut (.I0(\REG.mem_37_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n28), .I3(GND_net), .O(n5553));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4170_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1186_1260_add_4_22 (.CI(n10063), .I0(GND_net), 
            .I1(n5), .CO(n10064));
    SB_LUT4 i4171_3_lut (.I0(\REG.mem_38_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n27), .I3(GND_net), .O(n5554));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1186_1260_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6), .I3(n10062), .O(n111)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4172_3_lut (.I0(\REG.mem_38_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n27), .I3(GND_net), .O(n5555));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4173_3_lut (.I0(\REG.mem_38_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n27), .I3(GND_net), .O(n5556));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4173_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1186_1260_add_4_21 (.CI(n10062), .I0(GND_net), 
            .I1(n6), .CO(n10063));
    SB_LUT4 i4174_3_lut (.I0(\REG.mem_38_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n27), .I3(GND_net), .O(n5557));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1186_1260_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7), .I3(n10061), .O(n112)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4175_3_lut (.I0(\REG.mem_38_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n27), .I3(GND_net), .O(n5558));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4175_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1186_1260_add_4_20 (.CI(n10061), .I0(GND_net), 
            .I1(n7), .CO(n10062));
    SB_LUT4 i4176_3_lut (.I0(\REG.mem_38_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n27), .I3(GND_net), .O(n5559));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1186_1260_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_1238), .I3(n10060), .O(n113)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_19 (.CI(n10060), .I0(GND_net), 
            .I1(n8_adj_1238), .CO(n10061));
    SB_LUT4 led_counter_1186_1260_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9), .I3(n10059), .O(n114)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_18 (.CI(n10059), .I0(GND_net), 
            .I1(n9), .CO(n10060));
    SB_LUT4 led_counter_1186_1260_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_1237), .I3(n10058), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_17 (.CI(n10058), .I0(GND_net), 
            .I1(n10_adj_1237), .CO(n10059));
    SB_LUT4 led_counter_1186_1260_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_1236), .I3(n10057), .O(n116)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_16 (.CI(n10057), .I0(GND_net), 
            .I1(n11_adj_1236), .CO(n10058));
    SB_LUT4 led_counter_1186_1260_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12), .I3(n10056), .O(n117)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_15 (.CI(n10056), .I0(GND_net), 
            .I1(n12), .CO(n10057));
    SB_LUT4 led_counter_1186_1260_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13), .I3(n10055), .O(n118)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1186_1260_add_4_14 (.CI(n10055), .I0(GND_net), 
            .I1(n13), .CO(n10056));
    SB_LUT4 led_counter_1186_1260_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14), .I3(n10054), .O(n119)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_76 (.I0(reset_clk_counter[3]), .I1(reset_clk_counter[2]), 
            .I2(n9936), .I3(GND_net), .O(n10165));
    defparam i1_3_lut_adj_76.LUT_INIT = 16'ha9a9;
    SB_CARRY led_counter_1186_1260_add_4_13 (.CI(n10054), .I0(GND_net), 
            .I1(n14), .CO(n10055));
    SB_LUT4 i4177_3_lut (.I0(\REG.mem_38_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n27), .I3(GND_net), .O(n5560));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4177_3_lut.LUT_INIT = 16'hcaca;
    SB_IO FIFO_D1_pad (.PACKAGE_PIN(FIFO_D1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D1_c_1));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D1_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D1_pad.PULLUP = 1'b0;
    defparam FIFO_D1_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D2_pad (.PACKAGE_PIN(FIFO_D2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D2_c_2));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D2_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D2_pad.PULLUP = 1'b0;
    defparam FIFO_D2_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D3_pad (.PACKAGE_PIN(FIFO_D3), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D3_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D3_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D3_pad.PULLUP = 1'b0;
    defparam FIFO_D3_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 led_counter_1186_1260_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_1235), .I3(n10053), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_IO FIFO_D4_pad (.PACKAGE_PIN(FIFO_D4), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D4_c_4));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D4_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D4_pad.PULLUP = 1'b0;
    defparam FIFO_D4_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D5_pad (.PACKAGE_PIN(FIFO_D5), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D5_c_5));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D5_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D5_pad.PULLUP = 1'b0;
    defparam FIFO_D5_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D6_pad (.PACKAGE_PIN(FIFO_D6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D6_c_6));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D6_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D6_pad.PULLUP = 1'b0;
    defparam FIFO_D6_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D7_pad (.PACKAGE_PIN(FIFO_D7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D7_c_7));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D7_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D7_pad.PULLUP = 1'b0;
    defparam FIFO_D7_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D8_pad (.PACKAGE_PIN(FIFO_D8), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D8_c_8));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D8_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D8_pad.PULLUP = 1'b0;
    defparam FIFO_D8_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D9_pad (.PACKAGE_PIN(FIFO_D9), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D9_c_9));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D9_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D9_pad.PULLUP = 1'b0;
    defparam FIFO_D9_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D10_pad (.PACKAGE_PIN(FIFO_D10), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D10_c_10));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D10_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D10_pad.PULLUP = 1'b0;
    defparam FIFO_D10_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D11_pad (.PACKAGE_PIN(FIFO_D11), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D11_c_11));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D11_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D11_pad.PULLUP = 1'b0;
    defparam FIFO_D11_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D12_pad (.PACKAGE_PIN(FIFO_D12), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D12_c_12));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D12_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D12_pad.PULLUP = 1'b0;
    defparam FIFO_D12_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D13_pad (.PACKAGE_PIN(FIFO_D13), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D13_c_13));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D13_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D13_pad.PULLUP = 1'b0;
    defparam FIFO_D13_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D14_pad (.PACKAGE_PIN(FIFO_D14), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D14_c_14));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D14_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D14_pad.PULLUP = 1'b0;
    defparam FIFO_D14_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D15_pad (.PACKAGE_PIN(FIFO_D15), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D15_c_15));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D15_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D15_pad.PULLUP = 1'b0;
    defparam FIFO_D15_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO FIFO_CLK_pad (.PACKAGE_PIN(FIFO_CLK), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(FIFO_CLK_c));   // src/top.v(84[12:20])
    defparam FIFO_CLK_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_CLK_pad.PULLUP = 1'b0;
    defparam FIFO_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_1_c_pad (.PACKAGE_PIN(FR_RXF), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(DEBUG_1_c_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_1_c_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_1_c_pad.PULLUP = 1'b0;
    defparam DEBUG_1_c_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_1_c_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SOUT_pad (.PACKAGE_PIN(SOUT), .OUTPUT_ENABLE(VCC_net), .D_IN_0(SOUT_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SOUT_pad.PIN_TYPE = 6'b000001;
    defparam SOUT_pad.PULLUP = 1'b0;
    defparam SOUT_pad.NEG_TRIGGER = 1'b0;
    defparam SOUT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UART_RX_pad (.PACKAGE_PIN(UART_RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(UART_RX_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_RX_pad.PIN_TYPE = 6'b000001;
    defparam UART_RX_pad.PULLUP = 1'b0;
    defparam UART_RX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_SYSCLK_pad (.PACKAGE_PIN(ICE_SYSCLK), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ICE_SYSCLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_SYSCLK_pad.PIN_TYPE = 6'b000001;
    defparam ICE_SYSCLK_pad.PULLUP = 1'b0;
    defparam ICE_SYSCLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_SYSCLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CREST_pad (.PACKAGE_PIN(ICE_CREST), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CREST_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CREST_pad.PULLUP = 1'b0;
    defparam ICE_CREST_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CREST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4178_3_lut (.I0(\REG.mem_38_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n27), .I3(GND_net), .O(n5561));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4178_3_lut.LUT_INIT = 16'hcaca;
    SB_IO ICE_CDONE_pad (.PACKAGE_PIN(ICE_CDONE), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CDONE_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CDONE_pad.PULLUP = 1'b0;
    defparam ICE_CDONE_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CDONE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CLK_pad (.PACKAGE_PIN(ICE_CLK), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CLK_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CLK_pad.PULLUP = 1'b0;
    defparam ICE_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_9_pad (.PACKAGE_PIN(DEBUG_9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_9_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_9_pad.PULLUP = 1'b0;
    defparam DEBUG_9_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_8_pad (.PACKAGE_PIN(DEBUG_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_8_c_0_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_8_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_8_pad.PULLUP = 1'b0;
    defparam DEBUG_8_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_6_pad (.PACKAGE_PIN(DEBUG_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_6_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_6_pad.PULLUP = 1'b0;
    defparam DEBUG_6_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_5_pad (.PACKAGE_PIN(DEBUG_5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_5_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_5_pad.PULLUP = 1'b0;
    defparam DEBUG_5_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_3_pad (.PACKAGE_PIN(DEBUG_3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_3_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_3_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_3_pad.PULLUP = 1'b0;
    defparam DEBUG_3_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_2_pad (.PACKAGE_PIN(DEBUG_2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_2_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_2_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_2_pad.PULLUP = 1'b0;
    defparam DEBUG_2_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_1_pad (.PACKAGE_PIN(DEBUG_1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_1_c_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_1_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_1_pad.PULLUP = 1'b0;
    defparam DEBUG_1_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_0_pad (.PACKAGE_PIN(DEBUG_0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_0_c_24));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_0_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_0_pad.PULLUP = 1'b0;
    defparam DEBUG_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_SIWU_pad (.PACKAGE_PIN(FT_SIWU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_SIWU_pad.PIN_TYPE = 6'b011001;
    defparam FT_SIWU_pad.PULLUP = 1'b0;
    defparam FT_SIWU_pad.NEG_TRIGGER = 1'b0;
    defparam FT_SIWU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_WR_pad (.PACKAGE_PIN(FT_WR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_WR_pad.PIN_TYPE = 6'b011001;
    defparam FT_WR_pad.PULLUP = 1'b0;
    defparam FT_WR_pad.NEG_TRIGGER = 1'b0;
    defparam FT_WR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_RD_pad (.PACKAGE_PIN(FT_RD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_2_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_RD_pad.PIN_TYPE = 6'b011001;
    defparam FT_RD_pad.PULLUP = 1'b0;
    defparam FT_RD_pad.NEG_TRIGGER = 1'b0;
    defparam FT_RD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_OE_pad (.PACKAGE_PIN(FT_OE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_OE_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_OE_pad.PIN_TYPE = 6'b011001;
    defparam FT_OE_pad.PULLUP = 1'b0;
    defparam FT_OE_pad.NEG_TRIGGER = 1'b0;
    defparam FT_OE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA10_pad (.PACKAGE_PIN(DATA10), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA10_c_10));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA10_pad.PIN_TYPE = 6'b011001;
    defparam DATA10_pad.PULLUP = 1'b0;
    defparam DATA10_pad.NEG_TRIGGER = 1'b0;
    defparam DATA10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA9_pad (.PACKAGE_PIN(DATA9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA9_c_9));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA9_pad.PIN_TYPE = 6'b011001;
    defparam DATA9_pad.PULLUP = 1'b0;
    defparam DATA9_pad.NEG_TRIGGER = 1'b0;
    defparam DATA9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA11_pad (.PACKAGE_PIN(DATA11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA11_c_11));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA11_pad.PIN_TYPE = 6'b011001;
    defparam DATA11_pad.PULLUP = 1'b0;
    defparam DATA11_pad.NEG_TRIGGER = 1'b0;
    defparam DATA11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA12_pad (.PACKAGE_PIN(DATA12), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA12_c_12));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA12_pad.PIN_TYPE = 6'b011001;
    defparam DATA12_pad.PULLUP = 1'b0;
    defparam DATA12_pad.NEG_TRIGGER = 1'b0;
    defparam DATA12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA13_pad (.PACKAGE_PIN(DATA13), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA13_c_13));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA13_pad.PIN_TYPE = 6'b011001;
    defparam DATA13_pad.PULLUP = 1'b0;
    defparam DATA13_pad.NEG_TRIGGER = 1'b0;
    defparam DATA13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA14_pad (.PACKAGE_PIN(DATA14), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA14_c_14));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA14_pad.PIN_TYPE = 6'b011001;
    defparam DATA14_pad.PULLUP = 1'b0;
    defparam DATA14_pad.NEG_TRIGGER = 1'b0;
    defparam DATA14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA8_pad (.PACKAGE_PIN(DATA8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA8_c_8));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA8_pad.PIN_TYPE = 6'b011001;
    defparam DATA8_pad.PULLUP = 1'b0;
    defparam DATA8_pad.NEG_TRIGGER = 1'b0;
    defparam DATA8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA15_pad (.PACKAGE_PIN(DATA15), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA15_c_15));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA15_pad.PIN_TYPE = 6'b011001;
    defparam DATA15_pad.PULLUP = 1'b0;
    defparam DATA15_pad.NEG_TRIGGER = 1'b0;
    defparam DATA15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA16_pad (.PACKAGE_PIN(DATA16), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA16_pad.PIN_TYPE = 6'b011001;
    defparam DATA16_pad.PULLUP = 1'b0;
    defparam DATA16_pad.NEG_TRIGGER = 1'b0;
    defparam DATA16_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA7_pad (.PACKAGE_PIN(DATA7), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA7_c_7));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA7_pad.PIN_TYPE = 6'b011001;
    defparam DATA7_pad.PULLUP = 1'b0;
    defparam DATA7_pad.NEG_TRIGGER = 1'b0;
    defparam DATA7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA17_pad (.PACKAGE_PIN(DATA17), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA17_pad.PIN_TYPE = 6'b011001;
    defparam DATA17_pad.PULLUP = 1'b0;
    defparam DATA17_pad.NEG_TRIGGER = 1'b0;
    defparam DATA17_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA18_pad (.PACKAGE_PIN(DATA18), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA18_pad.PIN_TYPE = 6'b011001;
    defparam DATA18_pad.PULLUP = 1'b0;
    defparam DATA18_pad.NEG_TRIGGER = 1'b0;
    defparam DATA18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA6_pad (.PACKAGE_PIN(DATA6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA6_c_6));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA6_pad.PIN_TYPE = 6'b011001;
    defparam DATA6_pad.PULLUP = 1'b0;
    defparam DATA6_pad.NEG_TRIGGER = 1'b0;
    defparam DATA6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA19_pad (.PACKAGE_PIN(DATA19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA19_pad.PIN_TYPE = 6'b011001;
    defparam DATA19_pad.PULLUP = 1'b0;
    defparam DATA19_pad.NEG_TRIGGER = 1'b0;
    defparam DATA19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA20_pad (.PACKAGE_PIN(DATA20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA20_pad.PIN_TYPE = 6'b011001;
    defparam DATA20_pad.PULLUP = 1'b0;
    defparam DATA20_pad.NEG_TRIGGER = 1'b0;
    defparam DATA20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA5_pad (.PACKAGE_PIN(DATA5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA5_c_5));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA5_pad.PIN_TYPE = 6'b011001;
    defparam DATA5_pad.PULLUP = 1'b0;
    defparam DATA5_pad.NEG_TRIGGER = 1'b0;
    defparam DATA5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA21_pad (.PACKAGE_PIN(DATA21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA21_pad.PIN_TYPE = 6'b011001;
    defparam DATA21_pad.PULLUP = 1'b0;
    defparam DATA21_pad.NEG_TRIGGER = 1'b0;
    defparam DATA21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA22_pad (.PACKAGE_PIN(DATA22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA22_pad.PIN_TYPE = 6'b011001;
    defparam DATA22_pad.PULLUP = 1'b0;
    defparam DATA22_pad.NEG_TRIGGER = 1'b0;
    defparam DATA22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA4_pad (.PACKAGE_PIN(DATA4), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA4_c_4));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA4_pad.PIN_TYPE = 6'b011001;
    defparam DATA4_pad.PULLUP = 1'b0;
    defparam DATA4_pad.NEG_TRIGGER = 1'b0;
    defparam DATA4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA23_pad (.PACKAGE_PIN(DATA23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA23_pad.PIN_TYPE = 6'b011001;
    defparam DATA23_pad.PULLUP = 1'b0;
    defparam DATA23_pad.NEG_TRIGGER = 1'b0;
    defparam DATA23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA24_pad (.PACKAGE_PIN(DATA24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA24_pad.PIN_TYPE = 6'b011001;
    defparam DATA24_pad.PULLUP = 1'b0;
    defparam DATA24_pad.NEG_TRIGGER = 1'b0;
    defparam DATA24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA3_pad (.PACKAGE_PIN(DATA3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA3_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA3_pad.PIN_TYPE = 6'b011001;
    defparam DATA3_pad.PULLUP = 1'b0;
    defparam DATA3_pad.NEG_TRIGGER = 1'b0;
    defparam DATA3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_1186_1260_add_4_12 (.CI(n10053), .I0(GND_net), 
            .I1(n15_adj_1235), .CO(n10054));
    SB_IO DATA25_pad (.PACKAGE_PIN(DATA25), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA25_pad.PIN_TYPE = 6'b011001;
    defparam DATA25_pad.PULLUP = 1'b0;
    defparam DATA25_pad.NEG_TRIGGER = 1'b0;
    defparam DATA25_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA26_pad (.PACKAGE_PIN(DATA26), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA26_pad.PIN_TYPE = 6'b011001;
    defparam DATA26_pad.PULLUP = 1'b0;
    defparam DATA26_pad.NEG_TRIGGER = 1'b0;
    defparam DATA26_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA2_pad (.PACKAGE_PIN(DATA2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA2_c_2));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA2_pad.PIN_TYPE = 6'b011001;
    defparam DATA2_pad.PULLUP = 1'b0;
    defparam DATA2_pad.NEG_TRIGGER = 1'b0;
    defparam DATA2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA27_pad (.PACKAGE_PIN(DATA27), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA27_pad.PIN_TYPE = 6'b011001;
    defparam DATA27_pad.PULLUP = 1'b0;
    defparam DATA27_pad.NEG_TRIGGER = 1'b0;
    defparam DATA27_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA28_pad (.PACKAGE_PIN(DATA28), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA28_pad.PIN_TYPE = 6'b011001;
    defparam DATA28_pad.PULLUP = 1'b0;
    defparam DATA28_pad.NEG_TRIGGER = 1'b0;
    defparam DATA28_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA1_pad (.PACKAGE_PIN(DATA1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA1_c_1));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA1_pad.PIN_TYPE = 6'b011001;
    defparam DATA1_pad.PULLUP = 1'b0;
    defparam DATA1_pad.NEG_TRIGGER = 1'b0;
    defparam DATA1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA29_pad (.PACKAGE_PIN(DATA29), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA29_pad.PIN_TYPE = 6'b011001;
    defparam DATA29_pad.PULLUP = 1'b0;
    defparam DATA29_pad.NEG_TRIGGER = 1'b0;
    defparam DATA29_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA30_pad (.PACKAGE_PIN(DATA30), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA30_pad.PIN_TYPE = 6'b011001;
    defparam DATA30_pad.PULLUP = 1'b0;
    defparam DATA30_pad.NEG_TRIGGER = 1'b0;
    defparam DATA30_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA0_pad (.PACKAGE_PIN(DATA0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA0_pad.PIN_TYPE = 6'b011001;
    defparam DATA0_pad.PULLUP = 1'b0;
    defparam DATA0_pad.NEG_TRIGGER = 1'b0;
    defparam DATA0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 led_counter_1186_1260_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16), .I3(n10052), .O(n121)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_IO DATA31_pad (.PACKAGE_PIN(DATA31), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA31_pad.PIN_TYPE = 6'b011001;
    defparam DATA31_pad.PULLUP = 1'b0;
    defparam DATA31_pad.NEG_TRIGGER = 1'b0;
    defparam DATA31_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO VALID_pad (.PACKAGE_PIN(VALID), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam VALID_pad.PIN_TYPE = 6'b011001;
    defparam VALID_pad.PULLUP = 1'b0;
    defparam VALID_pad.NEG_TRIGGER = 1'b0;
    defparam VALID_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SYNC_pad (.PACKAGE_PIN(SYNC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SYNC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SYNC_pad.PIN_TYPE = 6'b011001;
    defparam SYNC_pad.PULLUP = 1'b0;
    defparam SYNC_pad.NEG_TRIGGER = 1'b0;
    defparam SYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INVERT_pad (.PACKAGE_PIN(INVERT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INVERT_c_3)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INVERT_pad.PIN_TYPE = 6'b011001;
    defparam INVERT_pad.PULLUP = 1'b0;
    defparam INVERT_pad.NEG_TRIGGER = 1'b0;
    defparam INVERT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SLM_CLK_pad (.PACKAGE_PIN(SLM_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SLM_CLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SLM_CLK_pad.PIN_TYPE = 6'b011001;
    defparam SLM_CLK_pad.PULLUP = 1'b0;
    defparam SLM_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam SLM_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO RESET_pad (.PACKAGE_PIN(RESET), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(RESET_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RESET_pad.PIN_TYPE = 6'b011001;
    defparam RESET_pad.PULLUP = 1'b0;
    defparam RESET_pad.NEG_TRIGGER = 1'b0;
    defparam RESET_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UPDATE_pad (.PACKAGE_PIN(UPDATE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UPDATE_c_2));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UPDATE_pad.PIN_TYPE = 6'b011001;
    defparam UPDATE_pad.PULLUP = 1'b0;
    defparam UPDATE_pad.NEG_TRIGGER = 1'b0;
    defparam UPDATE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SDAT_pad (.PACKAGE_PIN(SDAT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SDAT_c_15)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SDAT_pad.PIN_TYPE = 6'b011001;
    defparam SDAT_pad.PULLUP = 1'b0;
    defparam SDAT_pad.NEG_TRIGGER = 1'b0;
    defparam SDAT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SCK_pad (.PACKAGE_PIN(SCK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SCK_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SCK_pad.PIN_TYPE = 6'b011001;
    defparam SCK_pad.PULLUP = 1'b0;
    defparam SCK_pad.NEG_TRIGGER = 1'b0;
    defparam SCK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SEN_pad (.PACKAGE_PIN(SEN), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SEN_c_1)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SEN_pad.PIN_TYPE = 6'b011001;
    defparam SEN_pad.PULLUP = 1'b0;
    defparam SEN_pad.NEG_TRIGGER = 1'b0;
    defparam SEN_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UART_TX_pad (.PACKAGE_PIN(UART_TX), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UART_TX_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_TX_pad.PIN_TYPE = 6'b011001;
    defparam UART_TX_pad.PULLUP = 1'b0;
    defparam UART_TX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_TX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4179_3_lut (.I0(\REG.mem_38_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n27), .I3(GND_net), .O(n5562));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4180_3_lut (.I0(\REG.mem_38_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n27), .I3(GND_net), .O(n5563));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4181_3_lut (.I0(\REG.mem_38_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n27), .I3(GND_net), .O(n5564));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4182_3_lut (.I0(\REG.mem_38_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n27), .I3(GND_net), .O(n5565));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4182_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_addr_byte_r_i0_i0 (.Q(tx_addr_byte[0]), .C(SLM_CLK_c), .D(n4923));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i4183_3_lut (.I0(\REG.mem_38_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n27), .I3(GND_net), .O(n5566));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4184_3_lut (.I0(\REG.mem_38_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n27), .I3(GND_net), .O(n5567));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4185_3_lut (.I0(\REG.mem_38_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n27), .I3(GND_net), .O(n5568));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4186_3_lut (.I0(\REG.mem_38_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n27), .I3(GND_net), .O(n5569));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4187_3_lut (.I0(\REG.mem_39_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n26), .I3(GND_net), .O(n5570));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4189_3_lut (.I0(\REG.mem_39_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n26), .I3(GND_net), .O(n5572));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4190_3_lut (.I0(\REG.mem_39_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n26), .I3(GND_net), .O(n5573));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4191_3_lut (.I0(\REG.mem_39_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n26), .I3(GND_net), .O(n5574));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4192_3_lut (.I0(\REG.mem_39_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n26), .I3(GND_net), .O(n5575));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4193_3_lut (.I0(\REG.mem_39_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n26), .I3(GND_net), .O(n5576));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4194_3_lut (.I0(\REG.mem_39_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n26), .I3(GND_net), .O(n5577));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4195_3_lut (.I0(\REG.mem_39_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n26), .I3(GND_net), .O(n5578));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4196_3_lut (.I0(\REG.mem_39_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n26), .I3(GND_net), .O(n5579));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4197_3_lut (.I0(\REG.mem_39_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n26), .I3(GND_net), .O(n5580));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3514_3_lut (.I0(rx_buf_byte[0]), .I1(rx_shift_reg[0]), .I2(n3495), 
            .I3(GND_net), .O(n4897));   // src/spi.v(76[8] 221[4])
    defparam i3514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3515_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4898));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i3515_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4198_3_lut (.I0(\REG.mem_39_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n26), .I3(GND_net), .O(n5581));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4199_3_lut (.I0(\REG.mem_39_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n26), .I3(GND_net), .O(n5582));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4200_3_lut (.I0(\REG.mem_39_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n26), .I3(GND_net), .O(n5583));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4201_3_lut (.I0(\REG.mem_39_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n26), .I3(GND_net), .O(n5584));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4201_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1186_1260_add_4_11 (.CI(n10052), .I0(GND_net), 
            .I1(n16), .CO(n10053));
    SB_LUT4 led_counter_1186_1260_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_1234), .I3(n10051), .O(n122)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4434_3_lut (.I0(\REG.mem_54_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n11), .I3(GND_net), .O(n5817));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4434_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1186_1260_add_4_10 (.CI(n10051), .I0(GND_net), 
            .I1(n17_adj_1234), .CO(n10052));
    SB_LUT4 led_counter_1186_1260_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_1233), .I3(n10050), .O(n123)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4435_3_lut (.I0(\REG.mem_54_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n11), .I3(GND_net), .O(n5818));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4436_3_lut (.I0(\REG.mem_54_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n11), .I3(GND_net), .O(n5819));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4436_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF uart_rx_complete_rising_edge_82 (.Q(uart_rx_complete_rising_edge), 
           .C(SLM_CLK_c), .D(n4909));   // src/top.v(1065[8] 1071[4])
    SB_LUT4 i4437_3_lut (.I0(\REG.mem_54_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n11), .I3(GND_net), .O(n5820));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3559_2_lut (.I0(is_tx_fifo_full_flag), .I1(spi_rx_byte_ready), 
            .I2(GND_net), .I3(GND_net), .O(n4942));   // src/top.v(889[8] 898[4])
    defparam i3559_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY led_counter_1186_1260_add_4_9 (.CI(n10050), .I0(GND_net), .I1(n18_adj_1233), 
            .CO(n10051));
    SB_LUT4 i4438_3_lut (.I0(\REG.mem_54_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n11), .I3(GND_net), .O(n5821));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4439_3_lut (.I0(\REG.mem_54_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n11), .I3(GND_net), .O(n5822));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4440_3_lut (.I0(\REG.mem_54_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n11), .I3(GND_net), .O(n5823));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4441_3_lut (.I0(\REG.mem_54_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n11), .I3(GND_net), .O(n5824));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4442_3_lut (.I0(\REG.mem_54_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n11), .I3(GND_net), .O(n5825));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4442_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_addr_byte_r_i0_i1 (.Q(tx_addr_byte[1]), .C(SLM_CLK_c), .D(n5531));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_addr_byte_r_i0_i2 (.Q(tx_addr_byte[2]), .C(SLM_CLK_c), .D(n5530));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_addr_byte_r_i0_i3 (.Q(tx_addr_byte[3]), .C(SLM_CLK_c), .D(n5529));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_addr_byte_r_i0_i4 (.Q(tx_addr_byte[4]), .C(SLM_CLK_c), .D(n5528));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_addr_byte_r_i0_i5 (.Q(tx_addr_byte[5]), .C(SLM_CLK_c), .D(n5527));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_addr_byte_r_i0_i6 (.Q(tx_addr_byte[6]), .C(SLM_CLK_c), .D(n5526));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_addr_byte_r_i0_i7 (.Q(tx_addr_byte[7]), .C(SLM_CLK_c), .D(n5525));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 led_counter_1186_1260_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_1232), .I3(n10049), .O(n124)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF tx_data_byte_r_i0_i6 (.Q(tx_data_byte[6]), .C(SLM_CLK_c), .D(n5508));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i4443_3_lut (.I0(\REG.mem_54_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n11), .I3(GND_net), .O(n5826));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4444_3_lut (.I0(\REG.mem_54_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n11), .I3(GND_net), .O(n5827));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4445_3_lut (.I0(\REG.mem_54_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n11), .I3(GND_net), .O(n5828));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4446_3_lut (.I0(\REG.mem_54_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n11), .I3(GND_net), .O(n5829));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4447_3_lut (.I0(\REG.mem_54_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n11), .I3(GND_net), .O(n5830));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4448_3_lut (.I0(\REG.mem_54_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n11), .I3(GND_net), .O(n5831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i954_4_lut (.I0(n2034), .I1(n7440), .I2(state[3]), .I3(n63), 
            .O(n1879));   // src/timing_controller.v(48[11:16])
    defparam i954_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i3181_4_lut (.I0(n63), .I1(n4192), .I2(n7440), .I3(state[3]), 
            .O(n1774));   // src/timing_controller.v(48[11:16])
    defparam i3181_4_lut.LUT_INIT = 16'h0a88;
    SB_LUT4 i4449_3_lut (.I0(\REG.mem_54_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n11), .I3(GND_net), .O(n5832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4450_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n5833));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4450_2_lut.LUT_INIT = 16'h4444;
    SB_DFF reset_clk_counter_i3_1187__i0 (.Q(reset_clk_counter[0]), .C(SLM_CLK_c), 
           .D(n25_adj_1242));   // src/top.v(259[27:51])
    SB_LUT4 i4451_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5834));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4451_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4452_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5835));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4452_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4453_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5836));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4453_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4202_3_lut (.I0(\REG.mem_39_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n26), .I3(GND_net), .O(n5585));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3499_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[2]), .I2(\mem_LUT.data_raw_r [2]), 
            .I3(n4459), .O(n4882));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3499_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4455_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5838));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4455_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4456_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5839));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4456_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4457_3_lut (.I0(\REG.mem_55_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n10), .I3(GND_net), .O(n5840));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4458_3_lut (.I0(\REG.mem_55_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n10), .I3(GND_net), .O(n5841));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4459_3_lut (.I0(\REG.mem_55_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n10), .I3(GND_net), .O(n5842));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4460_3_lut (.I0(\REG.mem_55_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n10), .I3(GND_net), .O(n5843));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4461_3_lut (.I0(\REG.mem_55_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n10), .I3(GND_net), .O(n5844));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4203_3_lut (.I0(\REG.mem_39_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n26), .I3(GND_net), .O(n5586));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3562_3_lut (.I0(tx_data_byte[7]), .I1(pc_data_rx[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4945));   // src/top.v(1074[8] 1141[4])
    defparam i3562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4204_3_lut (.I0(\REG.mem_40_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n25), .I3(GND_net), .O(n5587));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4205_3_lut (.I0(\REG.mem_40_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n25), .I3(GND_net), .O(n5588));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4462_3_lut (.I0(\REG.mem_55_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n10), .I3(GND_net), .O(n5845));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4206_3_lut (.I0(\REG.mem_40_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n25), .I3(GND_net), .O(n5589));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4463_3_lut (.I0(\REG.mem_55_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n10), .I3(GND_net), .O(n5846));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4464_3_lut (.I0(\REG.mem_55_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n10), .I3(GND_net), .O(n5847));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4465_3_lut (.I0(\REG.mem_55_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n10), .I3(GND_net), .O(n5848));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4466_3_lut (.I0(\REG.mem_55_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n10), .I3(GND_net), .O(n5849));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4467_3_lut (.I0(\REG.mem_55_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n10), .I3(GND_net), .O(n5850));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4468_3_lut (.I0(\REG.mem_55_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n10), .I3(GND_net), .O(n5851));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4469_3_lut (.I0(\REG.mem_55_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n10), .I3(GND_net), .O(n5852));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5882_1_lut (.I0(n1774), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n7258));   // src/timing_controller.v(48[11:16])
    defparam i5882_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4470_3_lut (.I0(\REG.mem_55_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n10), .I3(GND_net), .O(n5853));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4471_3_lut (.I0(\REG.mem_55_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n10), .I3(GND_net), .O(n5854));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4472_3_lut (.I0(\REG.mem_55_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n10), .I3(GND_net), .O(n5855));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4473_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n5856));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4473_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4474_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5857));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4474_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4475_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5858));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4475_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4476_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5859));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4476_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4477_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5860));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4477_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4478_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5861));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4478_2_lut.LUT_INIT = 16'h4444;
    SB_DFF even_byte_flag_89 (.Q(even_byte_flag), .C(SLM_CLK_c), .D(n2944));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i4496_3_lut (.I0(\REG.mem_57_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4497_3_lut (.I0(\REG.mem_57_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5880));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4498_3_lut (.I0(\REG.mem_57_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5881));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4499_3_lut (.I0(\REG.mem_57_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5882));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4500_3_lut (.I0(\REG.mem_57_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5883));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4501_3_lut (.I0(\REG.mem_57_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4502_3_lut (.I0(\REG.mem_57_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5885));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4503_3_lut (.I0(\REG.mem_57_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5886));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4503_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1186_1260_add_4_8 (.CI(n10049), .I0(GND_net), .I1(n19_adj_1232), 
            .CO(n10050));
    SB_LUT4 i4504_3_lut (.I0(\REG.mem_57_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5887));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4505_3_lut (.I0(\REG.mem_57_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5888));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4506_3_lut (.I0(\REG.mem_57_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5889));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4507_3_lut (.I0(\REG.mem_57_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5890));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4508_3_lut (.I0(\REG.mem_57_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5891));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4509_3_lut (.I0(\REG.mem_57_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5892));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4510_3_lut (.I0(\REG.mem_57_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5893));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4511_3_lut (.I0(\REG.mem_57_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n8_adj_1223), .I3(GND_net), .O(n5894));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3930_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[5]), .I2(\mem_LUT.data_raw_r [5]), 
            .I3(n4459), .O(n5313));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3930_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i3927_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[4]), .I2(\mem_LUT.data_raw_r [4]), 
            .I3(n4459), .O(n5310));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3927_4_lut.LUT_INIT = 16'h5044;
    SB_DFFSR multi_byte_spi_trans_flag_r_86 (.Q(multi_byte_spi_trans_flag_r), 
            .C(SLM_CLK_c), .D(multi_byte_spi_trans_flag_r_N_72), .R(n4676));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_data_byte_r_i0_i1 (.Q(tx_data_byte[1]), .C(SLM_CLK_c), .D(n4860));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_data_byte_r_i0_i2 (.Q(tx_data_byte[2]), .C(SLM_CLK_c), .D(n4859));   // src/top.v(1074[8] 1141[4])
    SB_DFF tx_data_byte_r_i0_i3 (.Q(tx_data_byte[3]), .C(SLM_CLK_c), .D(n4855));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i4531_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_6__N_498[5]), 
            .I2(GND_net), .I3(GND_net), .O(n5914));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i4531_2_lut.LUT_INIT = 16'h4444;
    SB_DFF tx_data_byte_r_i0_i4 (.Q(tx_data_byte[4]), .C(SLM_CLK_c), .D(n4845));   // src/top.v(1074[8] 1141[4])
    SB_LUT4 i4533_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_6__N_498[3]), 
            .I2(GND_net), .I3(GND_net), .O(n5916));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i4533_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4534_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_6__N_498[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5917));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i4534_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4536_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n5919));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4536_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4537_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5920));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4537_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4538_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5921));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4538_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4555_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5938));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4555_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4556_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5939));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4556_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4557_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5940));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4557_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4558_2_lut (.I0(reset_per_frame), .I1(rd_addr_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n5941));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4558_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4559_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5942));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4559_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4560_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5943));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4560_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4561_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5944));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4561_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4562_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5945));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4562_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4563_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5946));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4563_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3555_4_lut_4_lut_4_lut (.I0(wr_fifo_en_w), .I1(reset_all_w), 
            .I2(wr_addr_r_adj_1284[0]), .I3(wr_addr_r_adj_1284[1]), .O(n4938));
    defparam i3555_4_lut_4_lut_4_lut.LUT_INIT = 16'h1320;
    SB_LUT4 i3558_4_lut_4_lut (.I0(wr_fifo_en_w), .I1(reset_all_w), .I2(wr_addr_p1_w_adj_1286[2]), 
            .I3(wr_addr_r_adj_1284[2]), .O(n4941));
    defparam i3558_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4580_3_lut (.I0(tx_data_byte[5]), .I1(pc_data_rx[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5963));   // src/top.v(1074[8] 1141[4])
    defparam i4580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[3]), 
            .I3(n10790), .O(n10662));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i3_4_lut (.I0(reset_clk_counter[0]), .I1(reset_clk_counter[2]), 
            .I2(reset_clk_counter[3]), .I3(reset_clk_counter[1]), .O(reset_all_w_N_61));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 led_counter_1186_1260_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_1231), .I3(n10048), .O(n125)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10160_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(n10681), .O(n11939));
    defparam i10160_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i6086_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(n63), 
            .I3(GND_net), .O(n7462));
    defparam i6086_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_DFF tx_data_byte_r_i0_i0 (.Q(tx_data_byte[0]), .C(SLM_CLK_c), .D(n4824));   // src/top.v(1074[8] 1141[4])
    SB_CARRY led_counter_1186_1260_add_4_7 (.CI(n10048), .I0(GND_net), .I1(n20_adj_1231), 
            .CO(n10049));
    SB_LUT4 led_counter_1186_1260_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_1230), .I3(n10047), .O(n126)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1186_1260_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF fifo_read_cmd_80 (.Q(fifo_read_cmd), .C(SLM_CLK_c), .D(start_tx_N_64));   // src/top.v(910[8] 928[4])
    SB_LUT4 i4598_3_lut (.I0(\REG.mem_62_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n3), .I3(GND_net), .O(n5981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4599_3_lut (.I0(\REG.mem_62_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n3), .I3(GND_net), .O(n5982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4600_3_lut (.I0(\REG.mem_62_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n3), .I3(GND_net), .O(n5983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4601_3_lut (.I0(\REG.mem_62_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n3), .I3(GND_net), .O(n5984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4602_3_lut (.I0(\REG.mem_62_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n3), .I3(GND_net), .O(n5985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4603_3_lut (.I0(\REG.mem_62_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n3), .I3(GND_net), .O(n5986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4269_3_lut (.I0(\REG.mem_44_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n21), .I3(GND_net), .O(n5652));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4604_3_lut (.I0(\REG.mem_62_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n3), .I3(GND_net), .O(n5987));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8227_2_lut_3_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(reset_clk_counter[1]), .I3(GND_net), .O(n9936));   // src/top.v(259[27:51])
    defparam i8227_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i4605_3_lut (.I0(\REG.mem_62_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n3), .I3(GND_net), .O(n5988));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4606_3_lut (.I0(\REG.mem_62_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n3), .I3(GND_net), .O(n5989));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3507_3_lut (.I0(r_Tx_Data[0]), .I1(fifo_temp_output[0]), .I2(n3794), 
            .I3(GND_net), .O(n4890));   // src/uart_tx.v(38[10] 141[8])
    defparam i3507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3505_3_lut (.I0(rx_shift_reg[1]), .I1(rx_shift_reg[0]), .I2(n4312), 
            .I3(GND_net), .O(n4888));   // src/spi.v(76[8] 221[4])
    defparam i3505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4057_3_lut (.I0(\REG.mem_31_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n34), .I3(GND_net), .O(n5440));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(reset_clk_counter[1]), .I3(GND_net), .O(n10163));   // src/top.v(259[27:51])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i4056_3_lut (.I0(\REG.mem_31_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n34), .I3(GND_net), .O(n5439));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4055_3_lut (.I0(\REG.mem_31_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n34), .I3(GND_net), .O(n5438));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4054_3_lut (.I0(\REG.mem_31_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n34), .I3(GND_net), .O(n5437));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4053_3_lut (.I0(\REG.mem_31_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n34), .I3(GND_net), .O(n5436));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4052_3_lut (.I0(\REG.mem_31_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n34), .I3(GND_net), .O(n5435));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4051_3_lut (.I0(\REG.mem_31_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n34), .I3(GND_net), .O(n5434));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4050_3_lut (.I0(\REG.mem_31_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n34), .I3(GND_net), .O(n5433));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4049_3_lut (.I0(\REG.mem_31_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n34), .I3(GND_net), .O(n5432));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4048_3_lut (.I0(\REG.mem_31_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n34), .I3(GND_net), .O(n5431));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4047_3_lut (.I0(\REG.mem_31_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n34), .I3(GND_net), .O(n5430));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4046_3_lut (.I0(\REG.mem_31_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n34), .I3(GND_net), .O(n5429));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4045_3_lut (.I0(\REG.mem_31_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n34), .I3(GND_net), .O(n5428));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4044_3_lut (.I0(\REG.mem_31_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n34), .I3(GND_net), .O(n5427));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4043_3_lut (.I0(\REG.mem_31_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n34), .I3(GND_net), .O(n5426));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4042_3_lut (.I0(\REG.mem_31_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n34), .I3(GND_net), .O(n5425));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4041_3_lut (.I0(\REG.mem_30_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n35), .I3(GND_net), .O(n5424));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4040_3_lut (.I0(\REG.mem_30_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n35), .I3(GND_net), .O(n5423));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4039_3_lut (.I0(\REG.mem_30_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n35), .I3(GND_net), .O(n5422));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4038_3_lut (.I0(\REG.mem_30_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n35), .I3(GND_net), .O(n5421));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4037_3_lut (.I0(\REG.mem_30_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n35), .I3(GND_net), .O(n5420));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4036_3_lut (.I0(\REG.mem_30_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n35), .I3(GND_net), .O(n5419));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4035_3_lut (.I0(\REG.mem_30_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n35), .I3(GND_net), .O(n5418));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4034_3_lut (.I0(\REG.mem_30_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n35), .I3(GND_net), .O(n5417));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4033_3_lut (.I0(\REG.mem_30_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n35), .I3(GND_net), .O(n5416));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4032_3_lut (.I0(\REG.mem_30_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n35), .I3(GND_net), .O(n5415));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4031_3_lut (.I0(\REG.mem_30_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n35), .I3(GND_net), .O(n5414));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4030_3_lut (.I0(\REG.mem_30_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n35), .I3(GND_net), .O(n5413));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4029_3_lut (.I0(\REG.mem_30_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n35), .I3(GND_net), .O(n5412));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4028_3_lut (.I0(\REG.mem_30_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n35), .I3(GND_net), .O(n5411));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4027_3_lut (.I0(\REG.mem_30_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n35), .I3(GND_net), .O(n5410));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4026_3_lut (.I0(\REG.mem_30_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n35), .I3(GND_net), .O(n5409));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_1242));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3500_3_lut (.I0(rx_shift_reg[2]), .I1(rx_shift_reg[1]), .I2(n4312), 
            .I3(GND_net), .O(n4883));   // src/spi.v(76[8] 221[4])
    defparam i3500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3961_3_lut (.I0(\REG.mem_25_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n40), .I3(GND_net), .O(n5344));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3960_3_lut (.I0(\REG.mem_25_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n40), .I3(GND_net), .O(n5343));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3959_3_lut (.I0(\REG.mem_25_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n40), .I3(GND_net), .O(n5342));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3958_3_lut (.I0(\REG.mem_25_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n40), .I3(GND_net), .O(n5341));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3957_3_lut (.I0(\REG.mem_25_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n40), .I3(GND_net), .O(n5340));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3956_3_lut (.I0(\REG.mem_25_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n40), .I3(GND_net), .O(n5339));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3955_3_lut (.I0(\REG.mem_25_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n40), .I3(GND_net), .O(n5338));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3954_3_lut (.I0(\REG.mem_25_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n40), .I3(GND_net), .O(n5337));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3953_3_lut (.I0(\REG.mem_25_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n40), .I3(GND_net), .O(n5336));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3952_3_lut (.I0(\REG.mem_25_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n40), .I3(GND_net), .O(n5335));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3951_3_lut (.I0(\REG.mem_25_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n40), .I3(GND_net), .O(n5334));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3950_3_lut (.I0(\REG.mem_25_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n40), .I3(GND_net), .O(n5333));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3949_3_lut (.I0(\REG.mem_25_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n40), .I3(GND_net), .O(n5332));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3948_3_lut (.I0(\REG.mem_25_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n40), .I3(GND_net), .O(n5331));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3947_3_lut (.I0(\REG.mem_25_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n40), .I3(GND_net), .O(n5330));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3946_3_lut (.I0(\REG.mem_25_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n40), .I3(GND_net), .O(n5329));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3923_3_lut (.I0(\REG.mem_23_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n42), .I3(GND_net), .O(n5306));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3922_3_lut (.I0(\REG.mem_23_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n42), .I3(GND_net), .O(n5305));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3921_3_lut (.I0(\REG.mem_23_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n42), .I3(GND_net), .O(n5304));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3920_3_lut (.I0(\REG.mem_23_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n42), .I3(GND_net), .O(n5303));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3919_3_lut (.I0(\REG.mem_23_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n42), .I3(GND_net), .O(n5302));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3918_3_lut (.I0(\REG.mem_23_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n42), .I3(GND_net), .O(n5301));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3917_3_lut (.I0(\REG.mem_23_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n42), .I3(GND_net), .O(n5300));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3916_3_lut (.I0(\REG.mem_23_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n42), .I3(GND_net), .O(n5299));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3915_3_lut (.I0(\REG.mem_23_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n42), .I3(GND_net), .O(n5298));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3914_3_lut (.I0(\REG.mem_23_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n42), .I3(GND_net), .O(n5297));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3913_3_lut (.I0(\REG.mem_23_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n42), .I3(GND_net), .O(n5296));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3912_3_lut (.I0(\REG.mem_23_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n42), .I3(GND_net), .O(n5295));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3911_3_lut (.I0(\REG.mem_23_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n42), .I3(GND_net), .O(n5294));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3910_3_lut (.I0(\REG.mem_23_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n42), .I3(GND_net), .O(n5293));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3909_3_lut (.I0(\REG.mem_23_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n42), .I3(GND_net), .O(n5292));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3908_3_lut (.I0(\REG.mem_23_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n42), .I3(GND_net), .O(n5291));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3907_3_lut (.I0(\REG.mem_22_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n43), .I3(GND_net), .O(n5290));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3906_3_lut (.I0(\REG.mem_22_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n43), .I3(GND_net), .O(n5289));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3905_3_lut (.I0(\REG.mem_22_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n43), .I3(GND_net), .O(n5288));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3904_3_lut (.I0(\REG.mem_22_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n43), .I3(GND_net), .O(n5287));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3903_3_lut (.I0(\REG.mem_22_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n43), .I3(GND_net), .O(n5286));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3902_3_lut (.I0(\REG.mem_22_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n43), .I3(GND_net), .O(n5285));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3901_3_lut (.I0(\REG.mem_22_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n43), .I3(GND_net), .O(n5284));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3900_3_lut (.I0(\REG.mem_22_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n43), .I3(GND_net), .O(n5283));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3899_3_lut (.I0(\REG.mem_22_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n43), .I3(GND_net), .O(n5282));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3898_3_lut (.I0(\REG.mem_22_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n43), .I3(GND_net), .O(n5281));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3897_3_lut (.I0(\REG.mem_22_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n43), .I3(GND_net), .O(n5280));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3896_3_lut (.I0(\REG.mem_22_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n43), .I3(GND_net), .O(n5279));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3895_3_lut (.I0(\REG.mem_22_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n43), .I3(GND_net), .O(n5278));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3894_3_lut (.I0(\REG.mem_22_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n43), .I3(GND_net), .O(n5277));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3893_3_lut (.I0(\REG.mem_22_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n43), .I3(GND_net), .O(n5276));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3892_3_lut (.I0(\REG.mem_22_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n43), .I3(GND_net), .O(n5275));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3843_3_lut (.I0(\REG.mem_18_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n47), .I3(GND_net), .O(n5226));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3842_3_lut (.I0(\REG.mem_18_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n47), .I3(GND_net), .O(n5225));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3841_3_lut (.I0(\REG.mem_18_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n47), .I3(GND_net), .O(n5224));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3840_3_lut (.I0(\REG.mem_18_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n47), .I3(GND_net), .O(n5223));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3839_3_lut (.I0(\REG.mem_18_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n47), .I3(GND_net), .O(n5222));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3838_3_lut (.I0(\REG.mem_18_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n47), .I3(GND_net), .O(n5221));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3837_3_lut (.I0(\REG.mem_18_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n47), .I3(GND_net), .O(n5220));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3836_3_lut (.I0(\REG.mem_18_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n47), .I3(GND_net), .O(n5219));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3835_3_lut (.I0(\REG.mem_18_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n47), .I3(GND_net), .O(n5218));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3834_3_lut (.I0(\REG.mem_18_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n47), .I3(GND_net), .O(n5217));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3833_3_lut (.I0(\REG.mem_18_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n47), .I3(GND_net), .O(n5216));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3832_3_lut (.I0(\REG.mem_18_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n47), .I3(GND_net), .O(n5215));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3831_3_lut (.I0(\REG.mem_18_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n47), .I3(GND_net), .O(n5214));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3830_3_lut (.I0(\REG.mem_18_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n47), .I3(GND_net), .O(n5213));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3829_3_lut (.I0(\REG.mem_18_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n47), .I3(GND_net), .O(n5212));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3828_3_lut (.I0(\REG.mem_18_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n47), .I3(GND_net), .O(n5211));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1590_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n2944));   // src/top.v(1074[8] 1141[4])
    defparam i1590_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3811_3_lut (.I0(r_Tx_Data[1]), .I1(fifo_temp_output[1]), .I2(n3794), 
            .I3(GND_net), .O(n5194));   // src/uart_tx.v(38[10] 141[8])
    defparam i3811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3810_3_lut (.I0(r_Tx_Data[2]), .I1(fifo_temp_output[2]), .I2(n3794), 
            .I3(GND_net), .O(n5193));   // src/uart_tx.v(38[10] 141[8])
    defparam i3810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3809_3_lut (.I0(r_Tx_Data[3]), .I1(fifo_temp_output[3]), .I2(n3794), 
            .I3(GND_net), .O(n5192));   // src/uart_tx.v(38[10] 141[8])
    defparam i3809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3808_3_lut (.I0(r_Tx_Data[4]), .I1(fifo_temp_output[4]), .I2(n3794), 
            .I3(GND_net), .O(n5191));   // src/uart_tx.v(38[10] 141[8])
    defparam i3808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3807_3_lut (.I0(\REG.mem_16_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n49), .I3(GND_net), .O(n5190));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3806_3_lut (.I0(r_Tx_Data[5]), .I1(fifo_temp_output[5]), .I2(n3794), 
            .I3(GND_net), .O(n5189));   // src/uart_tx.v(38[10] 141[8])
    defparam i3806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3805_3_lut (.I0(\REG.mem_16_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n49), .I3(GND_net), .O(n5188));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3804_3_lut (.I0(\REG.mem_16_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n49), .I3(GND_net), .O(n5187));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3803_3_lut (.I0(\REG.mem_16_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n49), .I3(GND_net), .O(n5186));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3802_3_lut (.I0(\REG.mem_16_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n49), .I3(GND_net), .O(n5185));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3801_3_lut (.I0(\REG.mem_16_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n49), .I3(GND_net), .O(n5184));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3800_3_lut (.I0(\REG.mem_16_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n49), .I3(GND_net), .O(n5183));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3799_3_lut (.I0(\REG.mem_16_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n49), .I3(GND_net), .O(n5182));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3798_3_lut (.I0(\REG.mem_16_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n49), .I3(GND_net), .O(n5181));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3797_3_lut (.I0(\REG.mem_16_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n49), .I3(GND_net), .O(n5180));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3796_3_lut (.I0(\REG.mem_16_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n49), .I3(GND_net), .O(n5179));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3795_3_lut (.I0(\REG.mem_16_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n49), .I3(GND_net), .O(n5178));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3794_3_lut (.I0(\REG.mem_16_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n49), .I3(GND_net), .O(n5177));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3793_3_lut (.I0(\REG.mem_16_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n49), .I3(GND_net), .O(n5176));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(rd_fifo_en_prev_r), .I1(fifo_read_cmd), 
            .I2(is_fifo_empty_flag), .I3(reset_all_w), .O(n4459));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hffae;
    SB_LUT4 i3792_3_lut (.I0(\REG.mem_16_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n49), .I3(GND_net), .O(n5175));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3791_3_lut (.I0(\REG.mem_16_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n49), .I3(GND_net), .O(n5174));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3790_3_lut (.I0(r_Tx_Data[6]), .I1(fifo_temp_output[6]), .I2(n3794), 
            .I3(GND_net), .O(n5173));   // src/uart_tx.v(38[10] 141[8])
    defparam i3790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3789_3_lut (.I0(r_Tx_Data[7]), .I1(fifo_temp_output[7]), .I2(n3794), 
            .I3(GND_net), .O(n5172));   // src/uart_tx.v(38[10] 141[8])
    defparam i3789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3788_3_lut (.I0(\REG.mem_15_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n50), .I3(GND_net), .O(n5171));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3787_3_lut (.I0(\REG.mem_15_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n50), .I3(GND_net), .O(n5170));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3786_3_lut (.I0(\REG.mem_15_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n50), .I3(GND_net), .O(n5169));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3785_3_lut (.I0(\REG.mem_15_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n50), .I3(GND_net), .O(n5168));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3293_1_lut_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n4676));   // src/top.v(1074[8] 1141[4])
    defparam i3293_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i3495_2_lut_3_lut (.I0(reset_all_w), .I1(fifo_read_cmd), .I2(is_fifo_empty_flag), 
            .I3(GND_net), .O(n4878));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    defparam i3495_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i3784_3_lut (.I0(\REG.mem_15_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n50), .I3(GND_net), .O(n5167));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3783_3_lut (.I0(\REG.mem_15_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n50), .I3(GND_net), .O(n5166));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3782_3_lut (.I0(\REG.mem_15_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n50), .I3(GND_net), .O(n5165));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3781_3_lut (.I0(\REG.mem_15_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n50), .I3(GND_net), .O(n5164));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3780_3_lut (.I0(\REG.mem_15_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n50), .I3(GND_net), .O(n5163));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3779_3_lut (.I0(\REG.mem_15_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n50), .I3(GND_net), .O(n5162));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3778_3_lut (.I0(\REG.mem_15_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n50), .I3(GND_net), .O(n5161));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3777_3_lut (.I0(\REG.mem_15_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n50), .I3(GND_net), .O(n5160));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3776_3_lut (.I0(\REG.mem_15_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n50), .I3(GND_net), .O(n5159));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3775_3_lut (.I0(\REG.mem_15_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n50), .I3(GND_net), .O(n5158));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3774_3_lut (.I0(\REG.mem_15_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n50), .I3(GND_net), .O(n5157));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3773_3_lut (.I0(\REG.mem_15_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n50), .I3(GND_net), .O(n5156));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3772_3_lut (.I0(\REG.mem_14_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n51), .I3(GND_net), .O(n5155));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3506_4_lut_4_lut (.I0(tx_uart_active_flag), .I1(r_SM_Main_adj_1261[1]), 
            .I2(r_SM_Main_adj_1261[2]), .I3(n10653), .O(n4889));   // src/uart_tx.v(38[10] 141[8])
    defparam i3506_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i3771_3_lut (.I0(\REG.mem_14_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n51), .I3(GND_net), .O(n5154));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3770_3_lut (.I0(\REG.mem_14_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n51), .I3(GND_net), .O(n5153));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3769_3_lut (.I0(\REG.mem_14_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n51), .I3(GND_net), .O(n5152));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3768_3_lut (.I0(\REG.mem_14_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n51), .I3(GND_net), .O(n5151));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3767_3_lut (.I0(\REG.mem_14_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n51), .I3(GND_net), .O(n5150));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3766_3_lut (.I0(\REG.mem_14_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n51), .I3(GND_net), .O(n5149));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3765_3_lut (.I0(\REG.mem_14_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n51), .I3(GND_net), .O(n5148));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3764_3_lut (.I0(\REG.mem_14_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n51), .I3(GND_net), .O(n5147));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3763_3_lut (.I0(\REG.mem_14_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n51), .I3(GND_net), .O(n5146));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3762_3_lut (.I0(\REG.mem_14_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n51), .I3(GND_net), .O(n5145));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3761_3_lut (.I0(\REG.mem_14_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n51), .I3(GND_net), .O(n5144));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3760_3_lut (.I0(\REG.mem_14_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n51), .I3(GND_net), .O(n5143));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3759_3_lut (.I0(\REG.mem_14_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n51), .I3(GND_net), .O(n5142));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3758_3_lut (.I0(\REG.mem_14_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n51), .I3(GND_net), .O(n5141));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3757_3_lut (.I0(\REG.mem_14_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n51), .I3(GND_net), .O(n5140));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3756_3_lut (.I0(\REG.mem_13_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n52), .I3(GND_net), .O(n5139));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3755_3_lut (.I0(\REG.mem_13_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n52), .I3(GND_net), .O(n5138));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3754_3_lut (.I0(\REG.mem_13_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n52), .I3(GND_net), .O(n5137));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3753_3_lut (.I0(\REG.mem_13_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n52), .I3(GND_net), .O(n5136));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3752_3_lut (.I0(\REG.mem_13_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n52), .I3(GND_net), .O(n5135));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3751_3_lut (.I0(\REG.mem_13_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n52), .I3(GND_net), .O(n5134));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3750_3_lut (.I0(\REG.mem_13_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n52), .I3(GND_net), .O(n5133));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3494_3_lut (.I0(rx_shift_reg[3]), .I1(rx_shift_reg[2]), .I2(n4312), 
            .I3(GND_net), .O(n4877));   // src/spi.v(76[8] 221[4])
    defparam i3494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3749_3_lut (.I0(\REG.mem_13_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n52), .I3(GND_net), .O(n5132));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3748_3_lut (.I0(\REG.mem_13_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n52), .I3(GND_net), .O(n5131));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_1261[1]), .I1(r_SM_Main_2__N_841[1]), 
            .I2(r_SM_Main_adj_1261[0]), .I3(r_SM_Main_adj_1261[2]), .O(n13737));   // src/uart_tx.v(38[10] 141[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i3747_3_lut (.I0(\REG.mem_13_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n52), .I3(GND_net), .O(n5130));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3746_3_lut (.I0(\REG.mem_13_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n52), .I3(GND_net), .O(n5129));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3745_3_lut (.I0(\REG.mem_13_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n52), .I3(GND_net), .O(n5128));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1601_2_lut_3_lut_4_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(reset_all_w), .I3(wr_addr_r_adj_1284[0]), .O(n8));
    defparam i1601_2_lut_3_lut_4_lut.LUT_INIT = 16'h0df2;
    SB_LUT4 i3744_3_lut (.I0(\REG.mem_13_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n52), .I3(GND_net), .O(n5127));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3743_3_lut (.I0(\REG.mem_13_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n52), .I3(GND_net), .O(n5126));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3742_3_lut (.I0(\REG.mem_13_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n52), .I3(GND_net), .O(n5125));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3741_3_lut (.I0(\REG.mem_13_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n52), .I3(GND_net), .O(n5124));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3740_3_lut (.I0(\REG.mem_12_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n53), .I3(GND_net), .O(n5123));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3739_3_lut (.I0(\REG.mem_12_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n53), .I3(GND_net), .O(n5122));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3738_3_lut (.I0(\REG.mem_12_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n53), .I3(GND_net), .O(n5121));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3737_3_lut (.I0(\REG.mem_12_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n53), .I3(GND_net), .O(n5120));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3736_3_lut (.I0(\REG.mem_12_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n53), .I3(GND_net), .O(n5119));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3735_3_lut (.I0(\REG.mem_12_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n53), .I3(GND_net), .O(n5118));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3734_3_lut (.I0(\REG.mem_12_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n53), .I3(GND_net), .O(n5117));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3733_3_lut (.I0(\REG.mem_12_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n53), .I3(GND_net), .O(n5116));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3486_3_lut (.I0(rx_shift_reg[4]), .I1(rx_shift_reg[3]), .I2(n4312), 
            .I3(GND_net), .O(n4869));   // src/spi.v(76[8] 221[4])
    defparam i3486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3732_3_lut (.I0(\REG.mem_12_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n53), .I3(GND_net), .O(n5115));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3731_3_lut (.I0(\REG.mem_12_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n53), .I3(GND_net), .O(n5114));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3730_3_lut (.I0(\REG.mem_12_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n53), .I3(GND_net), .O(n5113));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3729_3_lut (.I0(\REG.mem_12_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n53), .I3(GND_net), .O(n5112));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3728_3_lut (.I0(\REG.mem_12_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n53), .I3(GND_net), .O(n5111));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3727_3_lut (.I0(\REG.mem_12_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n53), .I3(GND_net), .O(n5110));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3726_3_lut (.I0(\REG.mem_12_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n53), .I3(GND_net), .O(n5109));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3725_3_lut (.I0(\REG.mem_12_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n53), .I3(GND_net), .O(n5108));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3724_3_lut (.I0(\REG.mem_11_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n54), .I3(GND_net), .O(n5107));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10191_4_lut (.I0(tx_data_byte[0]), .I1(tx_data_byte[1]), .I2(tx_data_byte[6]), 
            .I3(n10834), .O(multi_byte_spi_trans_flag_r_N_72));   // src/top.v(1123[10:31])
    defparam i10191_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i8984_4_lut (.I0(tx_data_byte[3]), .I1(tx_data_byte[2]), .I2(tx_data_byte[4]), 
            .I3(n10754), .O(n10834));
    defparam i8984_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8905_2_lut (.I0(tx_data_byte[5]), .I1(tx_data_byte[7]), .I2(GND_net), 
            .I3(GND_net), .O(n10754));
    defparam i8905_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3723_3_lut (.I0(\REG.mem_11_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n54), .I3(GND_net), .O(n5106));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3722_3_lut (.I0(\REG.mem_11_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n54), .I3(GND_net), .O(n5105));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3721_3_lut (.I0(\REG.mem_11_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n54), .I3(GND_net), .O(n5104));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3720_3_lut (.I0(\REG.mem_11_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n54), .I3(GND_net), .O(n5103));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3719_3_lut (.I0(\REG.mem_11_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n54), .I3(GND_net), .O(n5102));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3718_3_lut (.I0(\REG.mem_11_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n54), .I3(GND_net), .O(n5101));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3717_3_lut (.I0(\REG.mem_11_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n54), .I3(GND_net), .O(n5100));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3716_3_lut (.I0(\REG.mem_11_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n54), .I3(GND_net), .O(n5099));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3715_3_lut (.I0(\REG.mem_11_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n54), .I3(GND_net), .O(n5098));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3715_3_lut.LUT_INIT = 16'hcaca;
    fifo_dc_32_lut_gen2 fifo_dc_32_lut_gen_inst (.dc32_fifo_almost_full(dc32_fifo_almost_full), 
            .FIFO_CLK_c(FIFO_CLK_c), .reset_per_frame(reset_per_frame), 
            .\REG.mem_16_7 (\REG.mem_16_7 ), .\rd_addr_r[0] (rd_addr_r[0]), 
            .\REG.mem_6_2 (\REG.mem_6_2 ), .\REG.mem_7_2 (\REG.mem_7_2 ), 
            .\dc32_fifo_data_in[7] (dc32_fifo_data_in[7]), .\REG.mem_46_9 (\REG.mem_46_9 ), 
            .\REG.mem_47_9 (\REG.mem_47_9 ), .\REG.mem_25_5 (\REG.mem_25_5 ), 
            .GND_net(GND_net), .t_rd_fifo_en_w(t_rd_fifo_en_w), .\REG.out_raw[0] (\REG.out_raw [0]), 
            .SLM_CLK_c(SLM_CLK_c), .\REG.mem_45_9 (\REG.mem_45_9 ), .\REG.mem_44_9 (\REG.mem_44_9 ), 
            .\REG.mem_57_15 (\REG.mem_57_15 ), .\REG.mem_62_15 (\REG.mem_62_15 ), 
            .\REG.mem_63_15 (\REG.mem_63_15 ), .\REG.mem_6_1 (\REG.mem_6_1 ), 
            .\REG.mem_7_1 (\REG.mem_7_1 ), .\REG.mem_5_1 (\REG.mem_5_1 ), 
            .\REG.mem_4_1 (\REG.mem_4_1 ), .\REG.mem_57_1 (\REG.mem_57_1 ), 
            .\REG.mem_25_9 (\REG.mem_25_9 ), .\dc32_fifo_data_in[6] (dc32_fifo_data_in[6]), 
            .\dc32_fifo_data_in[15] (dc32_fifo_data_in[15]), .\REG.mem_46_3 (\REG.mem_46_3 ), 
            .\REG.mem_47_3 (\REG.mem_47_3 ), .\REG.mem_45_3 (\REG.mem_45_3 ), 
            .\REG.mem_44_3 (\REG.mem_44_3 ), .\REG.mem_54_13 (\REG.mem_54_13 ), 
            .\REG.mem_55_13 (\REG.mem_55_13 ), .\REG.mem_50_11 (\REG.mem_50_11 ), 
            .\REG.mem_48_11 (\REG.mem_48_11 ), .\dc32_fifo_data_in[5] (dc32_fifo_data_in[5]), 
            .\REG.mem_42_12 (\REG.mem_42_12 ), .\REG.mem_43_12 (\REG.mem_43_12 ), 
            .\REG.mem_41_12 (\REG.mem_41_12 ), .\REG.mem_40_12 (\REG.mem_40_12 ), 
            .\dc32_fifo_data_in[4] (dc32_fifo_data_in[4]), .\dc32_fifo_data_in[3] (dc32_fifo_data_in[3]), 
            .\dc32_fifo_data_in[2] (dc32_fifo_data_in[2]), .\rd_grey_sync_r[0] (rd_grey_sync_r[0]), 
            .\REG.mem_57_6 (\REG.mem_57_6 ), .DEBUG_3_c(DEBUG_3_c), .wr_grey_sync_r({wr_grey_sync_r}), 
            .\dc32_fifo_data_in[1] (dc32_fifo_data_in[1]), .\REG.mem_54_11 (\REG.mem_54_11 ), 
            .\REG.mem_55_11 (\REG.mem_55_11 ), .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .dc32_fifo_almost_empty(dc32_fifo_almost_empty), .\REG.mem_14_12 (\REG.mem_14_12 ), 
            .\REG.mem_15_12 (\REG.mem_15_12 ), .\REG.mem_30_0 (\REG.mem_30_0 ), 
            .\REG.mem_31_0 (\REG.mem_31_0 ), .\REG.mem_13_12 (\REG.mem_13_12 ), 
            .\REG.mem_12_12 (\REG.mem_12_12 ), .\REG.mem_3_5 (\REG.mem_3_5 ), 
            .\REG.mem_6_5 (\REG.mem_6_5 ), .\REG.mem_7_5 (\REG.mem_7_5 ), 
            .\REG.mem_4_5 (\REG.mem_4_5 ), .\REG.mem_5_5 (\REG.mem_5_5 ), 
            .\REG.mem_57_11 (\REG.mem_57_11 ), .n62(n62), .\REG.mem_62_13 (\REG.mem_62_13 ), 
            .\REG.mem_63_13 (\REG.mem_63_13 ), .\REG.mem_46_1 (\REG.mem_46_1 ), 
            .\REG.mem_47_1 (\REG.mem_47_1 ), .\REG.mem_45_1 (\REG.mem_45_1 ), 
            .\REG.mem_44_1 (\REG.mem_44_1 ), .\dc32_fifo_data_in[0] (dc32_fifo_data_in[0]), 
            .\REG.mem_3_11 (\REG.mem_3_11 ), .\REG.mem_6_11 (\REG.mem_6_11 ), 
            .\REG.mem_7_11 (\REG.mem_7_11 ), .n30(n30), .\REG.mem_5_2 (\REG.mem_5_2 ), 
            .\REG.mem_4_2 (\REG.mem_4_2 ), .\REG.mem_18_5 (\REG.mem_18_5 ), 
            .\REG.mem_62_1 (\REG.mem_62_1 ), .\REG.mem_63_1 (\REG.mem_63_1 ), 
            .\REG.mem_38_13 (\REG.mem_38_13 ), .\REG.mem_39_13 (\REG.mem_39_13 ), 
            .\REG.mem_5_11 (\REG.mem_5_11 ), .\REG.mem_4_11 (\REG.mem_4_11 ), 
            .\dc32_fifo_data_in[8] (dc32_fifo_data_in[8]), .\REG.mem_14_5 (\REG.mem_14_5 ), 
            .\REG.mem_15_5 (\REG.mem_15_5 ), .\REG.mem_13_5 (\REG.mem_13_5 ), 
            .\REG.mem_12_5 (\REG.mem_12_5 ), .\REG.mem_30_9 (\REG.mem_30_9 ), 
            .\REG.mem_31_9 (\REG.mem_31_9 ), .\wr_addr_nxt_c[5] (wr_addr_nxt_c[5]), 
            .\REG.mem_46_12 (\REG.mem_46_12 ), .\REG.mem_47_12 (\REG.mem_47_12 ), 
            .\REG.mem_45_12 (\REG.mem_45_12 ), .\REG.mem_44_12 (\REG.mem_44_12 ), 
            .\REG.mem_62_11 (\REG.mem_62_11 ), .\REG.mem_63_11 (\REG.mem_63_11 ), 
            .\REG.mem_57_8 (\REG.mem_57_8 ), .\REG.mem_62_6 (\REG.mem_62_6 ), 
            .\REG.mem_63_6 (\REG.mem_63_6 ), .\REG.mem_62_8 (\REG.mem_62_8 ), 
            .\REG.mem_63_8 (\REG.mem_63_8 ), .\REG.mem_35_0 (\REG.mem_35_0 ), 
            .\REG.mem_25_15 (\REG.mem_25_15 ), .\REG.mem_35_7 (\REG.mem_35_7 ), 
            .\REG.mem_35_9 (\REG.mem_35_9 ), .\REG.mem_18_12 (\REG.mem_18_12 ), 
            .\REG.mem_16_12 (\REG.mem_16_12 ), .\REG.mem_14_8 (\REG.mem_14_8 ), 
            .\REG.mem_15_8 (\REG.mem_15_8 ), .\REG.mem_13_8 (\REG.mem_13_8 ), 
            .\REG.mem_12_8 (\REG.mem_12_8 ), .\REG.mem_14_2 (\REG.mem_14_2 ), 
            .\REG.mem_15_2 (\REG.mem_15_2 ), .\REG.mem_13_2 (\REG.mem_13_2 ), 
            .\REG.mem_12_2 (\REG.mem_12_2 ), .\REG.mem_38_7 (\REG.mem_38_7 ), 
            .\REG.mem_39_7 (\REG.mem_39_7 ), .\REG.mem_36_7 (\REG.mem_36_7 ), 
            .\REG.mem_37_7 (\REG.mem_37_7 ), .\REG.mem_50_12 (\REG.mem_50_12 ), 
            .\REG.mem_48_12 (\REG.mem_48_12 ), .\REG.mem_62_9 (\REG.mem_62_9 ), 
            .\REG.mem_63_9 (\REG.mem_63_9 ), .\REG.mem_6_9 (\REG.mem_6_9 ), 
            .\REG.mem_7_9 (\REG.mem_7_9 ), .\REG.mem_35_6 (\REG.mem_35_6 ), 
            .\REG.mem_5_9 (\REG.mem_5_9 ), .\REG.mem_4_9 (\REG.mem_4_9 ), 
            .\REG.mem_37_13 (\REG.mem_37_13 ), .\REG.mem_36_13 (\REG.mem_36_13 ), 
            .\REG.mem_42_8 (\REG.mem_42_8 ), .\REG.mem_43_8 (\REG.mem_43_8 ), 
            .\REG.mem_41_8 (\REG.mem_41_8 ), .\REG.mem_40_8 (\REG.mem_40_8 ), 
            .\REG.mem_22_7 (\REG.mem_22_7 ), .\REG.mem_23_7 (\REG.mem_23_7 ), 
            .\REG.mem_10_11 (\REG.mem_10_11 ), .\REG.mem_11_11 (\REG.mem_11_11 ), 
            .\REG.mem_9_11 (\REG.mem_9_11 ), .\REG.mem_8_11 (\REG.mem_8_11 ), 
            .\REG.mem_3_15 (\REG.mem_3_15 ), .\REG.mem_46_8 (\REG.mem_46_8 ), 
            .\REG.mem_47_8 (\REG.mem_47_8 ), .\REG.mem_45_8 (\REG.mem_45_8 ), 
            .\REG.mem_44_8 (\REG.mem_44_8 ), .\REG.mem_46_5 (\REG.mem_46_5 ), 
            .\REG.mem_47_5 (\REG.mem_47_5 ), .\REG.mem_45_5 (\REG.mem_45_5 ), 
            .\REG.mem_44_5 (\REG.mem_44_5 ), .\REG.mem_10_2 (\REG.mem_10_2 ), 
            .\REG.mem_11_2 (\REG.mem_11_2 ), .\REG.mem_54_9 (\REG.mem_54_9 ), 
            .\REG.mem_55_9 (\REG.mem_55_9 ), .\REG.mem_57_9 (\REG.mem_57_9 ), 
            .\REG.mem_57_14 (\REG.mem_57_14 ), .\REG.mem_30_15 (\REG.mem_30_15 ), 
            .\REG.mem_31_15 (\REG.mem_31_15 ), .\REG.mem_42_15 (\REG.mem_42_15 ), 
            .\REG.mem_43_15 (\REG.mem_43_15 ), .\REG.mem_16_5 (\REG.mem_16_5 ), 
            .\REG.mem_9_2 (\REG.mem_9_2 ), .\REG.mem_8_2 (\REG.mem_8_2 ), 
            .\REG.mem_62_12 (\REG.mem_62_12 ), .\REG.mem_63_12 (\REG.mem_63_12 ), 
            .\wr_addr_nxt_c[3] (wr_addr_nxt_c[3]), .\REG.mem_18_8 (\REG.mem_18_8 ), 
            .\REG.mem_16_8 (\REG.mem_16_8 ), .\REG.mem_22_12 (\REG.mem_22_12 ), 
            .\REG.mem_23_12 (\REG.mem_23_12 ), .\REG.mem_25_2 (\REG.mem_25_2 ), 
            .\REG.mem_30_2 (\REG.mem_30_2 ), .\REG.mem_31_2 (\REG.mem_31_2 ), 
            .\dc32_fifo_data_in[14] (dc32_fifo_data_in[14]), .\REG.mem_48_10 (\REG.mem_48_10 ), 
            .\REG.mem_50_10 (\REG.mem_50_10 ), .\dc32_fifo_data_in[13] (dc32_fifo_data_in[13]), 
            .\REG.mem_54_10 (\REG.mem_54_10 ), .\REG.mem_55_10 (\REG.mem_55_10 ), 
            .\REG.mem_14_11 (\REG.mem_14_11 ), .\REG.mem_15_11 (\REG.mem_15_11 ), 
            .\dc32_fifo_data_in[12] (dc32_fifo_data_in[12]), .\REG.mem_54_12 (\REG.mem_54_12 ), 
            .\REG.mem_55_12 (\REG.mem_55_12 ), .\REG.mem_13_11 (\REG.mem_13_11 ), 
            .\REG.mem_12_11 (\REG.mem_12_11 ), .\REG.mem_35_15 (\REG.mem_35_15 ), 
            .\REG.mem_38_6 (\REG.mem_38_6 ), .\REG.mem_39_6 (\REG.mem_39_6 ), 
            .\dc32_fifo_data_in[11] (dc32_fifo_data_in[11]), .\REG.mem_37_6 (\REG.mem_37_6 ), 
            .\REG.mem_36_6 (\REG.mem_36_6 ), .\REG.mem_57_13 (\REG.mem_57_13 ), 
            .\dc32_fifo_data_in[10] (dc32_fifo_data_in[10]), .\dc32_fifo_data_in[9] (dc32_fifo_data_in[9]), 
            .\REG.mem_30_13 (\REG.mem_30_13 ), .\REG.mem_31_13 (\REG.mem_31_13 ), 
            .\REG.mem_30_5 (\REG.mem_30_5 ), .\REG.mem_31_5 (\REG.mem_31_5 ), 
            .\REG.mem_48_7 (\REG.mem_48_7 ), .\REG.mem_50_7 (\REG.mem_50_7 ), 
            .\REG.mem_54_7 (\REG.mem_54_7 ), .\REG.mem_55_7 (\REG.mem_55_7 ), 
            .n6106(n6106), .VCC_net(VCC_net), .\fifo_data_out[2] (fifo_data_out[2]), 
            .n6103(n6103), .\fifo_data_out[1] (fifo_data_out[1]), .\REG.mem_35_13 (\REG.mem_35_13 ), 
            .\REG.mem_3_3 (\REG.mem_3_3 ), .\rd_addr_r[6] (rd_addr_r[6]), 
            .n4827(n4827), .\fifo_data_out[3] (fifo_data_out[3]), .\REG.mem_50_1 (\REG.mem_50_1 ), 
            .n4830(n4830), .\fifo_data_out[4] (fifo_data_out[4]), .n4841(n4841), 
            .\fifo_data_out[5] (fifo_data_out[5]), .n4844(n4844), .\fifo_data_out[6] (fifo_data_out[6]), 
            .n4848(n4848), .\fifo_data_out[7] (fifo_data_out[7]), .n4851(n4851), 
            .\fifo_data_out[8] (fifo_data_out[8]), .n4854(n4854), .\fifo_data_out[9] (fifo_data_out[9]), 
            .n4858(n4858), .\fifo_data_out[10] (fifo_data_out[10]), .n4864(n4864), 
            .\fifo_data_out[11] (fifo_data_out[11]), .\REG.mem_62_14 (\REG.mem_62_14 ), 
            .\REG.mem_63_14 (\REG.mem_63_14 ), .\REG.mem_48_1 (\REG.mem_48_1 ), 
            .\REG.mem_18_11 (\REG.mem_18_11 ), .\REG.mem_16_11 (\REG.mem_16_11 ), 
            .\REG.mem_6_3 (\REG.mem_6_3 ), .\REG.mem_7_3 (\REG.mem_7_3 ), 
            .\REG.mem_5_3 (\REG.mem_5_3 ), .\REG.mem_4_3 (\REG.mem_4_3 ), 
            .\REG.mem_42_2 (\REG.mem_42_2 ), .\REG.mem_43_2 (\REG.mem_43_2 ), 
            .\REG.mem_41_2 (\REG.mem_41_2 ), .\REG.mem_40_2 (\REG.mem_40_2 ), 
            .n6070(n6070), .\fifo_data_out[0] (fifo_data_out[0]), .\REG.mem_46_2 (\REG.mem_46_2 ), 
            .\REG.mem_47_2 (\REG.mem_47_2 ), .\REG.mem_45_2 (\REG.mem_45_2 ), 
            .\REG.mem_44_2 (\REG.mem_44_2 ), .\REG.mem_14_7 (\REG.mem_14_7 ), 
            .\REG.mem_15_7 (\REG.mem_15_7 ), .n4872(n4872), .\fifo_data_out[12] (fifo_data_out[12]), 
            .n4875(n4875), .\fifo_data_out[13] (fifo_data_out[13]), .\REG.mem_13_7 (\REG.mem_13_7 ), 
            .\REG.mem_12_7 (\REG.mem_12_7 ), .n6034(n6034), .\REG.mem_25_13 (\REG.mem_25_13 ), 
            .n6032(n6032), .\REG.mem_10_3 (\REG.mem_10_3 ), .\REG.mem_11_3 (\REG.mem_11_3 ), 
            .\REG.mem_9_3 (\REG.mem_9_3 ), .\REG.mem_8_3 (\REG.mem_8_3 ), 
            .\REG.mem_50_9 (\REG.mem_50_9 ), .n6013(n6013), .n6012(n6012), 
            .n6011(n6011), .n6010(n6010), .n6009(n6009), .n6008(n6008), 
            .n6007(n6007), .\REG.mem_63_10 (\REG.mem_63_10 ), .n6006(n6006), 
            .n6005(n6005), .n6004(n6004), .\REG.mem_63_7 (\REG.mem_63_7 ), 
            .n6003(n6003), .n6002(n6002), .\REG.mem_63_5 (\REG.mem_63_5 ), 
            .\REG.mem_48_9 (\REG.mem_48_9 ), .\REG.mem_42_13 (\REG.mem_42_13 ), 
            .\REG.mem_43_13 (\REG.mem_43_13 ), .\REG.mem_38_0 (\REG.mem_38_0 ), 
            .\REG.mem_39_0 (\REG.mem_39_0 ), .n6001(n6001), .\REG.mem_63_4 (\REG.mem_63_4 ), 
            .n6000(n6000), .\REG.mem_63_3 (\REG.mem_63_3 ), .n5999(n5999), 
            .\REG.mem_63_2 (\REG.mem_63_2 ), .n5998(n5998), .n5997(n5997), 
            .\REG.mem_63_0 (\REG.mem_63_0 ), .n5996(n5996), .n5995(n5995), 
            .n5994(n5994), .n5993(n5993), .n5992(n5992), .n5991(n5991), 
            .\REG.mem_62_10 (\REG.mem_62_10 ), .n5990(n5990), .n5989(n5989), 
            .n5988(n5988), .\REG.mem_62_7 (\REG.mem_62_7 ), .n5987(n5987), 
            .n5986(n5986), .\REG.mem_62_5 (\REG.mem_62_5 ), .n5985(n5985), 
            .\REG.mem_62_4 (\REG.mem_62_4 ), .\REG.mem_41_13 (\REG.mem_41_13 ), 
            .\REG.mem_40_13 (\REG.mem_40_13 ), .\REG.mem_37_0 (\REG.mem_37_0 ), 
            .\REG.mem_36_0 (\REG.mem_36_0 ), .\REG.mem_10_6 (\REG.mem_10_6 ), 
            .\REG.mem_11_6 (\REG.mem_11_6 ), .n5984(n5984), .\REG.mem_62_3 (\REG.mem_62_3 ), 
            .n5983(n5983), .\REG.mem_62_2 (\REG.mem_62_2 ), .n5982(n5982), 
            .n5981(n5981), .\REG.mem_62_0 (\REG.mem_62_0 ), .\REG.mem_9_6 (\REG.mem_9_6 ), 
            .\REG.mem_8_6 (\REG.mem_8_6 ), .\REG.mem_42_0 (\REG.mem_42_0 ), 
            .\REG.mem_43_0 (\REG.mem_43_0 ), .\REG.mem_22_8 (\REG.mem_22_8 ), 
            .\REG.mem_23_8 (\REG.mem_23_8 ), .n5946(n5946), .rp_sync1_r({rp_sync1_r}), 
            .n5945(n5945), .n5944(n5944), .n5943(n5943), .n5942(n5942), 
            .n5941(n5941), .n5940(n5940), .n5939(n5939), .n5938(n5938), 
            .n5921(n5921), .n5920(n5920), .n5919(n5919), .\REG.mem_41_0 (\REG.mem_41_0 ), 
            .\REG.mem_40_0 (\REG.mem_40_0 ), .n5917(n5917), .n5916(n5916), 
            .n5914(n5914), .\REG.mem_8_14 (\REG.mem_8_14 ), .\REG.mem_9_14 (\REG.mem_9_14 ), 
            .\REG.mem_25_1 (\REG.mem_25_1 ), .\REG.mem_10_14 (\REG.mem_10_14 ), 
            .\REG.mem_11_14 (\REG.mem_11_14 ), .n5894(n5894), .n5893(n5893), 
            .n5892(n5892), .n5891(n5891), .\REG.mem_57_12 (\REG.mem_57_12 ), 
            .n5890(n5890), .n5889(n5889), .\REG.mem_57_10 (\REG.mem_57_10 ), 
            .n5888(n5888), .n5887(n5887), .n5886(n5886), .\REG.mem_57_7 (\REG.mem_57_7 ), 
            .\REG.mem_6_8 (\REG.mem_6_8 ), .\REG.mem_7_8 (\REG.mem_7_8 ), 
            .\REG.mem_38_15 (\REG.mem_38_15 ), .\REG.mem_39_15 (\REG.mem_39_15 ), 
            .n5885(n5885), .\REG.mem_5_8 (\REG.mem_5_8 ), .\REG.mem_4_8 (\REG.mem_4_8 ), 
            .\REG.mem_14_14 (\REG.mem_14_14 ), .\REG.mem_15_14 (\REG.mem_15_14 ), 
            .n5884(n5884), .\REG.mem_57_5 (\REG.mem_57_5 ), .n5883(n5883), 
            .\REG.mem_57_4 (\REG.mem_57_4 ), .n5882(n5882), .\REG.mem_57_3 (\REG.mem_57_3 ), 
            .n5881(n5881), .\REG.mem_57_2 (\REG.mem_57_2 ), .n5880(n5880), 
            .n5879(n5879), .\REG.mem_57_0 (\REG.mem_57_0 ), .\REG.mem_12_14 (\REG.mem_12_14 ), 
            .\REG.mem_13_14 (\REG.mem_13_14 ), .\REG.mem_37_15 (\REG.mem_37_15 ), 
            .\REG.mem_36_15 (\REG.mem_36_15 ), .n5861(n5861), .wp_sync1_r({wp_sync1_r}), 
            .n5860(n5860), .n5859(n5859), .n5858(n5858), .n5857(n5857), 
            .n5856(n5856), .n5855(n5855), .\REG.mem_55_15 (\REG.mem_55_15 ), 
            .n5854(n5854), .\REG.mem_55_14 (\REG.mem_55_14 ), .n5853(n5853), 
            .\rd_sig_diff0_w[0] (rd_sig_diff0_w[0]), .n5852(n5852), .n5851(n5851), 
            .n5850(n5850), .n5849(n5849), .n5848(n5848), .\REG.mem_55_8 (\REG.mem_55_8 ), 
            .n5847(n5847), .n5846(n5846), .\REG.mem_55_6 (\REG.mem_55_6 ), 
            .n5845(n5845), .\REG.mem_55_5 (\REG.mem_55_5 ), .n5844(n5844), 
            .\REG.mem_55_4 (\REG.mem_55_4 ), .n5843(n5843), .\REG.mem_55_3 (\REG.mem_55_3 ), 
            .n5842(n5842), .\REG.mem_55_2 (\REG.mem_55_2 ), .n5841(n5841), 
            .\REG.mem_55_1 (\REG.mem_55_1 ), .n5840(n5840), .\REG.mem_55_0 (\REG.mem_55_0 ), 
            .n5839(n5839), .n5838(n5838), .\REG.mem_40_4 (\REG.mem_40_4 ), 
            .\REG.mem_41_4 (\REG.mem_41_4 ), .\REG.mem_42_4 (\REG.mem_42_4 ), 
            .\REG.mem_43_4 (\REG.mem_43_4 ), .n5836(n5836), .n5835(n5835), 
            .n5834(n5834), .n5833(n5833), .n5832(n5832), .\REG.mem_54_15 (\REG.mem_54_15 ), 
            .n5831(n5831), .\REG.mem_54_14 (\REG.mem_54_14 ), .n5830(n5830), 
            .n5829(n5829), .n5828(n5828), .n5827(n5827), .n5826(n5826), 
            .n5825(n5825), .\REG.mem_54_8 (\REG.mem_54_8 ), .n5824(n5824), 
            .n5823(n5823), .\REG.mem_54_6 (\REG.mem_54_6 ), .n5822(n5822), 
            .\REG.mem_54_5 (\REG.mem_54_5 ), .n5821(n5821), .\REG.mem_54_4 (\REG.mem_54_4 ), 
            .\REG.mem_46_4 (\REG.mem_46_4 ), .\REG.mem_47_4 (\REG.mem_47_4 ), 
            .\REG.mem_44_4 (\REG.mem_44_4 ), .\REG.mem_45_4 (\REG.mem_45_4 ), 
            .n5820(n5820), .\REG.mem_54_3 (\REG.mem_54_3 ), .n5819(n5819), 
            .\REG.mem_54_2 (\REG.mem_54_2 ), .n5818(n5818), .\REG.mem_54_1 (\REG.mem_54_1 ), 
            .n5817(n5817), .\REG.mem_54_0 (\REG.mem_54_0 ), .\REG.mem_25_4 (\REG.mem_25_4 ), 
            .\REG.mem_30_4 (\REG.mem_30_4 ), .\REG.mem_31_4 (\REG.mem_31_4 ), 
            .\REG.mem_8_4 (\REG.mem_8_4 ), .\REG.mem_9_4 (\REG.mem_9_4 ), 
            .\REG.mem_10_4 (\REG.mem_10_4 ), .\REG.mem_11_4 (\REG.mem_11_4 ), 
            .\REG.mem_14_4 (\REG.mem_14_4 ), .\REG.mem_15_4 (\REG.mem_15_4 ), 
            .\REG.mem_12_4 (\REG.mem_12_4 ), .\REG.mem_13_4 (\REG.mem_13_4 ), 
            .n5768(n5768), .\REG.mem_50_15 (\REG.mem_50_15 ), .n5767(n5767), 
            .\REG.mem_50_14 (\REG.mem_50_14 ), .n5766(n5766), .\REG.mem_50_13 (\REG.mem_50_13 ), 
            .n5765(n5765), .n5764(n5764), .n5763(n5763), .n5762(n5762), 
            .n5761(n5761), .\REG.mem_50_8 (\REG.mem_50_8 ), .n5760(n5760), 
            .n5759(n5759), .\REG.mem_50_6 (\REG.mem_50_6 ), .n5758(n5758), 
            .\REG.mem_50_5 (\REG.mem_50_5 ), .n5757(n5757), .\REG.mem_50_4 (\REG.mem_50_4 ), 
            .n10700(n10700), .n5756(n5756), .\REG.mem_50_3 (\REG.mem_50_3 ), 
            .n5755(n5755), .\REG.mem_50_2 (\REG.mem_50_2 ), .n5754(n5754), 
            .n4893(n4893), .\fifo_data_out[14] (fifo_data_out[14]), .n4896(n4896), 
            .\fifo_data_out[15] (fifo_data_out[15]), .n5750(n5750), .\REG.mem_50_0 (\REG.mem_50_0 ), 
            .\REG.mem_38_5 (\REG.mem_38_5 ), .\REG.mem_39_5 (\REG.mem_39_5 ), 
            .n5733(n5733), .\REG.mem_48_15 (\REG.mem_48_15 ), .n5732(n5732), 
            .\REG.mem_48_14 (\REG.mem_48_14 ), .n5731(n5731), .\REG.mem_48_13 (\REG.mem_48_13 ), 
            .n5730(n5730), .n5729(n5729), .n5728(n5728), .n5727(n5727), 
            .n5726(n5726), .\REG.mem_48_8 (\REG.mem_48_8 ), .n5725(n5725), 
            .n5724(n5724), .\REG.mem_48_6 (\REG.mem_48_6 ), .n10748(n10748), 
            .n5723(n5723), .\REG.mem_48_5 (\REG.mem_48_5 ), .n5722(n5722), 
            .\REG.mem_48_4 (\REG.mem_48_4 ), .n5721(n5721), .\REG.mem_48_3 (\REG.mem_48_3 ), 
            .n5720(n5720), .\REG.mem_48_2 (\REG.mem_48_2 ), .n5719(n5719), 
            .\REG.mem_42_6 (\REG.mem_42_6 ), .\REG.mem_43_6 (\REG.mem_43_6 ), 
            .n5718(n5718), .\REG.mem_48_0 (\REG.mem_48_0 ), .n5717(n5717), 
            .\REG.mem_47_15 (\REG.mem_47_15 ), .\REG.mem_41_6 (\REG.mem_41_6 ), 
            .\REG.mem_40_6 (\REG.mem_40_6 ), .n5716(n5716), .\REG.mem_47_14 (\REG.mem_47_14 ), 
            .n5715(n5715), .\REG.mem_47_13 (\REG.mem_47_13 ), .n5714(n5714), 
            .n5713(n5713), .\REG.mem_47_11 (\REG.mem_47_11 ), .n5712(n5712), 
            .\REG.mem_47_10 (\REG.mem_47_10 ), .n5711(n5711), .n5710(n5710), 
            .n5709(n5709), .\REG.mem_47_7 (\REG.mem_47_7 ), .n5708(n5708), 
            .\REG.mem_47_6 (\REG.mem_47_6 ), .n5707(n5707), .n5706(n5706), 
            .n5705(n5705), .n5704(n5704), .n5703(n5703), .\REG.mem_25_12 (\REG.mem_25_12 ), 
            .\REG.mem_37_5 (\REG.mem_37_5 ), .\REG.mem_36_5 (\REG.mem_36_5 ), 
            .n5702(n5702), .\REG.mem_47_0 (\REG.mem_47_0 ), .n5701(n5701), 
            .\REG.mem_46_15 (\REG.mem_46_15 ), .n5700(n5700), .\REG.mem_46_14 (\REG.mem_46_14 ), 
            .n5699(n5699), .\REG.mem_46_13 (\REG.mem_46_13 ), .n5698(n5698), 
            .n5697(n5697), .\REG.mem_46_11 (\REG.mem_46_11 ), .n5696(n5696), 
            .\REG.mem_46_10 (\REG.mem_46_10 ), .n5695(n5695), .n5694(n5694), 
            .n5693(n5693), .\REG.mem_46_7 (\REG.mem_46_7 ), .n5692(n5692), 
            .\REG.mem_46_6 (\REG.mem_46_6 ), .n5691(n5691), .n5690(n5690), 
            .n5689(n5689), .n5688(n5688), .n5687(n5687), .n5686(n5686), 
            .\REG.mem_46_0 (\REG.mem_46_0 ), .n5685(n5685), .\REG.mem_45_15 (\REG.mem_45_15 ), 
            .n5684(n5684), .\REG.mem_45_14 (\REG.mem_45_14 ), .n5683(n5683), 
            .\REG.mem_45_13 (\REG.mem_45_13 ), .n5682(n5682), .n5681(n5681), 
            .\REG.mem_45_11 (\REG.mem_45_11 ), .n5680(n5680), .\REG.mem_45_10 (\REG.mem_45_10 ), 
            .n5679(n5679), .n5678(n5678), .\REG.mem_6_15 (\REG.mem_6_15 ), 
            .\REG.mem_7_15 (\REG.mem_7_15 ), .\REG.mem_3_1 (\REG.mem_3_1 ), 
            .n5677(n5677), .\REG.mem_45_7 (\REG.mem_45_7 ), .\REG.mem_5_15 (\REG.mem_5_15 ), 
            .\REG.mem_4_15 (\REG.mem_4_15 ), .n5676(n5676), .\REG.mem_45_6 (\REG.mem_45_6 ), 
            .n5675(n5675), .n5674(n5674), .n5673(n5673), .n5672(n5672), 
            .n5671(n5671), .n5670(n5670), .\REG.mem_45_0 (\REG.mem_45_0 ), 
            .n5668(n5668), .\REG.mem_44_15 (\REG.mem_44_15 ), .n5667(n5667), 
            .\REG.mem_44_14 (\REG.mem_44_14 ), .n5665(n5665), .\REG.mem_44_13 (\REG.mem_44_13 ), 
            .n5664(n5664), .n5663(n5663), .\REG.mem_44_11 (\REG.mem_44_11 ), 
            .n5661(n5661), .\REG.mem_44_10 (\REG.mem_44_10 ), .n5660(n5660), 
            .n5659(n5659), .n5658(n5658), .\REG.mem_44_7 (\REG.mem_44_7 ), 
            .n5657(n5657), .\REG.mem_44_6 (\REG.mem_44_6 ), .n5656(n5656), 
            .n5655(n5655), .n5654(n5654), .n5653(n5653), .n5652(n5652), 
            .n5651(n5651), .\REG.mem_44_0 (\REG.mem_44_0 ), .n5650(n5650), 
            .n5649(n5649), .\REG.mem_43_14 (\REG.mem_43_14 ), .n5648(n5648), 
            .n5647(n5647), .n5646(n5646), .\REG.mem_43_11 (\REG.mem_43_11 ), 
            .n5645(n5645), .\REG.mem_43_10 (\REG.mem_43_10 ), .n5644(n5644), 
            .\REG.mem_43_9 (\REG.mem_43_9 ), .\rd_addr_p1_w[0] (rd_addr_p1_w[0]), 
            .\REG.mem_18_7 (\REG.mem_18_7 ), .n5643(n5643), .n5642(n5642), 
            .\REG.mem_43_7 (\REG.mem_43_7 ), .n5641(n5641), .n5640(n5640), 
            .\REG.mem_43_5 (\REG.mem_43_5 ), .n5639(n5639), .n5638(n5638), 
            .\REG.mem_43_3 (\REG.mem_43_3 ), .n5637(n5637), .n5636(n5636), 
            .\REG.mem_43_1 (\REG.mem_43_1 ), .n5635(n5635), .n5634(n5634), 
            .n5633(n5633), .\REG.mem_42_14 (\REG.mem_42_14 ), .n5632(n5632), 
            .n5631(n5631), .n5630(n5630), .\REG.mem_42_11 (\REG.mem_42_11 ), 
            .n5629(n5629), .\REG.mem_42_10 (\REG.mem_42_10 ), .n4916(n4916), 
            .\REG.mem_22_11 (\REG.mem_22_11 ), .\REG.mem_23_11 (\REG.mem_23_11 ), 
            .n5628(n5628), .\REG.mem_42_9 (\REG.mem_42_9 ), .n5627(n5627), 
            .n5626(n5626), .\REG.mem_42_7 (\REG.mem_42_7 ), .n5625(n5625), 
            .n5624(n5624), .\REG.mem_42_5 (\REG.mem_42_5 ), .n5623(n5623), 
            .n5622(n5622), .\REG.mem_42_3 (\REG.mem_42_3 ), .n5621(n5621), 
            .n5620(n5620), .\REG.mem_42_1 (\REG.mem_42_1 ), .n5619(n5619), 
            .n5618(n5618), .\REG.mem_41_15 (\REG.mem_41_15 ), .n5617(n5617), 
            .\REG.mem_41_14 (\REG.mem_41_14 ), .n5616(n5616), .n5615(n5615), 
            .n5614(n5614), .\REG.mem_41_11 (\REG.mem_41_11 ), .n5613(n5613), 
            .\REG.mem_41_10 (\REG.mem_41_10 ), .\REG.mem_25_6 (\REG.mem_25_6 ), 
            .n5612(n5612), .\REG.mem_41_9 (\REG.mem_41_9 ), .n5611(n5611), 
            .n5610(n5610), .\REG.mem_41_7 (\REG.mem_41_7 ), .n5609(n5609), 
            .n5608(n5608), .\REG.mem_41_5 (\REG.mem_41_5 ), .n5607(n5607), 
            .n5606(n5606), .\REG.mem_41_3 (\REG.mem_41_3 ), .n5605(n5605), 
            .n5604(n5604), .\REG.mem_41_1 (\REG.mem_41_1 ), .n5603(n5603), 
            .n5602(n5602), .\REG.mem_40_15 (\REG.mem_40_15 ), .n5601(n5601), 
            .\REG.mem_40_14 (\REG.mem_40_14 ), .n5600(n5600), .n5599(n5599), 
            .n5598(n5598), .\REG.mem_40_11 (\REG.mem_40_11 ), .n5597(n5597), 
            .\REG.mem_40_10 (\REG.mem_40_10 ), .n4904(n4904), .n4903(n4903), 
            .n4901(n4901), .n4899(n4899), .n5596(n5596), .\REG.mem_40_9 (\REG.mem_40_9 ), 
            .n5595(n5595), .n5594(n5594), .\REG.mem_40_7 (\REG.mem_40_7 ), 
            .n5593(n5593), .n5592(n5592), .\REG.mem_40_5 (\REG.mem_40_5 ), 
            .n5591(n5591), .n5590(n5590), .\REG.mem_40_3 (\REG.mem_40_3 ), 
            .n5589(n5589), .n5588(n5588), .\REG.mem_40_1 (\REG.mem_40_1 ), 
            .n5587(n5587), .n5586(n5586), .n5585(n5585), .\REG.mem_39_14 (\REG.mem_39_14 ), 
            .n5584(n5584), .n5583(n5583), .\REG.mem_39_12 (\REG.mem_39_12 ), 
            .n5582(n5582), .\REG.mem_39_11 (\REG.mem_39_11 ), .n5581(n5581), 
            .\REG.mem_39_10 (\REG.mem_39_10 ), .n4898(n4898), .DEBUG_5_c(DEBUG_5_c), 
            .\REG.mem_3_4 (\REG.mem_3_4 ), .\REG.mem_6_4 (\REG.mem_6_4 ), 
            .\REG.mem_7_4 (\REG.mem_7_4 ), .n5580(n5580), .\REG.mem_39_9 (\REG.mem_39_9 ), 
            .n5579(n5579), .\REG.mem_39_8 (\REG.mem_39_8 ), .n5578(n5578), 
            .n5577(n5577), .n5576(n5576), .n5575(n5575), .\REG.mem_39_4 (\REG.mem_39_4 ), 
            .n5574(n5574), .\REG.mem_39_3 (\REG.mem_39_3 ), .n5573(n5573), 
            .\REG.mem_39_2 (\REG.mem_39_2 ), .n5572(n5572), .\REG.mem_39_1 (\REG.mem_39_1 ), 
            .n5570(n5570), .n5569(n5569), .n5568(n5568), .\REG.mem_38_14 (\REG.mem_38_14 ), 
            .n5567(n5567), .n5566(n5566), .\REG.mem_38_12 (\REG.mem_38_12 ), 
            .n5565(n5565), .\REG.mem_38_11 (\REG.mem_38_11 ), .n5564(n5564), 
            .\REG.mem_38_10 (\REG.mem_38_10 ), .\REG.mem_5_4 (\REG.mem_5_4 ), 
            .\REG.mem_4_4 (\REG.mem_4_4 ), .n5563(n5563), .\REG.mem_38_9 (\REG.mem_38_9 ), 
            .n5562(n5562), .\REG.mem_38_8 (\REG.mem_38_8 ), .n5561(n5561), 
            .n5560(n5560), .n5559(n5559), .n5558(n5558), .\REG.mem_38_4 (\REG.mem_38_4 ), 
            .n5557(n5557), .\REG.mem_38_3 (\REG.mem_38_3 ), .n5556(n5556), 
            .\REG.mem_38_2 (\REG.mem_38_2 ), .n5555(n5555), .\REG.mem_38_1 (\REG.mem_38_1 ), 
            .n5554(n5554), .n5553(n5553), .n5552(n5552), .\REG.mem_37_14 (\REG.mem_37_14 ), 
            .n5551(n5551), .n5550(n5550), .\REG.mem_37_12 (\REG.mem_37_12 ), 
            .n5549(n5549), .\REG.mem_37_11 (\REG.mem_37_11 ), .\REG.out_raw[15] (\REG.out_raw [15]), 
            .\REG.out_raw[14] (\REG.out_raw [14]), .\REG.out_raw[13] (\REG.out_raw [13]), 
            .\REG.out_raw[12] (\REG.out_raw [12]), .\REG.out_raw[11] (\REG.out_raw [11]), 
            .n5548(n5548), .\REG.mem_37_10 (\REG.mem_37_10 ), .n5547(n5547), 
            .\REG.mem_37_9 (\REG.mem_37_9 ), .n5546(n5546), .\REG.mem_37_8 (\REG.mem_37_8 ), 
            .n5545(n5545), .n5544(n5544), .n5543(n5543), .n5542(n5542), 
            .\REG.mem_37_4 (\REG.mem_37_4 ), .n5541(n5541), .\REG.mem_37_3 (\REG.mem_37_3 ), 
            .n5540(n5540), .\REG.mem_37_2 (\REG.mem_37_2 ), .n5539(n5539), 
            .\REG.mem_37_1 (\REG.mem_37_1 ), .n5538(n5538), .\REG.out_raw[10] (\REG.out_raw [10]), 
            .\REG.out_raw[9] (\REG.out_raw [9]), .\REG.out_raw[8] (\REG.out_raw [8]), 
            .\REG.out_raw[7] (\REG.out_raw [7]), .\REG.out_raw[6] (\REG.out_raw [6]), 
            .\REG.out_raw[5] (\REG.out_raw [5]), .\REG.out_raw[4] (\REG.out_raw [4]), 
            .\REG.out_raw[3] (\REG.out_raw [3]), .\REG.out_raw[2] (\REG.out_raw [2]), 
            .\REG.out_raw[1] (\REG.out_raw [1]), .n5524(n5524), .n5523(n5523), 
            .\REG.mem_36_14 (\REG.mem_36_14 ), .n5522(n5522), .n5521(n5521), 
            .\REG.mem_36_12 (\REG.mem_36_12 ), .n5520(n5520), .\REG.mem_36_11 (\REG.mem_36_11 ), 
            .n5519(n5519), .\REG.mem_36_10 (\REG.mem_36_10 ), .n5518(n5518), 
            .\REG.mem_36_9 (\REG.mem_36_9 ), .n5517(n5517), .\REG.mem_36_8 (\REG.mem_36_8 ), 
            .n5516(n5516), .\rd_sig_diff0_w[2] (rd_sig_diff0_w[2]), .n5515(n5515), 
            .n5514(n5514), .n5513(n5513), .\REG.mem_36_4 (\REG.mem_36_4 ), 
            .n5512(n5512), .\REG.mem_36_3 (\REG.mem_36_3 ), .n5511(n5511), 
            .\REG.mem_36_2 (\REG.mem_36_2 ), .n5510(n5510), .\REG.mem_36_1 (\REG.mem_36_1 ), 
            .n5509(n5509), .n5505(n5505), .n5504(n5504), .\REG.mem_35_14 (\REG.mem_35_14 ), 
            .n5503(n5503), .n5502(n5502), .\REG.mem_35_12 (\REG.mem_35_12 ), 
            .n5501(n5501), .\REG.mem_35_11 (\REG.mem_35_11 ), .n5500(n5500), 
            .\REG.mem_35_10 (\REG.mem_35_10 ), .\rd_sig_diff0_w[1] (rd_sig_diff0_w[1]), 
            .n5499(n5499), .n5498(n5498), .\REG.mem_35_8 (\REG.mem_35_8 ), 
            .n5497(n5497), .n5496(n5496), .n5495(n5495), .\REG.mem_35_5 (\REG.mem_35_5 ), 
            .n5494(n5494), .\REG.mem_35_4 (\REG.mem_35_4 ), .n5493(n5493), 
            .\REG.mem_35_3 (\REG.mem_35_3 ), .n5492(n5492), .\REG.mem_35_2 (\REG.mem_35_2 ), 
            .n5491(n5491), .\REG.mem_35_1 (\REG.mem_35_1 ), .n5490(n5490), 
            .\REG.mem_25_11 (\REG.mem_25_11 ), .\REG.mem_10_13 (\REG.mem_10_13 ), 
            .\REG.mem_11_13 (\REG.mem_11_13 ), .\REG.mem_9_13 (\REG.mem_9_13 ), 
            .\REG.mem_8_13 (\REG.mem_8_13 ), .n5440(n5440), .n5439(n5439), 
            .\REG.mem_31_14 (\REG.mem_31_14 ), .n5438(n5438), .n5437(n5437), 
            .\REG.mem_31_12 (\REG.mem_31_12 ), .n5436(n5436), .\REG.mem_31_11 (\REG.mem_31_11 ), 
            .n5435(n5435), .\REG.mem_31_10 (\REG.mem_31_10 ), .n5434(n5434), 
            .n5433(n5433), .\REG.mem_31_8 (\REG.mem_31_8 ), .n5432(n5432), 
            .\REG.mem_31_7 (\REG.mem_31_7 ), .n5431(n5431), .\REG.mem_31_6 (\REG.mem_31_6 ), 
            .n5430(n5430), .n5429(n5429), .n5428(n5428), .\REG.mem_31_3 (\REG.mem_31_3 ), 
            .n5427(n5427), .n5426(n5426), .\REG.mem_31_1 (\REG.mem_31_1 ), 
            .n5425(n5425), .n5424(n5424), .n5423(n5423), .\REG.mem_30_14 (\REG.mem_30_14 ), 
            .n5422(n5422), .n5421(n5421), .\REG.mem_30_12 (\REG.mem_30_12 ), 
            .n5420(n5420), .\REG.mem_30_11 (\REG.mem_30_11 ), .DEBUG_1_c_c(DEBUG_1_c_c), 
            .write_to_dc32_fifo_latched_N_425(write_to_dc32_fifo_latched_N_425), 
            .\REG.mem_18_6 (\REG.mem_18_6 ), .n5419(n5419), .\REG.mem_30_10 (\REG.mem_30_10 ), 
            .n5418(n5418), .n5417(n5417), .\REG.mem_30_8 (\REG.mem_30_8 ), 
            .n5416(n5416), .\REG.mem_30_7 (\REG.mem_30_7 ), .n5415(n5415), 
            .\REG.mem_30_6 (\REG.mem_30_6 ), .n5414(n5414), .n5413(n5413), 
            .n5412(n5412), .\REG.mem_30_3 (\REG.mem_30_3 ), .n5411(n5411), 
            .n5410(n5410), .\REG.mem_30_1 (\REG.mem_30_1 ), .n5409(n5409), 
            .\REG.mem_16_6 (\REG.mem_16_6 ), .\wr_addr_nxt_c[1] (wr_addr_nxt_c[1]), 
            .\REG.mem_10_9 (\REG.mem_10_9 ), .\REG.mem_11_9 (\REG.mem_11_9 ), 
            .\REG.mem_9_9 (\REG.mem_9_9 ), .\REG.mem_8_9 (\REG.mem_8_9 ), 
            .\REG.mem_14_13 (\REG.mem_14_13 ), .\REG.mem_15_13 (\REG.mem_15_13 ), 
            .\REG.mem_13_13 (\REG.mem_13_13 ), .\REG.mem_12_13 (\REG.mem_12_13 ), 
            .n56(n56), .\REG.mem_14_9 (\REG.mem_14_9 ), .\REG.mem_15_9 (\REG.mem_15_9 ), 
            .\REG.mem_10_15 (\REG.mem_10_15 ), .\REG.mem_11_15 (\REG.mem_11_15 ), 
            .\REG.mem_9_15 (\REG.mem_9_15 ), .\REG.mem_8_15 (\REG.mem_8_15 ), 
            .\REG.mem_10_7 (\REG.mem_10_7 ), .\REG.mem_11_7 (\REG.mem_11_7 ), 
            .\REG.mem_13_9 (\REG.mem_13_9 ), .\REG.mem_12_9 (\REG.mem_12_9 ), 
            .n5344(n5344), .n5343(n5343), .\REG.mem_25_14 (\REG.mem_25_14 ), 
            .n5342(n5342), .n5341(n5341), .n5340(n5340), .n5339(n5339), 
            .\REG.mem_25_10 (\REG.mem_25_10 ), .n5338(n5338), .n5337(n5337), 
            .\REG.mem_25_8 (\REG.mem_25_8 ), .n5336(n5336), .\REG.mem_25_7 (\REG.mem_25_7 ), 
            .\REG.mem_18_13 (\REG.mem_18_13 ), .\REG.mem_9_7 (\REG.mem_9_7 ), 
            .\REG.mem_8_7 (\REG.mem_8_7 ), .\REG.mem_16_13 (\REG.mem_16_13 ), 
            .n5335(n5335), .n5334(n5334), .n5333(n5333), .n5332(n5332), 
            .\REG.mem_25_3 (\REG.mem_25_3 ), .n5331(n5331), .n5330(n5330), 
            .n5329(n5329), .\REG.mem_25_0 (\REG.mem_25_0 ), .n52(n52), 
            .n20(n20), .n5306(n5306), .\REG.mem_23_15 (\REG.mem_23_15 ), 
            .n5305(n5305), .\REG.mem_23_14 (\REG.mem_23_14 ), .n5304(n5304), 
            .\REG.mem_23_13 (\REG.mem_23_13 ), .n5303(n5303), .n5302(n5302), 
            .n5301(n5301), .\REG.mem_23_10 (\REG.mem_23_10 ), .n5300(n5300), 
            .\REG.mem_23_9 (\REG.mem_23_9 ), .n5299(n5299), .n5298(n5298), 
            .n5297(n5297), .\REG.mem_23_6 (\REG.mem_23_6 ), .n5296(n5296), 
            .\REG.mem_23_5 (\REG.mem_23_5 ), .n5295(n5295), .\REG.mem_23_4 (\REG.mem_23_4 ), 
            .n5294(n5294), .\REG.mem_23_3 (\REG.mem_23_3 ), .n5293(n5293), 
            .\REG.mem_23_2 (\REG.mem_23_2 ), .n5292(n5292), .\REG.mem_23_1 (\REG.mem_23_1 ), 
            .n5291(n5291), .\REG.mem_23_0 (\REG.mem_23_0 ), .n5290(n5290), 
            .\REG.mem_22_15 (\REG.mem_22_15 ), .n5289(n5289), .\REG.mem_22_14 (\REG.mem_22_14 ), 
            .n5288(n5288), .\REG.mem_22_13 (\REG.mem_22_13 ), .n5287(n5287), 
            .n5286(n5286), .n5285(n5285), .\REG.mem_22_10 (\REG.mem_22_10 ), 
            .\rd_grey_sync_r[5] (rd_grey_sync_r[5]), .\rd_grey_sync_r[4] (rd_grey_sync_r[4]), 
            .\rd_grey_sync_r[3] (rd_grey_sync_r[3]), .\rd_grey_sync_r[2] (rd_grey_sync_r[2]), 
            .\rd_grey_sync_r[1] (rd_grey_sync_r[1]), .n5284(n5284), .\REG.mem_22_9 (\REG.mem_22_9 ), 
            .n5283(n5283), .n5282(n5282), .n5281(n5281), .\REG.mem_22_6 (\REG.mem_22_6 ), 
            .n5280(n5280), .\REG.mem_22_5 (\REG.mem_22_5 ), .n5279(n5279), 
            .\REG.mem_22_4 (\REG.mem_22_4 ), .n5278(n5278), .\REG.mem_22_3 (\REG.mem_22_3 ), 
            .n5277(n5277), .\REG.mem_22_2 (\REG.mem_22_2 ), .n5276(n5276), 
            .\REG.mem_22_1 (\REG.mem_22_1 ), .n5275(n5275), .\REG.mem_22_0 (\REG.mem_22_0 ), 
            .\REG.mem_14_3 (\REG.mem_14_3 ), .\REG.mem_15_3 (\REG.mem_15_3 ), 
            .\REG.mem_13_3 (\REG.mem_13_3 ), .\REG.mem_12_3 (\REG.mem_12_3 ), 
            .\REG.mem_10_8 (\REG.mem_10_8 ), .\REG.mem_11_8 (\REG.mem_11_8 ), 
            .\REG.mem_9_8 (\REG.mem_9_8 ), .\REG.mem_8_8 (\REG.mem_8_8 ), 
            .get_next_word(get_next_word), .\REG.mem_16_2 (\REG.mem_16_2 ), 
            .\REG.mem_18_2 (\REG.mem_18_2 ), .\REG.mem_18_3 (\REG.mem_18_3 ), 
            .n5226(n5226), .\REG.mem_18_15 (\REG.mem_18_15 ), .n5225(n5225), 
            .\REG.mem_18_14 (\REG.mem_18_14 ), .n5224(n5224), .n5223(n5223), 
            .n5222(n5222), .n5221(n5221), .\REG.mem_18_10 (\REG.mem_18_10 ), 
            .n5220(n5220), .\REG.mem_18_9 (\REG.mem_18_9 ), .rd_fifo_en_w(rd_fifo_en_w), 
            .\REG.mem_16_3 (\REG.mem_16_3 ), .\REG.mem_16_15 (\REG.mem_16_15 ), 
            .n5219(n5219), .n5218(n5218), .n5217(n5217), .n5216(n5216), 
            .n5215(n5215), .\REG.mem_18_4 (\REG.mem_18_4 ), .n5214(n5214), 
            .n5213(n5213), .n5212(n5212), .\REG.mem_18_1 (\REG.mem_18_1 ), 
            .n5211(n5211), .\REG.mem_18_0 (\REG.mem_18_0 ), .n5190(n5190), 
            .n5188(n5188), .\REG.mem_16_14 (\REG.mem_16_14 ), .n5187(n5187), 
            .n5186(n5186), .n5185(n5185), .n5184(n5184), .\REG.mem_16_10 (\REG.mem_16_10 ), 
            .\REG.mem_3_2 (\REG.mem_3_2 ), .\REG.mem_3_0 (\REG.mem_3_0 ), 
            .n5183(n5183), .\REG.mem_16_9 (\REG.mem_16_9 ), .n5182(n5182), 
            .n5181(n5181), .n5180(n5180), .n5179(n5179), .n5178(n5178), 
            .\REG.mem_16_4 (\REG.mem_16_4 ), .n5177(n5177), .n5176(n5176), 
            .\REG.mem_6_0 (\REG.mem_6_0 ), .\REG.mem_7_0 (\REG.mem_7_0 ), 
            .n5175(n5175), .\REG.mem_16_1 (\REG.mem_16_1 ), .n5174(n5174), 
            .\REG.mem_16_0 (\REG.mem_16_0 ), .n5171(n5171), .\REG.mem_15_15 (\REG.mem_15_15 ), 
            .n5170(n5170), .n5169(n5169), .n5168(n5168), .n5167(n5167), 
            .n5166(n5166), .\REG.mem_15_10 (\REG.mem_15_10 ), .n5165(n5165), 
            .n5164(n5164), .n5163(n5163), .n5162(n5162), .\REG.mem_15_6 (\REG.mem_15_6 ), 
            .\REG.mem_5_0 (\REG.mem_5_0 ), .\REG.mem_4_0 (\REG.mem_4_0 ), 
            .n5161(n5161), .n5160(n5160), .n5159(n5159), .n5158(n5158), 
            .n5157(n5157), .\REG.mem_15_1 (\REG.mem_15_1 ), .n5156(n5156), 
            .\REG.mem_15_0 (\REG.mem_15_0 ), .n5155(n5155), .\REG.mem_14_15 (\REG.mem_14_15 ), 
            .n5154(n5154), .n5153(n5153), .n5152(n5152), .n5151(n5151), 
            .n5150(n5150), .\REG.mem_14_10 (\REG.mem_14_10 ), .n5149(n5149), 
            .n5148(n5148), .n5147(n5147), .n5146(n5146), .\REG.mem_14_6 (\REG.mem_14_6 ), 
            .n5145(n5145), .n5144(n5144), .n5143(n5143), .n5142(n5142), 
            .n5141(n5141), .\REG.mem_14_1 (\REG.mem_14_1 ), .n5140(n5140), 
            .\REG.mem_14_0 (\REG.mem_14_0 ), .n5139(n5139), .\REG.mem_13_15 (\REG.mem_13_15 ), 
            .n5138(n5138), .n5137(n5137), .n5136(n5136), .n5135(n5135), 
            .n5134(n5134), .\REG.mem_13_10 (\REG.mem_13_10 ), .n5133(n5133), 
            .n5132(n5132), .n5131(n5131), .n47(n47), .n15(n15_adj_1224), 
            .n50(n50), .n5130(n5130), .\REG.mem_13_6 (\REG.mem_13_6 ), 
            .n18(n18), .n5129(n5129), .n5128(n5128), .n5127(n5127), 
            .n5126(n5126), .n5125(n5125), .\REG.mem_13_1 (\REG.mem_13_1 ), 
            .n5124(n5124), .\REG.mem_13_0 (\REG.mem_13_0 ), .n5123(n5123), 
            .\REG.mem_12_15 (\REG.mem_12_15 ), .n5122(n5122), .n5121(n5121), 
            .n5120(n5120), .n5119(n5119), .n5118(n5118), .\REG.mem_12_10 (\REG.mem_12_10 ), 
            .n5117(n5117), .n5116(n5116), .\REG.mem_3_12 (\REG.mem_3_12 ), 
            .\REG.mem_3_14 (\REG.mem_3_14 ), .n5115(n5115), .n5114(n5114), 
            .\REG.mem_12_6 (\REG.mem_12_6 ), .n5113(n5113), .n5112(n5112), 
            .n53(n53), .n21(n21), .\REG.mem_10_0 (\REG.mem_10_0 ), .\REG.mem_11_0 (\REG.mem_11_0 ), 
            .\REG.mem_9_0 (\REG.mem_9_0 ), .\REG.mem_8_0 (\REG.mem_8_0 ), 
            .n5111(n5111), .n5110(n5110), .n5109(n5109), .\REG.mem_12_1 (\REG.mem_12_1 ), 
            .n5108(n5108), .\REG.mem_12_0 (\REG.mem_12_0 ), .n51(n51), 
            .n19(n19), .n5107(n5107), .n54(n54), .n22(n22), .n5106(n5106), 
            .n5105(n5105), .n5104(n5104), .\REG.mem_11_12 (\REG.mem_11_12 ), 
            .n5103(n5103), .n5102(n5102), .\REG.mem_11_10 (\REG.mem_11_10 ), 
            .n5101(n5101), .n5100(n5100), .n5099(n5099), .n5098(n5098), 
            .n5097(n5097), .\REG.mem_11_5 (\REG.mem_11_5 ), .\rd_addr_nxt_c_6__N_498[5] (rd_addr_nxt_c_6__N_498[5]), 
            .n5096(n5096), .n5095(n5095), .n5094(n5094), .n5093(n5093), 
            .\REG.mem_11_1 (\REG.mem_11_1 ), .n5092(n5092), .n5091(n5091), 
            .n5090(n5090), .n5089(n5089), .n5088(n5088), .\REG.mem_10_12 (\REG.mem_10_12 ), 
            .n5087(n5087), .n5086(n5086), .\REG.mem_10_10 (\REG.mem_10_10 ), 
            .n5085(n5085), .n5084(n5084), .n5083(n5083), .n5082(n5082), 
            .n5081(n5081), .\REG.mem_10_5 (\REG.mem_10_5 ), .n5080(n5080), 
            .\rd_addr_nxt_c_6__N_498[3] (rd_addr_nxt_c_6__N_498[3]), .n5079(n5079), 
            .\rd_addr_nxt_c_6__N_498[2] (rd_addr_nxt_c_6__N_498[2]), .n49(n49), 
            .n17(n17), .\REG.mem_6_14 (\REG.mem_6_14 ), .\REG.mem_7_14 (\REG.mem_7_14 ), 
            .\REG.mem_4_14 (\REG.mem_4_14 ), .\REG.mem_5_14 (\REG.mem_5_14 ), 
            .n24(n24_adj_1225), .n5078(n5078), .\REG.mem_3_6 (\REG.mem_3_6 ), 
            .n5077(n5077), .\REG.mem_10_1 (\REG.mem_10_1 ), .n5076(n5076), 
            .n5075(n5075), .\REG.mem_3_9 (\REG.mem_3_9 ), .n5074(n5074), 
            .n5073(n5073), .n55(n55), .n23(n23), .n40(n40), .n8(n8_adj_1223), 
            .n5072(n5072), .\REG.mem_9_12 (\REG.mem_9_12 ), .n34(n34), 
            .n5071(n5071), .n5070(n5070), .\REG.mem_9_10 (\REG.mem_9_10 ), 
            .n5069(n5069), .n2(n2), .n5068(n5068), .n5067(n5067), .n5066(n5066), 
            .n5065(n5065), .\REG.mem_9_5 (\REG.mem_9_5 ), .n5064(n5064), 
            .n5063(n5063), .n5062(n5062), .n5061(n5061), .\REG.mem_9_1 (\REG.mem_9_1 ), 
            .n5060(n5060), .n5059(n5059), .n5058(n5058), .n5057(n5057), 
            .n5056(n5056), .\REG.mem_8_12 (\REG.mem_8_12 ), .n5055(n5055), 
            .n5054(n5054), .\REG.mem_8_10 (\REG.mem_8_10 ), .n5053(n5053), 
            .n5052(n5052), .n5051(n5051), .n5050(n5050), .n5049(n5049), 
            .\REG.mem_8_5 (\REG.mem_8_5 ), .n5048(n5048), .n5047(n5047), 
            .n5046(n5046), .n5045(n5045), .\REG.mem_8_1 (\REG.mem_8_1 ), 
            .n5044(n5044), .n5043(n5043), .n5042(n5042), .n5041(n5041), 
            .\REG.mem_7_13 (\REG.mem_7_13 ), .n5040(n5040), .\REG.mem_7_12 (\REG.mem_7_12 ), 
            .n5039(n5039), .n5038(n5038), .\REG.mem_7_10 (\REG.mem_7_10 ), 
            .n5037(n5037), .n5036(n5036), .n5035(n5035), .\REG.mem_7_7 (\REG.mem_7_7 ), 
            .n5034(n5034), .\REG.mem_7_6 (\REG.mem_7_6 ), .n5033(n5033), 
            .n5032(n5032), .n5031(n5031), .n5030(n5030), .n5029(n5029), 
            .n5028(n5028), .n5027(n5027), .n5026(n5026), .n5025(n5025), 
            .\REG.mem_6_13 (\REG.mem_6_13 ), .n5024(n5024), .\REG.mem_6_12 (\REG.mem_6_12 ), 
            .n5023(n5023), .n5022(n5022), .\REG.mem_6_10 (\REG.mem_6_10 ), 
            .n5021(n5021), .n5020(n5020), .n5019(n5019), .\REG.mem_6_7 (\REG.mem_6_7 ), 
            .n5018(n5018), .\REG.mem_6_6 (\REG.mem_6_6 ), .n5017(n5017), 
            .n5016(n5016), .n5015(n5015), .n5014(n5014), .n5013(n5013), 
            .n5012(n5012), .n5011(n5011), .n5010(n5010), .n5009(n5009), 
            .\REG.mem_5_13 (\REG.mem_5_13 ), .n5008(n5008), .\REG.mem_5_12 (\REG.mem_5_12 ), 
            .n5007(n5007), .n5006(n5006), .\REG.mem_5_10 (\REG.mem_5_10 ), 
            .n5005(n5005), .n5004(n5004), .n5003(n5003), .\REG.mem_5_7 (\REG.mem_5_7 ), 
            .n5002(n5002), .\REG.mem_5_6 (\REG.mem_5_6 ), .n5001(n5001), 
            .n5000(n5000), .n4999(n4999), .n4998(n4998), .n4997(n4997), 
            .n4996(n4996), .n4995(n4995), .n4994(n4994), .n4993(n4993), 
            .\REG.mem_4_13 (\REG.mem_4_13 ), .n4992(n4992), .\REG.mem_4_12 (\REG.mem_4_12 ), 
            .n4991(n4991), .n4990(n4990), .\REG.mem_4_10 (\REG.mem_4_10 ), 
            .n4989(n4989), .n4988(n4988), .n4987(n4987), .\REG.mem_4_7 (\REG.mem_4_7 ), 
            .n4986(n4986), .\REG.mem_4_6 (\REG.mem_4_6 ), .n4985(n4985), 
            .n4984(n4984), .n4983(n4983), .n4982(n4982), .n4981(n4981), 
            .n4980(n4980), .n4979(n4979), .n4978(n4978), .n4977(n4977), 
            .\REG.mem_3_13 (\REG.mem_3_13 ), .n4976(n4976), .n4975(n4975), 
            .n4974(n4974), .\REG.mem_3_10 (\REG.mem_3_10 ), .n4973(n4973), 
            .n4972(n4972), .\REG.mem_3_8 (\REG.mem_3_8 ), .n4971(n4971), 
            .\REG.mem_3_7 (\REG.mem_3_7 ), .n4970(n4970), .n4969(n4969), 
            .FT_OE_N_420(FT_OE_N_420), .n57(n57), .n25(n25), .n42(n42), 
            .n10(n10), .n58(n58), .n26(n26), .n43(n43), .n35(n35), 
            .n11(n11), .n3(n3), .n4968(n4968), .n4967(n4967), .n4966(n4966), 
            .n4965(n4965), .n4964(n4964), .n60(n60), .n28(n28), .n59(n59), 
            .n27(n27), .n61(n61), .n29(n29), .n4672(n4672), .n4671(n4671), 
            .n4670(n4670), .n4669(n4669), .n4668(n4668), .n4667(n4667), 
            .n4666(n4666), .n4665(n4665), .n4664(n4664), .n4663(n4663), 
            .n4662(n4662), .n4661(n4661), .n4660(n4660), .n4659(n4659), 
            .n4658(n4658)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(547[21] 562[2])
    SB_LUT4 i3477_3_lut (.I0(tx_data_byte[1]), .I1(pc_data_rx[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4860));   // src/top.v(1074[8] 1141[4])
    defparam i3477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3714_3_lut (.I0(\REG.mem_11_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n54), .I3(GND_net), .O(n5097));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3713_3_lut (.I0(\REG.mem_11_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n54), .I3(GND_net), .O(n5096));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3712_3_lut (.I0(\REG.mem_11_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n54), .I3(GND_net), .O(n5095));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3711_3_lut (.I0(\REG.mem_11_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n54), .I3(GND_net), .O(n5094));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3710_3_lut (.I0(\REG.mem_11_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n54), .I3(GND_net), .O(n5093));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3709_3_lut (.I0(\REG.mem_11_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n54), .I3(GND_net), .O(n5092));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3708_3_lut (.I0(\REG.mem_10_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n55), .I3(GND_net), .O(n5091));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3707_3_lut (.I0(\REG.mem_10_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n55), .I3(GND_net), .O(n5090));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3706_3_lut (.I0(\REG.mem_10_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n55), .I3(GND_net), .O(n5089));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3476_3_lut (.I0(tx_data_byte[2]), .I1(pc_data_rx[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4859));   // src/top.v(1074[8] 1141[4])
    defparam i3476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3472_3_lut (.I0(tx_data_byte[3]), .I1(pc_data_rx[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4855));   // src/top.v(1074[8] 1141[4])
    defparam i3472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3705_3_lut (.I0(\REG.mem_10_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n55), .I3(GND_net), .O(n5088));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3704_3_lut (.I0(\REG.mem_10_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n55), .I3(GND_net), .O(n5087));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3703_3_lut (.I0(\REG.mem_10_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n55), .I3(GND_net), .O(n5086));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3702_3_lut (.I0(\REG.mem_10_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n55), .I3(GND_net), .O(n5085));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3701_3_lut (.I0(\REG.mem_10_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n55), .I3(GND_net), .O(n5084));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3700_3_lut (.I0(\REG.mem_10_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n55), .I3(GND_net), .O(n5083));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3699_3_lut (.I0(\REG.mem_10_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n55), .I3(GND_net), .O(n5082));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3698_3_lut (.I0(\REG.mem_10_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n55), .I3(GND_net), .O(n5081));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3697_3_lut (.I0(\REG.mem_10_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n55), .I3(GND_net), .O(n5080));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3462_3_lut (.I0(tx_data_byte[4]), .I1(pc_data_rx[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4845));   // src/top.v(1074[8] 1141[4])
    defparam i3462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3696_3_lut (.I0(\REG.mem_10_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n55), .I3(GND_net), .O(n5079));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3695_3_lut (.I0(\REG.mem_10_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n55), .I3(GND_net), .O(n5078));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3694_3_lut (.I0(\REG.mem_10_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n55), .I3(GND_net), .O(n5077));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3694_3_lut.LUT_INIT = 16'hcaca;
    \uart_rx(CLKS_PER_BIT=20)  pc_rx (.SLM_CLK_c(SLM_CLK_c), .r_Rx_Data(r_Rx_Data), 
            .GND_net(GND_net), .debug_led3(debug_led3), .n4248(n4248), 
            .n4253(n4253), .n4(n4_adj_1220), .n4_adj_1(n4_adj_1244), .n7347(n7347), 
            .n6083(n6083), .pc_data_rx({pc_data_rx}), .VCC_net(VCC_net), 
            .n6067(n6067), .n6066(n6066), .n6064(n6064), .n6063(n6063), 
            .n6062(n6062), .n6060(n6060), .n4_adj_2(n4_adj_1243), .n10211(n10211), 
            .UART_RX_c(UART_RX_c), .n6030(n6030)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(699[42] 704[3])
    SB_LUT4 i3693_3_lut (.I0(\REG.mem_10_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n55), .I3(GND_net), .O(n5076));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3692_3_lut (.I0(\REG.mem_9_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n56), .I3(GND_net), .O(n5075));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3455_3_lut (.I0(rx_shift_reg[5]), .I1(rx_shift_reg[4]), .I2(n4312), 
            .I3(GND_net), .O(n4838));   // src/spi.v(76[8] 221[4])
    defparam i3455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3691_3_lut (.I0(\REG.mem_9_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n56), .I3(GND_net), .O(n5074));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3690_3_lut (.I0(\REG.mem_9_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n56), .I3(GND_net), .O(n5073));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3689_3_lut (.I0(\REG.mem_9_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n56), .I3(GND_net), .O(n5072));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3688_3_lut (.I0(\REG.mem_9_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n56), .I3(GND_net), .O(n5071));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3687_3_lut (.I0(\REG.mem_9_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n56), .I3(GND_net), .O(n5070));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3686_3_lut (.I0(\REG.mem_9_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n56), .I3(GND_net), .O(n5069));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3453_3_lut (.I0(rx_shift_reg[6]), .I1(rx_shift_reg[5]), .I2(n4312), 
            .I3(GND_net), .O(n4836));   // src/spi.v(76[8] 221[4])
    defparam i3453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3685_3_lut (.I0(\REG.mem_9_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n56), .I3(GND_net), .O(n5068));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3684_3_lut (.I0(\REG.mem_9_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n56), .I3(GND_net), .O(n5067));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3683_3_lut (.I0(\REG.mem_9_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n56), .I3(GND_net), .O(n5066));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3682_3_lut (.I0(\REG.mem_9_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n56), .I3(GND_net), .O(n5065));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3681_3_lut (.I0(\REG.mem_9_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n56), .I3(GND_net), .O(n5064));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3680_3_lut (.I0(\REG.mem_9_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n56), .I3(GND_net), .O(n5063));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3679_3_lut (.I0(\REG.mem_9_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n56), .I3(GND_net), .O(n5062));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3678_3_lut (.I0(\REG.mem_9_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n56), .I3(GND_net), .O(n5061));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3677_3_lut (.I0(\REG.mem_9_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n56), .I3(GND_net), .O(n5060));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3676_3_lut (.I0(\REG.mem_8_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n57), .I3(GND_net), .O(n5059));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3675_3_lut (.I0(\REG.mem_8_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n57), .I3(GND_net), .O(n5058));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3674_3_lut (.I0(\REG.mem_8_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n57), .I3(GND_net), .O(n5057));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3673_3_lut (.I0(\REG.mem_8_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n57), .I3(GND_net), .O(n5056));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3672_3_lut (.I0(\REG.mem_8_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n57), .I3(GND_net), .O(n5055));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3671_3_lut (.I0(\REG.mem_8_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n57), .I3(GND_net), .O(n5054));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3670_3_lut (.I0(\REG.mem_8_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n57), .I3(GND_net), .O(n5053));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3669_3_lut (.I0(\REG.mem_8_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n57), .I3(GND_net), .O(n5052));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3668_3_lut (.I0(\REG.mem_8_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n57), .I3(GND_net), .O(n5051));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3667_3_lut (.I0(\REG.mem_8_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n57), .I3(GND_net), .O(n5050));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3666_3_lut (.I0(\REG.mem_8_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n57), .I3(GND_net), .O(n5049));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3665_3_lut (.I0(\REG.mem_8_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n57), .I3(GND_net), .O(n5048));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3664_3_lut (.I0(\REG.mem_8_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n57), .I3(GND_net), .O(n5047));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3663_3_lut (.I0(\REG.mem_8_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n57), .I3(GND_net), .O(n5046));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3662_3_lut (.I0(\REG.mem_8_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n57), .I3(GND_net), .O(n5045));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3661_3_lut (.I0(\REG.mem_8_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n57), .I3(GND_net), .O(n5044));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3660_3_lut (.I0(\REG.mem_7_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n58), .I3(GND_net), .O(n5043));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3659_3_lut (.I0(\REG.mem_7_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n58), .I3(GND_net), .O(n5042));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3658_3_lut (.I0(\REG.mem_7_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n58), .I3(GND_net), .O(n5041));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3657_3_lut (.I0(\REG.mem_7_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n58), .I3(GND_net), .O(n5040));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3656_3_lut (.I0(\REG.mem_7_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n58), .I3(GND_net), .O(n5039));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3655_3_lut (.I0(\REG.mem_7_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n58), .I3(GND_net), .O(n5038));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3654_3_lut (.I0(\REG.mem_7_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n58), .I3(GND_net), .O(n5037));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3653_3_lut (.I0(\REG.mem_7_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n58), .I3(GND_net), .O(n5036));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3652_3_lut (.I0(\REG.mem_7_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n58), .I3(GND_net), .O(n5035));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3651_3_lut (.I0(\REG.mem_7_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n58), .I3(GND_net), .O(n5034));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3650_3_lut (.I0(\REG.mem_7_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n58), .I3(GND_net), .O(n5033));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3649_3_lut (.I0(\REG.mem_7_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n58), .I3(GND_net), .O(n5032));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3648_3_lut (.I0(\REG.mem_7_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n58), .I3(GND_net), .O(n5031));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3647_3_lut (.I0(\REG.mem_7_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n58), .I3(GND_net), .O(n5030));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3646_3_lut (.I0(\REG.mem_7_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n58), .I3(GND_net), .O(n5029));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3645_3_lut (.I0(\REG.mem_7_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n58), .I3(GND_net), .O(n5028));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3644_3_lut (.I0(\REG.mem_6_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n59), .I3(GND_net), .O(n5027));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3643_3_lut (.I0(\REG.mem_6_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n59), .I3(GND_net), .O(n5026));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3642_3_lut (.I0(\REG.mem_6_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n59), .I3(GND_net), .O(n5025));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3641_3_lut (.I0(\REG.mem_6_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n59), .I3(GND_net), .O(n5024));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3640_3_lut (.I0(\REG.mem_6_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n59), .I3(GND_net), .O(n5023));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3639_3_lut (.I0(\REG.mem_6_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n59), .I3(GND_net), .O(n5022));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3638_3_lut (.I0(\REG.mem_6_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n59), .I3(GND_net), .O(n5021));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3637_3_lut (.I0(\REG.mem_6_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n59), .I3(GND_net), .O(n5020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3636_3_lut (.I0(\REG.mem_6_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n59), .I3(GND_net), .O(n5019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3635_3_lut (.I0(\REG.mem_6_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n59), .I3(GND_net), .O(n5018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3634_3_lut (.I0(\REG.mem_6_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n59), .I3(GND_net), .O(n5017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3633_3_lut (.I0(\REG.mem_6_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n59), .I3(GND_net), .O(n5016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3632_3_lut (.I0(\REG.mem_6_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n59), .I3(GND_net), .O(n5015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3631_3_lut (.I0(\REG.mem_6_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n59), .I3(GND_net), .O(n5014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3630_3_lut (.I0(\REG.mem_6_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n59), .I3(GND_net), .O(n5013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3629_3_lut (.I0(\REG.mem_6_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n59), .I3(GND_net), .O(n5012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3628_3_lut (.I0(\REG.mem_5_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n60), .I3(GND_net), .O(n5011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3627_3_lut (.I0(\REG.mem_5_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n60), .I3(GND_net), .O(n5010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3626_3_lut (.I0(\REG.mem_5_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n60), .I3(GND_net), .O(n5009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3625_3_lut (.I0(\REG.mem_5_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n60), .I3(GND_net), .O(n5008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3624_3_lut (.I0(\REG.mem_5_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n60), .I3(GND_net), .O(n5007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3623_3_lut (.I0(\REG.mem_5_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n60), .I3(GND_net), .O(n5006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3622_3_lut (.I0(\REG.mem_5_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n60), .I3(GND_net), .O(n5005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3621_3_lut (.I0(\REG.mem_5_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n60), .I3(GND_net), .O(n5004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3620_3_lut (.I0(\REG.mem_5_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n60), .I3(GND_net), .O(n5003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3619_3_lut (.I0(\REG.mem_5_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n60), .I3(GND_net), .O(n5002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3618_3_lut (.I0(\REG.mem_5_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n60), .I3(GND_net), .O(n5001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3617_3_lut (.I0(\REG.mem_5_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n60), .I3(GND_net), .O(n5000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3616_3_lut (.I0(\REG.mem_5_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n60), .I3(GND_net), .O(n4999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3615_3_lut (.I0(\REG.mem_5_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n60), .I3(GND_net), .O(n4998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3614_3_lut (.I0(\REG.mem_5_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n60), .I3(GND_net), .O(n4997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3613_3_lut (.I0(\REG.mem_5_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n60), .I3(GND_net), .O(n4996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3612_3_lut (.I0(\REG.mem_4_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n61), .I3(GND_net), .O(n4995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1216_2_lut_3_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(reset_all_w), .I3(GND_net), .O(empty_o_N_1149));
    defparam i1216_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i3611_3_lut (.I0(\REG.mem_4_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n61), .I3(GND_net), .O(n4994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3610_3_lut (.I0(\REG.mem_4_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n61), .I3(GND_net), .O(n4993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3609_3_lut (.I0(\REG.mem_4_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n61), .I3(GND_net), .O(n4992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3608_3_lut (.I0(\REG.mem_4_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n61), .I3(GND_net), .O(n4991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3607_3_lut (.I0(\REG.mem_4_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n61), .I3(GND_net), .O(n4990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3606_3_lut (.I0(\REG.mem_4_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n61), .I3(GND_net), .O(n4989));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3605_3_lut (.I0(\REG.mem_4_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n61), .I3(GND_net), .O(n4988));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3604_3_lut (.I0(\REG.mem_4_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n61), .I3(GND_net), .O(n4987));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3603_3_lut (.I0(\REG.mem_4_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n61), .I3(GND_net), .O(n4986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3602_3_lut (.I0(\REG.mem_4_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n61), .I3(GND_net), .O(n4985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3601_3_lut (.I0(\REG.mem_4_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n61), .I3(GND_net), .O(n4984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3600_3_lut (.I0(\REG.mem_4_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n61), .I3(GND_net), .O(n4983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3599_3_lut (.I0(\REG.mem_4_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n61), .I3(GND_net), .O(n4982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3598_3_lut (.I0(\REG.mem_4_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n61), .I3(GND_net), .O(n4981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3597_3_lut (.I0(\REG.mem_4_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n61), .I3(GND_net), .O(n4980));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3596_3_lut (.I0(\REG.mem_3_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n62), .I3(GND_net), .O(n4979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3595_3_lut (.I0(\REG.mem_3_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n62), .I3(GND_net), .O(n4978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3594_3_lut (.I0(\REG.mem_3_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n62), .I3(GND_net), .O(n4977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3593_3_lut (.I0(\REG.mem_3_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n62), .I3(GND_net), .O(n4976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3592_3_lut (.I0(\REG.mem_3_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n62), .I3(GND_net), .O(n4975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3591_3_lut (.I0(\REG.mem_3_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n62), .I3(GND_net), .O(n4974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3590_3_lut (.I0(\REG.mem_3_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n62), .I3(GND_net), .O(n4973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3589_3_lut (.I0(\REG.mem_3_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n62), .I3(GND_net), .O(n4972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3588_3_lut (.I0(\REG.mem_3_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n62), .I3(GND_net), .O(n4971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3587_3_lut (.I0(\REG.mem_3_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n62), .I3(GND_net), .O(n4970));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3586_3_lut (.I0(\REG.mem_3_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n62), .I3(GND_net), .O(n4969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i949_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(n63), 
            .I3(state[2]), .O(n2034));   // src/timing_controller.v(48[11:16])
    defparam i949_4_lut_4_lut.LUT_INIT = 16'h0806;
    SB_LUT4 i4723_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [2]), .I3(fifo_data_out[2]), .O(n6106));
    defparam i4723_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3536_4_lut_4_lut (.I0(reset_all_w), .I1(rd_addr_r_adj_1287[1]), 
            .I2(rd_addr_r_adj_1287[0]), .I3(rd_fifo_en_w_adj_1221), .O(n4919));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i3536_4_lut_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i4720_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [1]), .I3(fifo_data_out[1]), .O(n6103));
    defparam i4720_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i1_2_lut_4_lut (.I0(reset_clk_counter[2]), .I1(reset_all_w_N_61), 
            .I2(reset_clk_counter[0]), .I3(reset_clk_counter[1]), .O(n10167));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'haaa6;
    SB_LUT4 i3444_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [3]), .I3(fifo_data_out[3]), .O(n4827));
    defparam i3444_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3447_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_per_frame), 
            .I2(\REG.out_raw [4]), .I3(fifo_data_out[4]), .O(n4830));
    defparam i3447_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4715_3_lut_4_lut (.I0(r_SM_Main_2__N_844[0]), .I1(fifo_read_cmd), 
            .I2(is_fifo_empty_flag), .I3(tx_uart_active_flag), .O(n6098));   // src/top.v(910[8] 928[4])
    defparam i4715_3_lut_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4704_2_lut_3_lut (.I0(fifo_data_out[0]), .I1(bluejay_data_out_31__N_736), 
            .I2(bluejay_data_out_31__N_737), .I3(GND_net), .O(n6087));   // src/bluejay_data.v(126[8] 148[4])
    defparam i4704_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i3451_3_lut (.I0(rx_shift_reg[7]), .I1(rx_shift_reg[6]), .I2(n4312), 
            .I3(GND_net), .O(n4834));   // src/spi.v(76[8] 221[4])
    defparam i3451_3_lut.LUT_INIT = 16'hcaca;
    FIFO_Quad_Word tx_fifo (.rd_fifo_en_w(rd_fifo_en_w_adj_1221), .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r [7]), 
            .SLM_CLK_c(SLM_CLK_c), .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r [6]), 
            .rd_addr_r({rd_addr_r_adj_1287}), .\rd_addr_p1_w[2] (rd_addr_p1_w_adj_1289[2]), 
            .GND_net(GND_net), .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r [5]), 
            .n13895(n13895), .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r [0]), 
            .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r [4]), .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r [3]), 
            .reset_all_w(reset_all_w), .n8(n8), .wr_addr_r({wr_addr_r_adj_1284}), 
            .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r [2]), .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r [1]), 
            .n4941(n4941), .VCC_net(VCC_net), .n4938(n4938), .rx_buf_byte({rx_buf_byte}), 
            .n6112(n6112), .\fifo_temp_output[1] (fifo_temp_output[1]), 
            .n10302(n10302), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .n6073(n6073), .\fifo_temp_output[0] (fifo_temp_output[0]), 
            .n1(n1), .\wr_addr_p1_w[2] (wr_addr_p1_w_adj_1286[2]), .n10098(n10098), 
            .n5310(n5310), .\fifo_temp_output[4] (fifo_temp_output[4]), 
            .n5313(n5313), .\fifo_temp_output[5] (fifo_temp_output[5]), 
            .n4882(n4882), .\fifo_temp_output[2] (fifo_temp_output[2]), 
            .n4887(n4887), .\fifo_temp_output[3] (fifo_temp_output[3]), 
            .n5534(n5534), .\fifo_temp_output[6] (fifo_temp_output[6]), 
            .n5537(n5537), .\fifo_temp_output[7] (fifo_temp_output[7]), 
            .n10632(n10632), .is_fifo_empty_flag(is_fifo_empty_flag), .n4919(n4919), 
            .n4922(n4922), .fifo_write_cmd(fifo_write_cmd), .wr_fifo_en_w(wr_fifo_en_w), 
            .n4878(n4878), .rd_fifo_en_prev_r(rd_fifo_en_prev_r), .fifo_read_cmd(fifo_read_cmd)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(933[16] 949[2])
    SB_LUT4 i1_4_lut_4_lut (.I0(is_tx_fifo_full_flag), .I1(n10712), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3585_3_lut (.I0(\REG.mem_3_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n62), .I3(GND_net), .O(n4968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3584_3_lut (.I0(\REG.mem_3_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n62), .I3(GND_net), .O(n4967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3583_3_lut (.I0(\REG.mem_3_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n62), .I3(GND_net), .O(n4966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3582_3_lut (.I0(\REG.mem_3_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n62), .I3(GND_net), .O(n4965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3581_3_lut (.I0(\REG.mem_3_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n62), .I3(GND_net), .O(n4964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3441_3_lut (.I0(tx_data_byte[0]), .I1(pc_data_rx[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4824));   // src/top.v(1074[8] 1141[4])
    defparam i3441_3_lut.LUT_INIT = 16'hcaca;
    clock clock_inst (.GND_net(GND_net), .VCC_net(VCC_net), .ICE_SYSCLK_c(ICE_SYSCLK_c), 
          .pll_clk_unbuf(pll_clk_unbuf)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(222[7] 228[3])
    SB_LUT4 i4151_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[6]), 
            .I2(\mem_LUT.data_raw_r [6]), .I3(n4459), .O(n5534));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4151_4_lut_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i3533_2_lut_3_lut (.I0(reset_per_frame), .I1(DEBUG_3_c), .I2(get_next_word), 
            .I3(GND_net), .O(n4916));   // src/fifo_dc_32_lut_gen.v(751[29] 761[32])
    defparam i3533_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i4154_4_lut_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[7]), 
            .I2(\mem_LUT.data_raw_r [7]), .I3(n4459), .O(n5537));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4154_4_lut_4_lut.LUT_INIT = 16'h5044;
    usb3_if usb3_if_inst (.reset_per_frame(reset_per_frame), .reset_per_frame_latched(reset_per_frame_latched), 
            .SLM_CLK_c(SLM_CLK_c), .write_to_dc32_fifo_latched_N_425(write_to_dc32_fifo_latched_N_425), 
            .n2352(n2352), .DEBUG_3_c(DEBUG_3_c), .DEBUG_2_c(DEBUG_2_c), 
            .FIFO_CLK_c(FIFO_CLK_c), .\dc32_fifo_data_in[0] (dc32_fifo_data_in[0]), 
            .DEBUG_5_c(DEBUG_5_c), .buffer_switch_done(buffer_switch_done), 
            .buffer_switch_done_latched(buffer_switch_done_latched), .n571(n571), 
            .n575(n575), .GND_net(GND_net), .VCC_net(VCC_net), .FT_OE_N_420(FT_OE_N_420), 
            .n4911(n4911), .n4910(n4910), .n4907(n4907), .dc32_fifo_almost_full(dc32_fifo_almost_full), 
            .FT_OE_c(FT_OE_c), .FIFO_D15_c_15(FIFO_D15_c_15), .FIFO_D14_c_14(FIFO_D14_c_14), 
            .FIFO_D13_c_13(FIFO_D13_c_13), .FIFO_D12_c_12(FIFO_D12_c_12), 
            .FIFO_D11_c_11(FIFO_D11_c_11), .FIFO_D10_c_10(FIFO_D10_c_10), 
            .FIFO_D9_c_9(FIFO_D9_c_9), .FIFO_D8_c_8(FIFO_D8_c_8), .FIFO_D7_c_7(FIFO_D7_c_7), 
            .FIFO_D6_c_6(FIFO_D6_c_6), .FIFO_D5_c_5(FIFO_D5_c_5), .FIFO_D4_c_4(FIFO_D4_c_4), 
            .FIFO_D3_c_3(FIFO_D3_c_3), .FIFO_D2_c_2(FIFO_D2_c_2), .FIFO_D1_c_1(FIFO_D1_c_1), 
            .\dc32_fifo_data_in[15] (dc32_fifo_data_in[15]), .\dc32_fifo_data_in[14] (dc32_fifo_data_in[14]), 
            .\dc32_fifo_data_in[13] (dc32_fifo_data_in[13]), .\dc32_fifo_data_in[12] (dc32_fifo_data_in[12]), 
            .\dc32_fifo_data_in[11] (dc32_fifo_data_in[11]), .\dc32_fifo_data_in[10] (dc32_fifo_data_in[10]), 
            .\dc32_fifo_data_in[9] (dc32_fifo_data_in[9]), .\dc32_fifo_data_in[8] (dc32_fifo_data_in[8]), 
            .\dc32_fifo_data_in[7] (dc32_fifo_data_in[7]), .\dc32_fifo_data_in[6] (dc32_fifo_data_in[6]), 
            .\dc32_fifo_data_in[5] (dc32_fifo_data_in[5]), .\dc32_fifo_data_in[4] (dc32_fifo_data_in[4]), 
            .\dc32_fifo_data_in[3] (dc32_fifo_data_in[3]), .\dc32_fifo_data_in[2] (dc32_fifo_data_in[2]), 
            .\dc32_fifo_data_in[1] (dc32_fifo_data_in[1]), .DEBUG_1_c_c(DEBUG_1_c_c)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(513[9] 530[3])
    \uart_tx(CLKS_PER_BIT=20)  pc_tx (.UART_TX_c(UART_TX_c), .SLM_CLK_c(SLM_CLK_c), 
            .r_SM_Main({r_SM_Main_adj_1261}), .GND_net(GND_net), .\r_SM_Main_2__N_841[1] (r_SM_Main_2__N_841[1]), 
            .\r_SM_Main_2__N_844[0] (r_SM_Main_2__N_844[0]), .n3794(n3794), 
            .VCC_net(VCC_net), .n13737(n13737), .n4890(n4890), .r_Tx_Data({r_Tx_Data}), 
            .n4889(n4889), .tx_uart_active_flag(tx_uart_active_flag), .n5194(n5194), 
            .n5193(n5193), .n5192(n5192), .n5191(n5191), .n5189(n5189), 
            .n5173(n5173), .n5172(n5172), .n10653(n10653)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(768[42] 777[3])
    SB_LUT4 i1_2_lut_4_lut_adj_77 (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(wr_addr_r_adj_1284[0]), .I3(rd_addr_r_adj_1287[0]), .O(n4));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_2_lut_4_lut_adj_77.LUT_INIT = 16'h0220;
    spi spi0 (.SEN_c_1(SEN_c_1), .SLM_CLK_c(SLM_CLK_c), .SOUT_c(SOUT_c), 
        .n4312(n4312), .\rx_shift_reg[0] (rx_shift_reg[0]), .\tx_data_byte[3] (tx_data_byte[3]), 
        .n2086(n2086), .GND_net(GND_net), .\tx_data_byte[4] (tx_data_byte[4]), 
        .\tx_data_byte[5] (tx_data_byte[5]), .n4319(n4319), .SDAT_c_15(SDAT_c_15), 
        .\tx_data_byte[6] (tx_data_byte[6]), .\tx_data_byte[7] (tx_data_byte[7]), 
        .tx_addr_byte({tx_addr_byte}), .VCC_net(VCC_net), .n10300(n10300), 
        .\tx_shift_reg[0] (tx_shift_reg[0]), .n6049(n6049), .rx_buf_byte({rx_buf_byte}), 
        .n6048(n6048), .n6047(n6047), .n6046(n6046), .n6045(n6045), 
        .n6044(n6044), .n6043(n6043), .spi_rx_byte_ready(spi_rx_byte_ready), 
        .SCK_c_0(SCK_c_0), .spi_start_transfer_r(spi_start_transfer_r), 
        .n4897(n4897), .n4888(n4888), .\rx_shift_reg[1] (rx_shift_reg[1]), 
        .n4883(n4883), .\rx_shift_reg[2] (rx_shift_reg[2]), .n4877(n4877), 
        .\rx_shift_reg[3] (rx_shift_reg[3]), .n4869(n4869), .\rx_shift_reg[4] (rx_shift_reg[4]), 
        .n4838(n4838), .\rx_shift_reg[5] (rx_shift_reg[5]), .n4836(n4836), 
        .\rx_shift_reg[6] (rx_shift_reg[6]), .n4834(n4834), .\rx_shift_reg[7] (rx_shift_reg[7]), 
        .multi_byte_spi_trans_flag_r(multi_byte_spi_trans_flag_r), .\tx_data_byte[2] (tx_data_byte[2]), 
        .\tx_data_byte[1] (tx_data_byte[1]), .n3495(n3495)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(833[5] 857[2])
    SB_LUT4 i3518_2_lut_4_lut (.I0(reset_per_frame), .I1(rd_addr_r[0]), 
            .I2(rd_addr_p1_w[0]), .I3(rd_fifo_en_w), .O(n4901));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i3518_2_lut_4_lut.LUT_INIT = 16'h5044;
    
endmodule
//
// Verilog Description of module timing_controller
//

module timing_controller (state, SLM_CLK_c, n1879, GND_net, n10384, 
            VCC_net, n10662, reset_per_frame, n1774, n7258, INVERT_c_3, 
            buffer_switch_done, n4245, n7440, n7462, n4192, n63, 
            n10681, UPDATE_c_2) /* synthesis syn_module_defined=1 */ ;
    output [3:0]state;
    input SLM_CLK_c;
    input n1879;
    input GND_net;
    input n10384;
    input VCC_net;
    input n10662;
    output reset_per_frame;
    input n1774;
    input n7258;
    output INVERT_c_3;
    output buffer_switch_done;
    output n4245;
    output n7440;
    input n7462;
    output n4192;
    output n63;
    output n10681;
    output UPDATE_c_2;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [3:0]state_3__N_80;
    
    wire n10683, n11902;
    wire [31:0]n1880;
    
    wire n11901;
    wire [31:0]n506;
    
    wire n4491;
    wire [31:0]state_timeout_counter;   // src/timing_controller.v(49[12:33])
    
    wire n4809, n13747, n10655, n1951;
    wire [31:0]n1952;
    
    wire n9993, n9994, n9977, n9978, n11900, n9976, n11893, n9992, 
        n9975, n11894, n9991, n9974, n9990, n11886, n9989, n10004, 
        n10003, n11895, n9988, n11896, n9987, n10002, n9986, n11897, 
        n9985, n10001, n10000, n9999, n9984, n11898, n9983, n9998, 
        n11899, n9982, n9981, n11889, n9997, n11890, n9996, n11891, 
        n9995, n9980;
    wire [3:0]n968;
    
    wire n9979, n4806, n11903, n10678, n11892, n11937, n2033, 
        n4496, n10687, n38, n52, n56, n54, n55, n53, n50, 
        n58, n62, n49, n12025, n5, n7442, n7;
    
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n10683), .D(state_3__N_80[0]));   // src/timing_controller.v(53[8] 129[4])
    SB_LUT4 mux_890_i2_3_lut (.I0(n11902), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[1]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i3_3_lut (.I0(n11901), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[2]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFESR state_timeout_counter_i0_i31 (.Q(state_timeout_counter[31]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[31]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i30 (.Q(state_timeout_counter[30]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[30]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_LUT4 i3_4_lut (.I0(state[3]), .I1(state[0]), .I2(state[1]), .I3(state[2]), 
            .O(n13747));
    defparam i3_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 mux_898_i25_3_lut_4_lut (.I0(state[1]), .I1(n10655), .I2(n1951), 
            .I3(n1880[24]), .O(n1952[24]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_898_i25_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i24_3_lut_4_lut (.I0(state[1]), .I1(n10655), .I2(n1951), 
            .I3(n1880[23]), .O(n1952[23]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_898_i24_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i23_3_lut_4_lut (.I0(state[1]), .I1(n10655), .I2(n1951), 
            .I3(n1880[22]), .O(n1952[22]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_898_i23_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i21_3_lut_4_lut (.I0(state[1]), .I1(n10655), .I2(n1951), 
            .I3(n1880[20]), .O(n1952[20]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_898_i21_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i20_3_lut_4_lut (.I0(state[1]), .I1(n10655), .I2(n1951), 
            .I3(n1880[19]), .O(n1952[19]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_898_i20_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i19_3_lut_4_lut (.I0(state[1]), .I1(n10655), .I2(n1951), 
            .I3(n1880[18]), .O(n1952[18]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_898_i19_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i16_3_lut_4_lut (.I0(state[1]), .I1(n10655), .I2(n1951), 
            .I3(n1880[15]), .O(n1952[15]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_898_i16_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i15_3_lut_4_lut (.I0(state[1]), .I1(n10655), .I2(n1951), 
            .I3(n1880[14]), .O(n1952[14]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_898_i15_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i13_3_lut_4_lut (.I0(state[1]), .I1(n10655), .I2(n1951), 
            .I3(n1880[12]), .O(n1952[12]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_898_i13_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i10_3_lut_4_lut (.I0(state[1]), .I1(n10655), .I2(n1951), 
            .I3(n1880[9]), .O(n1952[9]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_898_i10_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i11_3_lut_4_lut (.I0(state[1]), .I1(n10655), .I2(n1951), 
            .I3(n1880[10]), .O(n1952[10]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_898_i11_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_898_i4_3_lut_4_lut (.I0(state[1]), .I1(n10655), .I2(n1951), 
            .I3(n1880[3]), .O(n1952[3]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_898_i4_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(VCC_net), .D(n10384));   // src/timing_controller.v(53[8] 129[4])
    SB_DFF invert_55_i0 (.Q(reset_per_frame), .C(SLM_CLK_c), .D(n10662));   // src/timing_controller.v(59[5] 128[12])
    SB_DFFESR state_timeout_counter_i0_i29 (.Q(state_timeout_counter[29]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[29]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i28 (.Q(state_timeout_counter[28]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[28]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i27 (.Q(state_timeout_counter[27]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[27]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i26 (.Q(state_timeout_counter[26]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[26]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i25 (.Q(state_timeout_counter[25]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[25]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i21 (.Q(state_timeout_counter[21]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[21]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i17 (.Q(state_timeout_counter[17]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[17]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i16 (.Q(state_timeout_counter[16]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[16]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i13 (.Q(state_timeout_counter[13]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[13]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i11 (.Q(state_timeout_counter[11]), 
            .C(SLM_CLK_c), .E(n4491), .D(n506[11]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_CARRY sub_31_add_2_22 (.CI(n9993), .I0(state_timeout_counter[20]), 
            .I1(VCC_net), .CO(n9994));
    SB_CARRY sub_31_add_2_6 (.CI(n9977), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n9978));
    SB_LUT4 sub_31_add_2_5_lut (.I0(n1774), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n9976), .O(n11900)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_21_lut (.I0(n1774), .I1(state_timeout_counter[19]), 
            .I2(VCC_net), .I3(n9992), .O(n11893)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_21 (.CI(n9992), .I0(state_timeout_counter[19]), 
            .I1(VCC_net), .CO(n9993));
    SB_CARRY sub_31_add_2_5 (.CI(n9976), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n9977));
    SB_LUT4 sub_31_add_2_4_lut (.I0(n7258), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n9975), .O(n11901)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_31_add_2_20_lut (.I0(n1774), .I1(state_timeout_counter[18]), 
            .I2(VCC_net), .I3(n9991), .O(n11894)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_20 (.CI(n9991), .I0(state_timeout_counter[18]), 
            .I1(VCC_net), .CO(n9992));
    SB_CARRY sub_31_add_2_4 (.CI(n9975), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n9976));
    SB_LUT4 sub_31_add_2_3_lut (.I0(n1774), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n9974), .O(n11902)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_19_lut (.I0(GND_net), .I1(state_timeout_counter[17]), 
            .I2(VCC_net), .I3(n9990), .O(n506[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_19 (.CI(n9990), .I0(state_timeout_counter[17]), 
            .I1(VCC_net), .CO(n9991));
    SB_CARRY sub_31_add_2_3 (.CI(n9974), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n9975));
    SB_LUT4 sub_31_add_2_2_lut (.I0(n7258), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n11886)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_31_add_2_18_lut (.I0(GND_net), .I1(state_timeout_counter[16]), 
            .I2(VCC_net), .I3(n9989), .O(n506[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_33_lut (.I0(GND_net), .I1(state_timeout_counter[31]), 
            .I2(VCC_net), .I3(n10004), .O(n506[31])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_32_lut (.I0(GND_net), .I1(state_timeout_counter[30]), 
            .I2(VCC_net), .I3(n10003), .O(n506[30])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_18 (.CI(n9989), .I0(state_timeout_counter[16]), 
            .I1(VCC_net), .CO(n9990));
    SB_CARRY sub_31_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n9974));
    SB_LUT4 sub_31_add_2_17_lut (.I0(n1774), .I1(state_timeout_counter[15]), 
            .I2(VCC_net), .I3(n9988), .O(n11895)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_32 (.CI(n10003), .I0(state_timeout_counter[30]), 
            .I1(VCC_net), .CO(n10004));
    SB_CARRY sub_31_add_2_17 (.CI(n9988), .I0(state_timeout_counter[15]), 
            .I1(VCC_net), .CO(n9989));
    SB_LUT4 sub_31_add_2_16_lut (.I0(n1774), .I1(state_timeout_counter[14]), 
            .I2(VCC_net), .I3(n9987), .O(n11896)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_31_lut (.I0(GND_net), .I1(state_timeout_counter[29]), 
            .I2(VCC_net), .I3(n10002), .O(n506[29])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_16 (.CI(n9987), .I0(state_timeout_counter[14]), 
            .I1(VCC_net), .CO(n9988));
    SB_LUT4 sub_31_add_2_15_lut (.I0(GND_net), .I1(state_timeout_counter[13]), 
            .I2(VCC_net), .I3(n9986), .O(n506[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_31 (.CI(n10002), .I0(state_timeout_counter[29]), 
            .I1(VCC_net), .CO(n10003));
    SB_CARRY sub_31_add_2_15 (.CI(n9986), .I0(state_timeout_counter[13]), 
            .I1(VCC_net), .CO(n9987));
    SB_LUT4 sub_31_add_2_14_lut (.I0(n1774), .I1(state_timeout_counter[12]), 
            .I2(VCC_net), .I3(n9985), .O(n11897)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_30_lut (.I0(GND_net), .I1(state_timeout_counter[28]), 
            .I2(VCC_net), .I3(n10001), .O(n506[28])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_30 (.CI(n10001), .I0(state_timeout_counter[28]), 
            .I1(VCC_net), .CO(n10002));
    SB_LUT4 sub_31_add_2_29_lut (.I0(GND_net), .I1(state_timeout_counter[27]), 
            .I2(VCC_net), .I3(n10000), .O(n506[27])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_29 (.CI(n10000), .I0(state_timeout_counter[27]), 
            .I1(VCC_net), .CO(n10001));
    SB_LUT4 sub_31_add_2_28_lut (.I0(GND_net), .I1(state_timeout_counter[26]), 
            .I2(VCC_net), .I3(n9999), .O(n506[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_14 (.CI(n9985), .I0(state_timeout_counter[12]), 
            .I1(VCC_net), .CO(n9986));
    SB_LUT4 sub_31_add_2_13_lut (.I0(GND_net), .I1(state_timeout_counter[11]), 
            .I2(VCC_net), .I3(n9984), .O(n506[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_28 (.CI(n9999), .I0(state_timeout_counter[26]), 
            .I1(VCC_net), .CO(n10000));
    SB_CARRY sub_31_add_2_13 (.CI(n9984), .I0(state_timeout_counter[11]), 
            .I1(VCC_net), .CO(n9985));
    SB_LUT4 sub_31_add_2_12_lut (.I0(n1774), .I1(state_timeout_counter[10]), 
            .I2(VCC_net), .I3(n9983), .O(n11898)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_27_lut (.I0(GND_net), .I1(state_timeout_counter[25]), 
            .I2(VCC_net), .I3(n9998), .O(n506[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_12 (.CI(n9983), .I0(state_timeout_counter[10]), 
            .I1(VCC_net), .CO(n9984));
    SB_LUT4 sub_31_add_2_11_lut (.I0(n1774), .I1(state_timeout_counter[9]), 
            .I2(VCC_net), .I3(n9982), .O(n11899)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_27 (.CI(n9998), .I0(state_timeout_counter[25]), 
            .I1(VCC_net), .CO(n9999));
    SB_CARRY sub_31_add_2_11 (.CI(n9982), .I0(state_timeout_counter[9]), 
            .I1(VCC_net), .CO(n9983));
    SB_LUT4 sub_31_add_2_10_lut (.I0(GND_net), .I1(state_timeout_counter[8]), 
            .I2(VCC_net), .I3(n9981), .O(n506[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_26_lut (.I0(n1774), .I1(state_timeout_counter[24]), 
            .I2(VCC_net), .I3(n9997), .O(n11889)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_26 (.CI(n9997), .I0(state_timeout_counter[24]), 
            .I1(VCC_net), .CO(n9998));
    SB_LUT4 sub_31_add_2_25_lut (.I0(n1774), .I1(state_timeout_counter[23]), 
            .I2(VCC_net), .I3(n9996), .O(n11890)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_25 (.CI(n9996), .I0(state_timeout_counter[23]), 
            .I1(VCC_net), .CO(n9997));
    SB_LUT4 sub_31_add_2_24_lut (.I0(n1774), .I1(state_timeout_counter[22]), 
            .I2(VCC_net), .I3(n9995), .O(n11891)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_10 (.CI(n9981), .I0(state_timeout_counter[8]), 
            .I1(VCC_net), .CO(n9982));
    SB_LUT4 sub_31_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n9980), .O(n506[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_24 (.CI(n9995), .I0(state_timeout_counter[22]), 
            .I1(VCC_net), .CO(n9996));
    SB_DFFESR state_timeout_counter_i0_i8 (.Q(state_timeout_counter[8]), .C(SLM_CLK_c), 
            .E(n4491), .D(n506[8]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFF invert_55_i3 (.Q(INVERT_c_3), .C(SLM_CLK_c), .D(n968[3]));   // src/timing_controller.v(59[5] 128[12])
    SB_CARRY sub_31_add_2_9 (.CI(n9980), .I0(state_timeout_counter[7]), 
            .I1(VCC_net), .CO(n9981));
    SB_LUT4 sub_31_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n9979), .O(n506[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_23_lut (.I0(GND_net), .I1(state_timeout_counter[21]), 
            .I2(VCC_net), .I3(n9994), .O(n506[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_8 (.CI(n9979), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n9980));
    SB_DFFESR state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(SLM_CLK_c), 
            .E(n4491), .D(n506[7]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n4491), .D(n506[6]), .R(n4809));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1880[2]), .R(n4806));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1880[1]), .R(n4806));   // src/timing_controller.v(53[8] 129[4])
    SB_CARRY sub_31_add_2_23 (.CI(n9994), .I0(state_timeout_counter[21]), 
            .I1(VCC_net), .CO(n9995));
    SB_LUT4 sub_31_add_2_7_lut (.I0(n10678), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n9978), .O(n11903)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_DFF invert_55_i1 (.Q(buffer_switch_done), .C(SLM_CLK_c), .D(n13747));   // src/timing_controller.v(59[5] 128[12])
    SB_CARRY sub_31_add_2_7 (.CI(n9978), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n9979));
    SB_LUT4 sub_31_add_2_22_lut (.I0(n1774), .I1(state_timeout_counter[20]), 
            .I2(VCC_net), .I3(n9993), .O(n11892)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_6_lut (.I0(n1774), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n9977), .O(n11937)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n4245));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6064_3_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n7440));
    defparam i6064_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_69 (.I0(n1774), .I1(n1879), .I2(GND_net), .I3(GND_net), 
            .O(n10678));   // src/timing_controller.v(59[5] 128[12])
    defparam i1_2_lut_adj_69.LUT_INIT = 16'h2222;
    SB_LUT4 i959_4_lut (.I0(state[3]), .I1(n2033), .I2(n7462), .I3(state[2]), 
            .O(n1951));   // src/timing_controller.v(53[8] 129[4])
    defparam i959_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i10195_2_lut (.I0(state[3]), .I1(n4192), .I2(GND_net), .I3(GND_net), 
            .O(n4491));   // src/timing_controller.v(59[5] 128[12])
    defparam i10195_2_lut.LUT_INIT = 16'h7777;
    SB_DFFE state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[0]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n4496), .D(state_3__N_80[2]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n4496), .D(state_3__N_80[1]));   // src/timing_controller.v(53[8] 129[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(state[2]), .I1(state[0]), .I2(n63), .I3(GND_net), 
            .O(n10687));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_343_Mux_3_i15_4_lut_4_lut (.I0(state[2]), .I1(state[0]), 
            .I2(state[1]), .I3(state[3]), .O(n968[3]));
    defparam mux_343_Mux_3_i15_4_lut_4_lut.LUT_INIT = 16'h01a0;
    SB_DFFE state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[3]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[4]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[5]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i9 (.Q(state_timeout_counter[9]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[9]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i10 (.Q(state_timeout_counter[10]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[10]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i12 (.Q(state_timeout_counter[12]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[12]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i14 (.Q(state_timeout_counter[14]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[14]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i15 (.Q(state_timeout_counter[15]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[15]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i18 (.Q(state_timeout_counter[18]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[18]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i19 (.Q(state_timeout_counter[19]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[19]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i20 (.Q(state_timeout_counter[20]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[20]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i22 (.Q(state_timeout_counter[22]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[22]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i23 (.Q(state_timeout_counter[23]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[23]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i24 (.Q(state_timeout_counter[24]), .C(SLM_CLK_c), 
            .E(n4491), .D(n1952[24]));   // src/timing_controller.v(53[8] 129[4])
    SB_LUT4 i948_2_lut_3_lut (.I0(state[0]), .I1(n63), .I2(state[1]), 
            .I3(GND_net), .O(n2033));   // src/timing_controller.v(53[8] 129[4])
    defparam i948_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_adj_70 (.I0(state[3]), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n10681));
    defparam i1_2_lut_adj_70.LUT_INIT = 16'hbbbb;
    SB_LUT4 i6_2_lut (.I0(state_timeout_counter[9]), .I1(state_timeout_counter[12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // src/timing_controller.v(81[17:45])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut (.I0(state_timeout_counter[17]), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[24]), .I3(state_timeout_counter[4]), 
            .O(n52));   // src/timing_controller.v(81[17:45])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(state_timeout_counter[29]), .I1(state_timeout_counter[3]), 
            .I2(state_timeout_counter[13]), .I3(state_timeout_counter[31]), 
            .O(n56));   // src/timing_controller.v(81[17:45])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(state_timeout_counter[19]), .I1(state_timeout_counter[5]), 
            .I2(state_timeout_counter[22]), .I3(state_timeout_counter[6]), 
            .O(n54));   // src/timing_controller.v(81[17:45])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(state_timeout_counter[10]), .I1(state_timeout_counter[15]), 
            .I2(state_timeout_counter[20]), .I3(state_timeout_counter[23]), 
            .O(n55));   // src/timing_controller.v(81[17:45])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(state_timeout_counter[27]), .I1(state_timeout_counter[7]), 
            .I2(state_timeout_counter[30]), .I3(state_timeout_counter[14]), 
            .O(n53));   // src/timing_controller.v(81[17:45])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(state_timeout_counter[8]), .I1(state_timeout_counter[11]), 
            .I2(state_timeout_counter[16]), .I3(state_timeout_counter[21]), 
            .O(n50));   // src/timing_controller.v(81[17:45])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(state_timeout_counter[25]), .I1(n52), .I2(n38), 
            .I3(state_timeout_counter[26]), .O(n58));   // src/timing_controller.v(81[17:45])
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30_4_lut (.I0(n53), .I1(n55), .I2(n54), .I3(n56), .O(n62));   // src/timing_controller.v(81[17:45])
    defparam i30_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(state_timeout_counter[0]), .I1(state_timeout_counter[18]), 
            .I2(state_timeout_counter[28]), .I3(state_timeout_counter[2]), 
            .O(n49));   // src/timing_controller.v(81[17:45])
    defparam i17_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i31_4_lut (.I0(n49), .I1(n62), .I2(n58), .I3(n50), .O(n63));   // src/timing_controller.v(81[17:45])
    defparam i31_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR invert_55_i2 (.Q(UPDATE_c_2), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n12025), .R(n5));   // src/timing_controller.v(59[5] 128[12])
    SB_LUT4 i6066_3_lut (.I0(n63), .I1(state[1]), .I2(state[2]), .I3(GND_net), 
            .O(n7442));
    defparam i6066_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 state_3__I_0_59_Mux_0_i7_4_lut (.I0(state[1]), .I1(n63), .I2(state[2]), 
            .I3(state[0]), .O(n7));   // src/timing_controller.v(59[5] 128[12])
    defparam state_3__I_0_59_Mux_0_i7_4_lut.LUT_INIT = 16'hc535;
    SB_LUT4 state_3__I_0_59_Mux_0_i15_4_lut (.I0(n7), .I1(n7442), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_80[0]));   // src/timing_controller.v(59[5] 128[12])
    defparam state_3__I_0_59_Mux_0_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 state_3__I_0_59_Mux_1_i15_4_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[3]), .I3(n10687), .O(state_3__N_80[1]));   // src/timing_controller.v(59[5] 128[12])
    defparam state_3__I_0_59_Mux_1_i15_4_lut_4_lut.LUT_INIT = 16'hc6f6;
    SB_LUT4 mux_898_i1_4_lut (.I0(n1880[0]), .I1(state[1]), .I2(n1951), 
            .I3(n10655), .O(n1952[0]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_898_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 mux_890_i1_3_lut (.I0(n11886), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[0]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i1_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10246_2_lut (.I0(state[3]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // src/timing_controller.v(53[8] 129[4])
    defparam i10246_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_3__I_0_59_Mux_2_i15_4_lut (.I0(state[1]), .I1(state[2]), 
            .I2(state[3]), .I3(state[0]), .O(state_3__N_80[2]));   // src/timing_controller.v(59[5] 128[12])
    defparam state_3__I_0_59_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 i1_2_lut_3_lut_adj_71 (.I0(n7440), .I1(state[3]), .I2(n63), 
            .I3(GND_net), .O(n4496));
    defparam i1_2_lut_3_lut_adj_71.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[3]), .I1(n63), .I2(state[1]), .I3(state[2]), 
            .O(n10683));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[0]), .I1(n63), .I2(state[3]), 
            .I3(state[2]), .O(n10655));   // src/timing_controller.v(53[8] 129[4])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 mux_890_i4_3_lut (.I0(n11900), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[3]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8962_4_lut (.I0(n11937), .I1(state[1]), .I2(n1879), .I3(n1951), 
            .O(n1952[4]));   // src/timing_controller.v(59[5] 128[12])
    defparam i8962_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_898_i6_3_lut (.I0(n11903), .I1(state[1]), .I2(n1951), 
            .I3(GND_net), .O(n1952[5]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_898_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10250_3_lut_4_lut (.I0(state[3]), .I1(n4192), .I2(n1951), 
            .I3(n10678), .O(n4809));
    defparam i10250_3_lut_4_lut.LUT_INIT = 16'h7077;
    SB_LUT4 mux_890_i10_3_lut (.I0(n11899), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[9]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_2_lut_3_lut_adj_72 (.I0(state[2]), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n4192));
    defparam i1_2_lut_3_lut_adj_72.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_890_i11_3_lut (.I0(n11898), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[10]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i11_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i13_3_lut (.I0(n11897), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[12]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i13_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i15_3_lut (.I0(n11896), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[14]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i15_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i16_3_lut (.I0(n11895), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[15]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i19_3_lut (.I0(n11894), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[18]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i19_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i20_3_lut (.I0(n11893), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[19]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i21_3_lut (.I0(n11892), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[20]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i21_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i23_3_lut (.I0(n11891), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[22]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i23_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i24_3_lut (.I0(n11890), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[23]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_890_i25_3_lut (.I0(n11889), .I1(state[1]), .I2(n1879), 
            .I3(GND_net), .O(n1880[24]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_890_i25_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10175_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n12025));   // src/timing_controller.v(59[5] 128[12])
    defparam i10175_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i3423_2_lut_3_lut (.I0(state[3]), .I1(n4192), .I2(n1951), 
            .I3(GND_net), .O(n4806));   // src/timing_controller.v(53[8] 129[4])
    defparam i3423_2_lut_3_lut.LUT_INIT = 16'h7070;
    
endmodule
//
// Verilog Description of module bluejay_data
//

module bluejay_data (dc32_fifo_almost_full, n843, GND_net, DEBUG_9_c, 
            SLM_CLK_c, n771, buffer_switch_done_latched, dc32_fifo_almost_empty, 
            bluejay_data_out_31__N_736, buffer_switch_done, bluejay_data_out_31__N_737, 
            n6087, DEBUG_6_c, VCC_net, SYNC_c, n10149, \rd_sig_diff0_w[1] , 
            get_next_word, \rd_sig_diff0_w[0] , \rd_sig_diff0_w[2] , n10700, 
            n10748, \aempty_flag_impl.ae_flag_nxt_w , DATA10_c_10, n4672, 
            DATA9_c_9, n4671, DATA11_c_11, n4670, DATA12_c_12, n4669, 
            DATA13_c_13, n4668, DATA14_c_14, n4667, DATA8_c_8, n4666, 
            DATA15_c_15, n4665, DATA7_c_7, n4664, DATA6_c_6, n4663, 
            DATA5_c_5, n4662, DATA4_c_4, n4661, DATA3_c_3, n4660, 
            DATA2_c_2, n4659, DATA1_c_1, n4658) /* synthesis syn_module_defined=1 */ ;
    input dc32_fifo_almost_full;
    output n843;
    input GND_net;
    output DEBUG_9_c;
    input SLM_CLK_c;
    output n771;
    input buffer_switch_done_latched;
    input dc32_fifo_almost_empty;
    output bluejay_data_out_31__N_736;
    input buffer_switch_done;
    output bluejay_data_out_31__N_737;
    input n6087;
    output DEBUG_6_c;
    input VCC_net;
    output SYNC_c;
    input n10149;
    input \rd_sig_diff0_w[1] ;
    output get_next_word;
    input \rd_sig_diff0_w[0] ;
    input \rd_sig_diff0_w[2] ;
    input n10700;
    input n10748;
    output \aempty_flag_impl.ae_flag_nxt_w ;
    output DATA10_c_10;
    input n4672;
    output DATA9_c_9;
    input n4671;
    output DATA11_c_11;
    input n4670;
    output DATA12_c_12;
    input n4669;
    output DATA13_c_13;
    input n4668;
    output DATA14_c_14;
    input n4667;
    output DATA8_c_8;
    input n4666;
    output DATA15_c_15;
    input n4665;
    output DATA7_c_7;
    input n4664;
    output DATA6_c_6;
    input n4663;
    output DATA5_c_5;
    input n4662;
    output DATA4_c_4;
    input n4661;
    output DATA3_c_3;
    input n4660;
    output DATA2_c_2;
    input n4659;
    output DATA1_c_1;
    input n4658;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [10:0]v_counter;   // src/bluejay_data.v(51[12:21])
    
    wire n10806, n10804, n4, valid_N_740, n20, n10840;
    wire [7:0]state_timeout_counter;   // src/bluejay_data.v(52[11:32])
    
    wire n10742, n13, n10814;
    wire [15:0]n828;
    
    wire n27, n10440, n4228, n12, n10178, n10179, n10112, n3031, 
        n891, bluejay_data_out_31__N_735, n3033, n895;
    wire [10:0]v_counter_10__N_715;
    
    wire n4408, n1, n4370, n4694, n3035, n4_adj_1213, n4722, n1291, 
        n7310, bluejay_data_out_31__N_734, n3029, n10026, n10025, 
        n1_adj_1214, n4719, n10024, n10023, n10022, n1_adj_1215, 
        n10554, n10021, n10020, n10019, n1_adj_1216, n10018, n10017;
    wire [8:0]n62;
    
    wire n9961, n6564, n9960, n9957, n9955, n9956, n9958, n9959, 
        n1_adj_1217, n1_adj_1218, n15, n12_adj_1219, n4876;
    
    SB_LUT4 i8957_4_lut (.I0(v_counter[8]), .I1(v_counter[4]), .I2(v_counter[5]), 
            .I3(v_counter[3]), .O(n10806));
    defparam i8957_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8955_4_lut (.I0(v_counter[2]), .I1(v_counter[6]), .I2(v_counter[7]), 
            .I3(v_counter[9]), .O(n10804));
    defparam i8955_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(dc32_fifo_almost_full), .I1(n843), .I2(GND_net), 
            .I3(GND_net), .O(n4));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_DFFN valid_56 (.Q(DEBUG_9_c), .C(SLM_CLK_c), .D(valid_N_740));   // src/bluejay_data.v(126[8] 148[4])
    SB_LUT4 i8990_4_lut (.I0(n10804), .I1(n20), .I2(n10806), .I3(v_counter[10]), 
            .O(n10840));
    defparam i8990_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8893_2_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[5]), 
            .I2(GND_net), .I3(GND_net), .O(n10742));
    defparam i8893_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i8965_4_lut (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[2]), 
            .I2(state_timeout_counter[4]), .I3(n13), .O(n10814));
    defparam i8965_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(state_timeout_counter[0]), .I1(n10840), .I2(n4), 
            .I3(n828[9]), .O(n27));
    defparam i1_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1_4_lut_adj_55 (.I0(n828[2]), .I1(n27), .I2(n10814), .I3(n10742), 
            .O(n10440));
    defparam i1_4_lut_adj_55.LUT_INIT = 16'haaae;
    SB_LUT4 i1_3_lut (.I0(dc32_fifo_almost_full), .I1(n843), .I2(n771), 
            .I3(GND_net), .O(n4228));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 equal_1263_i20_2_lut (.I0(v_counter[0]), .I1(v_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n20));   // src/bluejay_data.v(106[21:49])
    defparam equal_1263_i20_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i5_4_lut (.I0(v_counter[8]), .I1(v_counter[7]), .I2(v_counter[4]), 
            .I3(v_counter[3]), .O(n12));   // src/bluejay_data.v(108[25:41])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(v_counter[5]), .I1(n12), .I2(v_counter[2]), 
            .I3(v_counter[6]), .O(n10178));   // src/bluejay_data.v(108[25:41])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n828[9]), .I1(n10178), .I2(n771), .I3(n10179), 
            .O(n10112));   // src/bluejay_data.v(66[9] 121[16])
    defparam i2_4_lut.LUT_INIT = 16'h0a08;
    SB_LUT4 i1664_4_lut (.I0(buffer_switch_done_latched), .I1(n10112), .I2(n828[5]), 
            .I3(dc32_fifo_almost_full), .O(n3031));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1664_4_lut.LUT_INIT = 16'hccdc;
    SB_LUT4 reduce_or_325_i1_4_lut (.I0(dc32_fifo_almost_full), .I1(n771), 
            .I2(n828[5]), .I3(n828[4]), .O(n891));   // src/bluejay_data.v(66[9] 121[16])
    defparam reduce_or_325_i1_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 i1_4_lut_adj_56 (.I0(dc32_fifo_almost_empty), .I1(bluejay_data_out_31__N_735), 
            .I2(bluejay_data_out_31__N_736), .I3(buffer_switch_done_latched), 
            .O(n3033));   // src/bluejay_data.v(43[15:31])
    defparam i1_4_lut_adj_56.LUT_INIT = 16'hccdc;
    SB_LUT4 i1_2_lut_adj_57 (.I0(bluejay_data_out_31__N_736), .I1(dc32_fifo_almost_empty), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_2_lut_adj_57.LUT_INIT = 16'h8888;
    SB_DFFESR v_counter_i1 (.Q(v_counter[1]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[1]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i2 (.Q(v_counter[2]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[2]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i3 (.Q(v_counter[3]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[3]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i4 (.Q(v_counter[4]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[4]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i5 (.Q(v_counter[5]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[5]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i6 (.Q(v_counter[6]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[6]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i7 (.Q(v_counter[7]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[7]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS v_counter_i8 (.Q(v_counter[8]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[8]), .S(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i9 (.Q(v_counter[9]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[9]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS v_counter_i10 (.Q(v_counter[10]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[10]), .S(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(SLM_CLK_c), 
            .E(n4370), .D(n1), .S(n4694));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 i1_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n771), 
            .I2(n828[9]), .I3(bluejay_data_out_31__N_737), .O(n3035));   // src/bluejay_data.v(62[9] 65[12])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hff40;
    SB_DFFESS state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n4370), .D(n4_adj_1213), .S(n4722));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 i10213_2_lut (.I0(n4370), .I1(n1291), .I2(GND_net), .I3(GND_net), 
            .O(n7310));
    defparam i10213_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1662_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n771), 
            .I2(bluejay_data_out_31__N_734), .I3(n828[4]), .O(n3029));   // src/bluejay_data.v(62[9] 65[12])
    defparam i1662_3_lut_4_lut.LUT_INIT = 16'hf4f0;
    SB_DFFN bluejay_data_out_i1 (.Q(DEBUG_6_c), .C(SLM_CLK_c), .D(n6087));   // src/bluejay_data.v(126[8] 148[4])
    SB_LUT4 i2_3_lut (.I0(n828[9]), .I1(n828[4]), .I2(n843), .I3(GND_net), 
            .O(n1291));   // src/bluejay_data.v(66[9] 121[16])
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 sub_118_add_2_12_lut (.I0(GND_net), .I1(v_counter[10]), .I2(VCC_net), 
            .I3(n10026), .O(v_counter_10__N_715[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_118_add_2_11_lut (.I0(GND_net), .I1(v_counter[9]), .I2(VCC_net), 
            .I3(n10025), .O(v_counter_10__N_715[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_11 (.CI(n10025), .I0(v_counter[9]), .I1(VCC_net), 
            .CO(n10026));
    SB_DFFESS state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(SLM_CLK_c), 
            .E(n4370), .D(n1_adj_1214), .S(n4719));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 sub_118_add_2_10_lut (.I0(GND_net), .I1(v_counter[8]), .I2(VCC_net), 
            .I3(n10024), .O(v_counter_10__N_715[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_10 (.CI(n10024), .I0(v_counter[8]), .I1(VCC_net), 
            .CO(n10025));
    SB_LUT4 sub_118_add_2_9_lut (.I0(GND_net), .I1(v_counter[7]), .I2(VCC_net), 
            .I3(n10023), .O(v_counter_10__N_715[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_9 (.CI(n10023), .I0(v_counter[7]), .I1(VCC_net), 
            .CO(n10024));
    SB_LUT4 sub_118_add_2_8_lut (.I0(GND_net), .I1(v_counter[6]), .I2(VCC_net), 
            .I3(n10022), .O(v_counter_10__N_715[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_8 (.CI(n10022), .I0(v_counter[6]), .I1(VCC_net), 
            .CO(n10023));
    SB_DFFESS state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(SLM_CLK_c), 
            .E(n4370), .D(n1_adj_1215), .S(n10554));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 sub_118_add_2_7_lut (.I0(GND_net), .I1(v_counter[5]), .I2(VCC_net), 
            .I3(n10021), .O(v_counter_10__N_715[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_7 (.CI(n10021), .I0(v_counter[5]), .I1(VCC_net), 
            .CO(n10022));
    SB_LUT4 sub_118_add_2_6_lut (.I0(GND_net), .I1(v_counter[4]), .I2(VCC_net), 
            .I3(n10020), .O(v_counter_10__N_715[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_6 (.CI(n10020), .I0(v_counter[4]), .I1(VCC_net), 
            .CO(n10021));
    SB_LUT4 sub_118_add_2_5_lut (.I0(GND_net), .I1(v_counter[3]), .I2(VCC_net), 
            .I3(n10019), .O(v_counter_10__N_715[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(SLM_CLK_c), 
            .E(n4370), .D(n1_adj_1216), .S(n4719));   // src/bluejay_data.v(56[8] 123[4])
    SB_CARRY sub_118_add_2_5 (.CI(n10019), .I0(v_counter[3]), .I1(VCC_net), 
            .CO(n10020));
    SB_LUT4 sub_118_add_2_4_lut (.I0(GND_net), .I1(v_counter[2]), .I2(VCC_net), 
            .I3(n10018), .O(v_counter_10__N_715[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_4 (.CI(n10018), .I0(v_counter[2]), .I1(VCC_net), 
            .CO(n10019));
    SB_LUT4 sub_118_add_2_3_lut (.I0(GND_net), .I1(v_counter[1]), .I2(VCC_net), 
            .I3(n10017), .O(v_counter_10__N_715[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_3 (.CI(n10017), .I0(v_counter[1]), .I1(VCC_net), 
            .CO(n10018));
    SB_LUT4 sub_118_add_2_2_lut (.I0(GND_net), .I1(v_counter[0]), .I2(n771), 
            .I3(VCC_net), .O(v_counter_10__N_715[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_2 (.CI(VCC_net), .I0(v_counter[0]), .I1(n771), 
            .CO(n10017));
    SB_LUT4 i1_2_lut_adj_58 (.I0(n4370), .I1(bluejay_data_out_31__N_737), 
            .I2(GND_net), .I3(GND_net), .O(n4722));   // src/bluejay_data.v(61[10] 122[8])
    defparam i1_2_lut_adj_58.LUT_INIT = 16'h8888;
    SB_LUT4 sub_116_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n9961), .O(n62[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_59 (.I0(n828[2]), .I1(n828[5]), .I2(bluejay_data_out_31__N_736), 
            .I3(GND_net), .O(n6564));   // src/bluejay_data.v(66[9] 121[16])
    defparam i2_3_lut_adj_59.LUT_INIT = 16'hfefe;
    SB_LUT4 i3311_2_lut (.I0(n4370), .I1(bluejay_data_out_31__N_734), .I2(GND_net), 
            .I3(GND_net), .O(n4694));   // src/bluejay_data.v(56[8] 123[4])
    defparam i3311_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10242_3_lut (.I0(buffer_switch_done_latched), .I1(buffer_switch_done), 
            .I2(n6564), .I3(GND_net), .O(n4370));   // src/bluejay_data.v(61[10] 122[8])
    defparam i10242_3_lut.LUT_INIT = 16'h2323;
    SB_LUT4 i1_2_lut_adj_60 (.I0(n828[9]), .I1(buffer_switch_done), .I2(GND_net), 
            .I3(GND_net), .O(n4408));
    defparam i1_2_lut_adj_60.LUT_INIT = 16'heeee;
    SB_LUT4 sub_116_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n9960), .O(n62[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_8 (.CI(n9960), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n9961));
    SB_LUT4 sub_116_add_2_5_lut (.I0(n1291), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n9957), .O(n1_adj_1214)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_116_add_2_3_lut (.I0(n1291), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n9955), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_116_add_2_3 (.CI(n9955), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n9956));
    SB_CARRY sub_116_add_2_6 (.CI(n9958), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n9959));
    SB_DFFESR state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n4370), .D(n62[6]), .R(n7310));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFN sync_58 (.Q(SYNC_c), .C(SLM_CLK_c), .D(bluejay_data_out_31__N_734));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFSR state_FSM_i10 (.Q(n828[9]), .C(SLM_CLK_c), .D(n3035), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i9 (.Q(bluejay_data_out_31__N_737), .C(SLM_CLK_c), 
            .D(n895), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i8 (.Q(bluejay_data_out_31__N_736), .C(SLM_CLK_c), 
            .D(n3033), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i7 (.Q(bluejay_data_out_31__N_735), .C(SLM_CLK_c), 
            .D(n891), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i6 (.Q(n828[5]), .C(SLM_CLK_c), .D(n3031), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i5 (.Q(n828[4]), .C(SLM_CLK_c), .D(n3029), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i4 (.Q(bluejay_data_out_31__N_734), .C(SLM_CLK_c), 
            .D(n4228), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i3 (.Q(n828[2]), .C(SLM_CLK_c), .D(n10440), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i2 (.Q(n843), .C(SLM_CLK_c), .D(n10149), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFESR state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(SLM_CLK_c), 
            .E(n4370), .D(n62[7]), .R(n7310));   // src/bluejay_data.v(56[8] 123[4])
    SB_CARRY sub_116_add_2_5 (.CI(n9957), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n9958));
    SB_LUT4 sub_116_add_2_7_lut (.I0(n1291), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n9959), .O(n1_adj_1216)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_116_add_2_7 (.CI(n9959), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n9960));
    SB_LUT4 sub_116_add_2_6_lut (.I0(n1291), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n9958), .O(n1_adj_1215)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_116_add_2_2_lut (.I0(n1291), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n1_adj_1217)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_116_add_2_4_lut (.I0(n1291), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n9956), .O(n1_adj_1218)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_116_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n9955));
    SB_CARRY sub_116_add_2_4 (.CI(n9956), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n9957));
    SB_LUT4 i1_3_lut_adj_61 (.I0(\rd_sig_diff0_w[1] ), .I1(get_next_word), 
            .I2(\rd_sig_diff0_w[0] ), .I3(GND_net), .O(n15));   // src/fifo_dc_32_lut_gen.v(233[30:44])
    defparam i1_3_lut_adj_61.LUT_INIT = 16'h5d5d;
    SB_LUT4 i5_4_lut_adj_62 (.I0(\rd_sig_diff0_w[2] ), .I1(n10700), .I2(n15), 
            .I3(n10748), .O(\aempty_flag_impl.ae_flag_nxt_w ));   // src/fifo_dc_32_lut_gen.v(233[30:44])
    defparam i5_4_lut_adj_62.LUT_INIT = 16'h0010;
    SB_LUT4 equal_117_i13_2_lut (.I0(state_timeout_counter[6]), .I1(state_timeout_counter[7]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // src/bluejay_data.v(106[21:49])
    defparam equal_117_i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_63 (.I0(state_timeout_counter[3]), .I1(n13), .I2(state_timeout_counter[1]), 
            .I3(state_timeout_counter[2]), .O(n12_adj_1219));   // src/bluejay_data.v(106[21:49])
    defparam i5_4_lut_adj_63.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_64 (.I0(state_timeout_counter[4]), .I1(n12_adj_1219), 
            .I2(state_timeout_counter[5]), .I3(state_timeout_counter[0]), 
            .O(n771));   // src/bluejay_data.v(106[21:49])
    defparam i6_4_lut_adj_64.LUT_INIT = 16'hfeff;
    SB_DFFN get_next_word_57 (.Q(get_next_word), .C(SLM_CLK_c), .D(n4876));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFESS state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(SLM_CLK_c), 
            .E(n4370), .D(n1_adj_1217), .S(n4694));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 i1_2_lut_adj_65 (.I0(buffer_switch_done_latched), .I1(buffer_switch_done), 
            .I2(GND_net), .I3(GND_net), .O(n10554));   // src/bluejay_data.v(61[10] 122[8])
    defparam i1_2_lut_adj_65.LUT_INIT = 16'h2222;
    SB_DFFESR v_counter_i0 (.Q(v_counter[0]), .C(SLM_CLK_c), .E(n4408), 
            .D(v_counter_10__N_715[0]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFNESR bluejay_data_out_i11 (.Q(DATA10_c_10), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4672));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i10 (.Q(DATA9_c_9), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4671));   // src/bluejay_data.v(126[8] 148[4])
    SB_LUT4 i1_2_lut_adj_66 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_737), 
            .I2(GND_net), .I3(GND_net), .O(valid_N_740));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_2_lut_adj_66.LUT_INIT = 16'heeee;
    SB_DFFNESR bluejay_data_out_i12 (.Q(DATA11_c_11), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4670));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i13 (.Q(DATA12_c_12), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4669));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i14 (.Q(DATA13_c_13), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4668));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i15 (.Q(DATA14_c_14), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4667));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i9 (.Q(DATA8_c_8), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4666));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i16 (.Q(DATA15_c_15), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4665));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i8 (.Q(DATA7_c_7), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4664));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i7 (.Q(DATA6_c_6), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4663));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i6 (.Q(DATA5_c_5), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4662));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i5 (.Q(DATA4_c_4), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4661));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i4 (.Q(DATA3_c_3), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4660));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i3 (.Q(DATA2_c_2), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4659));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFNESR bluejay_data_out_i2 (.Q(DATA1_c_1), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_740), .R(n4658));   // src/bluejay_data.v(126[8] 148[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(buffer_switch_done_latched), .I1(n6564), 
            .I2(n1_adj_1218), .I3(GND_net), .O(n4_adj_1213));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3336_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n6564), 
            .I2(bluejay_data_out_31__N_735), .I3(n4370), .O(n4719));   // src/bluejay_data.v(66[9] 121[16])
    defparam i3336_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_adj_67 (.I0(bluejay_data_out_31__N_736), .I1(bluejay_data_out_31__N_735), 
            .I2(GND_net), .I3(GND_net), .O(n4876));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_2_lut_adj_67.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_4_lut_adj_68 (.I0(v_counter[9]), .I1(v_counter[0]), 
            .I2(v_counter[1]), .I3(v_counter[10]), .O(n10179));   // src/bluejay_data.v(108[25:41])
    defparam i1_3_lut_4_lut_adj_68.LUT_INIT = 16'hfffb;
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen2
//

module fifo_dc_32_lut_gen2 (dc32_fifo_almost_full, FIFO_CLK_c, reset_per_frame, 
            \REG.mem_16_7 , \rd_addr_r[0] , \REG.mem_6_2 , \REG.mem_7_2 , 
            \dc32_fifo_data_in[7] , \REG.mem_46_9 , \REG.mem_47_9 , \REG.mem_25_5 , 
            GND_net, t_rd_fifo_en_w, \REG.out_raw[0] , SLM_CLK_c, \REG.mem_45_9 , 
            \REG.mem_44_9 , \REG.mem_57_15 , \REG.mem_62_15 , \REG.mem_63_15 , 
            \REG.mem_6_1 , \REG.mem_7_1 , \REG.mem_5_1 , \REG.mem_4_1 , 
            \REG.mem_57_1 , \REG.mem_25_9 , \dc32_fifo_data_in[6] , \dc32_fifo_data_in[15] , 
            \REG.mem_46_3 , \REG.mem_47_3 , \REG.mem_45_3 , \REG.mem_44_3 , 
            \REG.mem_54_13 , \REG.mem_55_13 , \REG.mem_50_11 , \REG.mem_48_11 , 
            \dc32_fifo_data_in[5] , \REG.mem_42_12 , \REG.mem_43_12 , 
            \REG.mem_41_12 , \REG.mem_40_12 , \dc32_fifo_data_in[4] , 
            \dc32_fifo_data_in[3] , \dc32_fifo_data_in[2] , \rd_grey_sync_r[0] , 
            \REG.mem_57_6 , DEBUG_3_c, wr_grey_sync_r, \dc32_fifo_data_in[1] , 
            \REG.mem_54_11 , \REG.mem_55_11 , \aempty_flag_impl.ae_flag_nxt_w , 
            dc32_fifo_almost_empty, \REG.mem_14_12 , \REG.mem_15_12 , 
            \REG.mem_30_0 , \REG.mem_31_0 , \REG.mem_13_12 , \REG.mem_12_12 , 
            \REG.mem_3_5 , \REG.mem_6_5 , \REG.mem_7_5 , \REG.mem_4_5 , 
            \REG.mem_5_5 , \REG.mem_57_11 , n62, \REG.mem_62_13 , \REG.mem_63_13 , 
            \REG.mem_46_1 , \REG.mem_47_1 , \REG.mem_45_1 , \REG.mem_44_1 , 
            \dc32_fifo_data_in[0] , \REG.mem_3_11 , \REG.mem_6_11 , \REG.mem_7_11 , 
            n30, \REG.mem_5_2 , \REG.mem_4_2 , \REG.mem_18_5 , \REG.mem_62_1 , 
            \REG.mem_63_1 , \REG.mem_38_13 , \REG.mem_39_13 , \REG.mem_5_11 , 
            \REG.mem_4_11 , \dc32_fifo_data_in[8] , \REG.mem_14_5 , \REG.mem_15_5 , 
            \REG.mem_13_5 , \REG.mem_12_5 , \REG.mem_30_9 , \REG.mem_31_9 , 
            \wr_addr_nxt_c[5] , \REG.mem_46_12 , \REG.mem_47_12 , \REG.mem_45_12 , 
            \REG.mem_44_12 , \REG.mem_62_11 , \REG.mem_63_11 , \REG.mem_57_8 , 
            \REG.mem_62_6 , \REG.mem_63_6 , \REG.mem_62_8 , \REG.mem_63_8 , 
            \REG.mem_35_0 , \REG.mem_25_15 , \REG.mem_35_7 , \REG.mem_35_9 , 
            \REG.mem_18_12 , \REG.mem_16_12 , \REG.mem_14_8 , \REG.mem_15_8 , 
            \REG.mem_13_8 , \REG.mem_12_8 , \REG.mem_14_2 , \REG.mem_15_2 , 
            \REG.mem_13_2 , \REG.mem_12_2 , \REG.mem_38_7 , \REG.mem_39_7 , 
            \REG.mem_36_7 , \REG.mem_37_7 , \REG.mem_50_12 , \REG.mem_48_12 , 
            \REG.mem_62_9 , \REG.mem_63_9 , \REG.mem_6_9 , \REG.mem_7_9 , 
            \REG.mem_35_6 , \REG.mem_5_9 , \REG.mem_4_9 , \REG.mem_37_13 , 
            \REG.mem_36_13 , \REG.mem_42_8 , \REG.mem_43_8 , \REG.mem_41_8 , 
            \REG.mem_40_8 , \REG.mem_22_7 , \REG.mem_23_7 , \REG.mem_10_11 , 
            \REG.mem_11_11 , \REG.mem_9_11 , \REG.mem_8_11 , \REG.mem_3_15 , 
            \REG.mem_46_8 , \REG.mem_47_8 , \REG.mem_45_8 , \REG.mem_44_8 , 
            \REG.mem_46_5 , \REG.mem_47_5 , \REG.mem_45_5 , \REG.mem_44_5 , 
            \REG.mem_10_2 , \REG.mem_11_2 , \REG.mem_54_9 , \REG.mem_55_9 , 
            \REG.mem_57_9 , \REG.mem_57_14 , \REG.mem_30_15 , \REG.mem_31_15 , 
            \REG.mem_42_15 , \REG.mem_43_15 , \REG.mem_16_5 , \REG.mem_9_2 , 
            \REG.mem_8_2 , \REG.mem_62_12 , \REG.mem_63_12 , \wr_addr_nxt_c[3] , 
            \REG.mem_18_8 , \REG.mem_16_8 , \REG.mem_22_12 , \REG.mem_23_12 , 
            \REG.mem_25_2 , \REG.mem_30_2 , \REG.mem_31_2 , \dc32_fifo_data_in[14] , 
            \REG.mem_48_10 , \REG.mem_50_10 , \dc32_fifo_data_in[13] , 
            \REG.mem_54_10 , \REG.mem_55_10 , \REG.mem_14_11 , \REG.mem_15_11 , 
            \dc32_fifo_data_in[12] , \REG.mem_54_12 , \REG.mem_55_12 , 
            \REG.mem_13_11 , \REG.mem_12_11 , \REG.mem_35_15 , \REG.mem_38_6 , 
            \REG.mem_39_6 , \dc32_fifo_data_in[11] , \REG.mem_37_6 , \REG.mem_36_6 , 
            \REG.mem_57_13 , \dc32_fifo_data_in[10] , \dc32_fifo_data_in[9] , 
            \REG.mem_30_13 , \REG.mem_31_13 , \REG.mem_30_5 , \REG.mem_31_5 , 
            \REG.mem_48_7 , \REG.mem_50_7 , \REG.mem_54_7 , \REG.mem_55_7 , 
            n6106, VCC_net, \fifo_data_out[2] , n6103, \fifo_data_out[1] , 
            \REG.mem_35_13 , \REG.mem_3_3 , \rd_addr_r[6] , n4827, \fifo_data_out[3] , 
            \REG.mem_50_1 , n4830, \fifo_data_out[4] , n4841, \fifo_data_out[5] , 
            n4844, \fifo_data_out[6] , n4848, \fifo_data_out[7] , n4851, 
            \fifo_data_out[8] , n4854, \fifo_data_out[9] , n4858, \fifo_data_out[10] , 
            n4864, \fifo_data_out[11] , \REG.mem_62_14 , \REG.mem_63_14 , 
            \REG.mem_48_1 , \REG.mem_18_11 , \REG.mem_16_11 , \REG.mem_6_3 , 
            \REG.mem_7_3 , \REG.mem_5_3 , \REG.mem_4_3 , \REG.mem_42_2 , 
            \REG.mem_43_2 , \REG.mem_41_2 , \REG.mem_40_2 , n6070, \fifo_data_out[0] , 
            \REG.mem_46_2 , \REG.mem_47_2 , \REG.mem_45_2 , \REG.mem_44_2 , 
            \REG.mem_14_7 , \REG.mem_15_7 , n4872, \fifo_data_out[12] , 
            n4875, \fifo_data_out[13] , \REG.mem_13_7 , \REG.mem_12_7 , 
            n6034, \REG.mem_25_13 , n6032, \REG.mem_10_3 , \REG.mem_11_3 , 
            \REG.mem_9_3 , \REG.mem_8_3 , \REG.mem_50_9 , n6013, n6012, 
            n6011, n6010, n6009, n6008, n6007, \REG.mem_63_10 , 
            n6006, n6005, n6004, \REG.mem_63_7 , n6003, n6002, \REG.mem_63_5 , 
            \REG.mem_48_9 , \REG.mem_42_13 , \REG.mem_43_13 , \REG.mem_38_0 , 
            \REG.mem_39_0 , n6001, \REG.mem_63_4 , n6000, \REG.mem_63_3 , 
            n5999, \REG.mem_63_2 , n5998, n5997, \REG.mem_63_0 , n5996, 
            n5995, n5994, n5993, n5992, n5991, \REG.mem_62_10 , 
            n5990, n5989, n5988, \REG.mem_62_7 , n5987, n5986, \REG.mem_62_5 , 
            n5985, \REG.mem_62_4 , \REG.mem_41_13 , \REG.mem_40_13 , 
            \REG.mem_37_0 , \REG.mem_36_0 , \REG.mem_10_6 , \REG.mem_11_6 , 
            n5984, \REG.mem_62_3 , n5983, \REG.mem_62_2 , n5982, n5981, 
            \REG.mem_62_0 , \REG.mem_9_6 , \REG.mem_8_6 , \REG.mem_42_0 , 
            \REG.mem_43_0 , \REG.mem_22_8 , \REG.mem_23_8 , n5946, rp_sync1_r, 
            n5945, n5944, n5943, n5942, n5941, n5940, n5939, n5938, 
            n5921, n5920, n5919, \REG.mem_41_0 , \REG.mem_40_0 , n5917, 
            n5916, n5914, \REG.mem_8_14 , \REG.mem_9_14 , \REG.mem_25_1 , 
            \REG.mem_10_14 , \REG.mem_11_14 , n5894, n5893, n5892, 
            n5891, \REG.mem_57_12 , n5890, n5889, \REG.mem_57_10 , 
            n5888, n5887, n5886, \REG.mem_57_7 , \REG.mem_6_8 , \REG.mem_7_8 , 
            \REG.mem_38_15 , \REG.mem_39_15 , n5885, \REG.mem_5_8 , 
            \REG.mem_4_8 , \REG.mem_14_14 , \REG.mem_15_14 , n5884, 
            \REG.mem_57_5 , n5883, \REG.mem_57_4 , n5882, \REG.mem_57_3 , 
            n5881, \REG.mem_57_2 , n5880, n5879, \REG.mem_57_0 , \REG.mem_12_14 , 
            \REG.mem_13_14 , \REG.mem_37_15 , \REG.mem_36_15 , n5861, 
            wp_sync1_r, n5860, n5859, n5858, n5857, n5856, n5855, 
            \REG.mem_55_15 , n5854, \REG.mem_55_14 , n5853, \rd_sig_diff0_w[0] , 
            n5852, n5851, n5850, n5849, n5848, \REG.mem_55_8 , n5847, 
            n5846, \REG.mem_55_6 , n5845, \REG.mem_55_5 , n5844, \REG.mem_55_4 , 
            n5843, \REG.mem_55_3 , n5842, \REG.mem_55_2 , n5841, \REG.mem_55_1 , 
            n5840, \REG.mem_55_0 , n5839, n5838, \REG.mem_40_4 , \REG.mem_41_4 , 
            \REG.mem_42_4 , \REG.mem_43_4 , n5836, n5835, n5834, n5833, 
            n5832, \REG.mem_54_15 , n5831, \REG.mem_54_14 , n5830, 
            n5829, n5828, n5827, n5826, n5825, \REG.mem_54_8 , n5824, 
            n5823, \REG.mem_54_6 , n5822, \REG.mem_54_5 , n5821, \REG.mem_54_4 , 
            \REG.mem_46_4 , \REG.mem_47_4 , \REG.mem_44_4 , \REG.mem_45_4 , 
            n5820, \REG.mem_54_3 , n5819, \REG.mem_54_2 , n5818, \REG.mem_54_1 , 
            n5817, \REG.mem_54_0 , \REG.mem_25_4 , \REG.mem_30_4 , \REG.mem_31_4 , 
            \REG.mem_8_4 , \REG.mem_9_4 , \REG.mem_10_4 , \REG.mem_11_4 , 
            \REG.mem_14_4 , \REG.mem_15_4 , \REG.mem_12_4 , \REG.mem_13_4 , 
            n5768, \REG.mem_50_15 , n5767, \REG.mem_50_14 , n5766, 
            \REG.mem_50_13 , n5765, n5764, n5763, n5762, n5761, 
            \REG.mem_50_8 , n5760, n5759, \REG.mem_50_6 , n5758, \REG.mem_50_5 , 
            n5757, \REG.mem_50_4 , n10700, n5756, \REG.mem_50_3 , 
            n5755, \REG.mem_50_2 , n5754, n4893, \fifo_data_out[14] , 
            n4896, \fifo_data_out[15] , n5750, \REG.mem_50_0 , \REG.mem_38_5 , 
            \REG.mem_39_5 , n5733, \REG.mem_48_15 , n5732, \REG.mem_48_14 , 
            n5731, \REG.mem_48_13 , n5730, n5729, n5728, n5727, 
            n5726, \REG.mem_48_8 , n5725, n5724, \REG.mem_48_6 , n10748, 
            n5723, \REG.mem_48_5 , n5722, \REG.mem_48_4 , n5721, \REG.mem_48_3 , 
            n5720, \REG.mem_48_2 , n5719, \REG.mem_42_6 , \REG.mem_43_6 , 
            n5718, \REG.mem_48_0 , n5717, \REG.mem_47_15 , \REG.mem_41_6 , 
            \REG.mem_40_6 , n5716, \REG.mem_47_14 , n5715, \REG.mem_47_13 , 
            n5714, n5713, \REG.mem_47_11 , n5712, \REG.mem_47_10 , 
            n5711, n5710, n5709, \REG.mem_47_7 , n5708, \REG.mem_47_6 , 
            n5707, n5706, n5705, n5704, n5703, \REG.mem_25_12 , 
            \REG.mem_37_5 , \REG.mem_36_5 , n5702, \REG.mem_47_0 , n5701, 
            \REG.mem_46_15 , n5700, \REG.mem_46_14 , n5699, \REG.mem_46_13 , 
            n5698, n5697, \REG.mem_46_11 , n5696, \REG.mem_46_10 , 
            n5695, n5694, n5693, \REG.mem_46_7 , n5692, \REG.mem_46_6 , 
            n5691, n5690, n5689, n5688, n5687, n5686, \REG.mem_46_0 , 
            n5685, \REG.mem_45_15 , n5684, \REG.mem_45_14 , n5683, 
            \REG.mem_45_13 , n5682, n5681, \REG.mem_45_11 , n5680, 
            \REG.mem_45_10 , n5679, n5678, \REG.mem_6_15 , \REG.mem_7_15 , 
            \REG.mem_3_1 , n5677, \REG.mem_45_7 , \REG.mem_5_15 , \REG.mem_4_15 , 
            n5676, \REG.mem_45_6 , n5675, n5674, n5673, n5672, n5671, 
            n5670, \REG.mem_45_0 , n5668, \REG.mem_44_15 , n5667, 
            \REG.mem_44_14 , n5665, \REG.mem_44_13 , n5664, n5663, 
            \REG.mem_44_11 , n5661, \REG.mem_44_10 , n5660, n5659, 
            n5658, \REG.mem_44_7 , n5657, \REG.mem_44_6 , n5656, n5655, 
            n5654, n5653, n5652, n5651, \REG.mem_44_0 , n5650, n5649, 
            \REG.mem_43_14 , n5648, n5647, n5646, \REG.mem_43_11 , 
            n5645, \REG.mem_43_10 , n5644, \REG.mem_43_9 , \rd_addr_p1_w[0] , 
            \REG.mem_18_7 , n5643, n5642, \REG.mem_43_7 , n5641, n5640, 
            \REG.mem_43_5 , n5639, n5638, \REG.mem_43_3 , n5637, n5636, 
            \REG.mem_43_1 , n5635, n5634, n5633, \REG.mem_42_14 , 
            n5632, n5631, n5630, \REG.mem_42_11 , n5629, \REG.mem_42_10 , 
            n4916, \REG.mem_22_11 , \REG.mem_23_11 , n5628, \REG.mem_42_9 , 
            n5627, n5626, \REG.mem_42_7 , n5625, n5624, \REG.mem_42_5 , 
            n5623, n5622, \REG.mem_42_3 , n5621, n5620, \REG.mem_42_1 , 
            n5619, n5618, \REG.mem_41_15 , n5617, \REG.mem_41_14 , 
            n5616, n5615, n5614, \REG.mem_41_11 , n5613, \REG.mem_41_10 , 
            \REG.mem_25_6 , n5612, \REG.mem_41_9 , n5611, n5610, \REG.mem_41_7 , 
            n5609, n5608, \REG.mem_41_5 , n5607, n5606, \REG.mem_41_3 , 
            n5605, n5604, \REG.mem_41_1 , n5603, n5602, \REG.mem_40_15 , 
            n5601, \REG.mem_40_14 , n5600, n5599, n5598, \REG.mem_40_11 , 
            n5597, \REG.mem_40_10 , n4904, n4903, n4901, n4899, 
            n5596, \REG.mem_40_9 , n5595, n5594, \REG.mem_40_7 , n5593, 
            n5592, \REG.mem_40_5 , n5591, n5590, \REG.mem_40_3 , n5589, 
            n5588, \REG.mem_40_1 , n5587, n5586, n5585, \REG.mem_39_14 , 
            n5584, n5583, \REG.mem_39_12 , n5582, \REG.mem_39_11 , 
            n5581, \REG.mem_39_10 , n4898, DEBUG_5_c, \REG.mem_3_4 , 
            \REG.mem_6_4 , \REG.mem_7_4 , n5580, \REG.mem_39_9 , n5579, 
            \REG.mem_39_8 , n5578, n5577, n5576, n5575, \REG.mem_39_4 , 
            n5574, \REG.mem_39_3 , n5573, \REG.mem_39_2 , n5572, \REG.mem_39_1 , 
            n5570, n5569, n5568, \REG.mem_38_14 , n5567, n5566, 
            \REG.mem_38_12 , n5565, \REG.mem_38_11 , n5564, \REG.mem_38_10 , 
            \REG.mem_5_4 , \REG.mem_4_4 , n5563, \REG.mem_38_9 , n5562, 
            \REG.mem_38_8 , n5561, n5560, n5559, n5558, \REG.mem_38_4 , 
            n5557, \REG.mem_38_3 , n5556, \REG.mem_38_2 , n5555, \REG.mem_38_1 , 
            n5554, n5553, n5552, \REG.mem_37_14 , n5551, n5550, 
            \REG.mem_37_12 , n5549, \REG.mem_37_11 , \REG.out_raw[15] , 
            \REG.out_raw[14] , \REG.out_raw[13] , \REG.out_raw[12] , \REG.out_raw[11] , 
            n5548, \REG.mem_37_10 , n5547, \REG.mem_37_9 , n5546, 
            \REG.mem_37_8 , n5545, n5544, n5543, n5542, \REG.mem_37_4 , 
            n5541, \REG.mem_37_3 , n5540, \REG.mem_37_2 , n5539, \REG.mem_37_1 , 
            n5538, \REG.out_raw[10] , \REG.out_raw[9] , \REG.out_raw[8] , 
            \REG.out_raw[7] , \REG.out_raw[6] , \REG.out_raw[5] , \REG.out_raw[4] , 
            \REG.out_raw[3] , \REG.out_raw[2] , \REG.out_raw[1] , n5524, 
            n5523, \REG.mem_36_14 , n5522, n5521, \REG.mem_36_12 , 
            n5520, \REG.mem_36_11 , n5519, \REG.mem_36_10 , n5518, 
            \REG.mem_36_9 , n5517, \REG.mem_36_8 , n5516, \rd_sig_diff0_w[2] , 
            n5515, n5514, n5513, \REG.mem_36_4 , n5512, \REG.mem_36_3 , 
            n5511, \REG.mem_36_2 , n5510, \REG.mem_36_1 , n5509, n5505, 
            n5504, \REG.mem_35_14 , n5503, n5502, \REG.mem_35_12 , 
            n5501, \REG.mem_35_11 , n5500, \REG.mem_35_10 , \rd_sig_diff0_w[1] , 
            n5499, n5498, \REG.mem_35_8 , n5497, n5496, n5495, \REG.mem_35_5 , 
            n5494, \REG.mem_35_4 , n5493, \REG.mem_35_3 , n5492, \REG.mem_35_2 , 
            n5491, \REG.mem_35_1 , n5490, \REG.mem_25_11 , \REG.mem_10_13 , 
            \REG.mem_11_13 , \REG.mem_9_13 , \REG.mem_8_13 , n5440, 
            n5439, \REG.mem_31_14 , n5438, n5437, \REG.mem_31_12 , 
            n5436, \REG.mem_31_11 , n5435, \REG.mem_31_10 , n5434, 
            n5433, \REG.mem_31_8 , n5432, \REG.mem_31_7 , n5431, \REG.mem_31_6 , 
            n5430, n5429, n5428, \REG.mem_31_3 , n5427, n5426, \REG.mem_31_1 , 
            n5425, n5424, n5423, \REG.mem_30_14 , n5422, n5421, 
            \REG.mem_30_12 , n5420, \REG.mem_30_11 , DEBUG_1_c_c, write_to_dc32_fifo_latched_N_425, 
            \REG.mem_18_6 , n5419, \REG.mem_30_10 , n5418, n5417, 
            \REG.mem_30_8 , n5416, \REG.mem_30_7 , n5415, \REG.mem_30_6 , 
            n5414, n5413, n5412, \REG.mem_30_3 , n5411, n5410, \REG.mem_30_1 , 
            n5409, \REG.mem_16_6 , \wr_addr_nxt_c[1] , \REG.mem_10_9 , 
            \REG.mem_11_9 , \REG.mem_9_9 , \REG.mem_8_9 , \REG.mem_14_13 , 
            \REG.mem_15_13 , \REG.mem_13_13 , \REG.mem_12_13 , n56, 
            \REG.mem_14_9 , \REG.mem_15_9 , \REG.mem_10_15 , \REG.mem_11_15 , 
            \REG.mem_9_15 , \REG.mem_8_15 , \REG.mem_10_7 , \REG.mem_11_7 , 
            \REG.mem_13_9 , \REG.mem_12_9 , n5344, n5343, \REG.mem_25_14 , 
            n5342, n5341, n5340, n5339, \REG.mem_25_10 , n5338, 
            n5337, \REG.mem_25_8 , n5336, \REG.mem_25_7 , \REG.mem_18_13 , 
            \REG.mem_9_7 , \REG.mem_8_7 , \REG.mem_16_13 , n5335, n5334, 
            n5333, n5332, \REG.mem_25_3 , n5331, n5330, n5329, \REG.mem_25_0 , 
            n52, n20, n5306, \REG.mem_23_15 , n5305, \REG.mem_23_14 , 
            n5304, \REG.mem_23_13 , n5303, n5302, n5301, \REG.mem_23_10 , 
            n5300, \REG.mem_23_9 , n5299, n5298, n5297, \REG.mem_23_6 , 
            n5296, \REG.mem_23_5 , n5295, \REG.mem_23_4 , n5294, \REG.mem_23_3 , 
            n5293, \REG.mem_23_2 , n5292, \REG.mem_23_1 , n5291, \REG.mem_23_0 , 
            n5290, \REG.mem_22_15 , n5289, \REG.mem_22_14 , n5288, 
            \REG.mem_22_13 , n5287, n5286, n5285, \REG.mem_22_10 , 
            \rd_grey_sync_r[5] , \rd_grey_sync_r[4] , \rd_grey_sync_r[3] , 
            \rd_grey_sync_r[2] , \rd_grey_sync_r[1] , n5284, \REG.mem_22_9 , 
            n5283, n5282, n5281, \REG.mem_22_6 , n5280, \REG.mem_22_5 , 
            n5279, \REG.mem_22_4 , n5278, \REG.mem_22_3 , n5277, \REG.mem_22_2 , 
            n5276, \REG.mem_22_1 , n5275, \REG.mem_22_0 , \REG.mem_14_3 , 
            \REG.mem_15_3 , \REG.mem_13_3 , \REG.mem_12_3 , \REG.mem_10_8 , 
            \REG.mem_11_8 , \REG.mem_9_8 , \REG.mem_8_8 , get_next_word, 
            \REG.mem_16_2 , \REG.mem_18_2 , \REG.mem_18_3 , n5226, \REG.mem_18_15 , 
            n5225, \REG.mem_18_14 , n5224, n5223, n5222, n5221, 
            \REG.mem_18_10 , n5220, \REG.mem_18_9 , rd_fifo_en_w, \REG.mem_16_3 , 
            \REG.mem_16_15 , n5219, n5218, n5217, n5216, n5215, 
            \REG.mem_18_4 , n5214, n5213, n5212, \REG.mem_18_1 , n5211, 
            \REG.mem_18_0 , n5190, n5188, \REG.mem_16_14 , n5187, 
            n5186, n5185, n5184, \REG.mem_16_10 , \REG.mem_3_2 , \REG.mem_3_0 , 
            n5183, \REG.mem_16_9 , n5182, n5181, n5180, n5179, n5178, 
            \REG.mem_16_4 , n5177, n5176, \REG.mem_6_0 , \REG.mem_7_0 , 
            n5175, \REG.mem_16_1 , n5174, \REG.mem_16_0 , n5171, \REG.mem_15_15 , 
            n5170, n5169, n5168, n5167, n5166, \REG.mem_15_10 , 
            n5165, n5164, n5163, n5162, \REG.mem_15_6 , \REG.mem_5_0 , 
            \REG.mem_4_0 , n5161, n5160, n5159, n5158, n5157, \REG.mem_15_1 , 
            n5156, \REG.mem_15_0 , n5155, \REG.mem_14_15 , n5154, 
            n5153, n5152, n5151, n5150, \REG.mem_14_10 , n5149, 
            n5148, n5147, n5146, \REG.mem_14_6 , n5145, n5144, n5143, 
            n5142, n5141, \REG.mem_14_1 , n5140, \REG.mem_14_0 , n5139, 
            \REG.mem_13_15 , n5138, n5137, n5136, n5135, n5134, 
            \REG.mem_13_10 , n5133, n5132, n5131, n47, n15, n50, 
            n5130, \REG.mem_13_6 , n18, n5129, n5128, n5127, n5126, 
            n5125, \REG.mem_13_1 , n5124, \REG.mem_13_0 , n5123, \REG.mem_12_15 , 
            n5122, n5121, n5120, n5119, n5118, \REG.mem_12_10 , 
            n5117, n5116, \REG.mem_3_12 , \REG.mem_3_14 , n5115, n5114, 
            \REG.mem_12_6 , n5113, n5112, n53, n21, \REG.mem_10_0 , 
            \REG.mem_11_0 , \REG.mem_9_0 , \REG.mem_8_0 , n5111, n5110, 
            n5109, \REG.mem_12_1 , n5108, \REG.mem_12_0 , n51, n19, 
            n5107, n54, n22, n5106, n5105, n5104, \REG.mem_11_12 , 
            n5103, n5102, \REG.mem_11_10 , n5101, n5100, n5099, 
            n5098, n5097, \REG.mem_11_5 , \rd_addr_nxt_c_6__N_498[5] , 
            n5096, n5095, n5094, n5093, \REG.mem_11_1 , n5092, n5091, 
            n5090, n5089, n5088, \REG.mem_10_12 , n5087, n5086, 
            \REG.mem_10_10 , n5085, n5084, n5083, n5082, n5081, 
            \REG.mem_10_5 , n5080, \rd_addr_nxt_c_6__N_498[3] , n5079, 
            \rd_addr_nxt_c_6__N_498[2] , n49, n17, \REG.mem_6_14 , \REG.mem_7_14 , 
            \REG.mem_4_14 , \REG.mem_5_14 , n24, n5078, \REG.mem_3_6 , 
            n5077, \REG.mem_10_1 , n5076, n5075, \REG.mem_3_9 , n5074, 
            n5073, n55, n23, n40, n8, n5072, \REG.mem_9_12 , n34, 
            n5071, n5070, \REG.mem_9_10 , n5069, n2, n5068, n5067, 
            n5066, n5065, \REG.mem_9_5 , n5064, n5063, n5062, n5061, 
            \REG.mem_9_1 , n5060, n5059, n5058, n5057, n5056, \REG.mem_8_12 , 
            n5055, n5054, \REG.mem_8_10 , n5053, n5052, n5051, n5050, 
            n5049, \REG.mem_8_5 , n5048, n5047, n5046, n5045, \REG.mem_8_1 , 
            n5044, n5043, n5042, n5041, \REG.mem_7_13 , n5040, \REG.mem_7_12 , 
            n5039, n5038, \REG.mem_7_10 , n5037, n5036, n5035, \REG.mem_7_7 , 
            n5034, \REG.mem_7_6 , n5033, n5032, n5031, n5030, n5029, 
            n5028, n5027, n5026, n5025, \REG.mem_6_13 , n5024, \REG.mem_6_12 , 
            n5023, n5022, \REG.mem_6_10 , n5021, n5020, n5019, \REG.mem_6_7 , 
            n5018, \REG.mem_6_6 , n5017, n5016, n5015, n5014, n5013, 
            n5012, n5011, n5010, n5009, \REG.mem_5_13 , n5008, \REG.mem_5_12 , 
            n5007, n5006, \REG.mem_5_10 , n5005, n5004, n5003, \REG.mem_5_7 , 
            n5002, \REG.mem_5_6 , n5001, n5000, n4999, n4998, n4997, 
            n4996, n4995, n4994, n4993, \REG.mem_4_13 , n4992, \REG.mem_4_12 , 
            n4991, n4990, \REG.mem_4_10 , n4989, n4988, n4987, \REG.mem_4_7 , 
            n4986, \REG.mem_4_6 , n4985, n4984, n4983, n4982, n4981, 
            n4980, n4979, n4978, n4977, \REG.mem_3_13 , n4976, n4975, 
            n4974, \REG.mem_3_10 , n4973, n4972, \REG.mem_3_8 , n4971, 
            \REG.mem_3_7 , n4970, n4969, FT_OE_N_420, n57, n25, 
            n42, n10, n58, n26, n43, n35, n11, n3, n4968, 
            n4967, n4966, n4965, n4964, n60, n28, n59, n27, 
            n61, n29, n4672, n4671, n4670, n4669, n4668, n4667, 
            n4666, n4665, n4664, n4663, n4662, n4661, n4660, n4659, 
            n4658) /* synthesis syn_module_defined=1 */ ;
    output dc32_fifo_almost_full;
    input FIFO_CLK_c;
    input reset_per_frame;
    output \REG.mem_16_7 ;
    output \rd_addr_r[0] ;
    output \REG.mem_6_2 ;
    output \REG.mem_7_2 ;
    input \dc32_fifo_data_in[7] ;
    output \REG.mem_46_9 ;
    output \REG.mem_47_9 ;
    output \REG.mem_25_5 ;
    input GND_net;
    output t_rd_fifo_en_w;
    output \REG.out_raw[0] ;
    input SLM_CLK_c;
    output \REG.mem_45_9 ;
    output \REG.mem_44_9 ;
    output \REG.mem_57_15 ;
    output \REG.mem_62_15 ;
    output \REG.mem_63_15 ;
    output \REG.mem_6_1 ;
    output \REG.mem_7_1 ;
    output \REG.mem_5_1 ;
    output \REG.mem_4_1 ;
    output \REG.mem_57_1 ;
    output \REG.mem_25_9 ;
    input \dc32_fifo_data_in[6] ;
    input \dc32_fifo_data_in[15] ;
    output \REG.mem_46_3 ;
    output \REG.mem_47_3 ;
    output \REG.mem_45_3 ;
    output \REG.mem_44_3 ;
    output \REG.mem_54_13 ;
    output \REG.mem_55_13 ;
    output \REG.mem_50_11 ;
    output \REG.mem_48_11 ;
    input \dc32_fifo_data_in[5] ;
    output \REG.mem_42_12 ;
    output \REG.mem_43_12 ;
    output \REG.mem_41_12 ;
    output \REG.mem_40_12 ;
    input \dc32_fifo_data_in[4] ;
    input \dc32_fifo_data_in[3] ;
    input \dc32_fifo_data_in[2] ;
    output \rd_grey_sync_r[0] ;
    output \REG.mem_57_6 ;
    output DEBUG_3_c;
    output [6:0]wr_grey_sync_r;
    input \dc32_fifo_data_in[1] ;
    output \REG.mem_54_11 ;
    output \REG.mem_55_11 ;
    input \aempty_flag_impl.ae_flag_nxt_w ;
    output dc32_fifo_almost_empty;
    output \REG.mem_14_12 ;
    output \REG.mem_15_12 ;
    output \REG.mem_30_0 ;
    output \REG.mem_31_0 ;
    output \REG.mem_13_12 ;
    output \REG.mem_12_12 ;
    output \REG.mem_3_5 ;
    output \REG.mem_6_5 ;
    output \REG.mem_7_5 ;
    output \REG.mem_4_5 ;
    output \REG.mem_5_5 ;
    output \REG.mem_57_11 ;
    output n62;
    output \REG.mem_62_13 ;
    output \REG.mem_63_13 ;
    output \REG.mem_46_1 ;
    output \REG.mem_47_1 ;
    output \REG.mem_45_1 ;
    output \REG.mem_44_1 ;
    input \dc32_fifo_data_in[0] ;
    output \REG.mem_3_11 ;
    output \REG.mem_6_11 ;
    output \REG.mem_7_11 ;
    output n30;
    output \REG.mem_5_2 ;
    output \REG.mem_4_2 ;
    output \REG.mem_18_5 ;
    output \REG.mem_62_1 ;
    output \REG.mem_63_1 ;
    output \REG.mem_38_13 ;
    output \REG.mem_39_13 ;
    output \REG.mem_5_11 ;
    output \REG.mem_4_11 ;
    input \dc32_fifo_data_in[8] ;
    output \REG.mem_14_5 ;
    output \REG.mem_15_5 ;
    output \REG.mem_13_5 ;
    output \REG.mem_12_5 ;
    output \REG.mem_30_9 ;
    output \REG.mem_31_9 ;
    output \wr_addr_nxt_c[5] ;
    output \REG.mem_46_12 ;
    output \REG.mem_47_12 ;
    output \REG.mem_45_12 ;
    output \REG.mem_44_12 ;
    output \REG.mem_62_11 ;
    output \REG.mem_63_11 ;
    output \REG.mem_57_8 ;
    output \REG.mem_62_6 ;
    output \REG.mem_63_6 ;
    output \REG.mem_62_8 ;
    output \REG.mem_63_8 ;
    output \REG.mem_35_0 ;
    output \REG.mem_25_15 ;
    output \REG.mem_35_7 ;
    output \REG.mem_35_9 ;
    output \REG.mem_18_12 ;
    output \REG.mem_16_12 ;
    output \REG.mem_14_8 ;
    output \REG.mem_15_8 ;
    output \REG.mem_13_8 ;
    output \REG.mem_12_8 ;
    output \REG.mem_14_2 ;
    output \REG.mem_15_2 ;
    output \REG.mem_13_2 ;
    output \REG.mem_12_2 ;
    output \REG.mem_38_7 ;
    output \REG.mem_39_7 ;
    output \REG.mem_36_7 ;
    output \REG.mem_37_7 ;
    output \REG.mem_50_12 ;
    output \REG.mem_48_12 ;
    output \REG.mem_62_9 ;
    output \REG.mem_63_9 ;
    output \REG.mem_6_9 ;
    output \REG.mem_7_9 ;
    output \REG.mem_35_6 ;
    output \REG.mem_5_9 ;
    output \REG.mem_4_9 ;
    output \REG.mem_37_13 ;
    output \REG.mem_36_13 ;
    output \REG.mem_42_8 ;
    output \REG.mem_43_8 ;
    output \REG.mem_41_8 ;
    output \REG.mem_40_8 ;
    output \REG.mem_22_7 ;
    output \REG.mem_23_7 ;
    output \REG.mem_10_11 ;
    output \REG.mem_11_11 ;
    output \REG.mem_9_11 ;
    output \REG.mem_8_11 ;
    output \REG.mem_3_15 ;
    output \REG.mem_46_8 ;
    output \REG.mem_47_8 ;
    output \REG.mem_45_8 ;
    output \REG.mem_44_8 ;
    output \REG.mem_46_5 ;
    output \REG.mem_47_5 ;
    output \REG.mem_45_5 ;
    output \REG.mem_44_5 ;
    output \REG.mem_10_2 ;
    output \REG.mem_11_2 ;
    output \REG.mem_54_9 ;
    output \REG.mem_55_9 ;
    output \REG.mem_57_9 ;
    output \REG.mem_57_14 ;
    output \REG.mem_30_15 ;
    output \REG.mem_31_15 ;
    output \REG.mem_42_15 ;
    output \REG.mem_43_15 ;
    output \REG.mem_16_5 ;
    output \REG.mem_9_2 ;
    output \REG.mem_8_2 ;
    output \REG.mem_62_12 ;
    output \REG.mem_63_12 ;
    output \wr_addr_nxt_c[3] ;
    output \REG.mem_18_8 ;
    output \REG.mem_16_8 ;
    output \REG.mem_22_12 ;
    output \REG.mem_23_12 ;
    output \REG.mem_25_2 ;
    output \REG.mem_30_2 ;
    output \REG.mem_31_2 ;
    input \dc32_fifo_data_in[14] ;
    output \REG.mem_48_10 ;
    output \REG.mem_50_10 ;
    input \dc32_fifo_data_in[13] ;
    output \REG.mem_54_10 ;
    output \REG.mem_55_10 ;
    output \REG.mem_14_11 ;
    output \REG.mem_15_11 ;
    input \dc32_fifo_data_in[12] ;
    output \REG.mem_54_12 ;
    output \REG.mem_55_12 ;
    output \REG.mem_13_11 ;
    output \REG.mem_12_11 ;
    output \REG.mem_35_15 ;
    output \REG.mem_38_6 ;
    output \REG.mem_39_6 ;
    input \dc32_fifo_data_in[11] ;
    output \REG.mem_37_6 ;
    output \REG.mem_36_6 ;
    output \REG.mem_57_13 ;
    input \dc32_fifo_data_in[10] ;
    input \dc32_fifo_data_in[9] ;
    output \REG.mem_30_13 ;
    output \REG.mem_31_13 ;
    output \REG.mem_30_5 ;
    output \REG.mem_31_5 ;
    output \REG.mem_48_7 ;
    output \REG.mem_50_7 ;
    output \REG.mem_54_7 ;
    output \REG.mem_55_7 ;
    input n6106;
    input VCC_net;
    output \fifo_data_out[2] ;
    input n6103;
    output \fifo_data_out[1] ;
    output \REG.mem_35_13 ;
    output \REG.mem_3_3 ;
    output \rd_addr_r[6] ;
    input n4827;
    output \fifo_data_out[3] ;
    output \REG.mem_50_1 ;
    input n4830;
    output \fifo_data_out[4] ;
    input n4841;
    output \fifo_data_out[5] ;
    input n4844;
    output \fifo_data_out[6] ;
    input n4848;
    output \fifo_data_out[7] ;
    input n4851;
    output \fifo_data_out[8] ;
    input n4854;
    output \fifo_data_out[9] ;
    input n4858;
    output \fifo_data_out[10] ;
    input n4864;
    output \fifo_data_out[11] ;
    output \REG.mem_62_14 ;
    output \REG.mem_63_14 ;
    output \REG.mem_48_1 ;
    output \REG.mem_18_11 ;
    output \REG.mem_16_11 ;
    output \REG.mem_6_3 ;
    output \REG.mem_7_3 ;
    output \REG.mem_5_3 ;
    output \REG.mem_4_3 ;
    output \REG.mem_42_2 ;
    output \REG.mem_43_2 ;
    output \REG.mem_41_2 ;
    output \REG.mem_40_2 ;
    input n6070;
    output \fifo_data_out[0] ;
    output \REG.mem_46_2 ;
    output \REG.mem_47_2 ;
    output \REG.mem_45_2 ;
    output \REG.mem_44_2 ;
    output \REG.mem_14_7 ;
    output \REG.mem_15_7 ;
    input n4872;
    output \fifo_data_out[12] ;
    input n4875;
    output \fifo_data_out[13] ;
    output \REG.mem_13_7 ;
    output \REG.mem_12_7 ;
    input n6034;
    output \REG.mem_25_13 ;
    input n6032;
    output \REG.mem_10_3 ;
    output \REG.mem_11_3 ;
    output \REG.mem_9_3 ;
    output \REG.mem_8_3 ;
    output \REG.mem_50_9 ;
    input n6013;
    input n6012;
    input n6011;
    input n6010;
    input n6009;
    input n6008;
    input n6007;
    output \REG.mem_63_10 ;
    input n6006;
    input n6005;
    input n6004;
    output \REG.mem_63_7 ;
    input n6003;
    input n6002;
    output \REG.mem_63_5 ;
    output \REG.mem_48_9 ;
    output \REG.mem_42_13 ;
    output \REG.mem_43_13 ;
    output \REG.mem_38_0 ;
    output \REG.mem_39_0 ;
    input n6001;
    output \REG.mem_63_4 ;
    input n6000;
    output \REG.mem_63_3 ;
    input n5999;
    output \REG.mem_63_2 ;
    input n5998;
    input n5997;
    output \REG.mem_63_0 ;
    input n5996;
    input n5995;
    input n5994;
    input n5993;
    input n5992;
    input n5991;
    output \REG.mem_62_10 ;
    input n5990;
    input n5989;
    input n5988;
    output \REG.mem_62_7 ;
    input n5987;
    input n5986;
    output \REG.mem_62_5 ;
    input n5985;
    output \REG.mem_62_4 ;
    output \REG.mem_41_13 ;
    output \REG.mem_40_13 ;
    output \REG.mem_37_0 ;
    output \REG.mem_36_0 ;
    output \REG.mem_10_6 ;
    output \REG.mem_11_6 ;
    input n5984;
    output \REG.mem_62_3 ;
    input n5983;
    output \REG.mem_62_2 ;
    input n5982;
    input n5981;
    output \REG.mem_62_0 ;
    output \REG.mem_9_6 ;
    output \REG.mem_8_6 ;
    output \REG.mem_42_0 ;
    output \REG.mem_43_0 ;
    output \REG.mem_22_8 ;
    output \REG.mem_23_8 ;
    input n5946;
    output [6:0]rp_sync1_r;
    input n5945;
    input n5944;
    input n5943;
    input n5942;
    input n5941;
    input n5940;
    input n5939;
    input n5938;
    input n5921;
    input n5920;
    input n5919;
    output \REG.mem_41_0 ;
    output \REG.mem_40_0 ;
    input n5917;
    input n5916;
    input n5914;
    output \REG.mem_8_14 ;
    output \REG.mem_9_14 ;
    output \REG.mem_25_1 ;
    output \REG.mem_10_14 ;
    output \REG.mem_11_14 ;
    input n5894;
    input n5893;
    input n5892;
    input n5891;
    output \REG.mem_57_12 ;
    input n5890;
    input n5889;
    output \REG.mem_57_10 ;
    input n5888;
    input n5887;
    input n5886;
    output \REG.mem_57_7 ;
    output \REG.mem_6_8 ;
    output \REG.mem_7_8 ;
    output \REG.mem_38_15 ;
    output \REG.mem_39_15 ;
    input n5885;
    output \REG.mem_5_8 ;
    output \REG.mem_4_8 ;
    output \REG.mem_14_14 ;
    output \REG.mem_15_14 ;
    input n5884;
    output \REG.mem_57_5 ;
    input n5883;
    output \REG.mem_57_4 ;
    input n5882;
    output \REG.mem_57_3 ;
    input n5881;
    output \REG.mem_57_2 ;
    input n5880;
    input n5879;
    output \REG.mem_57_0 ;
    output \REG.mem_12_14 ;
    output \REG.mem_13_14 ;
    output \REG.mem_37_15 ;
    output \REG.mem_36_15 ;
    input n5861;
    output [6:0]wp_sync1_r;
    input n5860;
    input n5859;
    input n5858;
    input n5857;
    input n5856;
    input n5855;
    output \REG.mem_55_15 ;
    input n5854;
    output \REG.mem_55_14 ;
    input n5853;
    output \rd_sig_diff0_w[0] ;
    input n5852;
    input n5851;
    input n5850;
    input n5849;
    input n5848;
    output \REG.mem_55_8 ;
    input n5847;
    input n5846;
    output \REG.mem_55_6 ;
    input n5845;
    output \REG.mem_55_5 ;
    input n5844;
    output \REG.mem_55_4 ;
    input n5843;
    output \REG.mem_55_3 ;
    input n5842;
    output \REG.mem_55_2 ;
    input n5841;
    output \REG.mem_55_1 ;
    input n5840;
    output \REG.mem_55_0 ;
    input n5839;
    input n5838;
    output \REG.mem_40_4 ;
    output \REG.mem_41_4 ;
    output \REG.mem_42_4 ;
    output \REG.mem_43_4 ;
    input n5836;
    input n5835;
    input n5834;
    input n5833;
    input n5832;
    output \REG.mem_54_15 ;
    input n5831;
    output \REG.mem_54_14 ;
    input n5830;
    input n5829;
    input n5828;
    input n5827;
    input n5826;
    input n5825;
    output \REG.mem_54_8 ;
    input n5824;
    input n5823;
    output \REG.mem_54_6 ;
    input n5822;
    output \REG.mem_54_5 ;
    input n5821;
    output \REG.mem_54_4 ;
    output \REG.mem_46_4 ;
    output \REG.mem_47_4 ;
    output \REG.mem_44_4 ;
    output \REG.mem_45_4 ;
    input n5820;
    output \REG.mem_54_3 ;
    input n5819;
    output \REG.mem_54_2 ;
    input n5818;
    output \REG.mem_54_1 ;
    input n5817;
    output \REG.mem_54_0 ;
    output \REG.mem_25_4 ;
    output \REG.mem_30_4 ;
    output \REG.mem_31_4 ;
    output \REG.mem_8_4 ;
    output \REG.mem_9_4 ;
    output \REG.mem_10_4 ;
    output \REG.mem_11_4 ;
    output \REG.mem_14_4 ;
    output \REG.mem_15_4 ;
    output \REG.mem_12_4 ;
    output \REG.mem_13_4 ;
    input n5768;
    output \REG.mem_50_15 ;
    input n5767;
    output \REG.mem_50_14 ;
    input n5766;
    output \REG.mem_50_13 ;
    input n5765;
    input n5764;
    input n5763;
    input n5762;
    input n5761;
    output \REG.mem_50_8 ;
    input n5760;
    input n5759;
    output \REG.mem_50_6 ;
    input n5758;
    output \REG.mem_50_5 ;
    input n5757;
    output \REG.mem_50_4 ;
    output n10700;
    input n5756;
    output \REG.mem_50_3 ;
    input n5755;
    output \REG.mem_50_2 ;
    input n5754;
    input n4893;
    output \fifo_data_out[14] ;
    input n4896;
    output \fifo_data_out[15] ;
    input n5750;
    output \REG.mem_50_0 ;
    output \REG.mem_38_5 ;
    output \REG.mem_39_5 ;
    input n5733;
    output \REG.mem_48_15 ;
    input n5732;
    output \REG.mem_48_14 ;
    input n5731;
    output \REG.mem_48_13 ;
    input n5730;
    input n5729;
    input n5728;
    input n5727;
    input n5726;
    output \REG.mem_48_8 ;
    input n5725;
    input n5724;
    output \REG.mem_48_6 ;
    output n10748;
    input n5723;
    output \REG.mem_48_5 ;
    input n5722;
    output \REG.mem_48_4 ;
    input n5721;
    output \REG.mem_48_3 ;
    input n5720;
    output \REG.mem_48_2 ;
    input n5719;
    output \REG.mem_42_6 ;
    output \REG.mem_43_6 ;
    input n5718;
    output \REG.mem_48_0 ;
    input n5717;
    output \REG.mem_47_15 ;
    output \REG.mem_41_6 ;
    output \REG.mem_40_6 ;
    input n5716;
    output \REG.mem_47_14 ;
    input n5715;
    output \REG.mem_47_13 ;
    input n5714;
    input n5713;
    output \REG.mem_47_11 ;
    input n5712;
    output \REG.mem_47_10 ;
    input n5711;
    input n5710;
    input n5709;
    output \REG.mem_47_7 ;
    input n5708;
    output \REG.mem_47_6 ;
    input n5707;
    input n5706;
    input n5705;
    input n5704;
    input n5703;
    output \REG.mem_25_12 ;
    output \REG.mem_37_5 ;
    output \REG.mem_36_5 ;
    input n5702;
    output \REG.mem_47_0 ;
    input n5701;
    output \REG.mem_46_15 ;
    input n5700;
    output \REG.mem_46_14 ;
    input n5699;
    output \REG.mem_46_13 ;
    input n5698;
    input n5697;
    output \REG.mem_46_11 ;
    input n5696;
    output \REG.mem_46_10 ;
    input n5695;
    input n5694;
    input n5693;
    output \REG.mem_46_7 ;
    input n5692;
    output \REG.mem_46_6 ;
    input n5691;
    input n5690;
    input n5689;
    input n5688;
    input n5687;
    input n5686;
    output \REG.mem_46_0 ;
    input n5685;
    output \REG.mem_45_15 ;
    input n5684;
    output \REG.mem_45_14 ;
    input n5683;
    output \REG.mem_45_13 ;
    input n5682;
    input n5681;
    output \REG.mem_45_11 ;
    input n5680;
    output \REG.mem_45_10 ;
    input n5679;
    input n5678;
    output \REG.mem_6_15 ;
    output \REG.mem_7_15 ;
    output \REG.mem_3_1 ;
    input n5677;
    output \REG.mem_45_7 ;
    output \REG.mem_5_15 ;
    output \REG.mem_4_15 ;
    input n5676;
    output \REG.mem_45_6 ;
    input n5675;
    input n5674;
    input n5673;
    input n5672;
    input n5671;
    input n5670;
    output \REG.mem_45_0 ;
    input n5668;
    output \REG.mem_44_15 ;
    input n5667;
    output \REG.mem_44_14 ;
    input n5665;
    output \REG.mem_44_13 ;
    input n5664;
    input n5663;
    output \REG.mem_44_11 ;
    input n5661;
    output \REG.mem_44_10 ;
    input n5660;
    input n5659;
    input n5658;
    output \REG.mem_44_7 ;
    input n5657;
    output \REG.mem_44_6 ;
    input n5656;
    input n5655;
    input n5654;
    input n5653;
    input n5652;
    input n5651;
    output \REG.mem_44_0 ;
    input n5650;
    input n5649;
    output \REG.mem_43_14 ;
    input n5648;
    input n5647;
    input n5646;
    output \REG.mem_43_11 ;
    input n5645;
    output \REG.mem_43_10 ;
    input n5644;
    output \REG.mem_43_9 ;
    output \rd_addr_p1_w[0] ;
    output \REG.mem_18_7 ;
    input n5643;
    input n5642;
    output \REG.mem_43_7 ;
    input n5641;
    input n5640;
    output \REG.mem_43_5 ;
    input n5639;
    input n5638;
    output \REG.mem_43_3 ;
    input n5637;
    input n5636;
    output \REG.mem_43_1 ;
    input n5635;
    input n5634;
    input n5633;
    output \REG.mem_42_14 ;
    input n5632;
    input n5631;
    input n5630;
    output \REG.mem_42_11 ;
    input n5629;
    output \REG.mem_42_10 ;
    input n4916;
    output \REG.mem_22_11 ;
    output \REG.mem_23_11 ;
    input n5628;
    output \REG.mem_42_9 ;
    input n5627;
    input n5626;
    output \REG.mem_42_7 ;
    input n5625;
    input n5624;
    output \REG.mem_42_5 ;
    input n5623;
    input n5622;
    output \REG.mem_42_3 ;
    input n5621;
    input n5620;
    output \REG.mem_42_1 ;
    input n5619;
    input n5618;
    output \REG.mem_41_15 ;
    input n5617;
    output \REG.mem_41_14 ;
    input n5616;
    input n5615;
    input n5614;
    output \REG.mem_41_11 ;
    input n5613;
    output \REG.mem_41_10 ;
    output \REG.mem_25_6 ;
    input n5612;
    output \REG.mem_41_9 ;
    input n5611;
    input n5610;
    output \REG.mem_41_7 ;
    input n5609;
    input n5608;
    output \REG.mem_41_5 ;
    input n5607;
    input n5606;
    output \REG.mem_41_3 ;
    input n5605;
    input n5604;
    output \REG.mem_41_1 ;
    input n5603;
    input n5602;
    output \REG.mem_40_15 ;
    input n5601;
    output \REG.mem_40_14 ;
    input n5600;
    input n5599;
    input n5598;
    output \REG.mem_40_11 ;
    input n5597;
    output \REG.mem_40_10 ;
    input n4904;
    input n4903;
    input n4901;
    input n4899;
    input n5596;
    output \REG.mem_40_9 ;
    input n5595;
    input n5594;
    output \REG.mem_40_7 ;
    input n5593;
    input n5592;
    output \REG.mem_40_5 ;
    input n5591;
    input n5590;
    output \REG.mem_40_3 ;
    input n5589;
    input n5588;
    output \REG.mem_40_1 ;
    input n5587;
    input n5586;
    input n5585;
    output \REG.mem_39_14 ;
    input n5584;
    input n5583;
    output \REG.mem_39_12 ;
    input n5582;
    output \REG.mem_39_11 ;
    input n5581;
    output \REG.mem_39_10 ;
    input n4898;
    input DEBUG_5_c;
    output \REG.mem_3_4 ;
    output \REG.mem_6_4 ;
    output \REG.mem_7_4 ;
    input n5580;
    output \REG.mem_39_9 ;
    input n5579;
    output \REG.mem_39_8 ;
    input n5578;
    input n5577;
    input n5576;
    input n5575;
    output \REG.mem_39_4 ;
    input n5574;
    output \REG.mem_39_3 ;
    input n5573;
    output \REG.mem_39_2 ;
    input n5572;
    output \REG.mem_39_1 ;
    input n5570;
    input n5569;
    input n5568;
    output \REG.mem_38_14 ;
    input n5567;
    input n5566;
    output \REG.mem_38_12 ;
    input n5565;
    output \REG.mem_38_11 ;
    input n5564;
    output \REG.mem_38_10 ;
    output \REG.mem_5_4 ;
    output \REG.mem_4_4 ;
    input n5563;
    output \REG.mem_38_9 ;
    input n5562;
    output \REG.mem_38_8 ;
    input n5561;
    input n5560;
    input n5559;
    input n5558;
    output \REG.mem_38_4 ;
    input n5557;
    output \REG.mem_38_3 ;
    input n5556;
    output \REG.mem_38_2 ;
    input n5555;
    output \REG.mem_38_1 ;
    input n5554;
    input n5553;
    input n5552;
    output \REG.mem_37_14 ;
    input n5551;
    input n5550;
    output \REG.mem_37_12 ;
    input n5549;
    output \REG.mem_37_11 ;
    output \REG.out_raw[15] ;
    output \REG.out_raw[14] ;
    output \REG.out_raw[13] ;
    output \REG.out_raw[12] ;
    output \REG.out_raw[11] ;
    input n5548;
    output \REG.mem_37_10 ;
    input n5547;
    output \REG.mem_37_9 ;
    input n5546;
    output \REG.mem_37_8 ;
    input n5545;
    input n5544;
    input n5543;
    input n5542;
    output \REG.mem_37_4 ;
    input n5541;
    output \REG.mem_37_3 ;
    input n5540;
    output \REG.mem_37_2 ;
    input n5539;
    output \REG.mem_37_1 ;
    input n5538;
    output \REG.out_raw[10] ;
    output \REG.out_raw[9] ;
    output \REG.out_raw[8] ;
    output \REG.out_raw[7] ;
    output \REG.out_raw[6] ;
    output \REG.out_raw[5] ;
    output \REG.out_raw[4] ;
    output \REG.out_raw[3] ;
    output \REG.out_raw[2] ;
    output \REG.out_raw[1] ;
    input n5524;
    input n5523;
    output \REG.mem_36_14 ;
    input n5522;
    input n5521;
    output \REG.mem_36_12 ;
    input n5520;
    output \REG.mem_36_11 ;
    input n5519;
    output \REG.mem_36_10 ;
    input n5518;
    output \REG.mem_36_9 ;
    input n5517;
    output \REG.mem_36_8 ;
    input n5516;
    output \rd_sig_diff0_w[2] ;
    input n5515;
    input n5514;
    input n5513;
    output \REG.mem_36_4 ;
    input n5512;
    output \REG.mem_36_3 ;
    input n5511;
    output \REG.mem_36_2 ;
    input n5510;
    output \REG.mem_36_1 ;
    input n5509;
    input n5505;
    input n5504;
    output \REG.mem_35_14 ;
    input n5503;
    input n5502;
    output \REG.mem_35_12 ;
    input n5501;
    output \REG.mem_35_11 ;
    input n5500;
    output \REG.mem_35_10 ;
    output \rd_sig_diff0_w[1] ;
    input n5499;
    input n5498;
    output \REG.mem_35_8 ;
    input n5497;
    input n5496;
    input n5495;
    output \REG.mem_35_5 ;
    input n5494;
    output \REG.mem_35_4 ;
    input n5493;
    output \REG.mem_35_3 ;
    input n5492;
    output \REG.mem_35_2 ;
    input n5491;
    output \REG.mem_35_1 ;
    input n5490;
    output \REG.mem_25_11 ;
    output \REG.mem_10_13 ;
    output \REG.mem_11_13 ;
    output \REG.mem_9_13 ;
    output \REG.mem_8_13 ;
    input n5440;
    input n5439;
    output \REG.mem_31_14 ;
    input n5438;
    input n5437;
    output \REG.mem_31_12 ;
    input n5436;
    output \REG.mem_31_11 ;
    input n5435;
    output \REG.mem_31_10 ;
    input n5434;
    input n5433;
    output \REG.mem_31_8 ;
    input n5432;
    output \REG.mem_31_7 ;
    input n5431;
    output \REG.mem_31_6 ;
    input n5430;
    input n5429;
    input n5428;
    output \REG.mem_31_3 ;
    input n5427;
    input n5426;
    output \REG.mem_31_1 ;
    input n5425;
    input n5424;
    input n5423;
    output \REG.mem_30_14 ;
    input n5422;
    input n5421;
    output \REG.mem_30_12 ;
    input n5420;
    output \REG.mem_30_11 ;
    input DEBUG_1_c_c;
    output write_to_dc32_fifo_latched_N_425;
    output \REG.mem_18_6 ;
    input n5419;
    output \REG.mem_30_10 ;
    input n5418;
    input n5417;
    output \REG.mem_30_8 ;
    input n5416;
    output \REG.mem_30_7 ;
    input n5415;
    output \REG.mem_30_6 ;
    input n5414;
    input n5413;
    input n5412;
    output \REG.mem_30_3 ;
    input n5411;
    input n5410;
    output \REG.mem_30_1 ;
    input n5409;
    output \REG.mem_16_6 ;
    output \wr_addr_nxt_c[1] ;
    output \REG.mem_10_9 ;
    output \REG.mem_11_9 ;
    output \REG.mem_9_9 ;
    output \REG.mem_8_9 ;
    output \REG.mem_14_13 ;
    output \REG.mem_15_13 ;
    output \REG.mem_13_13 ;
    output \REG.mem_12_13 ;
    output n56;
    output \REG.mem_14_9 ;
    output \REG.mem_15_9 ;
    output \REG.mem_10_15 ;
    output \REG.mem_11_15 ;
    output \REG.mem_9_15 ;
    output \REG.mem_8_15 ;
    output \REG.mem_10_7 ;
    output \REG.mem_11_7 ;
    output \REG.mem_13_9 ;
    output \REG.mem_12_9 ;
    input n5344;
    input n5343;
    output \REG.mem_25_14 ;
    input n5342;
    input n5341;
    input n5340;
    input n5339;
    output \REG.mem_25_10 ;
    input n5338;
    input n5337;
    output \REG.mem_25_8 ;
    input n5336;
    output \REG.mem_25_7 ;
    output \REG.mem_18_13 ;
    output \REG.mem_9_7 ;
    output \REG.mem_8_7 ;
    output \REG.mem_16_13 ;
    input n5335;
    input n5334;
    input n5333;
    input n5332;
    output \REG.mem_25_3 ;
    input n5331;
    input n5330;
    input n5329;
    output \REG.mem_25_0 ;
    output n52;
    output n20;
    input n5306;
    output \REG.mem_23_15 ;
    input n5305;
    output \REG.mem_23_14 ;
    input n5304;
    output \REG.mem_23_13 ;
    input n5303;
    input n5302;
    input n5301;
    output \REG.mem_23_10 ;
    input n5300;
    output \REG.mem_23_9 ;
    input n5299;
    input n5298;
    input n5297;
    output \REG.mem_23_6 ;
    input n5296;
    output \REG.mem_23_5 ;
    input n5295;
    output \REG.mem_23_4 ;
    input n5294;
    output \REG.mem_23_3 ;
    input n5293;
    output \REG.mem_23_2 ;
    input n5292;
    output \REG.mem_23_1 ;
    input n5291;
    output \REG.mem_23_0 ;
    input n5290;
    output \REG.mem_22_15 ;
    input n5289;
    output \REG.mem_22_14 ;
    input n5288;
    output \REG.mem_22_13 ;
    input n5287;
    input n5286;
    input n5285;
    output \REG.mem_22_10 ;
    output \rd_grey_sync_r[5] ;
    output \rd_grey_sync_r[4] ;
    output \rd_grey_sync_r[3] ;
    output \rd_grey_sync_r[2] ;
    output \rd_grey_sync_r[1] ;
    input n5284;
    output \REG.mem_22_9 ;
    input n5283;
    input n5282;
    input n5281;
    output \REG.mem_22_6 ;
    input n5280;
    output \REG.mem_22_5 ;
    input n5279;
    output \REG.mem_22_4 ;
    input n5278;
    output \REG.mem_22_3 ;
    input n5277;
    output \REG.mem_22_2 ;
    input n5276;
    output \REG.mem_22_1 ;
    input n5275;
    output \REG.mem_22_0 ;
    output \REG.mem_14_3 ;
    output \REG.mem_15_3 ;
    output \REG.mem_13_3 ;
    output \REG.mem_12_3 ;
    output \REG.mem_10_8 ;
    output \REG.mem_11_8 ;
    output \REG.mem_9_8 ;
    output \REG.mem_8_8 ;
    input get_next_word;
    output \REG.mem_16_2 ;
    output \REG.mem_18_2 ;
    output \REG.mem_18_3 ;
    input n5226;
    output \REG.mem_18_15 ;
    input n5225;
    output \REG.mem_18_14 ;
    input n5224;
    input n5223;
    input n5222;
    input n5221;
    output \REG.mem_18_10 ;
    input n5220;
    output \REG.mem_18_9 ;
    output rd_fifo_en_w;
    output \REG.mem_16_3 ;
    output \REG.mem_16_15 ;
    input n5219;
    input n5218;
    input n5217;
    input n5216;
    input n5215;
    output \REG.mem_18_4 ;
    input n5214;
    input n5213;
    input n5212;
    output \REG.mem_18_1 ;
    input n5211;
    output \REG.mem_18_0 ;
    input n5190;
    input n5188;
    output \REG.mem_16_14 ;
    input n5187;
    input n5186;
    input n5185;
    input n5184;
    output \REG.mem_16_10 ;
    output \REG.mem_3_2 ;
    output \REG.mem_3_0 ;
    input n5183;
    output \REG.mem_16_9 ;
    input n5182;
    input n5181;
    input n5180;
    input n5179;
    input n5178;
    output \REG.mem_16_4 ;
    input n5177;
    input n5176;
    output \REG.mem_6_0 ;
    output \REG.mem_7_0 ;
    input n5175;
    output \REG.mem_16_1 ;
    input n5174;
    output \REG.mem_16_0 ;
    input n5171;
    output \REG.mem_15_15 ;
    input n5170;
    input n5169;
    input n5168;
    input n5167;
    input n5166;
    output \REG.mem_15_10 ;
    input n5165;
    input n5164;
    input n5163;
    input n5162;
    output \REG.mem_15_6 ;
    output \REG.mem_5_0 ;
    output \REG.mem_4_0 ;
    input n5161;
    input n5160;
    input n5159;
    input n5158;
    input n5157;
    output \REG.mem_15_1 ;
    input n5156;
    output \REG.mem_15_0 ;
    input n5155;
    output \REG.mem_14_15 ;
    input n5154;
    input n5153;
    input n5152;
    input n5151;
    input n5150;
    output \REG.mem_14_10 ;
    input n5149;
    input n5148;
    input n5147;
    input n5146;
    output \REG.mem_14_6 ;
    input n5145;
    input n5144;
    input n5143;
    input n5142;
    input n5141;
    output \REG.mem_14_1 ;
    input n5140;
    output \REG.mem_14_0 ;
    input n5139;
    output \REG.mem_13_15 ;
    input n5138;
    input n5137;
    input n5136;
    input n5135;
    input n5134;
    output \REG.mem_13_10 ;
    input n5133;
    input n5132;
    input n5131;
    output n47;
    output n15;
    output n50;
    input n5130;
    output \REG.mem_13_6 ;
    output n18;
    input n5129;
    input n5128;
    input n5127;
    input n5126;
    input n5125;
    output \REG.mem_13_1 ;
    input n5124;
    output \REG.mem_13_0 ;
    input n5123;
    output \REG.mem_12_15 ;
    input n5122;
    input n5121;
    input n5120;
    input n5119;
    input n5118;
    output \REG.mem_12_10 ;
    input n5117;
    input n5116;
    output \REG.mem_3_12 ;
    output \REG.mem_3_14 ;
    input n5115;
    input n5114;
    output \REG.mem_12_6 ;
    input n5113;
    input n5112;
    output n53;
    output n21;
    output \REG.mem_10_0 ;
    output \REG.mem_11_0 ;
    output \REG.mem_9_0 ;
    output \REG.mem_8_0 ;
    input n5111;
    input n5110;
    input n5109;
    output \REG.mem_12_1 ;
    input n5108;
    output \REG.mem_12_0 ;
    output n51;
    output n19;
    input n5107;
    output n54;
    output n22;
    input n5106;
    input n5105;
    input n5104;
    output \REG.mem_11_12 ;
    input n5103;
    input n5102;
    output \REG.mem_11_10 ;
    input n5101;
    input n5100;
    input n5099;
    input n5098;
    input n5097;
    output \REG.mem_11_5 ;
    output \rd_addr_nxt_c_6__N_498[5] ;
    input n5096;
    input n5095;
    input n5094;
    input n5093;
    output \REG.mem_11_1 ;
    input n5092;
    input n5091;
    input n5090;
    input n5089;
    input n5088;
    output \REG.mem_10_12 ;
    input n5087;
    input n5086;
    output \REG.mem_10_10 ;
    input n5085;
    input n5084;
    input n5083;
    input n5082;
    input n5081;
    output \REG.mem_10_5 ;
    input n5080;
    output \rd_addr_nxt_c_6__N_498[3] ;
    input n5079;
    output \rd_addr_nxt_c_6__N_498[2] ;
    output n49;
    output n17;
    output \REG.mem_6_14 ;
    output \REG.mem_7_14 ;
    output \REG.mem_4_14 ;
    output \REG.mem_5_14 ;
    output n24;
    input n5078;
    output \REG.mem_3_6 ;
    input n5077;
    output \REG.mem_10_1 ;
    input n5076;
    input n5075;
    output \REG.mem_3_9 ;
    input n5074;
    input n5073;
    output n55;
    output n23;
    output n40;
    output n8;
    input n5072;
    output \REG.mem_9_12 ;
    output n34;
    input n5071;
    input n5070;
    output \REG.mem_9_10 ;
    input n5069;
    output n2;
    input n5068;
    input n5067;
    input n5066;
    input n5065;
    output \REG.mem_9_5 ;
    input n5064;
    input n5063;
    input n5062;
    input n5061;
    output \REG.mem_9_1 ;
    input n5060;
    input n5059;
    input n5058;
    input n5057;
    input n5056;
    output \REG.mem_8_12 ;
    input n5055;
    input n5054;
    output \REG.mem_8_10 ;
    input n5053;
    input n5052;
    input n5051;
    input n5050;
    input n5049;
    output \REG.mem_8_5 ;
    input n5048;
    input n5047;
    input n5046;
    input n5045;
    output \REG.mem_8_1 ;
    input n5044;
    input n5043;
    input n5042;
    input n5041;
    output \REG.mem_7_13 ;
    input n5040;
    output \REG.mem_7_12 ;
    input n5039;
    input n5038;
    output \REG.mem_7_10 ;
    input n5037;
    input n5036;
    input n5035;
    output \REG.mem_7_7 ;
    input n5034;
    output \REG.mem_7_6 ;
    input n5033;
    input n5032;
    input n5031;
    input n5030;
    input n5029;
    input n5028;
    input n5027;
    input n5026;
    input n5025;
    output \REG.mem_6_13 ;
    input n5024;
    output \REG.mem_6_12 ;
    input n5023;
    input n5022;
    output \REG.mem_6_10 ;
    input n5021;
    input n5020;
    input n5019;
    output \REG.mem_6_7 ;
    input n5018;
    output \REG.mem_6_6 ;
    input n5017;
    input n5016;
    input n5015;
    input n5014;
    input n5013;
    input n5012;
    input n5011;
    input n5010;
    input n5009;
    output \REG.mem_5_13 ;
    input n5008;
    output \REG.mem_5_12 ;
    input n5007;
    input n5006;
    output \REG.mem_5_10 ;
    input n5005;
    input n5004;
    input n5003;
    output \REG.mem_5_7 ;
    input n5002;
    output \REG.mem_5_6 ;
    input n5001;
    input n5000;
    input n4999;
    input n4998;
    input n4997;
    input n4996;
    input n4995;
    input n4994;
    input n4993;
    output \REG.mem_4_13 ;
    input n4992;
    output \REG.mem_4_12 ;
    input n4991;
    input n4990;
    output \REG.mem_4_10 ;
    input n4989;
    input n4988;
    input n4987;
    output \REG.mem_4_7 ;
    input n4986;
    output \REG.mem_4_6 ;
    input n4985;
    input n4984;
    input n4983;
    input n4982;
    input n4981;
    input n4980;
    input n4979;
    input n4978;
    input n4977;
    output \REG.mem_3_13 ;
    input n4976;
    input n4975;
    input n4974;
    output \REG.mem_3_10 ;
    input n4973;
    input n4972;
    output \REG.mem_3_8 ;
    input n4971;
    output \REG.mem_3_7 ;
    input n4970;
    input n4969;
    output FT_OE_N_420;
    output n57;
    output n25;
    output n42;
    output n10;
    output n58;
    output n26;
    output n43;
    output n35;
    output n11;
    output n3;
    input n4968;
    input n4967;
    input n4966;
    input n4965;
    input n4964;
    output n60;
    output n28;
    output n59;
    output n27;
    output n61;
    output n29;
    output n4672;
    output n4671;
    output n4670;
    output n4669;
    output n4668;
    output n4667;
    output n4666;
    output n4665;
    output n4664;
    output n4663;
    output n4662;
    output n4661;
    output n4660;
    output n4659;
    output n4658;
    
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 lscc_fifo_dc_inst (.dc32_fifo_almost_full(dc32_fifo_almost_full), 
            .FIFO_CLK_c(FIFO_CLK_c), .reset_per_frame(reset_per_frame), 
            .\REG.mem_16_7 (\REG.mem_16_7 ), .\rd_addr_r[0] (\rd_addr_r[0] ), 
            .\REG.mem_6_2 (\REG.mem_6_2 ), .\REG.mem_7_2 (\REG.mem_7_2 ), 
            .\dc32_fifo_data_in[7] (\dc32_fifo_data_in[7] ), .\REG.mem_46_9 (\REG.mem_46_9 ), 
            .\REG.mem_47_9 (\REG.mem_47_9 ), .\REG.mem_25_5 (\REG.mem_25_5 ), 
            .GND_net(GND_net), .t_rd_fifo_en_w(t_rd_fifo_en_w), .\REG.out_raw[0] (\REG.out_raw[0] ), 
            .SLM_CLK_c(SLM_CLK_c), .\REG.mem_45_9 (\REG.mem_45_9 ), .\REG.mem_44_9 (\REG.mem_44_9 ), 
            .\REG.mem_57_15 (\REG.mem_57_15 ), .\REG.mem_62_15 (\REG.mem_62_15 ), 
            .\REG.mem_63_15 (\REG.mem_63_15 ), .\REG.mem_6_1 (\REG.mem_6_1 ), 
            .\REG.mem_7_1 (\REG.mem_7_1 ), .\REG.mem_5_1 (\REG.mem_5_1 ), 
            .\REG.mem_4_1 (\REG.mem_4_1 ), .\REG.mem_57_1 (\REG.mem_57_1 ), 
            .\REG.mem_25_9 (\REG.mem_25_9 ), .\dc32_fifo_data_in[6] (\dc32_fifo_data_in[6] ), 
            .\dc32_fifo_data_in[15] (\dc32_fifo_data_in[15] ), .\REG.mem_46_3 (\REG.mem_46_3 ), 
            .\REG.mem_47_3 (\REG.mem_47_3 ), .\REG.mem_45_3 (\REG.mem_45_3 ), 
            .\REG.mem_44_3 (\REG.mem_44_3 ), .\REG.mem_54_13 (\REG.mem_54_13 ), 
            .\REG.mem_55_13 (\REG.mem_55_13 ), .\REG.mem_50_11 (\REG.mem_50_11 ), 
            .\REG.mem_48_11 (\REG.mem_48_11 ), .\dc32_fifo_data_in[5] (\dc32_fifo_data_in[5] ), 
            .\REG.mem_42_12 (\REG.mem_42_12 ), .\REG.mem_43_12 (\REG.mem_43_12 ), 
            .\REG.mem_41_12 (\REG.mem_41_12 ), .\REG.mem_40_12 (\REG.mem_40_12 ), 
            .\dc32_fifo_data_in[4] (\dc32_fifo_data_in[4] ), .\dc32_fifo_data_in[3] (\dc32_fifo_data_in[3] ), 
            .\dc32_fifo_data_in[2] (\dc32_fifo_data_in[2] ), .\rd_grey_sync_r[0] (\rd_grey_sync_r[0] ), 
            .\REG.mem_57_6 (\REG.mem_57_6 ), .DEBUG_3_c(DEBUG_3_c), .wr_grey_sync_r({wr_grey_sync_r}), 
            .\dc32_fifo_data_in[1] (\dc32_fifo_data_in[1] ), .\REG.mem_54_11 (\REG.mem_54_11 ), 
            .\REG.mem_55_11 (\REG.mem_55_11 ), .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .dc32_fifo_almost_empty(dc32_fifo_almost_empty), .\REG.mem_14_12 (\REG.mem_14_12 ), 
            .\REG.mem_15_12 (\REG.mem_15_12 ), .\REG.mem_30_0 (\REG.mem_30_0 ), 
            .\REG.mem_31_0 (\REG.mem_31_0 ), .\REG.mem_13_12 (\REG.mem_13_12 ), 
            .\REG.mem_12_12 (\REG.mem_12_12 ), .\REG.mem_3_5 (\REG.mem_3_5 ), 
            .\REG.mem_6_5 (\REG.mem_6_5 ), .\REG.mem_7_5 (\REG.mem_7_5 ), 
            .\REG.mem_4_5 (\REG.mem_4_5 ), .\REG.mem_5_5 (\REG.mem_5_5 ), 
            .\REG.mem_57_11 (\REG.mem_57_11 ), .n62(n62), .\REG.mem_62_13 (\REG.mem_62_13 ), 
            .\REG.mem_63_13 (\REG.mem_63_13 ), .\REG.mem_46_1 (\REG.mem_46_1 ), 
            .\REG.mem_47_1 (\REG.mem_47_1 ), .\REG.mem_45_1 (\REG.mem_45_1 ), 
            .\REG.mem_44_1 (\REG.mem_44_1 ), .\dc32_fifo_data_in[0] (\dc32_fifo_data_in[0] ), 
            .\REG.mem_3_11 (\REG.mem_3_11 ), .\REG.mem_6_11 (\REG.mem_6_11 ), 
            .\REG.mem_7_11 (\REG.mem_7_11 ), .n30(n30), .\REG.mem_5_2 (\REG.mem_5_2 ), 
            .\REG.mem_4_2 (\REG.mem_4_2 ), .\REG.mem_18_5 (\REG.mem_18_5 ), 
            .\REG.mem_62_1 (\REG.mem_62_1 ), .\REG.mem_63_1 (\REG.mem_63_1 ), 
            .\REG.mem_38_13 (\REG.mem_38_13 ), .\REG.mem_39_13 (\REG.mem_39_13 ), 
            .\REG.mem_5_11 (\REG.mem_5_11 ), .\REG.mem_4_11 (\REG.mem_4_11 ), 
            .\dc32_fifo_data_in[8] (\dc32_fifo_data_in[8] ), .\REG.mem_14_5 (\REG.mem_14_5 ), 
            .\REG.mem_15_5 (\REG.mem_15_5 ), .\REG.mem_13_5 (\REG.mem_13_5 ), 
            .\REG.mem_12_5 (\REG.mem_12_5 ), .\REG.mem_30_9 (\REG.mem_30_9 ), 
            .\REG.mem_31_9 (\REG.mem_31_9 ), .\wr_addr_nxt_c[5] (\wr_addr_nxt_c[5] ), 
            .\REG.mem_46_12 (\REG.mem_46_12 ), .\REG.mem_47_12 (\REG.mem_47_12 ), 
            .\REG.mem_45_12 (\REG.mem_45_12 ), .\REG.mem_44_12 (\REG.mem_44_12 ), 
            .\REG.mem_62_11 (\REG.mem_62_11 ), .\REG.mem_63_11 (\REG.mem_63_11 ), 
            .\REG.mem_57_8 (\REG.mem_57_8 ), .\REG.mem_62_6 (\REG.mem_62_6 ), 
            .\REG.mem_63_6 (\REG.mem_63_6 ), .\REG.mem_62_8 (\REG.mem_62_8 ), 
            .\REG.mem_63_8 (\REG.mem_63_8 ), .\REG.mem_35_0 (\REG.mem_35_0 ), 
            .\REG.mem_25_15 (\REG.mem_25_15 ), .\REG.mem_35_7 (\REG.mem_35_7 ), 
            .\REG.mem_35_9 (\REG.mem_35_9 ), .\REG.mem_18_12 (\REG.mem_18_12 ), 
            .\REG.mem_16_12 (\REG.mem_16_12 ), .\REG.mem_14_8 (\REG.mem_14_8 ), 
            .\REG.mem_15_8 (\REG.mem_15_8 ), .\REG.mem_13_8 (\REG.mem_13_8 ), 
            .\REG.mem_12_8 (\REG.mem_12_8 ), .\REG.mem_14_2 (\REG.mem_14_2 ), 
            .\REG.mem_15_2 (\REG.mem_15_2 ), .\REG.mem_13_2 (\REG.mem_13_2 ), 
            .\REG.mem_12_2 (\REG.mem_12_2 ), .\REG.mem_38_7 (\REG.mem_38_7 ), 
            .\REG.mem_39_7 (\REG.mem_39_7 ), .\REG.mem_36_7 (\REG.mem_36_7 ), 
            .\REG.mem_37_7 (\REG.mem_37_7 ), .\REG.mem_50_12 (\REG.mem_50_12 ), 
            .\REG.mem_48_12 (\REG.mem_48_12 ), .\REG.mem_62_9 (\REG.mem_62_9 ), 
            .\REG.mem_63_9 (\REG.mem_63_9 ), .\REG.mem_6_9 (\REG.mem_6_9 ), 
            .\REG.mem_7_9 (\REG.mem_7_9 ), .\REG.mem_35_6 (\REG.mem_35_6 ), 
            .\REG.mem_5_9 (\REG.mem_5_9 ), .\REG.mem_4_9 (\REG.mem_4_9 ), 
            .\REG.mem_37_13 (\REG.mem_37_13 ), .\REG.mem_36_13 (\REG.mem_36_13 ), 
            .\REG.mem_42_8 (\REG.mem_42_8 ), .\REG.mem_43_8 (\REG.mem_43_8 ), 
            .\REG.mem_41_8 (\REG.mem_41_8 ), .\REG.mem_40_8 (\REG.mem_40_8 ), 
            .\REG.mem_22_7 (\REG.mem_22_7 ), .\REG.mem_23_7 (\REG.mem_23_7 ), 
            .\REG.mem_10_11 (\REG.mem_10_11 ), .\REG.mem_11_11 (\REG.mem_11_11 ), 
            .\REG.mem_9_11 (\REG.mem_9_11 ), .\REG.mem_8_11 (\REG.mem_8_11 ), 
            .\REG.mem_3_15 (\REG.mem_3_15 ), .\REG.mem_46_8 (\REG.mem_46_8 ), 
            .\REG.mem_47_8 (\REG.mem_47_8 ), .\REG.mem_45_8 (\REG.mem_45_8 ), 
            .\REG.mem_44_8 (\REG.mem_44_8 ), .\REG.mem_46_5 (\REG.mem_46_5 ), 
            .\REG.mem_47_5 (\REG.mem_47_5 ), .\REG.mem_45_5 (\REG.mem_45_5 ), 
            .\REG.mem_44_5 (\REG.mem_44_5 ), .\REG.mem_10_2 (\REG.mem_10_2 ), 
            .\REG.mem_11_2 (\REG.mem_11_2 ), .\REG.mem_54_9 (\REG.mem_54_9 ), 
            .\REG.mem_55_9 (\REG.mem_55_9 ), .\REG.mem_57_9 (\REG.mem_57_9 ), 
            .\REG.mem_57_14 (\REG.mem_57_14 ), .\REG.mem_30_15 (\REG.mem_30_15 ), 
            .\REG.mem_31_15 (\REG.mem_31_15 ), .\REG.mem_42_15 (\REG.mem_42_15 ), 
            .\REG.mem_43_15 (\REG.mem_43_15 ), .\REG.mem_16_5 (\REG.mem_16_5 ), 
            .\REG.mem_9_2 (\REG.mem_9_2 ), .\REG.mem_8_2 (\REG.mem_8_2 ), 
            .\REG.mem_62_12 (\REG.mem_62_12 ), .\REG.mem_63_12 (\REG.mem_63_12 ), 
            .\wr_addr_nxt_c[3] (\wr_addr_nxt_c[3] ), .\REG.mem_18_8 (\REG.mem_18_8 ), 
            .\REG.mem_16_8 (\REG.mem_16_8 ), .\REG.mem_22_12 (\REG.mem_22_12 ), 
            .\REG.mem_23_12 (\REG.mem_23_12 ), .\REG.mem_25_2 (\REG.mem_25_2 ), 
            .\REG.mem_30_2 (\REG.mem_30_2 ), .\REG.mem_31_2 (\REG.mem_31_2 ), 
            .\dc32_fifo_data_in[14] (\dc32_fifo_data_in[14] ), .\REG.mem_48_10 (\REG.mem_48_10 ), 
            .\REG.mem_50_10 (\REG.mem_50_10 ), .\dc32_fifo_data_in[13] (\dc32_fifo_data_in[13] ), 
            .\REG.mem_54_10 (\REG.mem_54_10 ), .\REG.mem_55_10 (\REG.mem_55_10 ), 
            .\REG.mem_14_11 (\REG.mem_14_11 ), .\REG.mem_15_11 (\REG.mem_15_11 ), 
            .\dc32_fifo_data_in[12] (\dc32_fifo_data_in[12] ), .\REG.mem_54_12 (\REG.mem_54_12 ), 
            .\REG.mem_55_12 (\REG.mem_55_12 ), .\REG.mem_13_11 (\REG.mem_13_11 ), 
            .\REG.mem_12_11 (\REG.mem_12_11 ), .\REG.mem_35_15 (\REG.mem_35_15 ), 
            .\REG.mem_38_6 (\REG.mem_38_6 ), .\REG.mem_39_6 (\REG.mem_39_6 ), 
            .\dc32_fifo_data_in[11] (\dc32_fifo_data_in[11] ), .\REG.mem_37_6 (\REG.mem_37_6 ), 
            .\REG.mem_36_6 (\REG.mem_36_6 ), .\REG.mem_57_13 (\REG.mem_57_13 ), 
            .\dc32_fifo_data_in[10] (\dc32_fifo_data_in[10] ), .\dc32_fifo_data_in[9] (\dc32_fifo_data_in[9] ), 
            .\REG.mem_30_13 (\REG.mem_30_13 ), .\REG.mem_31_13 (\REG.mem_31_13 ), 
            .\REG.mem_30_5 (\REG.mem_30_5 ), .\REG.mem_31_5 (\REG.mem_31_5 ), 
            .\REG.mem_48_7 (\REG.mem_48_7 ), .\REG.mem_50_7 (\REG.mem_50_7 ), 
            .\REG.mem_54_7 (\REG.mem_54_7 ), .\REG.mem_55_7 (\REG.mem_55_7 ), 
            .n6106(n6106), .VCC_net(VCC_net), .\fifo_data_out[2] (\fifo_data_out[2] ), 
            .n6103(n6103), .\fifo_data_out[1] (\fifo_data_out[1] ), .\REG.mem_35_13 (\REG.mem_35_13 ), 
            .\REG.mem_3_3 (\REG.mem_3_3 ), .\rd_addr_r[6] (\rd_addr_r[6] ), 
            .n4827(n4827), .\fifo_data_out[3] (\fifo_data_out[3] ), .\REG.mem_50_1 (\REG.mem_50_1 ), 
            .n4830(n4830), .\fifo_data_out[4] (\fifo_data_out[4] ), .n4841(n4841), 
            .\fifo_data_out[5] (\fifo_data_out[5] ), .n4844(n4844), .\fifo_data_out[6] (\fifo_data_out[6] ), 
            .n4848(n4848), .\fifo_data_out[7] (\fifo_data_out[7] ), .n4851(n4851), 
            .\fifo_data_out[8] (\fifo_data_out[8] ), .n4854(n4854), .\fifo_data_out[9] (\fifo_data_out[9] ), 
            .n4858(n4858), .\fifo_data_out[10] (\fifo_data_out[10] ), .n4864(n4864), 
            .\fifo_data_out[11] (\fifo_data_out[11] ), .\REG.mem_62_14 (\REG.mem_62_14 ), 
            .\REG.mem_63_14 (\REG.mem_63_14 ), .\REG.mem_48_1 (\REG.mem_48_1 ), 
            .\REG.mem_18_11 (\REG.mem_18_11 ), .\REG.mem_16_11 (\REG.mem_16_11 ), 
            .\REG.mem_6_3 (\REG.mem_6_3 ), .\REG.mem_7_3 (\REG.mem_7_3 ), 
            .\REG.mem_5_3 (\REG.mem_5_3 ), .\REG.mem_4_3 (\REG.mem_4_3 ), 
            .\REG.mem_42_2 (\REG.mem_42_2 ), .\REG.mem_43_2 (\REG.mem_43_2 ), 
            .\REG.mem_41_2 (\REG.mem_41_2 ), .\REG.mem_40_2 (\REG.mem_40_2 ), 
            .n6070(n6070), .\fifo_data_out[0] (\fifo_data_out[0] ), .\REG.mem_46_2 (\REG.mem_46_2 ), 
            .\REG.mem_47_2 (\REG.mem_47_2 ), .\REG.mem_45_2 (\REG.mem_45_2 ), 
            .\REG.mem_44_2 (\REG.mem_44_2 ), .\REG.mem_14_7 (\REG.mem_14_7 ), 
            .\REG.mem_15_7 (\REG.mem_15_7 ), .n4872(n4872), .\fifo_data_out[12] (\fifo_data_out[12] ), 
            .n4875(n4875), .\fifo_data_out[13] (\fifo_data_out[13] ), .\REG.mem_13_7 (\REG.mem_13_7 ), 
            .\REG.mem_12_7 (\REG.mem_12_7 ), .n6034(n6034), .\REG.mem_25_13 (\REG.mem_25_13 ), 
            .n6032(n6032), .\REG.mem_10_3 (\REG.mem_10_3 ), .\REG.mem_11_3 (\REG.mem_11_3 ), 
            .\REG.mem_9_3 (\REG.mem_9_3 ), .\REG.mem_8_3 (\REG.mem_8_3 ), 
            .\REG.mem_50_9 (\REG.mem_50_9 ), .n6013(n6013), .n6012(n6012), 
            .n6011(n6011), .n6010(n6010), .n6009(n6009), .n6008(n6008), 
            .n6007(n6007), .\REG.mem_63_10 (\REG.mem_63_10 ), .n6006(n6006), 
            .n6005(n6005), .n6004(n6004), .\REG.mem_63_7 (\REG.mem_63_7 ), 
            .n6003(n6003), .n6002(n6002), .\REG.mem_63_5 (\REG.mem_63_5 ), 
            .\REG.mem_48_9 (\REG.mem_48_9 ), .\REG.mem_42_13 (\REG.mem_42_13 ), 
            .\REG.mem_43_13 (\REG.mem_43_13 ), .\REG.mem_38_0 (\REG.mem_38_0 ), 
            .\REG.mem_39_0 (\REG.mem_39_0 ), .n6001(n6001), .\REG.mem_63_4 (\REG.mem_63_4 ), 
            .n6000(n6000), .\REG.mem_63_3 (\REG.mem_63_3 ), .n5999(n5999), 
            .\REG.mem_63_2 (\REG.mem_63_2 ), .n5998(n5998), .n5997(n5997), 
            .\REG.mem_63_0 (\REG.mem_63_0 ), .n5996(n5996), .n5995(n5995), 
            .n5994(n5994), .n5993(n5993), .n5992(n5992), .n5991(n5991), 
            .\REG.mem_62_10 (\REG.mem_62_10 ), .n5990(n5990), .n5989(n5989), 
            .n5988(n5988), .\REG.mem_62_7 (\REG.mem_62_7 ), .n5987(n5987), 
            .n5986(n5986), .\REG.mem_62_5 (\REG.mem_62_5 ), .n5985(n5985), 
            .\REG.mem_62_4 (\REG.mem_62_4 ), .\REG.mem_41_13 (\REG.mem_41_13 ), 
            .\REG.mem_40_13 (\REG.mem_40_13 ), .\REG.mem_37_0 (\REG.mem_37_0 ), 
            .\REG.mem_36_0 (\REG.mem_36_0 ), .\REG.mem_10_6 (\REG.mem_10_6 ), 
            .\REG.mem_11_6 (\REG.mem_11_6 ), .n5984(n5984), .\REG.mem_62_3 (\REG.mem_62_3 ), 
            .n5983(n5983), .\REG.mem_62_2 (\REG.mem_62_2 ), .n5982(n5982), 
            .n5981(n5981), .\REG.mem_62_0 (\REG.mem_62_0 ), .\REG.mem_9_6 (\REG.mem_9_6 ), 
            .\REG.mem_8_6 (\REG.mem_8_6 ), .\REG.mem_42_0 (\REG.mem_42_0 ), 
            .\REG.mem_43_0 (\REG.mem_43_0 ), .\REG.mem_22_8 (\REG.mem_22_8 ), 
            .\REG.mem_23_8 (\REG.mem_23_8 ), .n5946(n5946), .rp_sync1_r({rp_sync1_r}), 
            .n5945(n5945), .n5944(n5944), .n5943(n5943), .n5942(n5942), 
            .n5941(n5941), .n5940(n5940), .n5939(n5939), .n5938(n5938), 
            .n5921(n5921), .n5920(n5920), .n5919(n5919), .\REG.mem_41_0 (\REG.mem_41_0 ), 
            .\REG.mem_40_0 (\REG.mem_40_0 ), .n5917(n5917), .n5916(n5916), 
            .n5914(n5914), .\REG.mem_8_14 (\REG.mem_8_14 ), .\REG.mem_9_14 (\REG.mem_9_14 ), 
            .\REG.mem_25_1 (\REG.mem_25_1 ), .\REG.mem_10_14 (\REG.mem_10_14 ), 
            .\REG.mem_11_14 (\REG.mem_11_14 ), .n5894(n5894), .n5893(n5893), 
            .n5892(n5892), .n5891(n5891), .\REG.mem_57_12 (\REG.mem_57_12 ), 
            .n5890(n5890), .n5889(n5889), .\REG.mem_57_10 (\REG.mem_57_10 ), 
            .n5888(n5888), .n5887(n5887), .n5886(n5886), .\REG.mem_57_7 (\REG.mem_57_7 ), 
            .\REG.mem_6_8 (\REG.mem_6_8 ), .\REG.mem_7_8 (\REG.mem_7_8 ), 
            .\REG.mem_38_15 (\REG.mem_38_15 ), .\REG.mem_39_15 (\REG.mem_39_15 ), 
            .n5885(n5885), .\REG.mem_5_8 (\REG.mem_5_8 ), .\REG.mem_4_8 (\REG.mem_4_8 ), 
            .\REG.mem_14_14 (\REG.mem_14_14 ), .\REG.mem_15_14 (\REG.mem_15_14 ), 
            .n5884(n5884), .\REG.mem_57_5 (\REG.mem_57_5 ), .n5883(n5883), 
            .\REG.mem_57_4 (\REG.mem_57_4 ), .n5882(n5882), .\REG.mem_57_3 (\REG.mem_57_3 ), 
            .n5881(n5881), .\REG.mem_57_2 (\REG.mem_57_2 ), .n5880(n5880), 
            .n5879(n5879), .\REG.mem_57_0 (\REG.mem_57_0 ), .\REG.mem_12_14 (\REG.mem_12_14 ), 
            .\REG.mem_13_14 (\REG.mem_13_14 ), .\REG.mem_37_15 (\REG.mem_37_15 ), 
            .\REG.mem_36_15 (\REG.mem_36_15 ), .n5861(n5861), .wp_sync1_r({wp_sync1_r}), 
            .n5860(n5860), .n5859(n5859), .n5858(n5858), .n5857(n5857), 
            .n5856(n5856), .n5855(n5855), .\REG.mem_55_15 (\REG.mem_55_15 ), 
            .n5854(n5854), .\REG.mem_55_14 (\REG.mem_55_14 ), .n5853(n5853), 
            .\rd_sig_diff0_w[0] (\rd_sig_diff0_w[0] ), .n5852(n5852), .n5851(n5851), 
            .n5850(n5850), .n5849(n5849), .n5848(n5848), .\REG.mem_55_8 (\REG.mem_55_8 ), 
            .n5847(n5847), .n5846(n5846), .\REG.mem_55_6 (\REG.mem_55_6 ), 
            .n5845(n5845), .\REG.mem_55_5 (\REG.mem_55_5 ), .n5844(n5844), 
            .\REG.mem_55_4 (\REG.mem_55_4 ), .n5843(n5843), .\REG.mem_55_3 (\REG.mem_55_3 ), 
            .n5842(n5842), .\REG.mem_55_2 (\REG.mem_55_2 ), .n5841(n5841), 
            .\REG.mem_55_1 (\REG.mem_55_1 ), .n5840(n5840), .\REG.mem_55_0 (\REG.mem_55_0 ), 
            .n5839(n5839), .n5838(n5838), .\REG.mem_40_4 (\REG.mem_40_4 ), 
            .\REG.mem_41_4 (\REG.mem_41_4 ), .\REG.mem_42_4 (\REG.mem_42_4 ), 
            .\REG.mem_43_4 (\REG.mem_43_4 ), .n5836(n5836), .n5835(n5835), 
            .n5834(n5834), .n5833(n5833), .n5832(n5832), .\REG.mem_54_15 (\REG.mem_54_15 ), 
            .n5831(n5831), .\REG.mem_54_14 (\REG.mem_54_14 ), .n5830(n5830), 
            .n5829(n5829), .n5828(n5828), .n5827(n5827), .n5826(n5826), 
            .n5825(n5825), .\REG.mem_54_8 (\REG.mem_54_8 ), .n5824(n5824), 
            .n5823(n5823), .\REG.mem_54_6 (\REG.mem_54_6 ), .n5822(n5822), 
            .\REG.mem_54_5 (\REG.mem_54_5 ), .n5821(n5821), .\REG.mem_54_4 (\REG.mem_54_4 ), 
            .\REG.mem_46_4 (\REG.mem_46_4 ), .\REG.mem_47_4 (\REG.mem_47_4 ), 
            .\REG.mem_44_4 (\REG.mem_44_4 ), .\REG.mem_45_4 (\REG.mem_45_4 ), 
            .n5820(n5820), .\REG.mem_54_3 (\REG.mem_54_3 ), .n5819(n5819), 
            .\REG.mem_54_2 (\REG.mem_54_2 ), .n5818(n5818), .\REG.mem_54_1 (\REG.mem_54_1 ), 
            .n5817(n5817), .\REG.mem_54_0 (\REG.mem_54_0 ), .\REG.mem_25_4 (\REG.mem_25_4 ), 
            .\REG.mem_30_4 (\REG.mem_30_4 ), .\REG.mem_31_4 (\REG.mem_31_4 ), 
            .\REG.mem_8_4 (\REG.mem_8_4 ), .\REG.mem_9_4 (\REG.mem_9_4 ), 
            .\REG.mem_10_4 (\REG.mem_10_4 ), .\REG.mem_11_4 (\REG.mem_11_4 ), 
            .\REG.mem_14_4 (\REG.mem_14_4 ), .\REG.mem_15_4 (\REG.mem_15_4 ), 
            .\REG.mem_12_4 (\REG.mem_12_4 ), .\REG.mem_13_4 (\REG.mem_13_4 ), 
            .n5768(n5768), .\REG.mem_50_15 (\REG.mem_50_15 ), .n5767(n5767), 
            .\REG.mem_50_14 (\REG.mem_50_14 ), .n5766(n5766), .\REG.mem_50_13 (\REG.mem_50_13 ), 
            .n5765(n5765), .n5764(n5764), .n5763(n5763), .n5762(n5762), 
            .n5761(n5761), .\REG.mem_50_8 (\REG.mem_50_8 ), .n5760(n5760), 
            .n5759(n5759), .\REG.mem_50_6 (\REG.mem_50_6 ), .n5758(n5758), 
            .\REG.mem_50_5 (\REG.mem_50_5 ), .n5757(n5757), .\REG.mem_50_4 (\REG.mem_50_4 ), 
            .n10700(n10700), .n5756(n5756), .\REG.mem_50_3 (\REG.mem_50_3 ), 
            .n5755(n5755), .\REG.mem_50_2 (\REG.mem_50_2 ), .n5754(n5754), 
            .n4893(n4893), .\fifo_data_out[14] (\fifo_data_out[14] ), .n4896(n4896), 
            .\fifo_data_out[15] (\fifo_data_out[15] ), .n5750(n5750), .\REG.mem_50_0 (\REG.mem_50_0 ), 
            .\REG.mem_38_5 (\REG.mem_38_5 ), .\REG.mem_39_5 (\REG.mem_39_5 ), 
            .n5733(n5733), .\REG.mem_48_15 (\REG.mem_48_15 ), .n5732(n5732), 
            .\REG.mem_48_14 (\REG.mem_48_14 ), .n5731(n5731), .\REG.mem_48_13 (\REG.mem_48_13 ), 
            .n5730(n5730), .n5729(n5729), .n5728(n5728), .n5727(n5727), 
            .n5726(n5726), .\REG.mem_48_8 (\REG.mem_48_8 ), .n5725(n5725), 
            .n5724(n5724), .\REG.mem_48_6 (\REG.mem_48_6 ), .n10748(n10748), 
            .n5723(n5723), .\REG.mem_48_5 (\REG.mem_48_5 ), .n5722(n5722), 
            .\REG.mem_48_4 (\REG.mem_48_4 ), .n5721(n5721), .\REG.mem_48_3 (\REG.mem_48_3 ), 
            .n5720(n5720), .\REG.mem_48_2 (\REG.mem_48_2 ), .n5719(n5719), 
            .\REG.mem_42_6 (\REG.mem_42_6 ), .\REG.mem_43_6 (\REG.mem_43_6 ), 
            .n5718(n5718), .\REG.mem_48_0 (\REG.mem_48_0 ), .n5717(n5717), 
            .\REG.mem_47_15 (\REG.mem_47_15 ), .\REG.mem_41_6 (\REG.mem_41_6 ), 
            .\REG.mem_40_6 (\REG.mem_40_6 ), .n5716(n5716), .\REG.mem_47_14 (\REG.mem_47_14 ), 
            .n5715(n5715), .\REG.mem_47_13 (\REG.mem_47_13 ), .n5714(n5714), 
            .n5713(n5713), .\REG.mem_47_11 (\REG.mem_47_11 ), .n5712(n5712), 
            .\REG.mem_47_10 (\REG.mem_47_10 ), .n5711(n5711), .n5710(n5710), 
            .n5709(n5709), .\REG.mem_47_7 (\REG.mem_47_7 ), .n5708(n5708), 
            .\REG.mem_47_6 (\REG.mem_47_6 ), .n5707(n5707), .n5706(n5706), 
            .n5705(n5705), .n5704(n5704), .n5703(n5703), .\REG.mem_25_12 (\REG.mem_25_12 ), 
            .\REG.mem_37_5 (\REG.mem_37_5 ), .\REG.mem_36_5 (\REG.mem_36_5 ), 
            .n5702(n5702), .\REG.mem_47_0 (\REG.mem_47_0 ), .n5701(n5701), 
            .\REG.mem_46_15 (\REG.mem_46_15 ), .n5700(n5700), .\REG.mem_46_14 (\REG.mem_46_14 ), 
            .n5699(n5699), .\REG.mem_46_13 (\REG.mem_46_13 ), .n5698(n5698), 
            .n5697(n5697), .\REG.mem_46_11 (\REG.mem_46_11 ), .n5696(n5696), 
            .\REG.mem_46_10 (\REG.mem_46_10 ), .n5695(n5695), .n5694(n5694), 
            .n5693(n5693), .\REG.mem_46_7 (\REG.mem_46_7 ), .n5692(n5692), 
            .\REG.mem_46_6 (\REG.mem_46_6 ), .n5691(n5691), .n5690(n5690), 
            .n5689(n5689), .n5688(n5688), .n5687(n5687), .n5686(n5686), 
            .\REG.mem_46_0 (\REG.mem_46_0 ), .n5685(n5685), .\REG.mem_45_15 (\REG.mem_45_15 ), 
            .n5684(n5684), .\REG.mem_45_14 (\REG.mem_45_14 ), .n5683(n5683), 
            .\REG.mem_45_13 (\REG.mem_45_13 ), .n5682(n5682), .n5681(n5681), 
            .\REG.mem_45_11 (\REG.mem_45_11 ), .n5680(n5680), .\REG.mem_45_10 (\REG.mem_45_10 ), 
            .n5679(n5679), .n5678(n5678), .\REG.mem_6_15 (\REG.mem_6_15 ), 
            .\REG.mem_7_15 (\REG.mem_7_15 ), .\REG.mem_3_1 (\REG.mem_3_1 ), 
            .n5677(n5677), .\REG.mem_45_7 (\REG.mem_45_7 ), .\REG.mem_5_15 (\REG.mem_5_15 ), 
            .\REG.mem_4_15 (\REG.mem_4_15 ), .n5676(n5676), .\REG.mem_45_6 (\REG.mem_45_6 ), 
            .n5675(n5675), .n5674(n5674), .n5673(n5673), .n5672(n5672), 
            .n5671(n5671), .n5670(n5670), .\REG.mem_45_0 (\REG.mem_45_0 ), 
            .n5668(n5668), .\REG.mem_44_15 (\REG.mem_44_15 ), .n5667(n5667), 
            .\REG.mem_44_14 (\REG.mem_44_14 ), .n5665(n5665), .\REG.mem_44_13 (\REG.mem_44_13 ), 
            .n5664(n5664), .n5663(n5663), .\REG.mem_44_11 (\REG.mem_44_11 ), 
            .n5661(n5661), .\REG.mem_44_10 (\REG.mem_44_10 ), .n5660(n5660), 
            .n5659(n5659), .n5658(n5658), .\REG.mem_44_7 (\REG.mem_44_7 ), 
            .n5657(n5657), .\REG.mem_44_6 (\REG.mem_44_6 ), .n5656(n5656), 
            .n5655(n5655), .n5654(n5654), .n5653(n5653), .n5652(n5652), 
            .n5651(n5651), .\REG.mem_44_0 (\REG.mem_44_0 ), .n5650(n5650), 
            .n5649(n5649), .\REG.mem_43_14 (\REG.mem_43_14 ), .n5648(n5648), 
            .n5647(n5647), .n5646(n5646), .\REG.mem_43_11 (\REG.mem_43_11 ), 
            .n5645(n5645), .\REG.mem_43_10 (\REG.mem_43_10 ), .n5644(n5644), 
            .\REG.mem_43_9 (\REG.mem_43_9 ), .\rd_addr_p1_w[0] (\rd_addr_p1_w[0] ), 
            .\REG.mem_18_7 (\REG.mem_18_7 ), .n5643(n5643), .n5642(n5642), 
            .\REG.mem_43_7 (\REG.mem_43_7 ), .n5641(n5641), .n5640(n5640), 
            .\REG.mem_43_5 (\REG.mem_43_5 ), .n5639(n5639), .n5638(n5638), 
            .\REG.mem_43_3 (\REG.mem_43_3 ), .n5637(n5637), .n5636(n5636), 
            .\REG.mem_43_1 (\REG.mem_43_1 ), .n5635(n5635), .n5634(n5634), 
            .n5633(n5633), .\REG.mem_42_14 (\REG.mem_42_14 ), .n5632(n5632), 
            .n5631(n5631), .n5630(n5630), .\REG.mem_42_11 (\REG.mem_42_11 ), 
            .n5629(n5629), .\REG.mem_42_10 (\REG.mem_42_10 ), .n4916(n4916), 
            .\REG.mem_22_11 (\REG.mem_22_11 ), .\REG.mem_23_11 (\REG.mem_23_11 ), 
            .n5628(n5628), .\REG.mem_42_9 (\REG.mem_42_9 ), .n5627(n5627), 
            .n5626(n5626), .\REG.mem_42_7 (\REG.mem_42_7 ), .n5625(n5625), 
            .n5624(n5624), .\REG.mem_42_5 (\REG.mem_42_5 ), .n5623(n5623), 
            .n5622(n5622), .\REG.mem_42_3 (\REG.mem_42_3 ), .n5621(n5621), 
            .n5620(n5620), .\REG.mem_42_1 (\REG.mem_42_1 ), .n5619(n5619), 
            .n5618(n5618), .\REG.mem_41_15 (\REG.mem_41_15 ), .n5617(n5617), 
            .\REG.mem_41_14 (\REG.mem_41_14 ), .n5616(n5616), .n5615(n5615), 
            .n5614(n5614), .\REG.mem_41_11 (\REG.mem_41_11 ), .n5613(n5613), 
            .\REG.mem_41_10 (\REG.mem_41_10 ), .\REG.mem_25_6 (\REG.mem_25_6 ), 
            .n5612(n5612), .\REG.mem_41_9 (\REG.mem_41_9 ), .n5611(n5611), 
            .n5610(n5610), .\REG.mem_41_7 (\REG.mem_41_7 ), .n5609(n5609), 
            .n5608(n5608), .\REG.mem_41_5 (\REG.mem_41_5 ), .n5607(n5607), 
            .n5606(n5606), .\REG.mem_41_3 (\REG.mem_41_3 ), .n5605(n5605), 
            .n5604(n5604), .\REG.mem_41_1 (\REG.mem_41_1 ), .n5603(n5603), 
            .n5602(n5602), .\REG.mem_40_15 (\REG.mem_40_15 ), .n5601(n5601), 
            .\REG.mem_40_14 (\REG.mem_40_14 ), .n5600(n5600), .n5599(n5599), 
            .n5598(n5598), .\REG.mem_40_11 (\REG.mem_40_11 ), .n5597(n5597), 
            .\REG.mem_40_10 (\REG.mem_40_10 ), .n4904(n4904), .n4903(n4903), 
            .n4901(n4901), .n4899(n4899), .n5596(n5596), .\REG.mem_40_9 (\REG.mem_40_9 ), 
            .n5595(n5595), .n5594(n5594), .\REG.mem_40_7 (\REG.mem_40_7 ), 
            .n5593(n5593), .n5592(n5592), .\REG.mem_40_5 (\REG.mem_40_5 ), 
            .n5591(n5591), .n5590(n5590), .\REG.mem_40_3 (\REG.mem_40_3 ), 
            .n5589(n5589), .n5588(n5588), .\REG.mem_40_1 (\REG.mem_40_1 ), 
            .n5587(n5587), .n5586(n5586), .n5585(n5585), .\REG.mem_39_14 (\REG.mem_39_14 ), 
            .n5584(n5584), .n5583(n5583), .\REG.mem_39_12 (\REG.mem_39_12 ), 
            .n5582(n5582), .\REG.mem_39_11 (\REG.mem_39_11 ), .n5581(n5581), 
            .\REG.mem_39_10 (\REG.mem_39_10 ), .n4898(n4898), .DEBUG_5_c(DEBUG_5_c), 
            .\REG.mem_3_4 (\REG.mem_3_4 ), .\REG.mem_6_4 (\REG.mem_6_4 ), 
            .\REG.mem_7_4 (\REG.mem_7_4 ), .n5580(n5580), .\REG.mem_39_9 (\REG.mem_39_9 ), 
            .n5579(n5579), .\REG.mem_39_8 (\REG.mem_39_8 ), .n5578(n5578), 
            .n5577(n5577), .n5576(n5576), .n5575(n5575), .\REG.mem_39_4 (\REG.mem_39_4 ), 
            .n5574(n5574), .\REG.mem_39_3 (\REG.mem_39_3 ), .n5573(n5573), 
            .\REG.mem_39_2 (\REG.mem_39_2 ), .n5572(n5572), .\REG.mem_39_1 (\REG.mem_39_1 ), 
            .n5570(n5570), .n5569(n5569), .n5568(n5568), .\REG.mem_38_14 (\REG.mem_38_14 ), 
            .n5567(n5567), .n5566(n5566), .\REG.mem_38_12 (\REG.mem_38_12 ), 
            .n5565(n5565), .\REG.mem_38_11 (\REG.mem_38_11 ), .n5564(n5564), 
            .\REG.mem_38_10 (\REG.mem_38_10 ), .\REG.mem_5_4 (\REG.mem_5_4 ), 
            .\REG.mem_4_4 (\REG.mem_4_4 ), .n5563(n5563), .\REG.mem_38_9 (\REG.mem_38_9 ), 
            .n5562(n5562), .\REG.mem_38_8 (\REG.mem_38_8 ), .n5561(n5561), 
            .n5560(n5560), .n5559(n5559), .n5558(n5558), .\REG.mem_38_4 (\REG.mem_38_4 ), 
            .n5557(n5557), .\REG.mem_38_3 (\REG.mem_38_3 ), .n5556(n5556), 
            .\REG.mem_38_2 (\REG.mem_38_2 ), .n5555(n5555), .\REG.mem_38_1 (\REG.mem_38_1 ), 
            .n5554(n5554), .n5553(n5553), .n5552(n5552), .\REG.mem_37_14 (\REG.mem_37_14 ), 
            .n5551(n5551), .n5550(n5550), .\REG.mem_37_12 (\REG.mem_37_12 ), 
            .n5549(n5549), .\REG.mem_37_11 (\REG.mem_37_11 ), .\REG.out_raw[15] (\REG.out_raw[15] ), 
            .\REG.out_raw[14] (\REG.out_raw[14] ), .\REG.out_raw[13] (\REG.out_raw[13] ), 
            .\REG.out_raw[12] (\REG.out_raw[12] ), .\REG.out_raw[11] (\REG.out_raw[11] ), 
            .n5548(n5548), .\REG.mem_37_10 (\REG.mem_37_10 ), .n5547(n5547), 
            .\REG.mem_37_9 (\REG.mem_37_9 ), .n5546(n5546), .\REG.mem_37_8 (\REG.mem_37_8 ), 
            .n5545(n5545), .n5544(n5544), .n5543(n5543), .n5542(n5542), 
            .\REG.mem_37_4 (\REG.mem_37_4 ), .n5541(n5541), .\REG.mem_37_3 (\REG.mem_37_3 ), 
            .n5540(n5540), .\REG.mem_37_2 (\REG.mem_37_2 ), .n5539(n5539), 
            .\REG.mem_37_1 (\REG.mem_37_1 ), .n5538(n5538), .\REG.out_raw[10] (\REG.out_raw[10] ), 
            .\REG.out_raw[9] (\REG.out_raw[9] ), .\REG.out_raw[8] (\REG.out_raw[8] ), 
            .\REG.out_raw[7] (\REG.out_raw[7] ), .\REG.out_raw[6] (\REG.out_raw[6] ), 
            .\REG.out_raw[5] (\REG.out_raw[5] ), .\REG.out_raw[4] (\REG.out_raw[4] ), 
            .\REG.out_raw[3] (\REG.out_raw[3] ), .\REG.out_raw[2] (\REG.out_raw[2] ), 
            .\REG.out_raw[1] (\REG.out_raw[1] ), .n5524(n5524), .n5523(n5523), 
            .\REG.mem_36_14 (\REG.mem_36_14 ), .n5522(n5522), .n5521(n5521), 
            .\REG.mem_36_12 (\REG.mem_36_12 ), .n5520(n5520), .\REG.mem_36_11 (\REG.mem_36_11 ), 
            .n5519(n5519), .\REG.mem_36_10 (\REG.mem_36_10 ), .n5518(n5518), 
            .\REG.mem_36_9 (\REG.mem_36_9 ), .n5517(n5517), .\REG.mem_36_8 (\REG.mem_36_8 ), 
            .n5516(n5516), .\rd_sig_diff0_w[2] (\rd_sig_diff0_w[2] ), .n5515(n5515), 
            .n5514(n5514), .n5513(n5513), .\REG.mem_36_4 (\REG.mem_36_4 ), 
            .n5512(n5512), .\REG.mem_36_3 (\REG.mem_36_3 ), .n5511(n5511), 
            .\REG.mem_36_2 (\REG.mem_36_2 ), .n5510(n5510), .\REG.mem_36_1 (\REG.mem_36_1 ), 
            .n5509(n5509), .n5505(n5505), .n5504(n5504), .\REG.mem_35_14 (\REG.mem_35_14 ), 
            .n5503(n5503), .n5502(n5502), .\REG.mem_35_12 (\REG.mem_35_12 ), 
            .n5501(n5501), .\REG.mem_35_11 (\REG.mem_35_11 ), .n5500(n5500), 
            .\REG.mem_35_10 (\REG.mem_35_10 ), .\rd_sig_diff0_w[1] (\rd_sig_diff0_w[1] ), 
            .n5499(n5499), .n5498(n5498), .\REG.mem_35_8 (\REG.mem_35_8 ), 
            .n5497(n5497), .n5496(n5496), .n5495(n5495), .\REG.mem_35_5 (\REG.mem_35_5 ), 
            .n5494(n5494), .\REG.mem_35_4 (\REG.mem_35_4 ), .n5493(n5493), 
            .\REG.mem_35_3 (\REG.mem_35_3 ), .n5492(n5492), .\REG.mem_35_2 (\REG.mem_35_2 ), 
            .n5491(n5491), .\REG.mem_35_1 (\REG.mem_35_1 ), .n5490(n5490), 
            .\REG.mem_25_11 (\REG.mem_25_11 ), .\REG.mem_10_13 (\REG.mem_10_13 ), 
            .\REG.mem_11_13 (\REG.mem_11_13 ), .\REG.mem_9_13 (\REG.mem_9_13 ), 
            .\REG.mem_8_13 (\REG.mem_8_13 ), .n5440(n5440), .n5439(n5439), 
            .\REG.mem_31_14 (\REG.mem_31_14 ), .n5438(n5438), .n5437(n5437), 
            .\REG.mem_31_12 (\REG.mem_31_12 ), .n5436(n5436), .\REG.mem_31_11 (\REG.mem_31_11 ), 
            .n5435(n5435), .\REG.mem_31_10 (\REG.mem_31_10 ), .n5434(n5434), 
            .n5433(n5433), .\REG.mem_31_8 (\REG.mem_31_8 ), .n5432(n5432), 
            .\REG.mem_31_7 (\REG.mem_31_7 ), .n5431(n5431), .\REG.mem_31_6 (\REG.mem_31_6 ), 
            .n5430(n5430), .n5429(n5429), .n5428(n5428), .\REG.mem_31_3 (\REG.mem_31_3 ), 
            .n5427(n5427), .n5426(n5426), .\REG.mem_31_1 (\REG.mem_31_1 ), 
            .n5425(n5425), .n5424(n5424), .n5423(n5423), .\REG.mem_30_14 (\REG.mem_30_14 ), 
            .n5422(n5422), .n5421(n5421), .\REG.mem_30_12 (\REG.mem_30_12 ), 
            .n5420(n5420), .\REG.mem_30_11 (\REG.mem_30_11 ), .DEBUG_1_c_c(DEBUG_1_c_c), 
            .write_to_dc32_fifo_latched_N_425(write_to_dc32_fifo_latched_N_425), 
            .\REG.mem_18_6 (\REG.mem_18_6 ), .n5419(n5419), .\REG.mem_30_10 (\REG.mem_30_10 ), 
            .n5418(n5418), .n5417(n5417), .\REG.mem_30_8 (\REG.mem_30_8 ), 
            .n5416(n5416), .\REG.mem_30_7 (\REG.mem_30_7 ), .n5415(n5415), 
            .\REG.mem_30_6 (\REG.mem_30_6 ), .n5414(n5414), .n5413(n5413), 
            .n5412(n5412), .\REG.mem_30_3 (\REG.mem_30_3 ), .n5411(n5411), 
            .n5410(n5410), .\REG.mem_30_1 (\REG.mem_30_1 ), .n5409(n5409), 
            .\REG.mem_16_6 (\REG.mem_16_6 ), .\wr_addr_nxt_c[1] (\wr_addr_nxt_c[1] ), 
            .\REG.mem_10_9 (\REG.mem_10_9 ), .\REG.mem_11_9 (\REG.mem_11_9 ), 
            .\REG.mem_9_9 (\REG.mem_9_9 ), .\REG.mem_8_9 (\REG.mem_8_9 ), 
            .\REG.mem_14_13 (\REG.mem_14_13 ), .\REG.mem_15_13 (\REG.mem_15_13 ), 
            .\REG.mem_13_13 (\REG.mem_13_13 ), .\REG.mem_12_13 (\REG.mem_12_13 ), 
            .n56(n56), .\REG.mem_14_9 (\REG.mem_14_9 ), .\REG.mem_15_9 (\REG.mem_15_9 ), 
            .\REG.mem_10_15 (\REG.mem_10_15 ), .\REG.mem_11_15 (\REG.mem_11_15 ), 
            .\REG.mem_9_15 (\REG.mem_9_15 ), .\REG.mem_8_15 (\REG.mem_8_15 ), 
            .\REG.mem_10_7 (\REG.mem_10_7 ), .\REG.mem_11_7 (\REG.mem_11_7 ), 
            .\REG.mem_13_9 (\REG.mem_13_9 ), .\REG.mem_12_9 (\REG.mem_12_9 ), 
            .n5344(n5344), .n5343(n5343), .\REG.mem_25_14 (\REG.mem_25_14 ), 
            .n5342(n5342), .n5341(n5341), .n5340(n5340), .n5339(n5339), 
            .\REG.mem_25_10 (\REG.mem_25_10 ), .n5338(n5338), .n5337(n5337), 
            .\REG.mem_25_8 (\REG.mem_25_8 ), .n5336(n5336), .\REG.mem_25_7 (\REG.mem_25_7 ), 
            .\REG.mem_18_13 (\REG.mem_18_13 ), .\REG.mem_9_7 (\REG.mem_9_7 ), 
            .\REG.mem_8_7 (\REG.mem_8_7 ), .\REG.mem_16_13 (\REG.mem_16_13 ), 
            .n5335(n5335), .n5334(n5334), .n5333(n5333), .n5332(n5332), 
            .\REG.mem_25_3 (\REG.mem_25_3 ), .n5331(n5331), .n5330(n5330), 
            .n5329(n5329), .\REG.mem_25_0 (\REG.mem_25_0 ), .n52(n52), 
            .n20(n20), .n5306(n5306), .\REG.mem_23_15 (\REG.mem_23_15 ), 
            .n5305(n5305), .\REG.mem_23_14 (\REG.mem_23_14 ), .n5304(n5304), 
            .\REG.mem_23_13 (\REG.mem_23_13 ), .n5303(n5303), .n5302(n5302), 
            .n5301(n5301), .\REG.mem_23_10 (\REG.mem_23_10 ), .n5300(n5300), 
            .\REG.mem_23_9 (\REG.mem_23_9 ), .n5299(n5299), .n5298(n5298), 
            .n5297(n5297), .\REG.mem_23_6 (\REG.mem_23_6 ), .n5296(n5296), 
            .\REG.mem_23_5 (\REG.mem_23_5 ), .n5295(n5295), .\REG.mem_23_4 (\REG.mem_23_4 ), 
            .n5294(n5294), .\REG.mem_23_3 (\REG.mem_23_3 ), .n5293(n5293), 
            .\REG.mem_23_2 (\REG.mem_23_2 ), .n5292(n5292), .\REG.mem_23_1 (\REG.mem_23_1 ), 
            .n5291(n5291), .\REG.mem_23_0 (\REG.mem_23_0 ), .n5290(n5290), 
            .\REG.mem_22_15 (\REG.mem_22_15 ), .n5289(n5289), .\REG.mem_22_14 (\REG.mem_22_14 ), 
            .n5288(n5288), .\REG.mem_22_13 (\REG.mem_22_13 ), .n5287(n5287), 
            .n5286(n5286), .n5285(n5285), .\REG.mem_22_10 (\REG.mem_22_10 ), 
            .\rd_grey_sync_r[5] (\rd_grey_sync_r[5] ), .\rd_grey_sync_r[4] (\rd_grey_sync_r[4] ), 
            .\rd_grey_sync_r[3] (\rd_grey_sync_r[3] ), .\rd_grey_sync_r[2] (\rd_grey_sync_r[2] ), 
            .\rd_grey_sync_r[1] (\rd_grey_sync_r[1] ), .n5284(n5284), .\REG.mem_22_9 (\REG.mem_22_9 ), 
            .n5283(n5283), .n5282(n5282), .n5281(n5281), .\REG.mem_22_6 (\REG.mem_22_6 ), 
            .n5280(n5280), .\REG.mem_22_5 (\REG.mem_22_5 ), .n5279(n5279), 
            .\REG.mem_22_4 (\REG.mem_22_4 ), .n5278(n5278), .\REG.mem_22_3 (\REG.mem_22_3 ), 
            .n5277(n5277), .\REG.mem_22_2 (\REG.mem_22_2 ), .n5276(n5276), 
            .\REG.mem_22_1 (\REG.mem_22_1 ), .n5275(n5275), .\REG.mem_22_0 (\REG.mem_22_0 ), 
            .\REG.mem_14_3 (\REG.mem_14_3 ), .\REG.mem_15_3 (\REG.mem_15_3 ), 
            .\REG.mem_13_3 (\REG.mem_13_3 ), .\REG.mem_12_3 (\REG.mem_12_3 ), 
            .\REG.mem_10_8 (\REG.mem_10_8 ), .\REG.mem_11_8 (\REG.mem_11_8 ), 
            .\REG.mem_9_8 (\REG.mem_9_8 ), .\REG.mem_8_8 (\REG.mem_8_8 ), 
            .get_next_word(get_next_word), .\REG.mem_16_2 (\REG.mem_16_2 ), 
            .\REG.mem_18_2 (\REG.mem_18_2 ), .\REG.mem_18_3 (\REG.mem_18_3 ), 
            .n5226(n5226), .\REG.mem_18_15 (\REG.mem_18_15 ), .n5225(n5225), 
            .\REG.mem_18_14 (\REG.mem_18_14 ), .n5224(n5224), .n5223(n5223), 
            .n5222(n5222), .n5221(n5221), .\REG.mem_18_10 (\REG.mem_18_10 ), 
            .n5220(n5220), .\REG.mem_18_9 (\REG.mem_18_9 ), .rd_fifo_en_w(rd_fifo_en_w), 
            .\REG.mem_16_3 (\REG.mem_16_3 ), .\REG.mem_16_15 (\REG.mem_16_15 ), 
            .n5219(n5219), .n5218(n5218), .n5217(n5217), .n5216(n5216), 
            .n5215(n5215), .\REG.mem_18_4 (\REG.mem_18_4 ), .n5214(n5214), 
            .n5213(n5213), .n5212(n5212), .\REG.mem_18_1 (\REG.mem_18_1 ), 
            .n5211(n5211), .\REG.mem_18_0 (\REG.mem_18_0 ), .n5190(n5190), 
            .n5188(n5188), .\REG.mem_16_14 (\REG.mem_16_14 ), .n5187(n5187), 
            .n5186(n5186), .n5185(n5185), .n5184(n5184), .\REG.mem_16_10 (\REG.mem_16_10 ), 
            .\REG.mem_3_2 (\REG.mem_3_2 ), .\REG.mem_3_0 (\REG.mem_3_0 ), 
            .n5183(n5183), .\REG.mem_16_9 (\REG.mem_16_9 ), .n5182(n5182), 
            .n5181(n5181), .n5180(n5180), .n5179(n5179), .n5178(n5178), 
            .\REG.mem_16_4 (\REG.mem_16_4 ), .n5177(n5177), .n5176(n5176), 
            .\REG.mem_6_0 (\REG.mem_6_0 ), .\REG.mem_7_0 (\REG.mem_7_0 ), 
            .n5175(n5175), .\REG.mem_16_1 (\REG.mem_16_1 ), .n5174(n5174), 
            .\REG.mem_16_0 (\REG.mem_16_0 ), .n5171(n5171), .\REG.mem_15_15 (\REG.mem_15_15 ), 
            .n5170(n5170), .n5169(n5169), .n5168(n5168), .n5167(n5167), 
            .n5166(n5166), .\REG.mem_15_10 (\REG.mem_15_10 ), .n5165(n5165), 
            .n5164(n5164), .n5163(n5163), .n5162(n5162), .\REG.mem_15_6 (\REG.mem_15_6 ), 
            .\REG.mem_5_0 (\REG.mem_5_0 ), .\REG.mem_4_0 (\REG.mem_4_0 ), 
            .n5161(n5161), .n5160(n5160), .n5159(n5159), .n5158(n5158), 
            .n5157(n5157), .\REG.mem_15_1 (\REG.mem_15_1 ), .n5156(n5156), 
            .\REG.mem_15_0 (\REG.mem_15_0 ), .n5155(n5155), .\REG.mem_14_15 (\REG.mem_14_15 ), 
            .n5154(n5154), .n5153(n5153), .n5152(n5152), .n5151(n5151), 
            .n5150(n5150), .\REG.mem_14_10 (\REG.mem_14_10 ), .n5149(n5149), 
            .n5148(n5148), .n5147(n5147), .n5146(n5146), .\REG.mem_14_6 (\REG.mem_14_6 ), 
            .n5145(n5145), .n5144(n5144), .n5143(n5143), .n5142(n5142), 
            .n5141(n5141), .\REG.mem_14_1 (\REG.mem_14_1 ), .n5140(n5140), 
            .\REG.mem_14_0 (\REG.mem_14_0 ), .n5139(n5139), .\REG.mem_13_15 (\REG.mem_13_15 ), 
            .n5138(n5138), .n5137(n5137), .n5136(n5136), .n5135(n5135), 
            .n5134(n5134), .\REG.mem_13_10 (\REG.mem_13_10 ), .n5133(n5133), 
            .n5132(n5132), .n5131(n5131), .n47(n47), .n15(n15), .n50(n50), 
            .n5130(n5130), .\REG.mem_13_6 (\REG.mem_13_6 ), .n18(n18), 
            .n5129(n5129), .n5128(n5128), .n5127(n5127), .n5126(n5126), 
            .n5125(n5125), .\REG.mem_13_1 (\REG.mem_13_1 ), .n5124(n5124), 
            .\REG.mem_13_0 (\REG.mem_13_0 ), .n5123(n5123), .\REG.mem_12_15 (\REG.mem_12_15 ), 
            .n5122(n5122), .n5121(n5121), .n5120(n5120), .n5119(n5119), 
            .n5118(n5118), .\REG.mem_12_10 (\REG.mem_12_10 ), .n5117(n5117), 
            .n5116(n5116), .\REG.mem_3_12 (\REG.mem_3_12 ), .\REG.mem_3_14 (\REG.mem_3_14 ), 
            .n5115(n5115), .n5114(n5114), .\REG.mem_12_6 (\REG.mem_12_6 ), 
            .n5113(n5113), .n5112(n5112), .n53(n53), .n21(n21), .\REG.mem_10_0 (\REG.mem_10_0 ), 
            .\REG.mem_11_0 (\REG.mem_11_0 ), .\REG.mem_9_0 (\REG.mem_9_0 ), 
            .\REG.mem_8_0 (\REG.mem_8_0 ), .n5111(n5111), .n5110(n5110), 
            .n5109(n5109), .\REG.mem_12_1 (\REG.mem_12_1 ), .n5108(n5108), 
            .\REG.mem_12_0 (\REG.mem_12_0 ), .n51(n51), .n19(n19), .n5107(n5107), 
            .n54(n54), .n22(n22), .n5106(n5106), .n5105(n5105), .n5104(n5104), 
            .\REG.mem_11_12 (\REG.mem_11_12 ), .n5103(n5103), .n5102(n5102), 
            .\REG.mem_11_10 (\REG.mem_11_10 ), .n5101(n5101), .n5100(n5100), 
            .n5099(n5099), .n5098(n5098), .n5097(n5097), .\REG.mem_11_5 (\REG.mem_11_5 ), 
            .\rd_addr_nxt_c_6__N_498[5] (\rd_addr_nxt_c_6__N_498[5] ), .n5096(n5096), 
            .n5095(n5095), .n5094(n5094), .n5093(n5093), .\REG.mem_11_1 (\REG.mem_11_1 ), 
            .n5092(n5092), .n5091(n5091), .n5090(n5090), .n5089(n5089), 
            .n5088(n5088), .\REG.mem_10_12 (\REG.mem_10_12 ), .n5087(n5087), 
            .n5086(n5086), .\REG.mem_10_10 (\REG.mem_10_10 ), .n5085(n5085), 
            .n5084(n5084), .n5083(n5083), .n5082(n5082), .n5081(n5081), 
            .\REG.mem_10_5 (\REG.mem_10_5 ), .n5080(n5080), .\rd_addr_nxt_c_6__N_498[3] (\rd_addr_nxt_c_6__N_498[3] ), 
            .n5079(n5079), .\rd_addr_nxt_c_6__N_498[2] (\rd_addr_nxt_c_6__N_498[2] ), 
            .n49(n49), .n17(n17), .\REG.mem_6_14 (\REG.mem_6_14 ), .\REG.mem_7_14 (\REG.mem_7_14 ), 
            .\REG.mem_4_14 (\REG.mem_4_14 ), .\REG.mem_5_14 (\REG.mem_5_14 ), 
            .n24(n24), .n5078(n5078), .\REG.mem_3_6 (\REG.mem_3_6 ), .n5077(n5077), 
            .\REG.mem_10_1 (\REG.mem_10_1 ), .n5076(n5076), .n5075(n5075), 
            .\REG.mem_3_9 (\REG.mem_3_9 ), .n5074(n5074), .n5073(n5073), 
            .n55(n55), .n23(n23), .n40(n40), .n8(n8), .n5072(n5072), 
            .\REG.mem_9_12 (\REG.mem_9_12 ), .n34(n34), .n5071(n5071), 
            .n5070(n5070), .\REG.mem_9_10 (\REG.mem_9_10 ), .n5069(n5069), 
            .n2(n2), .n5068(n5068), .n5067(n5067), .n5066(n5066), .n5065(n5065), 
            .\REG.mem_9_5 (\REG.mem_9_5 ), .n5064(n5064), .n5063(n5063), 
            .n5062(n5062), .n5061(n5061), .\REG.mem_9_1 (\REG.mem_9_1 ), 
            .n5060(n5060), .n5059(n5059), .n5058(n5058), .n5057(n5057), 
            .n5056(n5056), .\REG.mem_8_12 (\REG.mem_8_12 ), .n5055(n5055), 
            .n5054(n5054), .\REG.mem_8_10 (\REG.mem_8_10 ), .n5053(n5053), 
            .n5052(n5052), .n5051(n5051), .n5050(n5050), .n5049(n5049), 
            .\REG.mem_8_5 (\REG.mem_8_5 ), .n5048(n5048), .n5047(n5047), 
            .n5046(n5046), .n5045(n5045), .\REG.mem_8_1 (\REG.mem_8_1 ), 
            .n5044(n5044), .n5043(n5043), .n5042(n5042), .n5041(n5041), 
            .\REG.mem_7_13 (\REG.mem_7_13 ), .n5040(n5040), .\REG.mem_7_12 (\REG.mem_7_12 ), 
            .n5039(n5039), .n5038(n5038), .\REG.mem_7_10 (\REG.mem_7_10 ), 
            .n5037(n5037), .n5036(n5036), .n5035(n5035), .\REG.mem_7_7 (\REG.mem_7_7 ), 
            .n5034(n5034), .\REG.mem_7_6 (\REG.mem_7_6 ), .n5033(n5033), 
            .n5032(n5032), .n5031(n5031), .n5030(n5030), .n5029(n5029), 
            .n5028(n5028), .n5027(n5027), .n5026(n5026), .n5025(n5025), 
            .\REG.mem_6_13 (\REG.mem_6_13 ), .n5024(n5024), .\REG.mem_6_12 (\REG.mem_6_12 ), 
            .n5023(n5023), .n5022(n5022), .\REG.mem_6_10 (\REG.mem_6_10 ), 
            .n5021(n5021), .n5020(n5020), .n5019(n5019), .\REG.mem_6_7 (\REG.mem_6_7 ), 
            .n5018(n5018), .\REG.mem_6_6 (\REG.mem_6_6 ), .n5017(n5017), 
            .n5016(n5016), .n5015(n5015), .n5014(n5014), .n5013(n5013), 
            .n5012(n5012), .n5011(n5011), .n5010(n5010), .n5009(n5009), 
            .\REG.mem_5_13 (\REG.mem_5_13 ), .n5008(n5008), .\REG.mem_5_12 (\REG.mem_5_12 ), 
            .n5007(n5007), .n5006(n5006), .\REG.mem_5_10 (\REG.mem_5_10 ), 
            .n5005(n5005), .n5004(n5004), .n5003(n5003), .\REG.mem_5_7 (\REG.mem_5_7 ), 
            .n5002(n5002), .\REG.mem_5_6 (\REG.mem_5_6 ), .n5001(n5001), 
            .n5000(n5000), .n4999(n4999), .n4998(n4998), .n4997(n4997), 
            .n4996(n4996), .n4995(n4995), .n4994(n4994), .n4993(n4993), 
            .\REG.mem_4_13 (\REG.mem_4_13 ), .n4992(n4992), .\REG.mem_4_12 (\REG.mem_4_12 ), 
            .n4991(n4991), .n4990(n4990), .\REG.mem_4_10 (\REG.mem_4_10 ), 
            .n4989(n4989), .n4988(n4988), .n4987(n4987), .\REG.mem_4_7 (\REG.mem_4_7 ), 
            .n4986(n4986), .\REG.mem_4_6 (\REG.mem_4_6 ), .n4985(n4985), 
            .n4984(n4984), .n4983(n4983), .n4982(n4982), .n4981(n4981), 
            .n4980(n4980), .n4979(n4979), .n4978(n4978), .n4977(n4977), 
            .\REG.mem_3_13 (\REG.mem_3_13 ), .n4976(n4976), .n4975(n4975), 
            .n4974(n4974), .\REG.mem_3_10 (\REG.mem_3_10 ), .n4973(n4973), 
            .n4972(n4972), .\REG.mem_3_8 (\REG.mem_3_8 ), .n4971(n4971), 
            .\REG.mem_3_7 (\REG.mem_3_7 ), .n4970(n4970), .n4969(n4969), 
            .FT_OE_N_420(FT_OE_N_420), .n57(n57), .n25(n25), .n42(n42), 
            .n10(n10), .n58(n58), .n26(n26), .n43(n43), .n35(n35), 
            .n11(n11), .n3(n3), .n4968(n4968), .n4967(n4967), .n4966(n4966), 
            .n4965(n4965), .n4964(n4964), .n60(n60), .n28(n28), .n59(n59), 
            .n27(n27), .n61(n61), .n29(n29), .n4672(n4672), .n4671(n4671), 
            .n4670(n4670), .n4669(n4669), .n4668(n4668), .n4667(n4667), 
            .n4666(n4666), .n4665(n4665), .n4664(n4664), .n4663(n4663), 
            .n4662(n4662), .n4661(n4661), .n4660(n4660), .n4659(n4659), 
            .n4658(n4658)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_dc_32_lut_gen.v(53[33] 72[34])
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1
//

module fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 (dc32_fifo_almost_full, 
            FIFO_CLK_c, reset_per_frame, \REG.mem_16_7 , \rd_addr_r[0] , 
            \REG.mem_6_2 , \REG.mem_7_2 , \dc32_fifo_data_in[7] , \REG.mem_46_9 , 
            \REG.mem_47_9 , \REG.mem_25_5 , GND_net, t_rd_fifo_en_w, 
            \REG.out_raw[0] , SLM_CLK_c, \REG.mem_45_9 , \REG.mem_44_9 , 
            \REG.mem_57_15 , \REG.mem_62_15 , \REG.mem_63_15 , \REG.mem_6_1 , 
            \REG.mem_7_1 , \REG.mem_5_1 , \REG.mem_4_1 , \REG.mem_57_1 , 
            \REG.mem_25_9 , \dc32_fifo_data_in[6] , \dc32_fifo_data_in[15] , 
            \REG.mem_46_3 , \REG.mem_47_3 , \REG.mem_45_3 , \REG.mem_44_3 , 
            \REG.mem_54_13 , \REG.mem_55_13 , \REG.mem_50_11 , \REG.mem_48_11 , 
            \dc32_fifo_data_in[5] , \REG.mem_42_12 , \REG.mem_43_12 , 
            \REG.mem_41_12 , \REG.mem_40_12 , \dc32_fifo_data_in[4] , 
            \dc32_fifo_data_in[3] , \dc32_fifo_data_in[2] , \rd_grey_sync_r[0] , 
            \REG.mem_57_6 , DEBUG_3_c, wr_grey_sync_r, \dc32_fifo_data_in[1] , 
            \REG.mem_54_11 , \REG.mem_55_11 , \aempty_flag_impl.ae_flag_nxt_w , 
            dc32_fifo_almost_empty, \REG.mem_14_12 , \REG.mem_15_12 , 
            \REG.mem_30_0 , \REG.mem_31_0 , \REG.mem_13_12 , \REG.mem_12_12 , 
            \REG.mem_3_5 , \REG.mem_6_5 , \REG.mem_7_5 , \REG.mem_4_5 , 
            \REG.mem_5_5 , \REG.mem_57_11 , n62, \REG.mem_62_13 , \REG.mem_63_13 , 
            \REG.mem_46_1 , \REG.mem_47_1 , \REG.mem_45_1 , \REG.mem_44_1 , 
            \dc32_fifo_data_in[0] , \REG.mem_3_11 , \REG.mem_6_11 , \REG.mem_7_11 , 
            n30, \REG.mem_5_2 , \REG.mem_4_2 , \REG.mem_18_5 , \REG.mem_62_1 , 
            \REG.mem_63_1 , \REG.mem_38_13 , \REG.mem_39_13 , \REG.mem_5_11 , 
            \REG.mem_4_11 , \dc32_fifo_data_in[8] , \REG.mem_14_5 , \REG.mem_15_5 , 
            \REG.mem_13_5 , \REG.mem_12_5 , \REG.mem_30_9 , \REG.mem_31_9 , 
            \wr_addr_nxt_c[5] , \REG.mem_46_12 , \REG.mem_47_12 , \REG.mem_45_12 , 
            \REG.mem_44_12 , \REG.mem_62_11 , \REG.mem_63_11 , \REG.mem_57_8 , 
            \REG.mem_62_6 , \REG.mem_63_6 , \REG.mem_62_8 , \REG.mem_63_8 , 
            \REG.mem_35_0 , \REG.mem_25_15 , \REG.mem_35_7 , \REG.mem_35_9 , 
            \REG.mem_18_12 , \REG.mem_16_12 , \REG.mem_14_8 , \REG.mem_15_8 , 
            \REG.mem_13_8 , \REG.mem_12_8 , \REG.mem_14_2 , \REG.mem_15_2 , 
            \REG.mem_13_2 , \REG.mem_12_2 , \REG.mem_38_7 , \REG.mem_39_7 , 
            \REG.mem_36_7 , \REG.mem_37_7 , \REG.mem_50_12 , \REG.mem_48_12 , 
            \REG.mem_62_9 , \REG.mem_63_9 , \REG.mem_6_9 , \REG.mem_7_9 , 
            \REG.mem_35_6 , \REG.mem_5_9 , \REG.mem_4_9 , \REG.mem_37_13 , 
            \REG.mem_36_13 , \REG.mem_42_8 , \REG.mem_43_8 , \REG.mem_41_8 , 
            \REG.mem_40_8 , \REG.mem_22_7 , \REG.mem_23_7 , \REG.mem_10_11 , 
            \REG.mem_11_11 , \REG.mem_9_11 , \REG.mem_8_11 , \REG.mem_3_15 , 
            \REG.mem_46_8 , \REG.mem_47_8 , \REG.mem_45_8 , \REG.mem_44_8 , 
            \REG.mem_46_5 , \REG.mem_47_5 , \REG.mem_45_5 , \REG.mem_44_5 , 
            \REG.mem_10_2 , \REG.mem_11_2 , \REG.mem_54_9 , \REG.mem_55_9 , 
            \REG.mem_57_9 , \REG.mem_57_14 , \REG.mem_30_15 , \REG.mem_31_15 , 
            \REG.mem_42_15 , \REG.mem_43_15 , \REG.mem_16_5 , \REG.mem_9_2 , 
            \REG.mem_8_2 , \REG.mem_62_12 , \REG.mem_63_12 , \wr_addr_nxt_c[3] , 
            \REG.mem_18_8 , \REG.mem_16_8 , \REG.mem_22_12 , \REG.mem_23_12 , 
            \REG.mem_25_2 , \REG.mem_30_2 , \REG.mem_31_2 , \dc32_fifo_data_in[14] , 
            \REG.mem_48_10 , \REG.mem_50_10 , \dc32_fifo_data_in[13] , 
            \REG.mem_54_10 , \REG.mem_55_10 , \REG.mem_14_11 , \REG.mem_15_11 , 
            \dc32_fifo_data_in[12] , \REG.mem_54_12 , \REG.mem_55_12 , 
            \REG.mem_13_11 , \REG.mem_12_11 , \REG.mem_35_15 , \REG.mem_38_6 , 
            \REG.mem_39_6 , \dc32_fifo_data_in[11] , \REG.mem_37_6 , \REG.mem_36_6 , 
            \REG.mem_57_13 , \dc32_fifo_data_in[10] , \dc32_fifo_data_in[9] , 
            \REG.mem_30_13 , \REG.mem_31_13 , \REG.mem_30_5 , \REG.mem_31_5 , 
            \REG.mem_48_7 , \REG.mem_50_7 , \REG.mem_54_7 , \REG.mem_55_7 , 
            n6106, VCC_net, \fifo_data_out[2] , n6103, \fifo_data_out[1] , 
            \REG.mem_35_13 , \REG.mem_3_3 , \rd_addr_r[6] , n4827, \fifo_data_out[3] , 
            \REG.mem_50_1 , n4830, \fifo_data_out[4] , n4841, \fifo_data_out[5] , 
            n4844, \fifo_data_out[6] , n4848, \fifo_data_out[7] , n4851, 
            \fifo_data_out[8] , n4854, \fifo_data_out[9] , n4858, \fifo_data_out[10] , 
            n4864, \fifo_data_out[11] , \REG.mem_62_14 , \REG.mem_63_14 , 
            \REG.mem_48_1 , \REG.mem_18_11 , \REG.mem_16_11 , \REG.mem_6_3 , 
            \REG.mem_7_3 , \REG.mem_5_3 , \REG.mem_4_3 , \REG.mem_42_2 , 
            \REG.mem_43_2 , \REG.mem_41_2 , \REG.mem_40_2 , n6070, \fifo_data_out[0] , 
            \REG.mem_46_2 , \REG.mem_47_2 , \REG.mem_45_2 , \REG.mem_44_2 , 
            \REG.mem_14_7 , \REG.mem_15_7 , n4872, \fifo_data_out[12] , 
            n4875, \fifo_data_out[13] , \REG.mem_13_7 , \REG.mem_12_7 , 
            n6034, \REG.mem_25_13 , n6032, \REG.mem_10_3 , \REG.mem_11_3 , 
            \REG.mem_9_3 , \REG.mem_8_3 , \REG.mem_50_9 , n6013, n6012, 
            n6011, n6010, n6009, n6008, n6007, \REG.mem_63_10 , 
            n6006, n6005, n6004, \REG.mem_63_7 , n6003, n6002, \REG.mem_63_5 , 
            \REG.mem_48_9 , \REG.mem_42_13 , \REG.mem_43_13 , \REG.mem_38_0 , 
            \REG.mem_39_0 , n6001, \REG.mem_63_4 , n6000, \REG.mem_63_3 , 
            n5999, \REG.mem_63_2 , n5998, n5997, \REG.mem_63_0 , n5996, 
            n5995, n5994, n5993, n5992, n5991, \REG.mem_62_10 , 
            n5990, n5989, n5988, \REG.mem_62_7 , n5987, n5986, \REG.mem_62_5 , 
            n5985, \REG.mem_62_4 , \REG.mem_41_13 , \REG.mem_40_13 , 
            \REG.mem_37_0 , \REG.mem_36_0 , \REG.mem_10_6 , \REG.mem_11_6 , 
            n5984, \REG.mem_62_3 , n5983, \REG.mem_62_2 , n5982, n5981, 
            \REG.mem_62_0 , \REG.mem_9_6 , \REG.mem_8_6 , \REG.mem_42_0 , 
            \REG.mem_43_0 , \REG.mem_22_8 , \REG.mem_23_8 , n5946, rp_sync1_r, 
            n5945, n5944, n5943, n5942, n5941, n5940, n5939, n5938, 
            n5921, n5920, n5919, \REG.mem_41_0 , \REG.mem_40_0 , n5917, 
            n5916, n5914, \REG.mem_8_14 , \REG.mem_9_14 , \REG.mem_25_1 , 
            \REG.mem_10_14 , \REG.mem_11_14 , n5894, n5893, n5892, 
            n5891, \REG.mem_57_12 , n5890, n5889, \REG.mem_57_10 , 
            n5888, n5887, n5886, \REG.mem_57_7 , \REG.mem_6_8 , \REG.mem_7_8 , 
            \REG.mem_38_15 , \REG.mem_39_15 , n5885, \REG.mem_5_8 , 
            \REG.mem_4_8 , \REG.mem_14_14 , \REG.mem_15_14 , n5884, 
            \REG.mem_57_5 , n5883, \REG.mem_57_4 , n5882, \REG.mem_57_3 , 
            n5881, \REG.mem_57_2 , n5880, n5879, \REG.mem_57_0 , \REG.mem_12_14 , 
            \REG.mem_13_14 , \REG.mem_37_15 , \REG.mem_36_15 , n5861, 
            wp_sync1_r, n5860, n5859, n5858, n5857, n5856, n5855, 
            \REG.mem_55_15 , n5854, \REG.mem_55_14 , n5853, \rd_sig_diff0_w[0] , 
            n5852, n5851, n5850, n5849, n5848, \REG.mem_55_8 , n5847, 
            n5846, \REG.mem_55_6 , n5845, \REG.mem_55_5 , n5844, \REG.mem_55_4 , 
            n5843, \REG.mem_55_3 , n5842, \REG.mem_55_2 , n5841, \REG.mem_55_1 , 
            n5840, \REG.mem_55_0 , n5839, n5838, \REG.mem_40_4 , \REG.mem_41_4 , 
            \REG.mem_42_4 , \REG.mem_43_4 , n5836, n5835, n5834, n5833, 
            n5832, \REG.mem_54_15 , n5831, \REG.mem_54_14 , n5830, 
            n5829, n5828, n5827, n5826, n5825, \REG.mem_54_8 , n5824, 
            n5823, \REG.mem_54_6 , n5822, \REG.mem_54_5 , n5821, \REG.mem_54_4 , 
            \REG.mem_46_4 , \REG.mem_47_4 , \REG.mem_44_4 , \REG.mem_45_4 , 
            n5820, \REG.mem_54_3 , n5819, \REG.mem_54_2 , n5818, \REG.mem_54_1 , 
            n5817, \REG.mem_54_0 , \REG.mem_25_4 , \REG.mem_30_4 , \REG.mem_31_4 , 
            \REG.mem_8_4 , \REG.mem_9_4 , \REG.mem_10_4 , \REG.mem_11_4 , 
            \REG.mem_14_4 , \REG.mem_15_4 , \REG.mem_12_4 , \REG.mem_13_4 , 
            n5768, \REG.mem_50_15 , n5767, \REG.mem_50_14 , n5766, 
            \REG.mem_50_13 , n5765, n5764, n5763, n5762, n5761, 
            \REG.mem_50_8 , n5760, n5759, \REG.mem_50_6 , n5758, \REG.mem_50_5 , 
            n5757, \REG.mem_50_4 , n10700, n5756, \REG.mem_50_3 , 
            n5755, \REG.mem_50_2 , n5754, n4893, \fifo_data_out[14] , 
            n4896, \fifo_data_out[15] , n5750, \REG.mem_50_0 , \REG.mem_38_5 , 
            \REG.mem_39_5 , n5733, \REG.mem_48_15 , n5732, \REG.mem_48_14 , 
            n5731, \REG.mem_48_13 , n5730, n5729, n5728, n5727, 
            n5726, \REG.mem_48_8 , n5725, n5724, \REG.mem_48_6 , n10748, 
            n5723, \REG.mem_48_5 , n5722, \REG.mem_48_4 , n5721, \REG.mem_48_3 , 
            n5720, \REG.mem_48_2 , n5719, \REG.mem_42_6 , \REG.mem_43_6 , 
            n5718, \REG.mem_48_0 , n5717, \REG.mem_47_15 , \REG.mem_41_6 , 
            \REG.mem_40_6 , n5716, \REG.mem_47_14 , n5715, \REG.mem_47_13 , 
            n5714, n5713, \REG.mem_47_11 , n5712, \REG.mem_47_10 , 
            n5711, n5710, n5709, \REG.mem_47_7 , n5708, \REG.mem_47_6 , 
            n5707, n5706, n5705, n5704, n5703, \REG.mem_25_12 , 
            \REG.mem_37_5 , \REG.mem_36_5 , n5702, \REG.mem_47_0 , n5701, 
            \REG.mem_46_15 , n5700, \REG.mem_46_14 , n5699, \REG.mem_46_13 , 
            n5698, n5697, \REG.mem_46_11 , n5696, \REG.mem_46_10 , 
            n5695, n5694, n5693, \REG.mem_46_7 , n5692, \REG.mem_46_6 , 
            n5691, n5690, n5689, n5688, n5687, n5686, \REG.mem_46_0 , 
            n5685, \REG.mem_45_15 , n5684, \REG.mem_45_14 , n5683, 
            \REG.mem_45_13 , n5682, n5681, \REG.mem_45_11 , n5680, 
            \REG.mem_45_10 , n5679, n5678, \REG.mem_6_15 , \REG.mem_7_15 , 
            \REG.mem_3_1 , n5677, \REG.mem_45_7 , \REG.mem_5_15 , \REG.mem_4_15 , 
            n5676, \REG.mem_45_6 , n5675, n5674, n5673, n5672, n5671, 
            n5670, \REG.mem_45_0 , n5668, \REG.mem_44_15 , n5667, 
            \REG.mem_44_14 , n5665, \REG.mem_44_13 , n5664, n5663, 
            \REG.mem_44_11 , n5661, \REG.mem_44_10 , n5660, n5659, 
            n5658, \REG.mem_44_7 , n5657, \REG.mem_44_6 , n5656, n5655, 
            n5654, n5653, n5652, n5651, \REG.mem_44_0 , n5650, n5649, 
            \REG.mem_43_14 , n5648, n5647, n5646, \REG.mem_43_11 , 
            n5645, \REG.mem_43_10 , n5644, \REG.mem_43_9 , \rd_addr_p1_w[0] , 
            \REG.mem_18_7 , n5643, n5642, \REG.mem_43_7 , n5641, n5640, 
            \REG.mem_43_5 , n5639, n5638, \REG.mem_43_3 , n5637, n5636, 
            \REG.mem_43_1 , n5635, n5634, n5633, \REG.mem_42_14 , 
            n5632, n5631, n5630, \REG.mem_42_11 , n5629, \REG.mem_42_10 , 
            n4916, \REG.mem_22_11 , \REG.mem_23_11 , n5628, \REG.mem_42_9 , 
            n5627, n5626, \REG.mem_42_7 , n5625, n5624, \REG.mem_42_5 , 
            n5623, n5622, \REG.mem_42_3 , n5621, n5620, \REG.mem_42_1 , 
            n5619, n5618, \REG.mem_41_15 , n5617, \REG.mem_41_14 , 
            n5616, n5615, n5614, \REG.mem_41_11 , n5613, \REG.mem_41_10 , 
            \REG.mem_25_6 , n5612, \REG.mem_41_9 , n5611, n5610, \REG.mem_41_7 , 
            n5609, n5608, \REG.mem_41_5 , n5607, n5606, \REG.mem_41_3 , 
            n5605, n5604, \REG.mem_41_1 , n5603, n5602, \REG.mem_40_15 , 
            n5601, \REG.mem_40_14 , n5600, n5599, n5598, \REG.mem_40_11 , 
            n5597, \REG.mem_40_10 , n4904, n4903, n4901, n4899, 
            n5596, \REG.mem_40_9 , n5595, n5594, \REG.mem_40_7 , n5593, 
            n5592, \REG.mem_40_5 , n5591, n5590, \REG.mem_40_3 , n5589, 
            n5588, \REG.mem_40_1 , n5587, n5586, n5585, \REG.mem_39_14 , 
            n5584, n5583, \REG.mem_39_12 , n5582, \REG.mem_39_11 , 
            n5581, \REG.mem_39_10 , n4898, DEBUG_5_c, \REG.mem_3_4 , 
            \REG.mem_6_4 , \REG.mem_7_4 , n5580, \REG.mem_39_9 , n5579, 
            \REG.mem_39_8 , n5578, n5577, n5576, n5575, \REG.mem_39_4 , 
            n5574, \REG.mem_39_3 , n5573, \REG.mem_39_2 , n5572, \REG.mem_39_1 , 
            n5570, n5569, n5568, \REG.mem_38_14 , n5567, n5566, 
            \REG.mem_38_12 , n5565, \REG.mem_38_11 , n5564, \REG.mem_38_10 , 
            \REG.mem_5_4 , \REG.mem_4_4 , n5563, \REG.mem_38_9 , n5562, 
            \REG.mem_38_8 , n5561, n5560, n5559, n5558, \REG.mem_38_4 , 
            n5557, \REG.mem_38_3 , n5556, \REG.mem_38_2 , n5555, \REG.mem_38_1 , 
            n5554, n5553, n5552, \REG.mem_37_14 , n5551, n5550, 
            \REG.mem_37_12 , n5549, \REG.mem_37_11 , \REG.out_raw[15] , 
            \REG.out_raw[14] , \REG.out_raw[13] , \REG.out_raw[12] , \REG.out_raw[11] , 
            n5548, \REG.mem_37_10 , n5547, \REG.mem_37_9 , n5546, 
            \REG.mem_37_8 , n5545, n5544, n5543, n5542, \REG.mem_37_4 , 
            n5541, \REG.mem_37_3 , n5540, \REG.mem_37_2 , n5539, \REG.mem_37_1 , 
            n5538, \REG.out_raw[10] , \REG.out_raw[9] , \REG.out_raw[8] , 
            \REG.out_raw[7] , \REG.out_raw[6] , \REG.out_raw[5] , \REG.out_raw[4] , 
            \REG.out_raw[3] , \REG.out_raw[2] , \REG.out_raw[1] , n5524, 
            n5523, \REG.mem_36_14 , n5522, n5521, \REG.mem_36_12 , 
            n5520, \REG.mem_36_11 , n5519, \REG.mem_36_10 , n5518, 
            \REG.mem_36_9 , n5517, \REG.mem_36_8 , n5516, \rd_sig_diff0_w[2] , 
            n5515, n5514, n5513, \REG.mem_36_4 , n5512, \REG.mem_36_3 , 
            n5511, \REG.mem_36_2 , n5510, \REG.mem_36_1 , n5509, n5505, 
            n5504, \REG.mem_35_14 , n5503, n5502, \REG.mem_35_12 , 
            n5501, \REG.mem_35_11 , n5500, \REG.mem_35_10 , \rd_sig_diff0_w[1] , 
            n5499, n5498, \REG.mem_35_8 , n5497, n5496, n5495, \REG.mem_35_5 , 
            n5494, \REG.mem_35_4 , n5493, \REG.mem_35_3 , n5492, \REG.mem_35_2 , 
            n5491, \REG.mem_35_1 , n5490, \REG.mem_25_11 , \REG.mem_10_13 , 
            \REG.mem_11_13 , \REG.mem_9_13 , \REG.mem_8_13 , n5440, 
            n5439, \REG.mem_31_14 , n5438, n5437, \REG.mem_31_12 , 
            n5436, \REG.mem_31_11 , n5435, \REG.mem_31_10 , n5434, 
            n5433, \REG.mem_31_8 , n5432, \REG.mem_31_7 , n5431, \REG.mem_31_6 , 
            n5430, n5429, n5428, \REG.mem_31_3 , n5427, n5426, \REG.mem_31_1 , 
            n5425, n5424, n5423, \REG.mem_30_14 , n5422, n5421, 
            \REG.mem_30_12 , n5420, \REG.mem_30_11 , DEBUG_1_c_c, write_to_dc32_fifo_latched_N_425, 
            \REG.mem_18_6 , n5419, \REG.mem_30_10 , n5418, n5417, 
            \REG.mem_30_8 , n5416, \REG.mem_30_7 , n5415, \REG.mem_30_6 , 
            n5414, n5413, n5412, \REG.mem_30_3 , n5411, n5410, \REG.mem_30_1 , 
            n5409, \REG.mem_16_6 , \wr_addr_nxt_c[1] , \REG.mem_10_9 , 
            \REG.mem_11_9 , \REG.mem_9_9 , \REG.mem_8_9 , \REG.mem_14_13 , 
            \REG.mem_15_13 , \REG.mem_13_13 , \REG.mem_12_13 , n56, 
            \REG.mem_14_9 , \REG.mem_15_9 , \REG.mem_10_15 , \REG.mem_11_15 , 
            \REG.mem_9_15 , \REG.mem_8_15 , \REG.mem_10_7 , \REG.mem_11_7 , 
            \REG.mem_13_9 , \REG.mem_12_9 , n5344, n5343, \REG.mem_25_14 , 
            n5342, n5341, n5340, n5339, \REG.mem_25_10 , n5338, 
            n5337, \REG.mem_25_8 , n5336, \REG.mem_25_7 , \REG.mem_18_13 , 
            \REG.mem_9_7 , \REG.mem_8_7 , \REG.mem_16_13 , n5335, n5334, 
            n5333, n5332, \REG.mem_25_3 , n5331, n5330, n5329, \REG.mem_25_0 , 
            n52, n20, n5306, \REG.mem_23_15 , n5305, \REG.mem_23_14 , 
            n5304, \REG.mem_23_13 , n5303, n5302, n5301, \REG.mem_23_10 , 
            n5300, \REG.mem_23_9 , n5299, n5298, n5297, \REG.mem_23_6 , 
            n5296, \REG.mem_23_5 , n5295, \REG.mem_23_4 , n5294, \REG.mem_23_3 , 
            n5293, \REG.mem_23_2 , n5292, \REG.mem_23_1 , n5291, \REG.mem_23_0 , 
            n5290, \REG.mem_22_15 , n5289, \REG.mem_22_14 , n5288, 
            \REG.mem_22_13 , n5287, n5286, n5285, \REG.mem_22_10 , 
            \rd_grey_sync_r[5] , \rd_grey_sync_r[4] , \rd_grey_sync_r[3] , 
            \rd_grey_sync_r[2] , \rd_grey_sync_r[1] , n5284, \REG.mem_22_9 , 
            n5283, n5282, n5281, \REG.mem_22_6 , n5280, \REG.mem_22_5 , 
            n5279, \REG.mem_22_4 , n5278, \REG.mem_22_3 , n5277, \REG.mem_22_2 , 
            n5276, \REG.mem_22_1 , n5275, \REG.mem_22_0 , \REG.mem_14_3 , 
            \REG.mem_15_3 , \REG.mem_13_3 , \REG.mem_12_3 , \REG.mem_10_8 , 
            \REG.mem_11_8 , \REG.mem_9_8 , \REG.mem_8_8 , get_next_word, 
            \REG.mem_16_2 , \REG.mem_18_2 , \REG.mem_18_3 , n5226, \REG.mem_18_15 , 
            n5225, \REG.mem_18_14 , n5224, n5223, n5222, n5221, 
            \REG.mem_18_10 , n5220, \REG.mem_18_9 , rd_fifo_en_w, \REG.mem_16_3 , 
            \REG.mem_16_15 , n5219, n5218, n5217, n5216, n5215, 
            \REG.mem_18_4 , n5214, n5213, n5212, \REG.mem_18_1 , n5211, 
            \REG.mem_18_0 , n5190, n5188, \REG.mem_16_14 , n5187, 
            n5186, n5185, n5184, \REG.mem_16_10 , \REG.mem_3_2 , \REG.mem_3_0 , 
            n5183, \REG.mem_16_9 , n5182, n5181, n5180, n5179, n5178, 
            \REG.mem_16_4 , n5177, n5176, \REG.mem_6_0 , \REG.mem_7_0 , 
            n5175, \REG.mem_16_1 , n5174, \REG.mem_16_0 , n5171, \REG.mem_15_15 , 
            n5170, n5169, n5168, n5167, n5166, \REG.mem_15_10 , 
            n5165, n5164, n5163, n5162, \REG.mem_15_6 , \REG.mem_5_0 , 
            \REG.mem_4_0 , n5161, n5160, n5159, n5158, n5157, \REG.mem_15_1 , 
            n5156, \REG.mem_15_0 , n5155, \REG.mem_14_15 , n5154, 
            n5153, n5152, n5151, n5150, \REG.mem_14_10 , n5149, 
            n5148, n5147, n5146, \REG.mem_14_6 , n5145, n5144, n5143, 
            n5142, n5141, \REG.mem_14_1 , n5140, \REG.mem_14_0 , n5139, 
            \REG.mem_13_15 , n5138, n5137, n5136, n5135, n5134, 
            \REG.mem_13_10 , n5133, n5132, n5131, n47, n15, n50, 
            n5130, \REG.mem_13_6 , n18, n5129, n5128, n5127, n5126, 
            n5125, \REG.mem_13_1 , n5124, \REG.mem_13_0 , n5123, \REG.mem_12_15 , 
            n5122, n5121, n5120, n5119, n5118, \REG.mem_12_10 , 
            n5117, n5116, \REG.mem_3_12 , \REG.mem_3_14 , n5115, n5114, 
            \REG.mem_12_6 , n5113, n5112, n53, n21, \REG.mem_10_0 , 
            \REG.mem_11_0 , \REG.mem_9_0 , \REG.mem_8_0 , n5111, n5110, 
            n5109, \REG.mem_12_1 , n5108, \REG.mem_12_0 , n51, n19, 
            n5107, n54, n22, n5106, n5105, n5104, \REG.mem_11_12 , 
            n5103, n5102, \REG.mem_11_10 , n5101, n5100, n5099, 
            n5098, n5097, \REG.mem_11_5 , \rd_addr_nxt_c_6__N_498[5] , 
            n5096, n5095, n5094, n5093, \REG.mem_11_1 , n5092, n5091, 
            n5090, n5089, n5088, \REG.mem_10_12 , n5087, n5086, 
            \REG.mem_10_10 , n5085, n5084, n5083, n5082, n5081, 
            \REG.mem_10_5 , n5080, \rd_addr_nxt_c_6__N_498[3] , n5079, 
            \rd_addr_nxt_c_6__N_498[2] , n49, n17, \REG.mem_6_14 , \REG.mem_7_14 , 
            \REG.mem_4_14 , \REG.mem_5_14 , n24, n5078, \REG.mem_3_6 , 
            n5077, \REG.mem_10_1 , n5076, n5075, \REG.mem_3_9 , n5074, 
            n5073, n55, n23, n40, n8, n5072, \REG.mem_9_12 , n34, 
            n5071, n5070, \REG.mem_9_10 , n5069, n2, n5068, n5067, 
            n5066, n5065, \REG.mem_9_5 , n5064, n5063, n5062, n5061, 
            \REG.mem_9_1 , n5060, n5059, n5058, n5057, n5056, \REG.mem_8_12 , 
            n5055, n5054, \REG.mem_8_10 , n5053, n5052, n5051, n5050, 
            n5049, \REG.mem_8_5 , n5048, n5047, n5046, n5045, \REG.mem_8_1 , 
            n5044, n5043, n5042, n5041, \REG.mem_7_13 , n5040, \REG.mem_7_12 , 
            n5039, n5038, \REG.mem_7_10 , n5037, n5036, n5035, \REG.mem_7_7 , 
            n5034, \REG.mem_7_6 , n5033, n5032, n5031, n5030, n5029, 
            n5028, n5027, n5026, n5025, \REG.mem_6_13 , n5024, \REG.mem_6_12 , 
            n5023, n5022, \REG.mem_6_10 , n5021, n5020, n5019, \REG.mem_6_7 , 
            n5018, \REG.mem_6_6 , n5017, n5016, n5015, n5014, n5013, 
            n5012, n5011, n5010, n5009, \REG.mem_5_13 , n5008, \REG.mem_5_12 , 
            n5007, n5006, \REG.mem_5_10 , n5005, n5004, n5003, \REG.mem_5_7 , 
            n5002, \REG.mem_5_6 , n5001, n5000, n4999, n4998, n4997, 
            n4996, n4995, n4994, n4993, \REG.mem_4_13 , n4992, \REG.mem_4_12 , 
            n4991, n4990, \REG.mem_4_10 , n4989, n4988, n4987, \REG.mem_4_7 , 
            n4986, \REG.mem_4_6 , n4985, n4984, n4983, n4982, n4981, 
            n4980, n4979, n4978, n4977, \REG.mem_3_13 , n4976, n4975, 
            n4974, \REG.mem_3_10 , n4973, n4972, \REG.mem_3_8 , n4971, 
            \REG.mem_3_7 , n4970, n4969, FT_OE_N_420, n57, n25, 
            n42, n10, n58, n26, n43, n35, n11, n3, n4968, 
            n4967, n4966, n4965, n4964, n60, n28, n59, n27, 
            n61, n29, n4672, n4671, n4670, n4669, n4668, n4667, 
            n4666, n4665, n4664, n4663, n4662, n4661, n4660, n4659, 
            n4658) /* synthesis syn_module_defined=1 */ ;
    output dc32_fifo_almost_full;
    input FIFO_CLK_c;
    input reset_per_frame;
    output \REG.mem_16_7 ;
    output \rd_addr_r[0] ;
    output \REG.mem_6_2 ;
    output \REG.mem_7_2 ;
    input \dc32_fifo_data_in[7] ;
    output \REG.mem_46_9 ;
    output \REG.mem_47_9 ;
    output \REG.mem_25_5 ;
    input GND_net;
    output t_rd_fifo_en_w;
    output \REG.out_raw[0] ;
    input SLM_CLK_c;
    output \REG.mem_45_9 ;
    output \REG.mem_44_9 ;
    output \REG.mem_57_15 ;
    output \REG.mem_62_15 ;
    output \REG.mem_63_15 ;
    output \REG.mem_6_1 ;
    output \REG.mem_7_1 ;
    output \REG.mem_5_1 ;
    output \REG.mem_4_1 ;
    output \REG.mem_57_1 ;
    output \REG.mem_25_9 ;
    input \dc32_fifo_data_in[6] ;
    input \dc32_fifo_data_in[15] ;
    output \REG.mem_46_3 ;
    output \REG.mem_47_3 ;
    output \REG.mem_45_3 ;
    output \REG.mem_44_3 ;
    output \REG.mem_54_13 ;
    output \REG.mem_55_13 ;
    output \REG.mem_50_11 ;
    output \REG.mem_48_11 ;
    input \dc32_fifo_data_in[5] ;
    output \REG.mem_42_12 ;
    output \REG.mem_43_12 ;
    output \REG.mem_41_12 ;
    output \REG.mem_40_12 ;
    input \dc32_fifo_data_in[4] ;
    input \dc32_fifo_data_in[3] ;
    input \dc32_fifo_data_in[2] ;
    output \rd_grey_sync_r[0] ;
    output \REG.mem_57_6 ;
    output DEBUG_3_c;
    output [6:0]wr_grey_sync_r;
    input \dc32_fifo_data_in[1] ;
    output \REG.mem_54_11 ;
    output \REG.mem_55_11 ;
    input \aempty_flag_impl.ae_flag_nxt_w ;
    output dc32_fifo_almost_empty;
    output \REG.mem_14_12 ;
    output \REG.mem_15_12 ;
    output \REG.mem_30_0 ;
    output \REG.mem_31_0 ;
    output \REG.mem_13_12 ;
    output \REG.mem_12_12 ;
    output \REG.mem_3_5 ;
    output \REG.mem_6_5 ;
    output \REG.mem_7_5 ;
    output \REG.mem_4_5 ;
    output \REG.mem_5_5 ;
    output \REG.mem_57_11 ;
    output n62;
    output \REG.mem_62_13 ;
    output \REG.mem_63_13 ;
    output \REG.mem_46_1 ;
    output \REG.mem_47_1 ;
    output \REG.mem_45_1 ;
    output \REG.mem_44_1 ;
    input \dc32_fifo_data_in[0] ;
    output \REG.mem_3_11 ;
    output \REG.mem_6_11 ;
    output \REG.mem_7_11 ;
    output n30;
    output \REG.mem_5_2 ;
    output \REG.mem_4_2 ;
    output \REG.mem_18_5 ;
    output \REG.mem_62_1 ;
    output \REG.mem_63_1 ;
    output \REG.mem_38_13 ;
    output \REG.mem_39_13 ;
    output \REG.mem_5_11 ;
    output \REG.mem_4_11 ;
    input \dc32_fifo_data_in[8] ;
    output \REG.mem_14_5 ;
    output \REG.mem_15_5 ;
    output \REG.mem_13_5 ;
    output \REG.mem_12_5 ;
    output \REG.mem_30_9 ;
    output \REG.mem_31_9 ;
    output \wr_addr_nxt_c[5] ;
    output \REG.mem_46_12 ;
    output \REG.mem_47_12 ;
    output \REG.mem_45_12 ;
    output \REG.mem_44_12 ;
    output \REG.mem_62_11 ;
    output \REG.mem_63_11 ;
    output \REG.mem_57_8 ;
    output \REG.mem_62_6 ;
    output \REG.mem_63_6 ;
    output \REG.mem_62_8 ;
    output \REG.mem_63_8 ;
    output \REG.mem_35_0 ;
    output \REG.mem_25_15 ;
    output \REG.mem_35_7 ;
    output \REG.mem_35_9 ;
    output \REG.mem_18_12 ;
    output \REG.mem_16_12 ;
    output \REG.mem_14_8 ;
    output \REG.mem_15_8 ;
    output \REG.mem_13_8 ;
    output \REG.mem_12_8 ;
    output \REG.mem_14_2 ;
    output \REG.mem_15_2 ;
    output \REG.mem_13_2 ;
    output \REG.mem_12_2 ;
    output \REG.mem_38_7 ;
    output \REG.mem_39_7 ;
    output \REG.mem_36_7 ;
    output \REG.mem_37_7 ;
    output \REG.mem_50_12 ;
    output \REG.mem_48_12 ;
    output \REG.mem_62_9 ;
    output \REG.mem_63_9 ;
    output \REG.mem_6_9 ;
    output \REG.mem_7_9 ;
    output \REG.mem_35_6 ;
    output \REG.mem_5_9 ;
    output \REG.mem_4_9 ;
    output \REG.mem_37_13 ;
    output \REG.mem_36_13 ;
    output \REG.mem_42_8 ;
    output \REG.mem_43_8 ;
    output \REG.mem_41_8 ;
    output \REG.mem_40_8 ;
    output \REG.mem_22_7 ;
    output \REG.mem_23_7 ;
    output \REG.mem_10_11 ;
    output \REG.mem_11_11 ;
    output \REG.mem_9_11 ;
    output \REG.mem_8_11 ;
    output \REG.mem_3_15 ;
    output \REG.mem_46_8 ;
    output \REG.mem_47_8 ;
    output \REG.mem_45_8 ;
    output \REG.mem_44_8 ;
    output \REG.mem_46_5 ;
    output \REG.mem_47_5 ;
    output \REG.mem_45_5 ;
    output \REG.mem_44_5 ;
    output \REG.mem_10_2 ;
    output \REG.mem_11_2 ;
    output \REG.mem_54_9 ;
    output \REG.mem_55_9 ;
    output \REG.mem_57_9 ;
    output \REG.mem_57_14 ;
    output \REG.mem_30_15 ;
    output \REG.mem_31_15 ;
    output \REG.mem_42_15 ;
    output \REG.mem_43_15 ;
    output \REG.mem_16_5 ;
    output \REG.mem_9_2 ;
    output \REG.mem_8_2 ;
    output \REG.mem_62_12 ;
    output \REG.mem_63_12 ;
    output \wr_addr_nxt_c[3] ;
    output \REG.mem_18_8 ;
    output \REG.mem_16_8 ;
    output \REG.mem_22_12 ;
    output \REG.mem_23_12 ;
    output \REG.mem_25_2 ;
    output \REG.mem_30_2 ;
    output \REG.mem_31_2 ;
    input \dc32_fifo_data_in[14] ;
    output \REG.mem_48_10 ;
    output \REG.mem_50_10 ;
    input \dc32_fifo_data_in[13] ;
    output \REG.mem_54_10 ;
    output \REG.mem_55_10 ;
    output \REG.mem_14_11 ;
    output \REG.mem_15_11 ;
    input \dc32_fifo_data_in[12] ;
    output \REG.mem_54_12 ;
    output \REG.mem_55_12 ;
    output \REG.mem_13_11 ;
    output \REG.mem_12_11 ;
    output \REG.mem_35_15 ;
    output \REG.mem_38_6 ;
    output \REG.mem_39_6 ;
    input \dc32_fifo_data_in[11] ;
    output \REG.mem_37_6 ;
    output \REG.mem_36_6 ;
    output \REG.mem_57_13 ;
    input \dc32_fifo_data_in[10] ;
    input \dc32_fifo_data_in[9] ;
    output \REG.mem_30_13 ;
    output \REG.mem_31_13 ;
    output \REG.mem_30_5 ;
    output \REG.mem_31_5 ;
    output \REG.mem_48_7 ;
    output \REG.mem_50_7 ;
    output \REG.mem_54_7 ;
    output \REG.mem_55_7 ;
    input n6106;
    input VCC_net;
    output \fifo_data_out[2] ;
    input n6103;
    output \fifo_data_out[1] ;
    output \REG.mem_35_13 ;
    output \REG.mem_3_3 ;
    output \rd_addr_r[6] ;
    input n4827;
    output \fifo_data_out[3] ;
    output \REG.mem_50_1 ;
    input n4830;
    output \fifo_data_out[4] ;
    input n4841;
    output \fifo_data_out[5] ;
    input n4844;
    output \fifo_data_out[6] ;
    input n4848;
    output \fifo_data_out[7] ;
    input n4851;
    output \fifo_data_out[8] ;
    input n4854;
    output \fifo_data_out[9] ;
    input n4858;
    output \fifo_data_out[10] ;
    input n4864;
    output \fifo_data_out[11] ;
    output \REG.mem_62_14 ;
    output \REG.mem_63_14 ;
    output \REG.mem_48_1 ;
    output \REG.mem_18_11 ;
    output \REG.mem_16_11 ;
    output \REG.mem_6_3 ;
    output \REG.mem_7_3 ;
    output \REG.mem_5_3 ;
    output \REG.mem_4_3 ;
    output \REG.mem_42_2 ;
    output \REG.mem_43_2 ;
    output \REG.mem_41_2 ;
    output \REG.mem_40_2 ;
    input n6070;
    output \fifo_data_out[0] ;
    output \REG.mem_46_2 ;
    output \REG.mem_47_2 ;
    output \REG.mem_45_2 ;
    output \REG.mem_44_2 ;
    output \REG.mem_14_7 ;
    output \REG.mem_15_7 ;
    input n4872;
    output \fifo_data_out[12] ;
    input n4875;
    output \fifo_data_out[13] ;
    output \REG.mem_13_7 ;
    output \REG.mem_12_7 ;
    input n6034;
    output \REG.mem_25_13 ;
    input n6032;
    output \REG.mem_10_3 ;
    output \REG.mem_11_3 ;
    output \REG.mem_9_3 ;
    output \REG.mem_8_3 ;
    output \REG.mem_50_9 ;
    input n6013;
    input n6012;
    input n6011;
    input n6010;
    input n6009;
    input n6008;
    input n6007;
    output \REG.mem_63_10 ;
    input n6006;
    input n6005;
    input n6004;
    output \REG.mem_63_7 ;
    input n6003;
    input n6002;
    output \REG.mem_63_5 ;
    output \REG.mem_48_9 ;
    output \REG.mem_42_13 ;
    output \REG.mem_43_13 ;
    output \REG.mem_38_0 ;
    output \REG.mem_39_0 ;
    input n6001;
    output \REG.mem_63_4 ;
    input n6000;
    output \REG.mem_63_3 ;
    input n5999;
    output \REG.mem_63_2 ;
    input n5998;
    input n5997;
    output \REG.mem_63_0 ;
    input n5996;
    input n5995;
    input n5994;
    input n5993;
    input n5992;
    input n5991;
    output \REG.mem_62_10 ;
    input n5990;
    input n5989;
    input n5988;
    output \REG.mem_62_7 ;
    input n5987;
    input n5986;
    output \REG.mem_62_5 ;
    input n5985;
    output \REG.mem_62_4 ;
    output \REG.mem_41_13 ;
    output \REG.mem_40_13 ;
    output \REG.mem_37_0 ;
    output \REG.mem_36_0 ;
    output \REG.mem_10_6 ;
    output \REG.mem_11_6 ;
    input n5984;
    output \REG.mem_62_3 ;
    input n5983;
    output \REG.mem_62_2 ;
    input n5982;
    input n5981;
    output \REG.mem_62_0 ;
    output \REG.mem_9_6 ;
    output \REG.mem_8_6 ;
    output \REG.mem_42_0 ;
    output \REG.mem_43_0 ;
    output \REG.mem_22_8 ;
    output \REG.mem_23_8 ;
    input n5946;
    output [6:0]rp_sync1_r;
    input n5945;
    input n5944;
    input n5943;
    input n5942;
    input n5941;
    input n5940;
    input n5939;
    input n5938;
    input n5921;
    input n5920;
    input n5919;
    output \REG.mem_41_0 ;
    output \REG.mem_40_0 ;
    input n5917;
    input n5916;
    input n5914;
    output \REG.mem_8_14 ;
    output \REG.mem_9_14 ;
    output \REG.mem_25_1 ;
    output \REG.mem_10_14 ;
    output \REG.mem_11_14 ;
    input n5894;
    input n5893;
    input n5892;
    input n5891;
    output \REG.mem_57_12 ;
    input n5890;
    input n5889;
    output \REG.mem_57_10 ;
    input n5888;
    input n5887;
    input n5886;
    output \REG.mem_57_7 ;
    output \REG.mem_6_8 ;
    output \REG.mem_7_8 ;
    output \REG.mem_38_15 ;
    output \REG.mem_39_15 ;
    input n5885;
    output \REG.mem_5_8 ;
    output \REG.mem_4_8 ;
    output \REG.mem_14_14 ;
    output \REG.mem_15_14 ;
    input n5884;
    output \REG.mem_57_5 ;
    input n5883;
    output \REG.mem_57_4 ;
    input n5882;
    output \REG.mem_57_3 ;
    input n5881;
    output \REG.mem_57_2 ;
    input n5880;
    input n5879;
    output \REG.mem_57_0 ;
    output \REG.mem_12_14 ;
    output \REG.mem_13_14 ;
    output \REG.mem_37_15 ;
    output \REG.mem_36_15 ;
    input n5861;
    output [6:0]wp_sync1_r;
    input n5860;
    input n5859;
    input n5858;
    input n5857;
    input n5856;
    input n5855;
    output \REG.mem_55_15 ;
    input n5854;
    output \REG.mem_55_14 ;
    input n5853;
    output \rd_sig_diff0_w[0] ;
    input n5852;
    input n5851;
    input n5850;
    input n5849;
    input n5848;
    output \REG.mem_55_8 ;
    input n5847;
    input n5846;
    output \REG.mem_55_6 ;
    input n5845;
    output \REG.mem_55_5 ;
    input n5844;
    output \REG.mem_55_4 ;
    input n5843;
    output \REG.mem_55_3 ;
    input n5842;
    output \REG.mem_55_2 ;
    input n5841;
    output \REG.mem_55_1 ;
    input n5840;
    output \REG.mem_55_0 ;
    input n5839;
    input n5838;
    output \REG.mem_40_4 ;
    output \REG.mem_41_4 ;
    output \REG.mem_42_4 ;
    output \REG.mem_43_4 ;
    input n5836;
    input n5835;
    input n5834;
    input n5833;
    input n5832;
    output \REG.mem_54_15 ;
    input n5831;
    output \REG.mem_54_14 ;
    input n5830;
    input n5829;
    input n5828;
    input n5827;
    input n5826;
    input n5825;
    output \REG.mem_54_8 ;
    input n5824;
    input n5823;
    output \REG.mem_54_6 ;
    input n5822;
    output \REG.mem_54_5 ;
    input n5821;
    output \REG.mem_54_4 ;
    output \REG.mem_46_4 ;
    output \REG.mem_47_4 ;
    output \REG.mem_44_4 ;
    output \REG.mem_45_4 ;
    input n5820;
    output \REG.mem_54_3 ;
    input n5819;
    output \REG.mem_54_2 ;
    input n5818;
    output \REG.mem_54_1 ;
    input n5817;
    output \REG.mem_54_0 ;
    output \REG.mem_25_4 ;
    output \REG.mem_30_4 ;
    output \REG.mem_31_4 ;
    output \REG.mem_8_4 ;
    output \REG.mem_9_4 ;
    output \REG.mem_10_4 ;
    output \REG.mem_11_4 ;
    output \REG.mem_14_4 ;
    output \REG.mem_15_4 ;
    output \REG.mem_12_4 ;
    output \REG.mem_13_4 ;
    input n5768;
    output \REG.mem_50_15 ;
    input n5767;
    output \REG.mem_50_14 ;
    input n5766;
    output \REG.mem_50_13 ;
    input n5765;
    input n5764;
    input n5763;
    input n5762;
    input n5761;
    output \REG.mem_50_8 ;
    input n5760;
    input n5759;
    output \REG.mem_50_6 ;
    input n5758;
    output \REG.mem_50_5 ;
    input n5757;
    output \REG.mem_50_4 ;
    output n10700;
    input n5756;
    output \REG.mem_50_3 ;
    input n5755;
    output \REG.mem_50_2 ;
    input n5754;
    input n4893;
    output \fifo_data_out[14] ;
    input n4896;
    output \fifo_data_out[15] ;
    input n5750;
    output \REG.mem_50_0 ;
    output \REG.mem_38_5 ;
    output \REG.mem_39_5 ;
    input n5733;
    output \REG.mem_48_15 ;
    input n5732;
    output \REG.mem_48_14 ;
    input n5731;
    output \REG.mem_48_13 ;
    input n5730;
    input n5729;
    input n5728;
    input n5727;
    input n5726;
    output \REG.mem_48_8 ;
    input n5725;
    input n5724;
    output \REG.mem_48_6 ;
    output n10748;
    input n5723;
    output \REG.mem_48_5 ;
    input n5722;
    output \REG.mem_48_4 ;
    input n5721;
    output \REG.mem_48_3 ;
    input n5720;
    output \REG.mem_48_2 ;
    input n5719;
    output \REG.mem_42_6 ;
    output \REG.mem_43_6 ;
    input n5718;
    output \REG.mem_48_0 ;
    input n5717;
    output \REG.mem_47_15 ;
    output \REG.mem_41_6 ;
    output \REG.mem_40_6 ;
    input n5716;
    output \REG.mem_47_14 ;
    input n5715;
    output \REG.mem_47_13 ;
    input n5714;
    input n5713;
    output \REG.mem_47_11 ;
    input n5712;
    output \REG.mem_47_10 ;
    input n5711;
    input n5710;
    input n5709;
    output \REG.mem_47_7 ;
    input n5708;
    output \REG.mem_47_6 ;
    input n5707;
    input n5706;
    input n5705;
    input n5704;
    input n5703;
    output \REG.mem_25_12 ;
    output \REG.mem_37_5 ;
    output \REG.mem_36_5 ;
    input n5702;
    output \REG.mem_47_0 ;
    input n5701;
    output \REG.mem_46_15 ;
    input n5700;
    output \REG.mem_46_14 ;
    input n5699;
    output \REG.mem_46_13 ;
    input n5698;
    input n5697;
    output \REG.mem_46_11 ;
    input n5696;
    output \REG.mem_46_10 ;
    input n5695;
    input n5694;
    input n5693;
    output \REG.mem_46_7 ;
    input n5692;
    output \REG.mem_46_6 ;
    input n5691;
    input n5690;
    input n5689;
    input n5688;
    input n5687;
    input n5686;
    output \REG.mem_46_0 ;
    input n5685;
    output \REG.mem_45_15 ;
    input n5684;
    output \REG.mem_45_14 ;
    input n5683;
    output \REG.mem_45_13 ;
    input n5682;
    input n5681;
    output \REG.mem_45_11 ;
    input n5680;
    output \REG.mem_45_10 ;
    input n5679;
    input n5678;
    output \REG.mem_6_15 ;
    output \REG.mem_7_15 ;
    output \REG.mem_3_1 ;
    input n5677;
    output \REG.mem_45_7 ;
    output \REG.mem_5_15 ;
    output \REG.mem_4_15 ;
    input n5676;
    output \REG.mem_45_6 ;
    input n5675;
    input n5674;
    input n5673;
    input n5672;
    input n5671;
    input n5670;
    output \REG.mem_45_0 ;
    input n5668;
    output \REG.mem_44_15 ;
    input n5667;
    output \REG.mem_44_14 ;
    input n5665;
    output \REG.mem_44_13 ;
    input n5664;
    input n5663;
    output \REG.mem_44_11 ;
    input n5661;
    output \REG.mem_44_10 ;
    input n5660;
    input n5659;
    input n5658;
    output \REG.mem_44_7 ;
    input n5657;
    output \REG.mem_44_6 ;
    input n5656;
    input n5655;
    input n5654;
    input n5653;
    input n5652;
    input n5651;
    output \REG.mem_44_0 ;
    input n5650;
    input n5649;
    output \REG.mem_43_14 ;
    input n5648;
    input n5647;
    input n5646;
    output \REG.mem_43_11 ;
    input n5645;
    output \REG.mem_43_10 ;
    input n5644;
    output \REG.mem_43_9 ;
    output \rd_addr_p1_w[0] ;
    output \REG.mem_18_7 ;
    input n5643;
    input n5642;
    output \REG.mem_43_7 ;
    input n5641;
    input n5640;
    output \REG.mem_43_5 ;
    input n5639;
    input n5638;
    output \REG.mem_43_3 ;
    input n5637;
    input n5636;
    output \REG.mem_43_1 ;
    input n5635;
    input n5634;
    input n5633;
    output \REG.mem_42_14 ;
    input n5632;
    input n5631;
    input n5630;
    output \REG.mem_42_11 ;
    input n5629;
    output \REG.mem_42_10 ;
    input n4916;
    output \REG.mem_22_11 ;
    output \REG.mem_23_11 ;
    input n5628;
    output \REG.mem_42_9 ;
    input n5627;
    input n5626;
    output \REG.mem_42_7 ;
    input n5625;
    input n5624;
    output \REG.mem_42_5 ;
    input n5623;
    input n5622;
    output \REG.mem_42_3 ;
    input n5621;
    input n5620;
    output \REG.mem_42_1 ;
    input n5619;
    input n5618;
    output \REG.mem_41_15 ;
    input n5617;
    output \REG.mem_41_14 ;
    input n5616;
    input n5615;
    input n5614;
    output \REG.mem_41_11 ;
    input n5613;
    output \REG.mem_41_10 ;
    output \REG.mem_25_6 ;
    input n5612;
    output \REG.mem_41_9 ;
    input n5611;
    input n5610;
    output \REG.mem_41_7 ;
    input n5609;
    input n5608;
    output \REG.mem_41_5 ;
    input n5607;
    input n5606;
    output \REG.mem_41_3 ;
    input n5605;
    input n5604;
    output \REG.mem_41_1 ;
    input n5603;
    input n5602;
    output \REG.mem_40_15 ;
    input n5601;
    output \REG.mem_40_14 ;
    input n5600;
    input n5599;
    input n5598;
    output \REG.mem_40_11 ;
    input n5597;
    output \REG.mem_40_10 ;
    input n4904;
    input n4903;
    input n4901;
    input n4899;
    input n5596;
    output \REG.mem_40_9 ;
    input n5595;
    input n5594;
    output \REG.mem_40_7 ;
    input n5593;
    input n5592;
    output \REG.mem_40_5 ;
    input n5591;
    input n5590;
    output \REG.mem_40_3 ;
    input n5589;
    input n5588;
    output \REG.mem_40_1 ;
    input n5587;
    input n5586;
    input n5585;
    output \REG.mem_39_14 ;
    input n5584;
    input n5583;
    output \REG.mem_39_12 ;
    input n5582;
    output \REG.mem_39_11 ;
    input n5581;
    output \REG.mem_39_10 ;
    input n4898;
    input DEBUG_5_c;
    output \REG.mem_3_4 ;
    output \REG.mem_6_4 ;
    output \REG.mem_7_4 ;
    input n5580;
    output \REG.mem_39_9 ;
    input n5579;
    output \REG.mem_39_8 ;
    input n5578;
    input n5577;
    input n5576;
    input n5575;
    output \REG.mem_39_4 ;
    input n5574;
    output \REG.mem_39_3 ;
    input n5573;
    output \REG.mem_39_2 ;
    input n5572;
    output \REG.mem_39_1 ;
    input n5570;
    input n5569;
    input n5568;
    output \REG.mem_38_14 ;
    input n5567;
    input n5566;
    output \REG.mem_38_12 ;
    input n5565;
    output \REG.mem_38_11 ;
    input n5564;
    output \REG.mem_38_10 ;
    output \REG.mem_5_4 ;
    output \REG.mem_4_4 ;
    input n5563;
    output \REG.mem_38_9 ;
    input n5562;
    output \REG.mem_38_8 ;
    input n5561;
    input n5560;
    input n5559;
    input n5558;
    output \REG.mem_38_4 ;
    input n5557;
    output \REG.mem_38_3 ;
    input n5556;
    output \REG.mem_38_2 ;
    input n5555;
    output \REG.mem_38_1 ;
    input n5554;
    input n5553;
    input n5552;
    output \REG.mem_37_14 ;
    input n5551;
    input n5550;
    output \REG.mem_37_12 ;
    input n5549;
    output \REG.mem_37_11 ;
    output \REG.out_raw[15] ;
    output \REG.out_raw[14] ;
    output \REG.out_raw[13] ;
    output \REG.out_raw[12] ;
    output \REG.out_raw[11] ;
    input n5548;
    output \REG.mem_37_10 ;
    input n5547;
    output \REG.mem_37_9 ;
    input n5546;
    output \REG.mem_37_8 ;
    input n5545;
    input n5544;
    input n5543;
    input n5542;
    output \REG.mem_37_4 ;
    input n5541;
    output \REG.mem_37_3 ;
    input n5540;
    output \REG.mem_37_2 ;
    input n5539;
    output \REG.mem_37_1 ;
    input n5538;
    output \REG.out_raw[10] ;
    output \REG.out_raw[9] ;
    output \REG.out_raw[8] ;
    output \REG.out_raw[7] ;
    output \REG.out_raw[6] ;
    output \REG.out_raw[5] ;
    output \REG.out_raw[4] ;
    output \REG.out_raw[3] ;
    output \REG.out_raw[2] ;
    output \REG.out_raw[1] ;
    input n5524;
    input n5523;
    output \REG.mem_36_14 ;
    input n5522;
    input n5521;
    output \REG.mem_36_12 ;
    input n5520;
    output \REG.mem_36_11 ;
    input n5519;
    output \REG.mem_36_10 ;
    input n5518;
    output \REG.mem_36_9 ;
    input n5517;
    output \REG.mem_36_8 ;
    input n5516;
    output \rd_sig_diff0_w[2] ;
    input n5515;
    input n5514;
    input n5513;
    output \REG.mem_36_4 ;
    input n5512;
    output \REG.mem_36_3 ;
    input n5511;
    output \REG.mem_36_2 ;
    input n5510;
    output \REG.mem_36_1 ;
    input n5509;
    input n5505;
    input n5504;
    output \REG.mem_35_14 ;
    input n5503;
    input n5502;
    output \REG.mem_35_12 ;
    input n5501;
    output \REG.mem_35_11 ;
    input n5500;
    output \REG.mem_35_10 ;
    output \rd_sig_diff0_w[1] ;
    input n5499;
    input n5498;
    output \REG.mem_35_8 ;
    input n5497;
    input n5496;
    input n5495;
    output \REG.mem_35_5 ;
    input n5494;
    output \REG.mem_35_4 ;
    input n5493;
    output \REG.mem_35_3 ;
    input n5492;
    output \REG.mem_35_2 ;
    input n5491;
    output \REG.mem_35_1 ;
    input n5490;
    output \REG.mem_25_11 ;
    output \REG.mem_10_13 ;
    output \REG.mem_11_13 ;
    output \REG.mem_9_13 ;
    output \REG.mem_8_13 ;
    input n5440;
    input n5439;
    output \REG.mem_31_14 ;
    input n5438;
    input n5437;
    output \REG.mem_31_12 ;
    input n5436;
    output \REG.mem_31_11 ;
    input n5435;
    output \REG.mem_31_10 ;
    input n5434;
    input n5433;
    output \REG.mem_31_8 ;
    input n5432;
    output \REG.mem_31_7 ;
    input n5431;
    output \REG.mem_31_6 ;
    input n5430;
    input n5429;
    input n5428;
    output \REG.mem_31_3 ;
    input n5427;
    input n5426;
    output \REG.mem_31_1 ;
    input n5425;
    input n5424;
    input n5423;
    output \REG.mem_30_14 ;
    input n5422;
    input n5421;
    output \REG.mem_30_12 ;
    input n5420;
    output \REG.mem_30_11 ;
    input DEBUG_1_c_c;
    output write_to_dc32_fifo_latched_N_425;
    output \REG.mem_18_6 ;
    input n5419;
    output \REG.mem_30_10 ;
    input n5418;
    input n5417;
    output \REG.mem_30_8 ;
    input n5416;
    output \REG.mem_30_7 ;
    input n5415;
    output \REG.mem_30_6 ;
    input n5414;
    input n5413;
    input n5412;
    output \REG.mem_30_3 ;
    input n5411;
    input n5410;
    output \REG.mem_30_1 ;
    input n5409;
    output \REG.mem_16_6 ;
    output \wr_addr_nxt_c[1] ;
    output \REG.mem_10_9 ;
    output \REG.mem_11_9 ;
    output \REG.mem_9_9 ;
    output \REG.mem_8_9 ;
    output \REG.mem_14_13 ;
    output \REG.mem_15_13 ;
    output \REG.mem_13_13 ;
    output \REG.mem_12_13 ;
    output n56;
    output \REG.mem_14_9 ;
    output \REG.mem_15_9 ;
    output \REG.mem_10_15 ;
    output \REG.mem_11_15 ;
    output \REG.mem_9_15 ;
    output \REG.mem_8_15 ;
    output \REG.mem_10_7 ;
    output \REG.mem_11_7 ;
    output \REG.mem_13_9 ;
    output \REG.mem_12_9 ;
    input n5344;
    input n5343;
    output \REG.mem_25_14 ;
    input n5342;
    input n5341;
    input n5340;
    input n5339;
    output \REG.mem_25_10 ;
    input n5338;
    input n5337;
    output \REG.mem_25_8 ;
    input n5336;
    output \REG.mem_25_7 ;
    output \REG.mem_18_13 ;
    output \REG.mem_9_7 ;
    output \REG.mem_8_7 ;
    output \REG.mem_16_13 ;
    input n5335;
    input n5334;
    input n5333;
    input n5332;
    output \REG.mem_25_3 ;
    input n5331;
    input n5330;
    input n5329;
    output \REG.mem_25_0 ;
    output n52;
    output n20;
    input n5306;
    output \REG.mem_23_15 ;
    input n5305;
    output \REG.mem_23_14 ;
    input n5304;
    output \REG.mem_23_13 ;
    input n5303;
    input n5302;
    input n5301;
    output \REG.mem_23_10 ;
    input n5300;
    output \REG.mem_23_9 ;
    input n5299;
    input n5298;
    input n5297;
    output \REG.mem_23_6 ;
    input n5296;
    output \REG.mem_23_5 ;
    input n5295;
    output \REG.mem_23_4 ;
    input n5294;
    output \REG.mem_23_3 ;
    input n5293;
    output \REG.mem_23_2 ;
    input n5292;
    output \REG.mem_23_1 ;
    input n5291;
    output \REG.mem_23_0 ;
    input n5290;
    output \REG.mem_22_15 ;
    input n5289;
    output \REG.mem_22_14 ;
    input n5288;
    output \REG.mem_22_13 ;
    input n5287;
    input n5286;
    input n5285;
    output \REG.mem_22_10 ;
    output \rd_grey_sync_r[5] ;
    output \rd_grey_sync_r[4] ;
    output \rd_grey_sync_r[3] ;
    output \rd_grey_sync_r[2] ;
    output \rd_grey_sync_r[1] ;
    input n5284;
    output \REG.mem_22_9 ;
    input n5283;
    input n5282;
    input n5281;
    output \REG.mem_22_6 ;
    input n5280;
    output \REG.mem_22_5 ;
    input n5279;
    output \REG.mem_22_4 ;
    input n5278;
    output \REG.mem_22_3 ;
    input n5277;
    output \REG.mem_22_2 ;
    input n5276;
    output \REG.mem_22_1 ;
    input n5275;
    output \REG.mem_22_0 ;
    output \REG.mem_14_3 ;
    output \REG.mem_15_3 ;
    output \REG.mem_13_3 ;
    output \REG.mem_12_3 ;
    output \REG.mem_10_8 ;
    output \REG.mem_11_8 ;
    output \REG.mem_9_8 ;
    output \REG.mem_8_8 ;
    input get_next_word;
    output \REG.mem_16_2 ;
    output \REG.mem_18_2 ;
    output \REG.mem_18_3 ;
    input n5226;
    output \REG.mem_18_15 ;
    input n5225;
    output \REG.mem_18_14 ;
    input n5224;
    input n5223;
    input n5222;
    input n5221;
    output \REG.mem_18_10 ;
    input n5220;
    output \REG.mem_18_9 ;
    output rd_fifo_en_w;
    output \REG.mem_16_3 ;
    output \REG.mem_16_15 ;
    input n5219;
    input n5218;
    input n5217;
    input n5216;
    input n5215;
    output \REG.mem_18_4 ;
    input n5214;
    input n5213;
    input n5212;
    output \REG.mem_18_1 ;
    input n5211;
    output \REG.mem_18_0 ;
    input n5190;
    input n5188;
    output \REG.mem_16_14 ;
    input n5187;
    input n5186;
    input n5185;
    input n5184;
    output \REG.mem_16_10 ;
    output \REG.mem_3_2 ;
    output \REG.mem_3_0 ;
    input n5183;
    output \REG.mem_16_9 ;
    input n5182;
    input n5181;
    input n5180;
    input n5179;
    input n5178;
    output \REG.mem_16_4 ;
    input n5177;
    input n5176;
    output \REG.mem_6_0 ;
    output \REG.mem_7_0 ;
    input n5175;
    output \REG.mem_16_1 ;
    input n5174;
    output \REG.mem_16_0 ;
    input n5171;
    output \REG.mem_15_15 ;
    input n5170;
    input n5169;
    input n5168;
    input n5167;
    input n5166;
    output \REG.mem_15_10 ;
    input n5165;
    input n5164;
    input n5163;
    input n5162;
    output \REG.mem_15_6 ;
    output \REG.mem_5_0 ;
    output \REG.mem_4_0 ;
    input n5161;
    input n5160;
    input n5159;
    input n5158;
    input n5157;
    output \REG.mem_15_1 ;
    input n5156;
    output \REG.mem_15_0 ;
    input n5155;
    output \REG.mem_14_15 ;
    input n5154;
    input n5153;
    input n5152;
    input n5151;
    input n5150;
    output \REG.mem_14_10 ;
    input n5149;
    input n5148;
    input n5147;
    input n5146;
    output \REG.mem_14_6 ;
    input n5145;
    input n5144;
    input n5143;
    input n5142;
    input n5141;
    output \REG.mem_14_1 ;
    input n5140;
    output \REG.mem_14_0 ;
    input n5139;
    output \REG.mem_13_15 ;
    input n5138;
    input n5137;
    input n5136;
    input n5135;
    input n5134;
    output \REG.mem_13_10 ;
    input n5133;
    input n5132;
    input n5131;
    output n47;
    output n15;
    output n50;
    input n5130;
    output \REG.mem_13_6 ;
    output n18;
    input n5129;
    input n5128;
    input n5127;
    input n5126;
    input n5125;
    output \REG.mem_13_1 ;
    input n5124;
    output \REG.mem_13_0 ;
    input n5123;
    output \REG.mem_12_15 ;
    input n5122;
    input n5121;
    input n5120;
    input n5119;
    input n5118;
    output \REG.mem_12_10 ;
    input n5117;
    input n5116;
    output \REG.mem_3_12 ;
    output \REG.mem_3_14 ;
    input n5115;
    input n5114;
    output \REG.mem_12_6 ;
    input n5113;
    input n5112;
    output n53;
    output n21;
    output \REG.mem_10_0 ;
    output \REG.mem_11_0 ;
    output \REG.mem_9_0 ;
    output \REG.mem_8_0 ;
    input n5111;
    input n5110;
    input n5109;
    output \REG.mem_12_1 ;
    input n5108;
    output \REG.mem_12_0 ;
    output n51;
    output n19;
    input n5107;
    output n54;
    output n22;
    input n5106;
    input n5105;
    input n5104;
    output \REG.mem_11_12 ;
    input n5103;
    input n5102;
    output \REG.mem_11_10 ;
    input n5101;
    input n5100;
    input n5099;
    input n5098;
    input n5097;
    output \REG.mem_11_5 ;
    output \rd_addr_nxt_c_6__N_498[5] ;
    input n5096;
    input n5095;
    input n5094;
    input n5093;
    output \REG.mem_11_1 ;
    input n5092;
    input n5091;
    input n5090;
    input n5089;
    input n5088;
    output \REG.mem_10_12 ;
    input n5087;
    input n5086;
    output \REG.mem_10_10 ;
    input n5085;
    input n5084;
    input n5083;
    input n5082;
    input n5081;
    output \REG.mem_10_5 ;
    input n5080;
    output \rd_addr_nxt_c_6__N_498[3] ;
    input n5079;
    output \rd_addr_nxt_c_6__N_498[2] ;
    output n49;
    output n17;
    output \REG.mem_6_14 ;
    output \REG.mem_7_14 ;
    output \REG.mem_4_14 ;
    output \REG.mem_5_14 ;
    output n24;
    input n5078;
    output \REG.mem_3_6 ;
    input n5077;
    output \REG.mem_10_1 ;
    input n5076;
    input n5075;
    output \REG.mem_3_9 ;
    input n5074;
    input n5073;
    output n55;
    output n23;
    output n40;
    output n8;
    input n5072;
    output \REG.mem_9_12 ;
    output n34;
    input n5071;
    input n5070;
    output \REG.mem_9_10 ;
    input n5069;
    output n2;
    input n5068;
    input n5067;
    input n5066;
    input n5065;
    output \REG.mem_9_5 ;
    input n5064;
    input n5063;
    input n5062;
    input n5061;
    output \REG.mem_9_1 ;
    input n5060;
    input n5059;
    input n5058;
    input n5057;
    input n5056;
    output \REG.mem_8_12 ;
    input n5055;
    input n5054;
    output \REG.mem_8_10 ;
    input n5053;
    input n5052;
    input n5051;
    input n5050;
    input n5049;
    output \REG.mem_8_5 ;
    input n5048;
    input n5047;
    input n5046;
    input n5045;
    output \REG.mem_8_1 ;
    input n5044;
    input n5043;
    input n5042;
    input n5041;
    output \REG.mem_7_13 ;
    input n5040;
    output \REG.mem_7_12 ;
    input n5039;
    input n5038;
    output \REG.mem_7_10 ;
    input n5037;
    input n5036;
    input n5035;
    output \REG.mem_7_7 ;
    input n5034;
    output \REG.mem_7_6 ;
    input n5033;
    input n5032;
    input n5031;
    input n5030;
    input n5029;
    input n5028;
    input n5027;
    input n5026;
    input n5025;
    output \REG.mem_6_13 ;
    input n5024;
    output \REG.mem_6_12 ;
    input n5023;
    input n5022;
    output \REG.mem_6_10 ;
    input n5021;
    input n5020;
    input n5019;
    output \REG.mem_6_7 ;
    input n5018;
    output \REG.mem_6_6 ;
    input n5017;
    input n5016;
    input n5015;
    input n5014;
    input n5013;
    input n5012;
    input n5011;
    input n5010;
    input n5009;
    output \REG.mem_5_13 ;
    input n5008;
    output \REG.mem_5_12 ;
    input n5007;
    input n5006;
    output \REG.mem_5_10 ;
    input n5005;
    input n5004;
    input n5003;
    output \REG.mem_5_7 ;
    input n5002;
    output \REG.mem_5_6 ;
    input n5001;
    input n5000;
    input n4999;
    input n4998;
    input n4997;
    input n4996;
    input n4995;
    input n4994;
    input n4993;
    output \REG.mem_4_13 ;
    input n4992;
    output \REG.mem_4_12 ;
    input n4991;
    input n4990;
    output \REG.mem_4_10 ;
    input n4989;
    input n4988;
    input n4987;
    output \REG.mem_4_7 ;
    input n4986;
    output \REG.mem_4_6 ;
    input n4985;
    input n4984;
    input n4983;
    input n4982;
    input n4981;
    input n4980;
    input n4979;
    input n4978;
    input n4977;
    output \REG.mem_3_13 ;
    input n4976;
    input n4975;
    input n4974;
    output \REG.mem_3_10 ;
    input n4973;
    input n4972;
    output \REG.mem_3_8 ;
    input n4971;
    output \REG.mem_3_7 ;
    input n4970;
    input n4969;
    output FT_OE_N_420;
    output n57;
    output n25;
    output n42;
    output n10;
    output n58;
    output n26;
    output n43;
    output n35;
    output n11;
    output n3;
    input n4968;
    input n4967;
    input n4966;
    input n4965;
    input n4964;
    output n60;
    output n28;
    output n59;
    output n27;
    output n61;
    output n29;
    output n4672;
    output n4671;
    output n4670;
    output n4669;
    output n4668;
    output n4667;
    output n4666;
    output n4665;
    output n4664;
    output n4663;
    output n4662;
    output n4661;
    output n4660;
    output n4659;
    output n4658;
    
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [6:0]rd_addr_r;   // src/fifo_dc_32_lut_gen.v(217[29:38])
    
    wire n11123, n12192, n12567, \afull_flag_impl.af_flag_nxt_w , n11048, 
        n10961, n11555, n12255, \REG.mem_17_7 , n12258, n11316, 
        n11317, n13161, n11296, n11295, n11434, n12129, \REG.mem_26_5 , 
        \REG.mem_27_5 , n13155, n4950, \REG.mem_2_2 , n40_c;
    wire [6:0]wr_addr_r;   // src/fifo_dc_32_lut_gen.v(196[29:38])
    
    wire \REG.mem_1_7 , n4905, n12561, \REG.mem_24_5 , n13158, n12678, 
        n12402, n11229, full_nxt_c_N_626, full_o, n12216, n13476, 
        n11230, n13140, n13080, n11233;
    wire [31:0]\REG.out_raw_31__N_559 ;
    
    wire n11388, n11389, n13149, n11386, n11385, n11437, n12564, 
        n4949, \REG.mem_2_1 , n12510, n10864, n12555, n10861, n10860, 
        n12558, \REG.mem_56_15 , n11766, \REG.mem_58_15 , \REG.mem_59_15 , 
        n11767, n11776, \REG.mem_60_15 , \REG.mem_61_15 , n11775, 
        n4948, \REG.mem_2_0 , n13143, n11081, \REG.mem_58_1 , \REG.mem_59_1 , 
        n12549, \REG.mem_56_1 , n12552, n11700, n11701, n12543, 
        n4947, \REG.mem_0_0 , \REG.mem_26_9 , \REG.mem_27_9 , n13137, 
        \REG.mem_24_9 , n11615, n11618, n12249, \REG.mem_1_6 , n4914, 
        n11698, n11697, n12546, n11606, n11594, n11796, n11797, 
        n12537, n11791, n11790, n12540, \REG.mem_1_15 , n4832, n13131, 
        n10955, n11757, n11758, n12531, n11755, n11754, n12534, 
        n13125, \REG.mem_51_11 , n12525, \REG.mem_49_11 , n11561, 
        \REG.mem_1_5 , n4835, n12519, n12522, \REG.mem_1_4 , n4837, 
        n11565, n11566, n12513, \REG.mem_53_13 , \REG.mem_52_13 , 
        n13128, \REG.mem_1_3 , n4861, \REG.mem_1_2 , n4868, n11545, 
        n11544, n12516, \REG.mem_58_6 , \REG.mem_59_6 , n13119;
    wire [6:0]rd_grey_w;   // src/fifo_dc_32_lut_gen.v(224[38:47])
    
    wire \REG.mem_56_6 , n11444, n4946, \REG.mem_0_1 , n11727, n11728, 
        n12507, n11686, n11685, n11532, n11533, n12501, empty_nxt_c_N_629, 
        n11488, n11487, n12504, n11382, n11383, n13113, n11362, 
        n11361, n11446;
    wire [6:0]wr_grey_w;   // src/fifo_dc_32_lut_gen.v(203[38:47])
    
    wire \REG.mem_1_1 , n4879, n4944, \REG.mem_0_2 , n12495, n4943, 
        \REG.mem_0_3 , \REG.mem_53_11 , \REG.mem_52_11 , n11570, n13107, 
        n12489, n13110, \REG.mem_29_0 , \REG.mem_28_0 , n12492, \REG.mem_0_5 , 
        n10887, \REG.mem_2_5 , n10888, n10924, n10923, \REG.mem_58_11 , 
        \REG.mem_59_11 , n12483, n12948, n13101, n11413, n12936, 
        n13104, \REG.mem_56_11 , n11573, n20_c, n12477, n13095, 
        \REG.mem_61_13 , \REG.mem_60_13 , n12480, n13098, \REG.mem_1_0 , 
        n4884, \REG.mem_2_11 , n13089, \REG.mem_1_11 , \REG.mem_0_11 , 
        n11459, n11315, n11336, n12471, n11258, n11219, n11579, 
        n13083, n12132, \REG.mem_19_5 , n12135, n12465, n12123, 
        \REG.mem_61_1 , \REG.mem_60_1 , n12468, n11462, \REG.mem_1_8 , 
        n4900, n12459, n12462, n13077;
    wire [6:0]wr_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(200[30:42])
    
    wire wr_sig_mv_w, \REG.mem_29_9 , \REG.mem_28_9 , n12453, n11022, 
        n11023, n13071, n12456;
    wire [6:0]n1;
    
    wire n11020, n11019, n11101, n12447, \REG.mem_61_11 , \REG.mem_60_11 , 
        n11588, \REG.mem_56_8 , n11721, n13065, \REG.mem_58_8 , \REG.mem_59_8 , 
        n11722, n11785, \REG.mem_60_8 , \REG.mem_61_8 , n11784, \REG.mem_61_6 , 
        \REG.mem_60_6 , n11465, \REG.mem_34_0 , n12441, \REG.mem_33_0 , 
        \REG.mem_32_0 , n11171, \REG.mem_26_15 , \REG.mem_27_15 , n12435, 
        \REG.mem_24_15 , n12438, n12954, n13059, n12942, n13062, 
        \REG.mem_32_7 , \REG.mem_33_7 , n11262, \REG.mem_34_7 , n11263, 
        \REG.mem_34_9 , n13053, \REG.mem_33_9 , \REG.mem_32_9 , n13056, 
        n11049, n11050, n13047, n10919, n10928, n12429, n10916, 
        n10910, n10988, n11474, n11483, n12423, n11044, n11043, 
        n11107, \REG.mem_19_12 , n13041, n10844, n10847, n12417, 
        n11867, n11861, n12420, \REG.mem_17_12 , n13044, n12411, 
        n12414, n13731, n13734, n11281, n11070, n11071, n13035, 
        n11280, \REG.mem_51_12 , n12405, n11068, n11067, n11110, 
        \REG.mem_49_12 , n12408, n13725, n12399, \REG.mem_61_9 , \REG.mem_60_9 , 
        n13728, \REG.mem_34_6 , n13719, n12126, \REG.mem_33_6 , \REG.mem_32_6 , 
        n12393, n12396, n13713, n13029, \REG.mem_21_7 , \REG.mem_20_7 , 
        n13716, n10940, n12387, \REG.mem_2_15 , n13023, n13707, 
        n13710, \REG.mem_0_15 , n13026, n4935, \REG.mem_0_4 , n13701, 
        n13704, n10937, n10931, n10997, n12117, n12159, \REG.mem_61_12 , 
        \REG.mem_60_12 , n12162, n11633, n12153, n12231, n12147, 
        \REG.mem_56_9 , n12150, \REG.mem_58_14 , \REG.mem_59_14 , n13695, 
        \REG.mem_56_14 , n11091, n11092, n13017, n12381, \REG.mem_29_15 , 
        \REG.mem_28_15 , n12384, n12141, \REG.mem_17_5 , n12138, n11089, 
        n11088, n11113, n12120, \REG.mem_19_8 , n13689, n11507, 
        n11519, n12375, n39, \REG.mem_17_15 , n5210, \REG.mem_17_8 , 
        n13692, n11510, n11504, n11495, n13011, \REG.mem_26_2 , 
        \REG.mem_27_2 , n13683, \REG.mem_21_12 , \REG.mem_20_12 , n13014, 
        \REG.mem_24_2 , n13686, n13677, n10976, n10979, n12369, 
        n10970, n10964, n11000, \REG.mem_17_14 , n5209, \REG.mem_49_10 , 
        n11367, \REG.mem_51_10 , n11368, \REG.mem_29_2 , \REG.mem_28_2 , 
        n13680, n13662, \REG.mem_17_13 , n5208, n11371, \REG.mem_52_10 , 
        \REG.mem_53_10 , n11370, n12756, n12870, n13005, n5207, 
        n12363, n11709, n11710, n13671, \REG.mem_53_12 , \REG.mem_52_12 , 
        n12366, n11707, n11706, n10876, n12912, n13386, \REG.mem_34_15 , 
        n12357, n13665, n12966, \REG.mem_58_13 , \REG.mem_59_13 , 
        n12999, \REG.mem_33_15 , \REG.mem_32_15 , n12360, n12672, 
        n13224, \REG.mem_17_11 , n5206, n12858, n13656, \REG.mem_56_13 , 
        n13002, \REG.mem_17_10 , n5205, n10873, n13659, n11543, 
        n11552, n12351, n11528, n11525, \REG.mem_17_9 , n5204, n5203, 
        n12960, n5202, n10870, \REG.mem_17_6 , n5201, n5200, n12993, 
        \REG.mem_17_4 , n5199, n11250, n11251, n13653, \REG.mem_17_3 , 
        n5198, \REG.mem_29_13 , \REG.mem_28_13 , n12996, \REG.mem_17_2 , 
        n5197, \REG.mem_17_1 , n5196, \REG.mem_17_0 , n5195, n43_c, 
        \REG.mem_19_15 , n5242, n11242, n11241, \REG.mem_19_14 , n5241, 
        n13398, n13608, \REG.mem_53_9 , \REG.mem_52_9 , n12234, n12684, 
        n12780, n10967, \REG.mem_19_13 , n5240, n11035, n4934, n12726, 
        n12606, n13434, n12345, n4933, \REG.mem_0_6 , n13170, n13647, 
        n5239, n13326, n13392, n11753, n12987, \REG.mem_19_11 , 
        n5238, n10982, \REG.mem_19_10 , n5237, \REG.mem_19_9 , n5236, 
        n5235, \REG.mem_19_7 , n5234, \REG.mem_19_6 , n5233, \REG.mem_49_7 , 
        n11325, \REG.mem_51_7 , n11326, n11356, \REG.mem_52_7 , \REG.mem_53_7 , 
        n11355, n5232, n13602, n13641, \REG.mem_19_4 , n5231, \REG.mem_19_3 , 
        n5230, \REG.mem_29_5 , \REG.mem_28_5 , n12990, \REG.mem_19_2 , 
        n5229, \REG.mem_19_1 , n5228, \REG.mem_19_0 , n5227, n45, 
        \REG.mem_20_15 , n5258, n13182, n13470, n11762, \REG.mem_20_14 , 
        n5257, n12339, \REG.mem_34_13 , n12981, \REG.mem_2_3 , n13635, 
        \REG.mem_33_13 , \REG.mem_32_13 , n12984, \REG.mem_49_15 , n5749, 
        n10886;
    wire [6:0]wp_sync2_r;   // src/fifo_dc_32_lut_gen.v(223[37:47])
    wire [6:0]wp_sync_w;   // src/fifo_dc_32_lut_gen.v(226[30:39])
    
    wire \REG.mem_49_14 , n5748, \REG.mem_51_1 , n12975, n13629, \REG.mem_49_13 , 
        n5747, n12708, n12630, n11748, \REG.mem_49_1 , n12978, \REG.mem_61_14 , 
        \REG.mem_60_14 , n11749, n12969, n12270, n11770, \REG.mem_20_13 , 
        n5256, n13623, n11769, n5255, n11418, n11419, n12963, 
        n10892, n11404, n12924, n13617, n13620, \REG.mem_20_11 , 
        n5254, \REG.mem_20_10 , n5253, n5746, n12930, n11410, n12957, 
        n5745, \REG.mem_20_9 , n5252, n13611, n11401, n12918, n13614, 
        n12327, n5744, \REG.mem_20_8 , n5251, n13605, \REG.mem_49_9 , 
        n5743, n4932, \REG.mem_0_7 , n5250, n12828, n12330, n12951, 
        \REG.mem_26_13 , \REG.mem_27_13 , n13599, \REG.mem_20_6 , n5249, 
        \REG.mem_20_5 , n5248, \REG.mem_20_4 , n5247, \REG.mem_49_8 , 
        n5742, \REG.mem_20_3 , n5246, n5741, \REG.mem_49_6 , n5740, 
        \REG.mem_20_2 , n5245, \REG.mem_49_5 , n5739, n12945, \REG.mem_24_13 , 
        n6033, \REG.mem_20_1 , n5244, n6031, n4931, \REG.mem_0_8 , 
        n13593, \REG.mem_20_0 , n5243, n47_c, \REG.mem_21_15 , n5274, 
        n10895, n12939, \REG.mem_21_14 , n5273, \REG.mem_21_13 , n5272, 
        n5271, \REG.mem_21_11 , n5270, \REG.mem_51_9 , n12309, \REG.mem_21_10 , 
        n5269, n4930, \REG.mem_0_9 , n12312, n13587, \REG.mem_21_9 , 
        n5268, \REG.mem_21_8 , n5267, n12303, n5266, \REG.mem_21_6 , 
        n5265, n4929, \REG.mem_0_10 , n4928, \REG.mem_21_5 , n5264, 
        \REG.mem_21_4 , n5263, n11291, n11340, n11341, n12933, n11329, 
        n11328, \REG.mem_21_3 , n5262, n11183, n13581, n11301, n11302, 
        n12927, n12294, n11807, n12297, n12300, n5979, n5978, 
        n5977, n5976, n5975, n5974, \REG.mem_61_10 , n5973, n5972, 
        n5971, \REG.mem_61_7 , n5970, n5969, \REG.mem_61_5 , n10853, 
        n11299, n11298, \REG.mem_21_2 , n5261, \REG.mem_21_1 , n5260, 
        n12291, \REG.mem_21_0 , n5259, n13575, n11094, n11095, n12921, 
        n53_c, n5328, n11053, n11052, \REG.mem_24_14 , n5327, \REG.mem_49_4 , 
        n5738, n11274, n11275, n12915, n5968, \REG.mem_61_4 , n5967, 
        \REG.mem_61_3 , n5966, \REG.mem_61_2 , n5965, n5964, \REG.mem_61_0 , 
        n5962, n5961, n5960, n5959, n5958, n5957, \REG.mem_60_10 , 
        n5956, n5955, n5954, \REG.mem_60_7 , n5953, n13578, n11266, 
        n11265, n5952, \REG.mem_60_5 , n5951, \REG.mem_60_4 , n5950, 
        \REG.mem_60_3 , n5949, \REG.mem_60_2 , n5948, n5947, \REG.mem_60_0 ;
    wire [6:0]rp_sync2_r;   // src/fifo_dc_32_lut_gen.v(202[37:47])
    
    wire n5937, n5326, \REG.mem_24_12 , n5325, n13569, n5936, n12804, 
        n11789, n12816, n5935, n5934, \REG.mem_59_12 , n5933, n5932, 
        \REG.mem_59_10 , n5931, \REG.mem_59_9 , n5930, n5929, \REG.mem_59_7 , 
        n5928, n5927, \REG.mem_59_5 , n5926, \REG.mem_59_4 , n5925, 
        \REG.mem_59_3 , n5924, \REG.mem_59_2 , n5923, n5922, \REG.mem_59_0 , 
        n5918, n4927, \REG.mem_0_12 , n12720, \REG.mem_26_1 , \REG.mem_27_1 , 
        n13563, n5915, n5913, n5912, n5911, n5910, n5909, \REG.mem_58_12 , 
        n5908, n5907, \REG.mem_58_10 , n5906, \REG.mem_58_9 , n5905, 
        n5904, \REG.mem_58_7 , n5903, n5902, \REG.mem_58_5 , n11322, 
        n11323, n12909, n13548, n13524, \REG.mem_24_11 , n5324, 
        \REG.mem_49_3 , n5737, n12285, \REG.mem_24_1 , n13566, \REG.mem_24_10 , 
        n5323, n5901, \REG.mem_58_4 , n5900, \REG.mem_58_3 , n5899, 
        \REG.mem_58_2 , n5898, n5897, \REG.mem_58_0 , n5322, \REG.mem_24_8 , 
        n5321, n11311, n12888, n11396, n11381, n13557, n12279, 
        n13560, \REG.mem_24_7 , n5320, n5878, n5877, n5876, n5875, 
        \REG.mem_56_12 , n5874, n5873, \REG.mem_56_10 , n5872, n5871, 
        n5870, \REG.mem_56_7 , n5869, \REG.mem_56_4 , n11253, n11254, 
        n12903, n12282, n5868, \REG.mem_56_5 , n5867, n5866, \REG.mem_56_3 , 
        n5865, \REG.mem_56_2 , n5864, n5862, \REG.mem_56_0 , n10009, 
        n10010, n10008, n10007, n9962, n9963, n10006, n10005;
    wire [6:0]rd_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(221[30:42])
    
    wire n10016, n10015;
    wire [6:0]n1_adj_1212;
    
    wire n9973, n10828;
    wire [6:0]rp_sync_w;   // src/fifo_dc_32_lut_gen.v(205[30:39])
    
    wire n9972, n10798, n10014, n10778, n9971, n2_adj_1188;
    wire [6:0]wr_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(212[30:44])
    
    wire n9970, n11236, n11235, n12906, n5816, \REG.mem_53_15 , 
        n5815, \REG.mem_53_14 , n5814, n5813, n5812, n5811, n5810, 
        n5809, \REG.mem_53_8 , n5808, n5807, \REG.mem_53_6 , n5806, 
        \REG.mem_53_5 , n5805, \REG.mem_53_4 , n5472, \REG.mem_24_4 , 
        n10013, \REG.mem_26_4 , \REG.mem_27_4 , n5804, \REG.mem_53_3 , 
        n5803, \REG.mem_53_2 , n5802, \REG.mem_53_1 , n5801, \REG.mem_53_0 , 
        n5800, \REG.mem_52_15 , n5799, \REG.mem_52_14 , n5798, n5797, 
        n5796, n5795, n5794, n5793, \REG.mem_52_8 , n5792, n5791, 
        \REG.mem_52_6 , n5790, \REG.mem_52_5 , n5789, \REG.mem_52_4 , 
        \REG.mem_24_6 , n5319, \REG.mem_28_4 , \REG.mem_29_4 , n9969, 
        n5788, \REG.mem_52_3 , n5787, \REG.mem_52_2 , n5786, \REG.mem_52_1 , 
        n5785, \REG.mem_52_0 , n5784, \REG.mem_51_15 , n5783, \REG.mem_51_14 , 
        n5782, \REG.mem_51_13 , n5781, n5780, n5779, n5778, n5777, 
        \REG.mem_51_8 , n5776, n5775, \REG.mem_51_6 , n5774, \REG.mem_51_5 , 
        n5773, \REG.mem_51_4 , n9968, n10012, n5772, \REG.mem_51_3 , 
        n5771, \REG.mem_51_2 , n5770, n5769, \REG.mem_51_0 , n9967;
    wire [6:0]rd_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(233[30:44])
    
    wire n9966, n5318, n10011, n5317, n12273, n5736, \REG.mem_49_2 , 
        n5735, n5734, \REG.mem_49_0 , \REG.mem_24_3 , n5316, n9965, 
        n4926, \REG.mem_0_13 , n4925, \REG.mem_0_14 , n13551, \REG.mem_26_12 , 
        \REG.mem_27_12 , n12897, n12900, n4924, n12276, n13545, 
        n5315, n5314, \REG.mem_24_0 , n5307, n12267, n57_c, n5360, 
        n12891, n12261, n12894, n5669, n11006, \REG.mem_26_14 , 
        n5359, n5358, n5357, n13539, \REG.mem_26_11 , n5356, n10900, 
        n9964, \REG.mem_26_10 , n5355, n5354, \REG.mem_26_8 , n5353, 
        \REG.mem_26_7 , n5352, \genblk16.rd_prev_r , n11153, n12174, 
        n12219, \REG.mem_26_6 , n5351, n13533, n12885, n5350, n12879, 
        n4915, n5349, \REG.mem_27_6 , n12873, n13527, n10903, \REG.mem_26_3 , 
        n5348, n4912, \REG.mem_1_12 , \REG.mem_33_14 , n5471, n5347, 
        n5346, n4902, \REG.mem_1_13 , \REG.mem_26_0 , n5345, n5470, 
        n12222, n59_c, n5376, n6_adj_1189, \REG.mem_27_14 , n5375, 
        n13521, n10126, n12750, n12867, \REG.mem_2_4 , n12165, n5374, 
        n12744, n5373, \REG.mem_27_11 , n5372, n13515, n12861, \REG.mem_27_10 , 
        n5371, n5370, n13518, \REG.mem_27_8 , n5369, \REG.mem_27_7 , 
        n5368, n5367, n5366, n5365, \REG.mem_27_3 , n5364, n12168, 
        n5363, n5362, \REG.mem_33_12 , n5469, \REG.mem_27_0 , n5361, 
        n61_c, n5392, \REG.mem_28_14 , n5391, n5390, \REG.mem_28_12 , 
        n5389, \REG.mem_28_11 , n5388, \REG.mem_28_10 , n5387, n5386, 
        \REG.mem_28_8 , n5385, \REG.mem_28_7 , n5384, \REG.mem_28_6 , 
        n5383, n5382, n5488, n5487, \REG.mem_34_14 , n5486, n5485, 
        \REG.mem_34_12 , n5484, \REG.mem_34_11 , n5381, n13509, n13512, 
        n5483, \REG.mem_34_10 , n5482, n5481, \REG.mem_34_8 , n5480, 
        n5479, n5478, \REG.mem_34_5 , n5477, \REG.mem_34_4 , n5476, 
        \REG.mem_34_3 , n5475, \REG.mem_34_2 , n5474, \REG.mem_34_1 , 
        n5473, n5468, \REG.mem_33_11 , n12840, n12855, \REG.mem_28_3 , 
        n5380, n13503, n5467, \REG.mem_33_10 , n5466, n5465, \REG.mem_33_8 , 
        n5464, n5463, n5462, \REG.mem_33_5 , n5461, \REG.mem_33_4 , 
        n5460, \REG.mem_33_3 , n5459, \REG.mem_33_2 , n5458, \REG.mem_33_1 , 
        n5457, n5456, n5455, \REG.mem_32_14 , n5454, n5453, \REG.mem_32_12 , 
        n5379, \REG.mem_28_1 , n5378, n5377, n5452, \REG.mem_32_11 , 
        n63, n5408, n5451, \REG.mem_32_10 , n5450, n5449, \REG.mem_32_8 , 
        n5448, n5447, n5446, \REG.mem_32_5 , n5445, \REG.mem_32_4 , 
        n5444, \REG.mem_32_3 , n5443, \REG.mem_32_2 , n5442, \REG.mem_32_1 , 
        n5441, n10946, n12849, n11876, n11864, n11819, \REG.mem_29_14 , 
        n5407, n5406, \REG.mem_29_12 , n5405, \REG.mem_29_11 , n5404, 
        \REG.mem_29_10 , n5403, n13497, n11333, n5402, n12843, n12111, 
        \REG.mem_29_8 , n5401, \REG.mem_29_7 , n5400, \REG.mem_29_6 , 
        n5399, n5398, n5397, \REG.mem_29_3 , n5396, n5395, \REG.mem_29_1 , 
        n5394, n12213, n5393, n13491, n38, n11061, n11062, n12837, 
        n13485, n13488, n11038, n11037, n13479, n23_c, n13482, 
        n13473, n12831, n12834, n12825, n13467, n15_c, n12819, 
        n13461, n11828, n42_c, n12822, n13455, n12813, n4274, 
        n10772, n10907, n12807, n13449, n13452, n10722, n4298, 
        n10_c, n8_adj_1191, n12, n12801, n10766, n10838, n10130, 
        n4963, n13443, n11351, n12795, n13437;
    wire [6:0]rd_addr_nxt_c_6__N_498;
    
    wire \REG.mem_2_14 , n4962, \REG.mem_2_13 , n4961, \REG.mem_2_12 , 
        n4960, n4959, \REG.mem_2_10 , n4958, \REG.mem_2_9 , n4957, 
        n12600, n13431, \REG.mem_2_8 , n4956, \REG.mem_2_7 , n4955, 
        \REG.mem_2_6 , n4954, n12789, n10879, n10878, n4953, n12114, 
        n12783, n13425, n13428, n13242, n12210, n13419, n11847, 
        n11848, n12777, n12207, n11834, n12201, n11842, n11841, 
        n13413, n4952, n12771, n11283, n11284, n13407, n12774, 
        n11272, n11271, n11365, n4951, n13401, n12765, n11840, 
        n11736, n11737, n13395, n11725, n11724, n12768, n13206, 
        n13389, n12576, n12759, n12588, n12654, n12762, n18_c, 
        n13383, n11344, n11343, n35_c, n12738, n12753, n13377, 
        n11100, n11085, n11086, n12747, n13371, n11077, n11076, 
        n12204, n11064, n11065, n12741, n11059, n11058, n13365, 
        n11846, \REG.mem_1_14 , n13359, n13344, n13362, n12195, 
        n11040, n11041, n12735, n13, n11029, n11028, n12198, n13353, 
        n12729, n13188, n12732, n14, n12636, n10921, n12723, n12717, 
        n12189, n33, n13347, n12711, n12714, n13341, n4867, n4866, 
        n13335, n12705, n13329, n11690, n13323, n12699, n13317, 
        n11286, n11287, n13311, n11278, n11277, n12693, n13305, 
        n11835, n11836, n12681, n11830, n11829, n11268, n11269, 
        n13299, n11239, n11238, n13302, n12675, n11763, n11764, 
        n13293, n11740, n11739, \REG.mem_1_9 , n11_c, n11871, n11872, 
        n12669, n11854, n11853, n12_adj_1199, n13287, n12663, n11811, 
        n11812, n13281, n36, n12657, n12660, n11794, n11793, n13284, 
        n12144, n13275, n12651, n13269, \REG.mem_1_10 , n13263, 
        full_max_w, n10760, n10724, n12_adj_1201, n10746, n10736, 
        n11883, n10744, n10836, n12645, n13266, n4833, n12639, 
        n13257, n11319, n11320, n13251, n11308, n11307, n4831, 
        n13245, n11718, n11719, n12633, n11716, n11715, n13239, 
        n12627, n9, n13233, n12621, n34_adj_1205, n13227, n13230, 
        n12615, n12594, n13221, n12618, n10855, n12609, n11358, 
        n11359, n13215, n11696, n11347, n11346, n10867, n12603, 
        n11800, n11799, n13209, n13203, n11742, n11743, n12597, 
        n11731, n11730, n11247, n11248, n13197, n11227, n11226, 
        n11712, n11713, n12591, n11704, n11703, n12171, n12585, 
        n13191, n13194, n12579, n13185, n13179, n13173, n12573, 
        n13176, n13167, n11689, n11695;
    
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10698 (.I0(rd_addr_r[2]), .I1(n11123), 
            .I2(n12192), .I3(rd_addr_r[3]), .O(n12567));
    defparam rd_addr_r_2__bdd_4_lut_10698.LUT_INIT = 16'he4aa;
    SB_DFFSR \afull_flag_impl.af_flag_ext_r_121  (.Q(dc32_fifo_almost_full), 
            .C(FIFO_CLK_c), .D(\afull_flag_impl.af_flag_nxt_w ), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    SB_LUT4 n12567_bdd_4_lut (.I0(n12567), .I1(n11048), .I2(n10961), .I3(rd_addr_r[3]), 
            .O(n11555));
    defparam n12567_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12255_bdd_4_lut (.I0(n12255), .I1(\REG.mem_17_7 ), .I2(\REG.mem_16_7 ), 
            .I3(rd_addr_r[1]), .O(n12258));
    defparam n12255_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11162 (.I0(rd_addr_r[1]), .I1(n11316), 
            .I2(n11317), .I3(rd_addr_r[2]), .O(n13161));
    defparam rd_addr_r_1__bdd_4_lut_11162.LUT_INIT = 16'he4aa;
    SB_LUT4 n13161_bdd_4_lut (.I0(n13161), .I1(n11296), .I2(n11295), .I3(rd_addr_r[2]), 
            .O(n11434));
    defparam n13161_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10283 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_6_2 ), 
            .I2(\REG.mem_7_2 ), .I3(rd_addr_r[1]), .O(n12129));
    defparam rd_addr_r_0__bdd_4_lut_10283.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11137 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_26_5 ), 
            .I2(\REG.mem_27_5 ), .I3(rd_addr_r[1]), .O(n13155));
    defparam rd_addr_r_0__bdd_4_lut_11137.LUT_INIT = 16'he4aa;
    SB_DFF i236_237 (.Q(\REG.mem_2_2 ), .C(FIFO_CLK_c), .D(n4950));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3522_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_1_7 ), .O(n4905));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3522_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10643 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_46_9 ), 
            .I2(\REG.mem_47_9 ), .I3(rd_addr_r[1]), .O(n12561));
    defparam rd_addr_r_0__bdd_4_lut_10643.LUT_INIT = 16'he4aa;
    SB_LUT4 n13155_bdd_4_lut (.I0(n13155), .I1(\REG.mem_25_5 ), .I2(\REG.mem_24_5 ), 
            .I3(rd_addr_r[1]), .O(n13158));
    defparam n13155_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9379_3_lut (.I0(n12678), .I1(n12402), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11229));
    defparam i9379_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR full_ext_r_117 (.Q(full_o), .C(FIFO_CLK_c), .D(full_nxt_c_N_626), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 i9380_3_lut (.I0(n12216), .I1(n13476), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11230));
    defparam i9380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9383_3_lut (.I0(n13140), .I1(n13080), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11233));
    defparam i9383_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE \REG.out_raw__i1  (.Q(\REG.out_raw[0] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [0]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11132 (.I0(rd_addr_r[1]), .I1(n11388), 
            .I2(n11389), .I3(rd_addr_r[2]), .O(n13149));
    defparam rd_addr_r_1__bdd_4_lut_11132.LUT_INIT = 16'he4aa;
    SB_LUT4 n13149_bdd_4_lut (.I0(n13149), .I1(n11386), .I2(n11385), .I3(rd_addr_r[2]), 
            .O(n11437));
    defparam n13149_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12561_bdd_4_lut (.I0(n12561), .I1(\REG.mem_45_9 ), .I2(\REG.mem_44_9 ), 
            .I3(rd_addr_r[1]), .O(n12564));
    defparam n12561_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i233_234 (.Q(\REG.mem_2_1 ), .C(FIFO_CLK_c), .D(n4949));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10668 (.I0(rd_addr_r[3]), .I1(n12510), 
            .I2(n10864), .I3(rd_addr_r[4]), .O(n12555));
    defparam rd_addr_r_3__bdd_4_lut_10668.LUT_INIT = 16'he4aa;
    SB_LUT4 n12555_bdd_4_lut (.I0(n12555), .I1(n10861), .I2(n10860), .I3(rd_addr_r[4]), 
            .O(n12558));
    defparam n12555_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9916_3_lut (.I0(\REG.mem_56_15 ), .I1(\REG.mem_57_15 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11766));
    defparam i9916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9917_3_lut (.I0(\REG.mem_58_15 ), .I1(\REG.mem_59_15 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11767));
    defparam i9917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9926_3_lut (.I0(\REG.mem_62_15 ), .I1(\REG.mem_63_15 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11776));
    defparam i9926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9925_3_lut (.I0(\REG.mem_60_15 ), .I1(\REG.mem_61_15 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11775));
    defparam i9925_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i230_231 (.Q(\REG.mem_2_0 ), .C(FIFO_CLK_c), .D(n4948));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11127 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_6_1 ), 
            .I2(\REG.mem_7_1 ), .I3(rd_addr_r[1]), .O(n13143));
    defparam rd_addr_r_0__bdd_4_lut_11127.LUT_INIT = 16'he4aa;
    SB_LUT4 n13143_bdd_4_lut (.I0(n13143), .I1(\REG.mem_5_1 ), .I2(\REG.mem_4_1 ), 
            .I3(rd_addr_r[1]), .O(n11081));
    defparam n13143_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10633 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_58_1 ), 
            .I2(\REG.mem_59_1 ), .I3(rd_addr_r[1]), .O(n12549));
    defparam rd_addr_r_0__bdd_4_lut_10633.LUT_INIT = 16'he4aa;
    SB_LUT4 n12549_bdd_4_lut (.I0(n12549), .I1(\REG.mem_57_1 ), .I2(\REG.mem_56_1 ), 
            .I3(rd_addr_r[1]), .O(n12552));
    defparam n12549_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10658 (.I0(rd_addr_r[1]), .I1(n11700), 
            .I2(n11701), .I3(rd_addr_r[2]), .O(n12543));
    defparam rd_addr_r_1__bdd_4_lut_10658.LUT_INIT = 16'he4aa;
    SB_DFF i38_39 (.Q(\REG.mem_0_0 ), .C(FIFO_CLK_c), .D(n4947));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11117 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_26_9 ), 
            .I2(\REG.mem_27_9 ), .I3(rd_addr_r[1]), .O(n13137));
    defparam rd_addr_r_0__bdd_4_lut_11117.LUT_INIT = 16'he4aa;
    SB_LUT4 n13137_bdd_4_lut (.I0(n13137), .I1(\REG.mem_25_9 ), .I2(\REG.mem_24_9 ), 
            .I3(rd_addr_r[1]), .O(n13140));
    defparam n13137_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10455 (.I0(rd_addr_r[4]), .I1(n11615), 
            .I2(n11618), .I3(rd_addr_r[5]), .O(n12249));
    defparam rd_addr_r_4__bdd_4_lut_10455.LUT_INIT = 16'he4aa;
    SB_LUT4 i3531_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_1_6 ), .O(n4914));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3531_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12543_bdd_4_lut (.I0(n12543), .I1(n11698), .I2(n11697), .I3(rd_addr_r[2]), 
            .O(n12546));
    defparam n12543_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12249_bdd_4_lut (.I0(n12249), .I1(n11606), .I2(n11594), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_559 [11]));
    defparam n12249_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10619 (.I0(rd_addr_r[1]), .I1(n11796), 
            .I2(n11797), .I3(rd_addr_r[2]), .O(n12537));
    defparam rd_addr_r_1__bdd_4_lut_10619.LUT_INIT = 16'he4aa;
    SB_LUT4 n12537_bdd_4_lut (.I0(n12537), .I1(n11791), .I2(n11790), .I3(rd_addr_r[2]), 
            .O(n12540));
    defparam n12537_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3449_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_1_15 ), .O(n4832));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3449_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11112 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_46_3 ), 
            .I2(\REG.mem_47_3 ), .I3(rd_addr_r[1]), .O(n13131));
    defparam rd_addr_r_0__bdd_4_lut_11112.LUT_INIT = 16'he4aa;
    SB_LUT4 n13131_bdd_4_lut (.I0(n13131), .I1(\REG.mem_45_3 ), .I2(\REG.mem_44_3 ), 
            .I3(rd_addr_r[1]), .O(n10955));
    defparam n13131_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10614 (.I0(rd_addr_r[1]), .I1(n11757), 
            .I2(n11758), .I3(rd_addr_r[2]), .O(n12531));
    defparam rd_addr_r_1__bdd_4_lut_10614.LUT_INIT = 16'he4aa;
    SB_LUT4 n12531_bdd_4_lut (.I0(n12531), .I1(n11755), .I2(n11754), .I3(rd_addr_r[2]), 
            .O(n12534));
    defparam n12531_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11107 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_54_13 ), 
            .I2(\REG.mem_55_13 ), .I3(rd_addr_r[1]), .O(n13125));
    defparam rd_addr_r_0__bdd_4_lut_11107.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10624 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_50_11 ), 
            .I2(\REG.mem_51_11 ), .I3(rd_addr_r[1]), .O(n12525));
    defparam rd_addr_r_0__bdd_4_lut_10624.LUT_INIT = 16'he4aa;
    SB_LUT4 n12525_bdd_4_lut (.I0(n12525), .I1(\REG.mem_49_11 ), .I2(\REG.mem_48_11 ), 
            .I3(rd_addr_r[1]), .O(n11561));
    defparam n12525_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3452_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_1_5 ), .O(n4835));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3452_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10604 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_42_12 ), 
            .I2(\REG.mem_43_12 ), .I3(rd_addr_r[1]), .O(n12519));
    defparam rd_addr_r_0__bdd_4_lut_10604.LUT_INIT = 16'he4aa;
    SB_LUT4 n12519_bdd_4_lut (.I0(n12519), .I1(\REG.mem_41_12 ), .I2(\REG.mem_40_12 ), 
            .I3(rd_addr_r[1]), .O(n12522));
    defparam n12519_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3454_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_1_4 ), .O(n4837));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3454_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10609 (.I0(rd_addr_r[1]), .I1(n11565), 
            .I2(n11566), .I3(rd_addr_r[2]), .O(n12513));
    defparam rd_addr_r_1__bdd_4_lut_10609.LUT_INIT = 16'he4aa;
    SB_LUT4 n13125_bdd_4_lut (.I0(n13125), .I1(\REG.mem_53_13 ), .I2(\REG.mem_52_13 ), 
            .I3(rd_addr_r[1]), .O(n13128));
    defparam n13125_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3478_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_1_3 ), .O(n4861));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3478_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3485_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_1_2 ), .O(n4868));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3485_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12513_bdd_4_lut (.I0(n12513), .I1(n11545), .I2(n11544), .I3(rd_addr_r[2]), 
            .O(n12516));
    defparam n12513_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11102 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_58_6 ), 
            .I2(\REG.mem_59_6 ), .I3(rd_addr_r[1]), .O(n13119));
    defparam rd_addr_r_0__bdd_4_lut_11102.LUT_INIT = 16'he4aa;
    SB_DFFSR rd_grey_sync_r__i0 (.Q(\rd_grey_sync_r[0] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[0]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 n13119_bdd_4_lut (.I0(n13119), .I1(\REG.mem_57_6 ), .I2(\REG.mem_56_6 ), 
            .I3(rd_addr_r[1]), .O(n11444));
    defparam n13119_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i41_42 (.Q(\REG.mem_0_1 ), .C(FIFO_CLK_c), .D(n4946));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10594 (.I0(rd_addr_r[1]), .I1(n11727), 
            .I2(n11728), .I3(rd_addr_r[2]), .O(n12507));
    defparam rd_addr_r_1__bdd_4_lut_10594.LUT_INIT = 16'he4aa;
    SB_LUT4 n12507_bdd_4_lut (.I0(n12507), .I1(n11686), .I2(n11685), .I3(rd_addr_r[2]), 
            .O(n12510));
    defparam n12507_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10589 (.I0(rd_addr_r[1]), .I1(n11532), 
            .I2(n11533), .I3(rd_addr_r[2]), .O(n12501));
    defparam rd_addr_r_1__bdd_4_lut_10589.LUT_INIT = 16'he4aa;
    SB_DFFSS empty_ext_r_124 (.Q(DEBUG_3_c), .C(SLM_CLK_c), .D(empty_nxt_c_N_629), 
            .S(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_LUT4 n12501_bdd_4_lut (.I0(n12501), .I1(n11488), .I2(n11487), .I3(rd_addr_r[2]), 
            .O(n12504));
    defparam n12501_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11122 (.I0(rd_addr_r[1]), .I1(n11382), 
            .I2(n11383), .I3(rd_addr_r[2]), .O(n13113));
    defparam rd_addr_r_1__bdd_4_lut_11122.LUT_INIT = 16'he4aa;
    SB_LUT4 n13113_bdd_4_lut (.I0(n13113), .I1(n11362), .I2(n11361), .I3(rd_addr_r[2]), 
            .O(n11446));
    defparam n13113_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR wr_grey_sync_r__i0 (.Q(wr_grey_sync_r[0]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[0]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_LUT4 i3496_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_1_1 ), .O(n4879));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3496_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i44_45 (.Q(\REG.mem_0_2 ), .C(FIFO_CLK_c), .D(n4944));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10599 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_54_11 ), 
            .I2(\REG.mem_55_11 ), .I3(rd_addr_r[1]), .O(n12495));
    defparam rd_addr_r_0__bdd_4_lut_10599.LUT_INIT = 16'he4aa;
    SB_DFF i47_48 (.Q(\REG.mem_0_3 ), .C(FIFO_CLK_c), .D(n4943));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFS \aempty_flag_impl.ae_flag_ext_r_130  (.Q(dc32_fifo_almost_empty), 
            .C(SLM_CLK_c), .D(\aempty_flag_impl.ae_flag_nxt_w ), .S(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(669[37] 672[40])
    SB_LUT4 n12495_bdd_4_lut (.I0(n12495), .I1(\REG.mem_53_11 ), .I2(\REG.mem_52_11 ), 
            .I3(rd_addr_r[1]), .O(n11570));
    defparam n12495_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11097 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_12 ), 
            .I2(\REG.mem_15_12 ), .I3(rd_addr_r[1]), .O(n13107));
    defparam rd_addr_r_0__bdd_4_lut_11097.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10580 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_30_0 ), 
            .I2(\REG.mem_31_0 ), .I3(rd_addr_r[1]), .O(n12489));
    defparam rd_addr_r_0__bdd_4_lut_10580.LUT_INIT = 16'he4aa;
    SB_LUT4 n13107_bdd_4_lut (.I0(n13107), .I1(\REG.mem_13_12 ), .I2(\REG.mem_12_12 ), 
            .I3(rd_addr_r[1]), .O(n13110));
    defparam n13107_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12489_bdd_4_lut (.I0(n12489), .I1(\REG.mem_29_0 ), .I2(\REG.mem_28_0 ), 
            .I3(rd_addr_r[1]), .O(n12492));
    defparam n12489_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9037_3_lut (.I0(\REG.mem_0_5 ), .I1(\REG.mem_1_5 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n10887));
    defparam i9037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9038_3_lut (.I0(\REG.mem_2_5 ), .I1(\REG.mem_3_5 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n10888));
    defparam i9038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9074_3_lut (.I0(\REG.mem_6_5 ), .I1(\REG.mem_7_5 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n10924));
    defparam i9074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9073_3_lut (.I0(\REG.mem_4_5 ), .I1(\REG.mem_5_5 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n10923));
    defparam i9073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10575 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_58_11 ), 
            .I2(\REG.mem_59_11 ), .I3(rd_addr_r[1]), .O(n12483));
    defparam rd_addr_r_0__bdd_4_lut_10575.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11182 (.I0(rd_addr_r[3]), .I1(n12948), 
            .I2(n11437), .I3(rd_addr_r[4]), .O(n13101));
    defparam rd_addr_r_3__bdd_4_lut_11182.LUT_INIT = 16'he4aa;
    SB_LUT4 n13101_bdd_4_lut (.I0(n13101), .I1(n11413), .I2(n12936), .I3(rd_addr_r[4]), 
            .O(n13104));
    defparam n13101_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12483_bdd_4_lut (.I0(n12483), .I1(\REG.mem_57_11 ), .I2(\REG.mem_56_11 ), 
            .I3(rd_addr_r[1]), .O(n11573));
    defparam n12483_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i76_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n62));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i76_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10570 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_62_13 ), 
            .I2(\REG.mem_63_13 ), .I3(rd_addr_r[1]), .O(n12477));
    defparam rd_addr_r_0__bdd_4_lut_10570.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11087 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_46_1 ), 
            .I2(\REG.mem_47_1 ), .I3(rd_addr_r[1]), .O(n13095));
    defparam rd_addr_r_0__bdd_4_lut_11087.LUT_INIT = 16'he4aa;
    SB_LUT4 n12477_bdd_4_lut (.I0(n12477), .I1(\REG.mem_61_13 ), .I2(\REG.mem_60_13 ), 
            .I3(rd_addr_r[1]), .O(n12480));
    defparam n12477_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13095_bdd_4_lut (.I0(n13095), .I1(\REG.mem_45_1 ), .I2(\REG.mem_44_1 ), 
            .I3(rd_addr_r[1]), .O(n13098));
    defparam n13095_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3501_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_1_0 ), .O(n4884));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3501_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11077 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_2_11 ), 
            .I2(\REG.mem_3_11 ), .I3(rd_addr_r[1]), .O(n13089));
    defparam rd_addr_r_0__bdd_4_lut_11077.LUT_INIT = 16'he4aa;
    SB_LUT4 n13089_bdd_4_lut (.I0(n13089), .I1(\REG.mem_1_11 ), .I2(\REG.mem_0_11 ), 
            .I3(rd_addr_r[1]), .O(n11459));
    defparam n13089_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10638 (.I0(rd_addr_r[2]), .I1(n11315), 
            .I2(n11336), .I3(rd_addr_r[3]), .O(n12471));
    defparam rd_addr_r_2__bdd_4_lut_10638.LUT_INIT = 16'he4aa;
    SB_LUT4 n12471_bdd_4_lut (.I0(n12471), .I1(n11258), .I2(n11219), .I3(rd_addr_r[3]), 
            .O(n11579));
    defparam n12471_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11072 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_6_11 ), 
            .I2(\REG.mem_7_11 ), .I3(rd_addr_r[1]), .O(n13083));
    defparam rd_addr_r_0__bdd_4_lut_11072.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i75_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n30));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i75_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 n12129_bdd_4_lut (.I0(n12129), .I1(\REG.mem_5_2 ), .I2(\REG.mem_4_2 ), 
            .I3(rd_addr_r[1]), .O(n12132));
    defparam n12129_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10288 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_18_5 ), 
            .I2(\REG.mem_19_5 ), .I3(rd_addr_r[1]), .O(n12135));
    defparam rd_addr_r_0__bdd_4_lut_10288.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10565 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_62_1 ), 
            .I2(\REG.mem_63_1 ), .I3(rd_addr_r[1]), .O(n12465));
    defparam rd_addr_r_0__bdd_4_lut_10565.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10278 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_38_13 ), 
            .I2(\REG.mem_39_13 ), .I3(rd_addr_r[1]), .O(n12123));
    defparam rd_addr_r_0__bdd_4_lut_10278.LUT_INIT = 16'he4aa;
    SB_LUT4 n12465_bdd_4_lut (.I0(n12465), .I1(\REG.mem_61_1 ), .I2(\REG.mem_60_1 ), 
            .I3(rd_addr_r[1]), .O(n12468));
    defparam n12465_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13083_bdd_4_lut (.I0(n13083), .I1(\REG.mem_5_11 ), .I2(\REG.mem_4_11 ), 
            .I3(rd_addr_r[1]), .O(n11462));
    defparam n13083_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3517_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_1_8 ), .O(n4900));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3517_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10555 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_5 ), 
            .I2(\REG.mem_15_5 ), .I3(rd_addr_r[1]), .O(n12459));
    defparam rd_addr_r_0__bdd_4_lut_10555.LUT_INIT = 16'he4aa;
    SB_LUT4 n12459_bdd_4_lut (.I0(n12459), .I1(\REG.mem_13_5 ), .I2(\REG.mem_12_5 ), 
            .I3(rd_addr_r[1]), .O(n12462));
    defparam n12459_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11067 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_30_9 ), 
            .I2(\REG.mem_31_9 ), .I3(rd_addr_r[1]), .O(n13077));
    defparam rd_addr_r_0__bdd_4_lut_11067.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_r_6__I_0_135_i6_3_lut (.I0(wr_addr_r[5]), .I1(wr_addr_p1_w[5]), 
            .I2(wr_sig_mv_w), .I3(GND_net), .O(\wr_addr_nxt_c[5] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13077_bdd_4_lut (.I0(n13077), .I1(\REG.mem_29_9 ), .I2(\REG.mem_28_9 ), 
            .I3(rd_addr_r[1]), .O(n13080));
    defparam n13077_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10550 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_46_12 ), 
            .I2(\REG.mem_47_12 ), .I3(rd_addr_r[1]), .O(n12453));
    defparam rd_addr_r_0__bdd_4_lut_10550.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11092 (.I0(rd_addr_r[1]), .I1(n11022), 
            .I2(n11023), .I3(rd_addr_r[2]), .O(n13071));
    defparam rd_addr_r_1__bdd_4_lut_11092.LUT_INIT = 16'he4aa;
    SB_LUT4 n12453_bdd_4_lut (.I0(n12453), .I1(\REG.mem_45_12 ), .I2(\REG.mem_44_12 ), 
            .I3(rd_addr_r[1]), .O(n12456));
    defparam n12453_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i4_1_lut (.I0(rd_addr_r[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n13071_bdd_4_lut (.I0(n13071), .I1(n11020), .I2(n11019), .I3(rd_addr_r[2]), 
            .O(n11101));
    defparam n13071_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10545 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_62_11 ), 
            .I2(\REG.mem_63_11 ), .I3(rd_addr_r[1]), .O(n12447));
    defparam rd_addr_r_0__bdd_4_lut_10545.LUT_INIT = 16'he4aa;
    SB_LUT4 n12447_bdd_4_lut (.I0(n12447), .I1(\REG.mem_61_11 ), .I2(\REG.mem_60_11 ), 
            .I3(rd_addr_r[1]), .O(n11588));
    defparam n12447_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9871_3_lut (.I0(\REG.mem_56_8 ), .I1(\REG.mem_57_8 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11721));
    defparam i9871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11062 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_62_6 ), 
            .I2(\REG.mem_63_6 ), .I3(rd_addr_r[1]), .O(n13065));
    defparam rd_addr_r_0__bdd_4_lut_11062.LUT_INIT = 16'he4aa;
    SB_LUT4 i9872_3_lut (.I0(\REG.mem_58_8 ), .I1(\REG.mem_59_8 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11722));
    defparam i9872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9935_3_lut (.I0(\REG.mem_62_8 ), .I1(\REG.mem_63_8 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11785));
    defparam i9935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9934_3_lut (.I0(\REG.mem_60_8 ), .I1(\REG.mem_61_8 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11784));
    defparam i9934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13065_bdd_4_lut (.I0(n13065), .I1(\REG.mem_61_6 ), .I2(\REG.mem_60_6 ), 
            .I3(rd_addr_r[1]), .O(n11465));
    defparam n13065_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10540 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_34_0 ), 
            .I2(\REG.mem_35_0 ), .I3(rd_addr_r[1]), .O(n12441));
    defparam rd_addr_r_0__bdd_4_lut_10540.LUT_INIT = 16'he4aa;
    SB_LUT4 n12441_bdd_4_lut (.I0(n12441), .I1(\REG.mem_33_0 ), .I2(\REG.mem_32_0 ), 
            .I3(rd_addr_r[1]), .O(n11171));
    defparam n12441_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10535 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_26_15 ), 
            .I2(\REG.mem_27_15 ), .I3(rd_addr_r[1]), .O(n12435));
    defparam rd_addr_r_0__bdd_4_lut_10535.LUT_INIT = 16'he4aa;
    SB_LUT4 n12435_bdd_4_lut (.I0(n12435), .I1(\REG.mem_25_15 ), .I2(\REG.mem_24_15 ), 
            .I3(rd_addr_r[1]), .O(n12438));
    defparam n12435_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11082 (.I0(rd_addr_r[3]), .I1(n12954), 
            .I2(n11446), .I3(rd_addr_r[4]), .O(n13059));
    defparam rd_addr_r_3__bdd_4_lut_11082.LUT_INIT = 16'he4aa;
    SB_LUT4 n13059_bdd_4_lut (.I0(n13059), .I1(n11434), .I2(n12942), .I3(rd_addr_r[4]), 
            .O(n13062));
    defparam n13059_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9412_3_lut (.I0(\REG.mem_32_7 ), .I1(\REG.mem_33_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11262));
    defparam i9412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9413_3_lut (.I0(\REG.mem_34_7 ), .I1(\REG.mem_35_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11263));
    defparam i9413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11052 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_34_9 ), 
            .I2(\REG.mem_35_9 ), .I3(rd_addr_r[1]), .O(n13053));
    defparam rd_addr_r_0__bdd_4_lut_11052.LUT_INIT = 16'he4aa;
    SB_LUT4 n13053_bdd_4_lut (.I0(n13053), .I1(\REG.mem_33_9 ), .I2(\REG.mem_32_9 ), 
            .I3(rd_addr_r[1]), .O(n13056));
    defparam n13053_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11057 (.I0(rd_addr_r[1]), .I1(n11049), 
            .I2(n11050), .I3(rd_addr_r[2]), .O(n13047));
    defparam rd_addr_r_1__bdd_4_lut_11057.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10560 (.I0(rd_addr_r[2]), .I1(n10919), 
            .I2(n10928), .I3(rd_addr_r[3]), .O(n12429));
    defparam rd_addr_r_2__bdd_4_lut_10560.LUT_INIT = 16'he4aa;
    SB_LUT4 n12429_bdd_4_lut (.I0(n12429), .I1(n10916), .I2(n10910), .I3(rd_addr_r[3]), 
            .O(n10988));
    defparam n12429_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10525 (.I0(rd_addr_r[2]), .I1(n11474), 
            .I2(n11483), .I3(rd_addr_r[3]), .O(n12423));
    defparam rd_addr_r_2__bdd_4_lut_10525.LUT_INIT = 16'he4aa;
    SB_LUT4 n12423_bdd_4_lut (.I0(n12423), .I1(n11462), .I2(n11459), .I3(rd_addr_r[3]), 
            .O(n11594));
    defparam n12423_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13047_bdd_4_lut (.I0(n13047), .I1(n11044), .I2(n11043), .I3(rd_addr_r[2]), 
            .O(n11107));
    defparam n13047_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11042 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_18_12 ), 
            .I2(\REG.mem_19_12 ), .I3(rd_addr_r[1]), .O(n13041));
    defparam rd_addr_r_0__bdd_4_lut_11042.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10520 (.I0(rd_addr_r[2]), .I1(n10844), 
            .I2(n10847), .I3(rd_addr_r[3]), .O(n12417));
    defparam rd_addr_r_2__bdd_4_lut_10520.LUT_INIT = 16'he4aa;
    SB_LUT4 n12417_bdd_4_lut (.I0(n12417), .I1(n11867), .I2(n11861), .I3(rd_addr_r[3]), 
            .O(n12420));
    defparam n12417_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13041_bdd_4_lut (.I0(n13041), .I1(\REG.mem_17_12 ), .I2(\REG.mem_16_12 ), 
            .I3(rd_addr_r[1]), .O(n13044));
    defparam n13041_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10530 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_8 ), 
            .I2(\REG.mem_15_8 ), .I3(rd_addr_r[1]), .O(n12411));
    defparam rd_addr_r_0__bdd_4_lut_10530.LUT_INIT = 16'he4aa;
    SB_LUT4 n12411_bdd_4_lut (.I0(n12411), .I1(\REG.mem_13_8 ), .I2(\REG.mem_12_8 ), 
            .I3(rd_addr_r[1]), .O(n12414));
    defparam n12411_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_2 ), 
            .I2(\REG.mem_15_2 ), .I3(rd_addr_r[1]), .O(n13731));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n13731_bdd_4_lut (.I0(n13731), .I1(\REG.mem_13_2 ), .I2(\REG.mem_12_2 ), 
            .I3(rd_addr_r[1]), .O(n13734));
    defparam n13731_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9431_3_lut (.I0(\REG.mem_38_7 ), .I1(\REG.mem_39_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11281));
    defparam i9431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11037 (.I0(rd_addr_r[1]), .I1(n11070), 
            .I2(n11071), .I3(rd_addr_r[2]), .O(n13035));
    defparam rd_addr_r_1__bdd_4_lut_11037.LUT_INIT = 16'he4aa;
    SB_LUT4 i9430_3_lut (.I0(\REG.mem_36_7 ), .I1(\REG.mem_37_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11280));
    defparam i9430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10510 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_50_12 ), 
            .I2(\REG.mem_51_12 ), .I3(rd_addr_r[1]), .O(n12405));
    defparam rd_addr_r_0__bdd_4_lut_10510.LUT_INIT = 16'he4aa;
    SB_LUT4 n13035_bdd_4_lut (.I0(n13035), .I1(n11068), .I2(n11067), .I3(rd_addr_r[2]), 
            .O(n11110));
    defparam n13035_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12405_bdd_4_lut (.I0(n12405), .I1(\REG.mem_49_12 ), .I2(\REG.mem_48_12 ), 
            .I3(rd_addr_r[1]), .O(n12408));
    defparam n12405_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11607 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_62_9 ), 
            .I2(\REG.mem_63_9 ), .I3(rd_addr_r[1]), .O(n13725));
    defparam rd_addr_r_0__bdd_4_lut_11607.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10505 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_6_9 ), 
            .I2(\REG.mem_7_9 ), .I3(rd_addr_r[1]), .O(n12399));
    defparam rd_addr_r_0__bdd_4_lut_10505.LUT_INIT = 16'he4aa;
    SB_LUT4 n13725_bdd_4_lut (.I0(n13725), .I1(\REG.mem_61_9 ), .I2(\REG.mem_60_9 ), 
            .I3(rd_addr_r[1]), .O(n13728));
    defparam n13725_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11602 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_34_6 ), 
            .I2(\REG.mem_35_6 ), .I3(rd_addr_r[1]), .O(n13719));
    defparam rd_addr_r_0__bdd_4_lut_11602.LUT_INIT = 16'he4aa;
    SB_LUT4 n12399_bdd_4_lut (.I0(n12399), .I1(\REG.mem_5_9 ), .I2(\REG.mem_4_9 ), 
            .I3(rd_addr_r[1]), .O(n12402));
    defparam n12399_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12123_bdd_4_lut (.I0(n12123), .I1(\REG.mem_37_13 ), .I2(\REG.mem_36_13 ), 
            .I3(rd_addr_r[1]), .O(n12126));
    defparam n12123_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13719_bdd_4_lut (.I0(n13719), .I1(\REG.mem_33_6 ), .I2(\REG.mem_32_6 ), 
            .I3(rd_addr_r[1]), .O(n11219));
    defparam n13719_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10500 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_42_8 ), 
            .I2(\REG.mem_43_8 ), .I3(rd_addr_r[1]), .O(n12393));
    defparam rd_addr_r_0__bdd_4_lut_10500.LUT_INIT = 16'he4aa;
    SB_LUT4 n12393_bdd_4_lut (.I0(n12393), .I1(\REG.mem_41_8 ), .I2(\REG.mem_40_8 ), 
            .I3(rd_addr_r[1]), .O(n12396));
    defparam n12393_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11597 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_22_7 ), 
            .I2(\REG.mem_23_7 ), .I3(rd_addr_r[1]), .O(n13713));
    defparam rd_addr_r_0__bdd_4_lut_11597.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11032 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_11 ), 
            .I2(\REG.mem_11_11 ), .I3(rd_addr_r[1]), .O(n13029));
    defparam rd_addr_r_0__bdd_4_lut_11032.LUT_INIT = 16'he4aa;
    SB_LUT4 n13713_bdd_4_lut (.I0(n13713), .I1(\REG.mem_21_7 ), .I2(\REG.mem_20_7 ), 
            .I3(rd_addr_r[1]), .O(n13716));
    defparam n13713_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i3_1_lut (.I0(rd_addr_r[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n13029_bdd_4_lut (.I0(n13029), .I1(\REG.mem_9_11 ), .I2(\REG.mem_8_11 ), 
            .I3(rd_addr_r[1]), .O(n11474));
    defparam n13029_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10515 (.I0(rd_addr_r[2]), .I1(n10940), 
            .I2(n10955), .I3(rd_addr_r[3]), .O(n12387));
    defparam rd_addr_r_2__bdd_4_lut_10515.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11022 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_2_15 ), 
            .I2(\REG.mem_3_15 ), .I3(rd_addr_r[1]), .O(n13023));
    defparam rd_addr_r_0__bdd_4_lut_11022.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11592 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_46_8 ), 
            .I2(\REG.mem_47_8 ), .I3(rd_addr_r[1]), .O(n13707));
    defparam rd_addr_r_0__bdd_4_lut_11592.LUT_INIT = 16'he4aa;
    SB_LUT4 n13707_bdd_4_lut (.I0(n13707), .I1(\REG.mem_45_8 ), .I2(\REG.mem_44_8 ), 
            .I3(rd_addr_r[1]), .O(n13710));
    defparam n13707_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13023_bdd_4_lut (.I0(n13023), .I1(\REG.mem_1_15 ), .I2(\REG.mem_0_15 ), 
            .I3(rd_addr_r[1]), .O(n13026));
    defparam n13023_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i50_51 (.Q(\REG.mem_0_4 ), .C(FIFO_CLK_c), .D(n4935));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11587 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_46_5 ), 
            .I2(\REG.mem_47_5 ), .I3(rd_addr_r[1]), .O(n13701));
    defparam rd_addr_r_0__bdd_4_lut_11587.LUT_INIT = 16'he4aa;
    SB_LUT4 n13701_bdd_4_lut (.I0(n13701), .I1(\REG.mem_45_5 ), .I2(\REG.mem_44_5 ), 
            .I3(rd_addr_r[1]), .O(n13704));
    defparam n13701_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12387_bdd_4_lut (.I0(n12387), .I1(n10937), .I2(n10931), .I3(rd_addr_r[3]), 
            .O(n10997));
    defparam n12387_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10273 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_2 ), 
            .I2(\REG.mem_11_2 ), .I3(rd_addr_r[1]), .O(n12117));
    defparam rd_addr_r_0__bdd_4_lut_10273.LUT_INIT = 16'he4aa;
    SB_LUT4 n12159_bdd_4_lut (.I0(n12159), .I1(\REG.mem_61_12 ), .I2(\REG.mem_60_12 ), 
            .I3(rd_addr_r[1]), .O(n12162));
    defparam n12159_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10375 (.I0(rd_addr_r[4]), .I1(n11579), 
            .I2(n11633), .I3(rd_addr_r[5]), .O(n12153));
    defparam rd_addr_r_4__bdd_4_lut_10375.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10380 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_54_9 ), 
            .I2(\REG.mem_55_9 ), .I3(rd_addr_r[1]), .O(n12231));
    defparam rd_addr_r_0__bdd_4_lut_10380.LUT_INIT = 16'he4aa;
    SB_LUT4 n12147_bdd_4_lut (.I0(n12147), .I1(\REG.mem_57_9 ), .I2(\REG.mem_56_9 ), 
            .I3(rd_addr_r[1]), .O(n12150));
    defparam n12147_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11582 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_58_14 ), 
            .I2(\REG.mem_59_14 ), .I3(rd_addr_r[1]), .O(n13695));
    defparam rd_addr_r_0__bdd_4_lut_11582.LUT_INIT = 16'he4aa;
    SB_LUT4 n13695_bdd_4_lut (.I0(n13695), .I1(\REG.mem_57_14 ), .I2(\REG.mem_56_14 ), 
            .I3(rd_addr_r[1]), .O(n10844));
    defparam n13695_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11027 (.I0(rd_addr_r[1]), .I1(n11091), 
            .I2(n11092), .I3(rd_addr_r[2]), .O(n13017));
    defparam rd_addr_r_1__bdd_4_lut_11027.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10495 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_30_15 ), 
            .I2(\REG.mem_31_15 ), .I3(rd_addr_r[1]), .O(n12381));
    defparam rd_addr_r_0__bdd_4_lut_10495.LUT_INIT = 16'he4aa;
    SB_LUT4 n12381_bdd_4_lut (.I0(n12381), .I1(\REG.mem_29_15 ), .I2(\REG.mem_28_15 ), 
            .I3(rd_addr_r[1]), .O(n12384));
    defparam n12381_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10293 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_42_15 ), 
            .I2(\REG.mem_43_15 ), .I3(rd_addr_r[1]), .O(n12141));
    defparam rd_addr_r_0__bdd_4_lut_10293.LUT_INIT = 16'he4aa;
    SB_LUT4 n12135_bdd_4_lut (.I0(n12135), .I1(\REG.mem_17_5 ), .I2(\REG.mem_16_5 ), 
            .I3(rd_addr_r[1]), .O(n12138));
    defparam n12135_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13017_bdd_4_lut (.I0(n13017), .I1(n11089), .I2(n11088), .I3(rd_addr_r[2]), 
            .O(n11113));
    defparam n13017_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12117_bdd_4_lut (.I0(n12117), .I1(\REG.mem_9_2 ), .I2(\REG.mem_8_2 ), 
            .I3(rd_addr_r[1]), .O(n12120));
    defparam n12117_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10307 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_62_12 ), 
            .I2(\REG.mem_63_12 ), .I3(rd_addr_r[1]), .O(n12159));
    defparam rd_addr_r_0__bdd_4_lut_10307.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_r_6__I_0_135_i4_3_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(wr_sig_mv_w), .I3(GND_net), .O(\wr_addr_nxt_c[3] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11577 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_18_8 ), 
            .I2(\REG.mem_19_8 ), .I3(rd_addr_r[1]), .O(n13689));
    defparam rd_addr_r_0__bdd_4_lut_11577.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10490 (.I0(rd_addr_r[2]), .I1(n11507), 
            .I2(n11519), .I3(rd_addr_r[3]), .O(n12375));
    defparam rd_addr_r_2__bdd_4_lut_10490.LUT_INIT = 16'he4aa;
    SB_LUT4 i3827_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_17_15 ), .O(n5210));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3827_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i5_1_lut (.I0(rd_addr_r[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n13689_bdd_4_lut (.I0(n13689), .I1(\REG.mem_17_8 ), .I2(\REG.mem_16_8 ), 
            .I3(rd_addr_r[1]), .O(n13692));
    defparam n13689_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12153_bdd_4_lut (.I0(n12153), .I1(n11555), .I2(n11510), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_559 [6]));
    defparam n12153_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12375_bdd_4_lut (.I0(n12375), .I1(n11504), .I2(n11495), .I3(rd_addr_r[3]), 
            .O(n11606));
    defparam n12375_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11017 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_22_12 ), 
            .I2(\REG.mem_23_12 ), .I3(rd_addr_r[1]), .O(n13011));
    defparam rd_addr_r_0__bdd_4_lut_11017.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11572 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_26_2 ), 
            .I2(\REG.mem_27_2 ), .I3(rd_addr_r[1]), .O(n13683));
    defparam rd_addr_r_0__bdd_4_lut_11572.LUT_INIT = 16'he4aa;
    SB_LUT4 n13011_bdd_4_lut (.I0(n13011), .I1(\REG.mem_21_12 ), .I2(\REG.mem_20_12 ), 
            .I3(rd_addr_r[1]), .O(n13014));
    defparam n13011_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13683_bdd_4_lut (.I0(n13683), .I1(\REG.mem_25_2 ), .I2(\REG.mem_24_2 ), 
            .I3(rd_addr_r[1]), .O(n13686));
    defparam n13683_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11567 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_30_2 ), 
            .I2(\REG.mem_31_2 ), .I3(rd_addr_r[1]), .O(n13677));
    defparam rd_addr_r_0__bdd_4_lut_11567.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10480 (.I0(rd_addr_r[2]), .I1(n10976), 
            .I2(n10979), .I3(rd_addr_r[3]), .O(n12369));
    defparam rd_addr_r_2__bdd_4_lut_10480.LUT_INIT = 16'he4aa;
    SB_LUT4 n12369_bdd_4_lut (.I0(n12369), .I1(n10970), .I2(n10964), .I3(rd_addr_r[3]), 
            .O(n11000));
    defparam n12369_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3826_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_17_14 ), .O(n5209));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3826_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9517_3_lut (.I0(\REG.mem_48_10 ), .I1(\REG.mem_49_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11367));
    defparam i9517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9518_3_lut (.I0(\REG.mem_50_10 ), .I1(\REG.mem_51_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11368));
    defparam i9518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13677_bdd_4_lut (.I0(n13677), .I1(\REG.mem_29_2 ), .I2(\REG.mem_28_2 ), 
            .I3(rd_addr_r[1]), .O(n13680));
    defparam n13677_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9033_3_lut (.I0(n12558), .I1(n13662), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [2]));
    defparam i9033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3825_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_17_13 ), .O(n5208));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3825_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9521_3_lut (.I0(\REG.mem_54_10 ), .I1(\REG.mem_55_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11371));
    defparam i9521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9520_3_lut (.I0(\REG.mem_52_10 ), .I1(\REG.mem_53_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11370));
    defparam i9520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9276_3_lut (.I0(n12756), .I1(n12870), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [4]));
    defparam i9276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11007 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_11 ), 
            .I2(\REG.mem_15_11 ), .I3(rd_addr_r[1]), .O(n13005));
    defparam rd_addr_r_0__bdd_4_lut_11007.LUT_INIT = 16'he4aa;
    SB_LUT4 i3824_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_17_12 ), .O(n5207));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3824_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10485 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_54_12 ), 
            .I2(\REG.mem_55_12 ), .I3(rd_addr_r[1]), .O(n12363));
    defparam rd_addr_r_0__bdd_4_lut_10485.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut (.I0(rd_addr_r[1]), .I1(n11709), .I2(n11710), 
            .I3(rd_addr_r[2]), .O(n13671));
    defparam rd_addr_r_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n13005_bdd_4_lut (.I0(n13005), .I1(\REG.mem_13_11 ), .I2(\REG.mem_12_11 ), 
            .I3(rd_addr_r[1]), .O(n11483));
    defparam n13005_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12363_bdd_4_lut (.I0(n12363), .I1(\REG.mem_53_12 ), .I2(\REG.mem_52_12 ), 
            .I3(rd_addr_r[1]), .O(n12366));
    defparam n12363_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13671_bdd_4_lut (.I0(n13671), .I1(n11707), .I2(n11706), .I3(rd_addr_r[2]), 
            .O(n10876));
    defparam n13671_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9528_3_lut (.I0(n12912), .I1(n13386), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [5]));
    defparam i9528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10470 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_34_15 ), 
            .I2(\REG.mem_35_15 ), .I3(rd_addr_r[1]), .O(n12357));
    defparam rd_addr_r_0__bdd_4_lut_10470.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11562 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_38_6 ), 
            .I2(\REG.mem_39_6 ), .I3(rd_addr_r[1]), .O(n13665));
    defparam rd_addr_r_0__bdd_4_lut_11562.LUT_INIT = 16'he4aa;
    SB_LUT4 i9618_3_lut (.I0(n12966), .I1(n13062), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [7]));
    defparam i9618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11002 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_58_13 ), 
            .I2(\REG.mem_59_13 ), .I3(rd_addr_r[1]), .O(n12999));
    defparam rd_addr_r_0__bdd_4_lut_11002.LUT_INIT = 16'he4aa;
    SB_LUT4 n12357_bdd_4_lut (.I0(n12357), .I1(\REG.mem_33_15 ), .I2(\REG.mem_32_15 ), 
            .I3(rd_addr_r[1]), .O(n12360));
    defparam n12357_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9099_3_lut (.I0(n12672), .I1(n13224), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [8]));
    defparam i9099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3823_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_17_11 ), .O(n5206));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3823_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9411_3_lut (.I0(n12858), .I1(n13656), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [9]));
    defparam i9411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13665_bdd_4_lut (.I0(n13665), .I1(\REG.mem_37_6 ), .I2(\REG.mem_36_6 ), 
            .I3(rd_addr_r[1]), .O(n11258));
    defparam n13665_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12999_bdd_4_lut (.I0(n12999), .I1(\REG.mem_57_13 ), .I2(\REG.mem_56_13 ), 
            .I3(rd_addr_r[1]), .O(n13002));
    defparam n12999_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3822_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_17_10 ), .O(n5205));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3822_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut (.I0(rd_addr_r[3]), .I1(n12540), .I2(n10873), 
            .I3(rd_addr_r[4]), .O(n13659));
    defparam rd_addr_r_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10475 (.I0(rd_addr_r[2]), .I1(n11543), 
            .I2(n11552), .I3(rd_addr_r[3]), .O(n12351));
    defparam rd_addr_r_2__bdd_4_lut_10475.LUT_INIT = 16'he4aa;
    SB_LUT4 n12351_bdd_4_lut (.I0(n12351), .I1(n11528), .I2(n11525), .I3(rd_addr_r[3]), 
            .O(n11615));
    defparam n12351_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3821_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_17_9 ), .O(n5204));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3821_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3820_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_17_8 ), .O(n5203));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3820_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9603_3_lut (.I0(n12960), .I1(n13104), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [10]));
    defparam i9603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3819_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_17_7 ), .O(n5202));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3819_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13659_bdd_4_lut (.I0(n13659), .I1(n10870), .I2(n12534), .I3(rd_addr_r[4]), 
            .O(n13662));
    defparam n13659_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3818_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_17_6 ), .O(n5201));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3818_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3817_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_17_5 ), .O(n5200));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3817_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10997 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_30_13 ), 
            .I2(\REG.mem_31_13 ), .I3(rd_addr_r[1]), .O(n12993));
    defparam rd_addr_r_0__bdd_4_lut_10997.LUT_INIT = 16'he4aa;
    SB_LUT4 i3816_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_17_4 ), .O(n5199));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3816_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11547 (.I0(rd_addr_r[3]), .I1(n11250), 
            .I2(n11251), .I3(rd_addr_r[4]), .O(n13653));
    defparam rd_addr_r_3__bdd_4_lut_11547.LUT_INIT = 16'he4aa;
    SB_LUT4 i3815_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_17_3 ), .O(n5198));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3815_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12993_bdd_4_lut (.I0(n12993), .I1(\REG.mem_29_13 ), .I2(\REG.mem_28_13 ), 
            .I3(rd_addr_r[1]), .O(n12996));
    defparam n12993_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3814_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_17_2 ), .O(n5197));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3814_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3813_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_17_1 ), .O(n5196));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3813_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3812_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_17_0 ), .O(n5195));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3812_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3859_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_19_15 ), .O(n5242));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3859_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13653_bdd_4_lut (.I0(n13653), .I1(n11242), .I2(n11241), .I3(rd_addr_r[4]), 
            .O(n13656));
    defparam n13653_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3858_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_19_14 ), .O(n5241));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3858_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9933_3_lut (.I0(n13398), .I1(n13608), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [12]));
    defparam i9933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12231_bdd_4_lut (.I0(n12231), .I1(\REG.mem_53_9 ), .I2(\REG.mem_52_9 ), 
            .I3(rd_addr_r[1]), .O(n12234));
    defparam n12231_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9117_3_lut (.I0(n12684), .I1(n12780), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n10967));
    defparam i9117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3857_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_19_13 ), .O(n5240));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3857_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9185_3_lut (.I0(n10967), .I1(n12420), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(n11035));
    defparam i9185_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i53_54 (.Q(\REG.mem_0_5 ), .C(FIFO_CLK_c), .D(n4934));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9186_3_lut (.I0(n12726), .I1(n11035), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [14]));
    defparam i9186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9063_3_lut (.I0(n12606), .I1(n13434), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_559 [15]));
    defparam i9063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10673 (.I0(rd_addr_r[4]), .I1(n10997), 
            .I2(n11000), .I3(rd_addr_r[5]), .O(n12345));
    defparam rd_addr_r_4__bdd_4_lut_10673.LUT_INIT = 16'he4aa;
    SB_DFF i56_57 (.Q(\REG.mem_0_6 ), .C(FIFO_CLK_c), .D(n4933));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut (.I0(rd_addr_r[2]), .I1(n13170), .I2(n13098), 
            .I3(rd_addr_r[3]), .O(n13647));
    defparam rd_addr_r_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i3856_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_19_12 ), .O(n5239));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3856_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13647_bdd_4_lut (.I0(n13647), .I1(n13326), .I2(n13392), .I3(rd_addr_r[3]), 
            .O(n11753));
    defparam n13647_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10992 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_30_5 ), 
            .I2(\REG.mem_31_5 ), .I3(rd_addr_r[1]), .O(n12987));
    defparam rd_addr_r_0__bdd_4_lut_10992.LUT_INIT = 16'he4aa;
    SB_LUT4 i3855_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_19_11 ), .O(n5238));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3855_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12345_bdd_4_lut (.I0(n12345), .I1(n10988), .I2(n10982), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_559 [3]));
    defparam n12345_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3854_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_19_10 ), .O(n5237));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3854_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3853_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_19_9 ), .O(n5236));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3853_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3852_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_19_8 ), .O(n5235));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3852_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3851_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_19_7 ), .O(n5234));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3851_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3850_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_19_6 ), .O(n5233));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3850_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9475_3_lut (.I0(\REG.mem_48_7 ), .I1(\REG.mem_49_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11325));
    defparam i9475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9476_3_lut (.I0(\REG.mem_50_7 ), .I1(\REG.mem_51_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11326));
    defparam i9476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9506_3_lut (.I0(\REG.mem_54_7 ), .I1(\REG.mem_55_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11356));
    defparam i9506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9505_3_lut (.I0(\REG.mem_52_7 ), .I1(\REG.mem_53_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11355));
    defparam i9505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3849_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_19_5 ), .O(n5232));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3849_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11537 (.I0(rd_addr_r[2]), .I1(n13602), 
            .I2(n12996), .I3(rd_addr_r[3]), .O(n13641));
    defparam rd_addr_r_2__bdd_4_lut_11537.LUT_INIT = 16'he4aa;
    SB_LUT4 i3848_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_19_4 ), .O(n5231));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3848_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3847_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_19_3 ), .O(n5230));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3847_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12987_bdd_4_lut (.I0(n12987), .I1(\REG.mem_29_5 ), .I2(\REG.mem_28_5 ), 
            .I3(rd_addr_r[1]), .O(n12990));
    defparam n12987_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3846_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_19_2 ), .O(n5229));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3846_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3845_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_19_1 ), .O(n5228));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3845_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3844_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_19_0 ), .O(n5227));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3844_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3875_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_20_15 ), .O(n5258));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3875_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_buffer__i2  (.Q(\fifo_data_out[2] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6106));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 n13641_bdd_4_lut (.I0(n13641), .I1(n13182), .I2(n13470), .I3(rd_addr_r[3]), 
            .O(n11762));
    defparam n13641_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3874_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_20_14 ), .O(n5257));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3874_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_buffer__i1  (.Q(\fifo_data_out[1] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6103));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10460 (.I0(rd_addr_r[2]), .I1(n11573), 
            .I2(n11588), .I3(rd_addr_r[3]), .O(n12339));
    defparam rd_addr_r_2__bdd_4_lut_10460.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10987 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_34_13 ), 
            .I2(\REG.mem_35_13 ), .I3(rd_addr_r[1]), .O(n12981));
    defparam rd_addr_r_0__bdd_4_lut_10987.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11552 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_2_3 ), 
            .I2(\REG.mem_3_3 ), .I3(rd_addr_r[1]), .O(n13635));
    defparam rd_addr_r_0__bdd_4_lut_11552.LUT_INIT = 16'he4aa;
    SB_LUT4 n12981_bdd_4_lut (.I0(n12981), .I1(\REG.mem_33_13 ), .I2(\REG.mem_32_13 ), 
            .I3(rd_addr_r[1]), .O(n12984));
    defparam n12981_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4366_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_49_15 ), .O(n5749));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4366_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13635_bdd_4_lut (.I0(n13635), .I1(\REG.mem_1_3 ), .I2(\REG.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(n10886));
    defparam n13635_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12339_bdd_4_lut (.I0(n12339), .I1(n11570), .I2(n11561), .I3(rd_addr_r[3]), 
            .O(n11618));
    defparam n12339_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i6_1_lut (.I0(rd_addr_r[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 wp_sync2_r_6__I_0_143_i1_2_lut (.I0(wp_sync2_r[5]), .I1(wp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(wp_sync_w[5]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam wp_sync2_r_6__I_0_143_i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i7_1_lut (.I0(\rd_addr_r[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4365_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_49_14 ), .O(n5748));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4365_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF \REG.out_buffer__i3  (.Q(\fifo_data_out[3] ), .C(SLM_CLK_c), 
           .D(n4827));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10982 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_50_1 ), 
            .I2(\REG.mem_51_1 ), .I3(rd_addr_r[1]), .O(n12975));
    defparam rd_addr_r_0__bdd_4_lut_10982.LUT_INIT = 16'he4aa;
    SB_DFF \REG.out_buffer__i4  (.Q(\fifo_data_out[4] ), .C(SLM_CLK_c), 
           .D(n4830));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i5  (.Q(\fifo_data_out[5] ), .C(SLM_CLK_c), 
           .D(n4841));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i6  (.Q(\fifo_data_out[6] ), .C(SLM_CLK_c), 
           .D(n4844));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i7  (.Q(\fifo_data_out[7] ), .C(SLM_CLK_c), 
           .D(n4848));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i8  (.Q(\fifo_data_out[8] ), .C(SLM_CLK_c), 
           .D(n4851));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i9  (.Q(\fifo_data_out[9] ), .C(SLM_CLK_c), 
           .D(n4854));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i10  (.Q(\fifo_data_out[10] ), .C(SLM_CLK_c), 
           .D(n4858));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i11  (.Q(\fifo_data_out[11] ), .C(SLM_CLK_c), 
           .D(n4864));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11527 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_62_14 ), 
            .I2(\REG.mem_63_14 ), .I3(rd_addr_r[1]), .O(n13629));
    defparam rd_addr_r_0__bdd_4_lut_11527.LUT_INIT = 16'he4aa;
    SB_LUT4 i4364_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_49_13 ), .O(n5747));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4364_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9898_3_lut (.I0(n12708), .I1(n12630), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11748));
    defparam i9898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12975_bdd_4_lut (.I0(n12975), .I1(\REG.mem_49_1 ), .I2(\REG.mem_48_1 ), 
            .I3(rd_addr_r[1]), .O(n12978));
    defparam n12975_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13629_bdd_4_lut (.I0(n13629), .I1(\REG.mem_61_14 ), .I2(\REG.mem_60_14 ), 
            .I3(rd_addr_r[1]), .O(n10847));
    defparam n13629_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9899_3_lut (.I0(n12522), .I1(n12456), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11749));
    defparam i9899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10977 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_18_11 ), 
            .I2(\REG.mem_19_11 ), .I3(rd_addr_r[1]), .O(n12969));
    defparam rd_addr_r_0__bdd_4_lut_10977.LUT_INIT = 16'he4aa;
    SB_LUT4 i9920_3_lut (.I0(n12270), .I1(n12162), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11770));
    defparam i9920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3873_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_20_13 ), .O(n5256));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3873_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12969_bdd_4_lut (.I0(n12969), .I1(\REG.mem_17_11 ), .I2(\REG.mem_16_11 ), 
            .I3(rd_addr_r[1]), .O(n11495));
    defparam n12969_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11522 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_6_3 ), 
            .I2(\REG.mem_7_3 ), .I3(rd_addr_r[1]), .O(n13623));
    defparam rd_addr_r_0__bdd_4_lut_11522.LUT_INIT = 16'he4aa;
    SB_LUT4 i9919_3_lut (.I0(n12408), .I1(n12366), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11769));
    defparam i9919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3872_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_20_12 ), .O(n5255));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3872_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11047 (.I0(rd_addr_r[3]), .I1(n11418), 
            .I2(n11419), .I3(rd_addr_r[4]), .O(n12963));
    defparam rd_addr_r_3__bdd_4_lut_11047.LUT_INIT = 16'he4aa;
    SB_LUT4 n13623_bdd_4_lut (.I0(n13623), .I1(\REG.mem_5_3 ), .I2(\REG.mem_4_3 ), 
            .I3(rd_addr_r[1]), .O(n10892));
    defparam n13623_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12963_bdd_4_lut (.I0(n12963), .I1(n11404), .I2(n12924), .I3(rd_addr_r[4]), 
            .O(n12966));
    defparam n12963_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11517 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_42_2 ), 
            .I2(\REG.mem_43_2 ), .I3(rd_addr_r[1]), .O(n13617));
    defparam rd_addr_r_0__bdd_4_lut_11517.LUT_INIT = 16'he4aa;
    SB_LUT4 n13617_bdd_4_lut (.I0(n13617), .I1(\REG.mem_41_2 ), .I2(\REG.mem_40_2 ), 
            .I3(rd_addr_r[1]), .O(n13620));
    defparam n13617_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3871_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_20_11 ), .O(n5254));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3871_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_buffer__i0  (.Q(\fifo_data_out[0] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6070));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 i3870_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_20_10 ), .O(n5253));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3870_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4363_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_49_12 ), .O(n5746));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4363_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10967 (.I0(rd_addr_r[3]), .I1(n12930), 
            .I2(n11410), .I3(rd_addr_r[4]), .O(n12957));
    defparam rd_addr_r_3__bdd_4_lut_10967.LUT_INIT = 16'he4aa;
    SB_LUT4 i4362_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_49_11 ), .O(n5745));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4362_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3869_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_20_9 ), .O(n5252));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3869_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11512 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_46_2 ), 
            .I2(\REG.mem_47_2 ), .I3(rd_addr_r[1]), .O(n13611));
    defparam rd_addr_r_0__bdd_4_lut_11512.LUT_INIT = 16'he4aa;
    SB_LUT4 n12957_bdd_4_lut (.I0(n12957), .I1(n11401), .I2(n12918), .I3(rd_addr_r[4]), 
            .O(n12960));
    defparam n12957_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13611_bdd_4_lut (.I0(n13611), .I1(\REG.mem_45_2 ), .I2(\REG.mem_44_2 ), 
            .I3(rd_addr_r[1]), .O(n13614));
    defparam n13611_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10465 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_7 ), 
            .I2(\REG.mem_15_7 ), .I3(rd_addr_r[1]), .O(n12327));
    defparam rd_addr_r_0__bdd_4_lut_10465.LUT_INIT = 16'he4aa;
    SB_LUT4 i4361_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_49_10 ), .O(n5744));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4361_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3868_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_20_8 ), .O(n5251));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3868_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11542 (.I0(rd_addr_r[3]), .I1(n11769), 
            .I2(n11770), .I3(rd_addr_r[4]), .O(n13605));
    defparam rd_addr_r_3__bdd_4_lut_11542.LUT_INIT = 16'he4aa;
    SB_LUT4 i4360_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_49_9 ), .O(n5743));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4360_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13605_bdd_4_lut (.I0(n13605), .I1(n11749), .I2(n11748), .I3(rd_addr_r[4]), 
            .O(n13608));
    defparam n13605_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF \REG.out_buffer__i12  (.Q(\fifo_data_out[12] ), .C(SLM_CLK_c), 
           .D(n4872));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i13  (.Q(\fifo_data_out[13] ), .C(SLM_CLK_c), 
           .D(n4875));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF i59_60 (.Q(\REG.mem_0_7 ), .C(FIFO_CLK_c), .D(n4932));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3867_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_20_7 ), .O(n5250));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3867_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9554_3_lut (.I0(n12828), .I1(n12330), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11404));
    defparam i9554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11012 (.I0(rd_addr_r[1]), .I1(n11355), 
            .I2(n11356), .I3(rd_addr_r[2]), .O(n12951));
    defparam rd_addr_r_1__bdd_4_lut_11012.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11507 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_26_13 ), 
            .I2(\REG.mem_27_13 ), .I3(rd_addr_r[1]), .O(n13599));
    defparam rd_addr_r_0__bdd_4_lut_11507.LUT_INIT = 16'he4aa;
    SB_LUT4 i3866_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_20_6 ), .O(n5249));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3866_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3865_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_20_5 ), .O(n5248));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3865_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12951_bdd_4_lut (.I0(n12951), .I1(n11326), .I2(n11325), .I3(rd_addr_r[2]), 
            .O(n12954));
    defparam n12951_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3864_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_20_4 ), .O(n5247));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3864_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12327_bdd_4_lut (.I0(n12327), .I1(\REG.mem_13_7 ), .I2(\REG.mem_12_7 ), 
            .I3(rd_addr_r[1]), .O(n12330));
    defparam n12327_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4359_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_49_8 ), .O(n5742));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4359_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3863_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_20_3 ), .O(n5246));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3863_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4358_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_49_7 ), .O(n5741));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4358_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4357_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_49_6 ), .O(n5740));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4357_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3862_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_20_2 ), .O(n5245));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3862_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4356_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_49_5 ), .O(n5739));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4356_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10957 (.I0(rd_addr_r[1]), .I1(n11370), 
            .I2(n11371), .I3(rd_addr_r[2]), .O(n12945));
    defparam rd_addr_r_1__bdd_4_lut_10957.LUT_INIT = 16'he4aa;
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(FIFO_CLK_c), .D(n6034));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 i9568_3_lut (.I0(n12258), .I1(n13716), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11418));
    defparam i9568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13599_bdd_4_lut (.I0(n13599), .I1(\REG.mem_25_13 ), .I2(\REG.mem_24_13 ), 
            .I3(rd_addr_r[1]), .O(n13602));
    defparam n13599_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12945_bdd_4_lut (.I0(n12945), .I1(n11368), .I2(n11367), .I3(rd_addr_r[2]), 
            .O(n12948));
    defparam n12945_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(FIFO_CLK_c), .D(n6033));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 i3861_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_20_1 ), .O(n5244));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3861_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wr_addr_r__i3 (.Q(wr_addr_r[3]), .C(FIFO_CLK_c), .D(n6032));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i4 (.Q(wr_addr_r[4]), .C(FIFO_CLK_c), .D(n6031));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i62_63 (.Q(\REG.mem_0_8 ), .C(FIFO_CLK_c), .D(n4931));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11497 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_3 ), 
            .I2(\REG.mem_11_3 ), .I3(rd_addr_r[1]), .O(n13593));
    defparam rd_addr_r_0__bdd_4_lut_11497.LUT_INIT = 16'he4aa;
    SB_LUT4 i3860_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_20_0 ), .O(n5243));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3860_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3891_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_21_15 ), .O(n5274));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3891_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13593_bdd_4_lut (.I0(n13593), .I1(\REG.mem_9_3 ), .I2(\REG.mem_8_3 ), 
            .I3(rd_addr_r[1]), .O(n10895));
    defparam n13593_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10952 (.I0(rd_addr_r[1]), .I1(n11280), 
            .I2(n11281), .I3(rd_addr_r[2]), .O(n12939));
    defparam rd_addr_r_1__bdd_4_lut_10952.LUT_INIT = 16'he4aa;
    SB_LUT4 i3890_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_21_14 ), .O(n5273));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3890_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3889_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_21_13 ), .O(n5272));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3889_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3888_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_21_12 ), .O(n5271));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3888_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3887_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_21_11 ), .O(n5270));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3887_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10440 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_50_9 ), 
            .I2(\REG.mem_51_9 ), .I3(rd_addr_r[1]), .O(n12309));
    defparam rd_addr_r_0__bdd_4_lut_10440.LUT_INIT = 16'he4aa;
    SB_LUT4 n12939_bdd_4_lut (.I0(n12939), .I1(n11263), .I2(n11262), .I3(rd_addr_r[2]), 
            .O(n12942));
    defparam n12939_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3886_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_21_10 ), .O(n5269));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3886_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wr_addr_r__i5 (.Q(wr_addr_r[5]), .C(FIFO_CLK_c), .D(n6013));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i6131_6132 (.Q(\REG.mem_63_15 ), .C(FIFO_CLK_c), .D(n6012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6128_6129 (.Q(\REG.mem_63_14 ), .C(FIFO_CLK_c), .D(n6011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6125_6126 (.Q(\REG.mem_63_13 ), .C(FIFO_CLK_c), .D(n6010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6122_6123 (.Q(\REG.mem_63_12 ), .C(FIFO_CLK_c), .D(n6009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6119_6120 (.Q(\REG.mem_63_11 ), .C(FIFO_CLK_c), .D(n6008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6116_6117 (.Q(\REG.mem_63_10 ), .C(FIFO_CLK_c), .D(n6007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6113_6114 (.Q(\REG.mem_63_9 ), .C(FIFO_CLK_c), .D(n6006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6110_6111 (.Q(\REG.mem_63_8 ), .C(FIFO_CLK_c), .D(n6005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6107_6108 (.Q(\REG.mem_63_7 ), .C(FIFO_CLK_c), .D(n6004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6104_6105 (.Q(\REG.mem_63_6 ), .C(FIFO_CLK_c), .D(n6003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6101_6102 (.Q(\REG.mem_63_5 ), .C(FIFO_CLK_c), .D(n6002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i65_66 (.Q(\REG.mem_0_9 ), .C(FIFO_CLK_c), .D(n4930));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12309_bdd_4_lut (.I0(n12309), .I1(\REG.mem_49_9 ), .I2(\REG.mem_48_9 ), 
            .I3(rd_addr_r[1]), .O(n12312));
    defparam n12309_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11492 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_42_13 ), 
            .I2(\REG.mem_43_13 ), .I3(rd_addr_r[1]), .O(n13587));
    defparam rd_addr_r_0__bdd_4_lut_11492.LUT_INIT = 16'he4aa;
    SB_LUT4 i3885_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_21_9 ), .O(n5268));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3885_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3884_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_21_8 ), .O(n5267));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3884_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10425 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_38_0 ), 
            .I2(\REG.mem_39_0 ), .I3(rd_addr_r[1]), .O(n12303));
    defparam rd_addr_r_0__bdd_4_lut_10425.LUT_INIT = 16'he4aa;
    SB_LUT4 i3883_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_21_7 ), .O(n5266));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3883_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3882_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_21_6 ), .O(n5265));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3882_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i68_69 (.Q(\REG.mem_0_10 ), .C(FIFO_CLK_c), .D(n4929));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i71_72 (.Q(\REG.mem_0_11 ), .C(FIFO_CLK_c), .D(n4928));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3881_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_21_5 ), .O(n5264));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3881_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i6098_6099 (.Q(\REG.mem_63_4 ), .C(FIFO_CLK_c), .D(n6001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6095_6096 (.Q(\REG.mem_63_3 ), .C(FIFO_CLK_c), .D(n6000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6092_6093 (.Q(\REG.mem_63_2 ), .C(FIFO_CLK_c), .D(n5999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6089_6090 (.Q(\REG.mem_63_1 ), .C(FIFO_CLK_c), .D(n5998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6086_6087 (.Q(\REG.mem_63_0 ), .C(FIFO_CLK_c), .D(n5997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6035_6036 (.Q(\REG.mem_62_15 ), .C(FIFO_CLK_c), .D(n5996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6032_6033 (.Q(\REG.mem_62_14 ), .C(FIFO_CLK_c), .D(n5995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6029_6030 (.Q(\REG.mem_62_13 ), .C(FIFO_CLK_c), .D(n5994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6026_6027 (.Q(\REG.mem_62_12 ), .C(FIFO_CLK_c), .D(n5993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6023_6024 (.Q(\REG.mem_62_11 ), .C(FIFO_CLK_c), .D(n5992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6020_6021 (.Q(\REG.mem_62_10 ), .C(FIFO_CLK_c), .D(n5991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6017_6018 (.Q(\REG.mem_62_9 ), .C(FIFO_CLK_c), .D(n5990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6014_6015 (.Q(\REG.mem_62_8 ), .C(FIFO_CLK_c), .D(n5989));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6011_6012 (.Q(\REG.mem_62_7 ), .C(FIFO_CLK_c), .D(n5988));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6008_6009 (.Q(\REG.mem_62_6 ), .C(FIFO_CLK_c), .D(n5987));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6005_6006 (.Q(\REG.mem_62_5 ), .C(FIFO_CLK_c), .D(n5986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6002_6003 (.Q(\REG.mem_62_4 ), .C(FIFO_CLK_c), .D(n5985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3880_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_21_4 ), .O(n5263));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3880_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13587_bdd_4_lut (.I0(n13587), .I1(\REG.mem_41_13 ), .I2(\REG.mem_40_13 ), 
            .I3(rd_addr_r[1]), .O(n11291));
    defparam n13587_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10947 (.I0(rd_addr_r[1]), .I1(n11340), 
            .I2(n11341), .I3(rd_addr_r[2]), .O(n12933));
    defparam rd_addr_r_1__bdd_4_lut_10947.LUT_INIT = 16'he4aa;
    SB_LUT4 n12933_bdd_4_lut (.I0(n12933), .I1(n11329), .I2(n11328), .I3(rd_addr_r[2]), 
            .O(n12936));
    defparam n12933_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3879_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_21_3 ), .O(n5262));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3879_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12303_bdd_4_lut (.I0(n12303), .I1(\REG.mem_37_0 ), .I2(\REG.mem_36_0 ), 
            .I3(rd_addr_r[1]), .O(n11183));
    defparam n12303_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11487 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_6 ), 
            .I2(\REG.mem_11_6 ), .I3(rd_addr_r[1]), .O(n13581));
    defparam rd_addr_r_0__bdd_4_lut_11487.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10942 (.I0(rd_addr_r[1]), .I1(n11301), 
            .I2(n11302), .I3(rd_addr_r[2]), .O(n12927));
    defparam rd_addr_r_1__bdd_4_lut_10942.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10450 (.I0(rd_addr_r[2]), .I1(n12294), 
            .I2(n11807), .I3(rd_addr_r[3]), .O(n12297));
    defparam rd_addr_r_2__bdd_4_lut_10450.LUT_INIT = 16'he4aa;
    SB_LUT4 n12297_bdd_4_lut (.I0(n12297), .I1(n11183), .I2(n11171), .I3(rd_addr_r[3]), 
            .O(n12300));
    defparam n12297_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5999_6000 (.Q(\REG.mem_62_3 ), .C(FIFO_CLK_c), .D(n5984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5996_5997 (.Q(\REG.mem_62_2 ), .C(FIFO_CLK_c), .D(n5983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5993_5994 (.Q(\REG.mem_62_1 ), .C(FIFO_CLK_c), .D(n5982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5990_5991 (.Q(\REG.mem_62_0 ), .C(FIFO_CLK_c), .D(n5981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5939_5940 (.Q(\REG.mem_61_15 ), .C(FIFO_CLK_c), .D(n5979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5936_5937 (.Q(\REG.mem_61_14 ), .C(FIFO_CLK_c), .D(n5978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5933_5934 (.Q(\REG.mem_61_13 ), .C(FIFO_CLK_c), .D(n5977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5930_5931 (.Q(\REG.mem_61_12 ), .C(FIFO_CLK_c), .D(n5976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5927_5928 (.Q(\REG.mem_61_11 ), .C(FIFO_CLK_c), .D(n5975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5924_5925 (.Q(\REG.mem_61_10 ), .C(FIFO_CLK_c), .D(n5974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5921_5922 (.Q(\REG.mem_61_9 ), .C(FIFO_CLK_c), .D(n5973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5918_5919 (.Q(\REG.mem_61_8 ), .C(FIFO_CLK_c), .D(n5972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5915_5916 (.Q(\REG.mem_61_7 ), .C(FIFO_CLK_c), .D(n5971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5912_5913 (.Q(\REG.mem_61_6 ), .C(FIFO_CLK_c), .D(n5970));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5909_5910 (.Q(\REG.mem_61_5 ), .C(FIFO_CLK_c), .D(n5969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13581_bdd_4_lut (.I0(n13581), .I1(\REG.mem_9_6 ), .I2(\REG.mem_8_6 ), 
            .I3(rd_addr_r[1]), .O(n10853));
    defparam n13581_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12927_bdd_4_lut (.I0(n12927), .I1(n11299), .I2(n11298), .I3(rd_addr_r[2]), 
            .O(n12930));
    defparam n12927_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3878_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_21_2 ), .O(n5261));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3878_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3877_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_21_1 ), .O(n5260));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3877_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10420 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_42_0 ), 
            .I2(\REG.mem_43_0 ), .I3(rd_addr_r[1]), .O(n12291));
    defparam rd_addr_r_0__bdd_4_lut_10420.LUT_INIT = 16'he4aa;
    SB_LUT4 i3876_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_21_0 ), .O(n5259));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3876_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11482 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_22_8 ), 
            .I2(\REG.mem_23_8 ), .I3(rd_addr_r[1]), .O(n13575));
    defparam rd_addr_r_0__bdd_4_lut_11482.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10937 (.I0(rd_addr_r[1]), .I1(n11094), 
            .I2(n11095), .I3(rd_addr_r[2]), .O(n12921));
    defparam rd_addr_r_1__bdd_4_lut_10937.LUT_INIT = 16'he4aa;
    SB_LUT4 i3945_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_24_15 ), .O(n5328));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3945_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12921_bdd_4_lut (.I0(n12921), .I1(n11053), .I2(n11052), .I3(rd_addr_r[2]), 
            .O(n12924));
    defparam n12921_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3944_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_24_14 ), .O(n5327));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3944_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4355_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_49_4 ), .O(n5738));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4355_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10932 (.I0(rd_addr_r[1]), .I1(n11274), 
            .I2(n11275), .I3(rd_addr_r[2]), .O(n12915));
    defparam rd_addr_r_1__bdd_4_lut_10932.LUT_INIT = 16'he4aa;
    SB_DFF i5906_5907 (.Q(\REG.mem_61_4 ), .C(FIFO_CLK_c), .D(n5968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5903_5904 (.Q(\REG.mem_61_3 ), .C(FIFO_CLK_c), .D(n5967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5900_5901 (.Q(\REG.mem_61_2 ), .C(FIFO_CLK_c), .D(n5966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5897_5898 (.Q(\REG.mem_61_1 ), .C(FIFO_CLK_c), .D(n5965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5894_5895 (.Q(\REG.mem_61_0 ), .C(FIFO_CLK_c), .D(n5964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5843_5844 (.Q(\REG.mem_60_15 ), .C(FIFO_CLK_c), .D(n5962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5840_5841 (.Q(\REG.mem_60_14 ), .C(FIFO_CLK_c), .D(n5961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5837_5838 (.Q(\REG.mem_60_13 ), .C(FIFO_CLK_c), .D(n5960));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5834_5835 (.Q(\REG.mem_60_12 ), .C(FIFO_CLK_c), .D(n5959));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5831_5832 (.Q(\REG.mem_60_11 ), .C(FIFO_CLK_c), .D(n5958));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5828_5829 (.Q(\REG.mem_60_10 ), .C(FIFO_CLK_c), .D(n5957));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5825_5826 (.Q(\REG.mem_60_9 ), .C(FIFO_CLK_c), .D(n5956));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5822_5823 (.Q(\REG.mem_60_8 ), .C(FIFO_CLK_c), .D(n5955));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5819_5820 (.Q(\REG.mem_60_7 ), .C(FIFO_CLK_c), .D(n5954));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5816_5817 (.Q(\REG.mem_60_6 ), .C(FIFO_CLK_c), .D(n5953));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13575_bdd_4_lut (.I0(n13575), .I1(\REG.mem_21_8 ), .I2(\REG.mem_20_8 ), 
            .I3(rd_addr_r[1]), .O(n13578));
    defparam n13575_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12915_bdd_4_lut (.I0(n12915), .I1(n11266), .I2(n11265), .I3(rd_addr_r[2]), 
            .O(n12918));
    defparam n12915_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5813_5814 (.Q(\REG.mem_60_5 ), .C(FIFO_CLK_c), .D(n5952));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5810_5811 (.Q(\REG.mem_60_4 ), .C(FIFO_CLK_c), .D(n5951));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5807_5808 (.Q(\REG.mem_60_3 ), .C(FIFO_CLK_c), .D(n5950));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5804_5805 (.Q(\REG.mem_60_2 ), .C(FIFO_CLK_c), .D(n5949));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5801_5802 (.Q(\REG.mem_60_1 ), .C(FIFO_CLK_c), .D(n5948));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5798_5799 (.Q(\REG.mem_60_0 ), .C(FIFO_CLK_c), .D(n5947));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync1_r__i1 (.Q(rp_sync1_r[1]), .C(FIFO_CLK_c), .D(n5946));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i2 (.Q(rp_sync1_r[2]), .C(FIFO_CLK_c), .D(n5945));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i3 (.Q(rp_sync1_r[3]), .C(FIFO_CLK_c), .D(n5944));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i4 (.Q(rp_sync1_r[4]), .C(FIFO_CLK_c), .D(n5943));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i5 (.Q(rp_sync1_r[5]), .C(FIFO_CLK_c), .D(n5942));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i6 (.Q(rp_sync1_r[6]), .C(FIFO_CLK_c), .D(n5941));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i1 (.Q(rp_sync2_r[1]), .C(FIFO_CLK_c), .D(n5940));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i2 (.Q(rp_sync2_r[2]), .C(FIFO_CLK_c), .D(n5939));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i3 (.Q(rp_sync2_r[3]), .C(FIFO_CLK_c), .D(n5938));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i5747_5748 (.Q(\REG.mem_59_15 ), .C(FIFO_CLK_c), .D(n5937));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3943_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_24_13 ), .O(n5326));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3943_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3942_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_24_12 ), .O(n5325));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3942_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11532 (.I0(rd_addr_r[2]), .I1(n12552), 
            .I2(n12468), .I3(rd_addr_r[3]), .O(n13569));
    defparam rd_addr_r_2__bdd_4_lut_11532.LUT_INIT = 16'he4aa;
    SB_DFF i5744_5745 (.Q(\REG.mem_59_14 ), .C(FIFO_CLK_c), .D(n5936));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13569_bdd_4_lut (.I0(n13569), .I1(n12804), .I2(n12978), .I3(rd_addr_r[3]), 
            .O(n11789));
    defparam n13569_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9391_3_lut (.I0(n13056), .I1(n12816), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11241));
    defparam i9391_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5741_5742 (.Q(\REG.mem_59_13 ), .C(FIFO_CLK_c), .D(n5935));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5738_5739 (.Q(\REG.mem_59_12 ), .C(FIFO_CLK_c), .D(n5934));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5735_5736 (.Q(\REG.mem_59_11 ), .C(FIFO_CLK_c), .D(n5933));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5732_5733 (.Q(\REG.mem_59_10 ), .C(FIFO_CLK_c), .D(n5932));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5729_5730 (.Q(\REG.mem_59_9 ), .C(FIFO_CLK_c), .D(n5931));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5726_5727 (.Q(\REG.mem_59_8 ), .C(FIFO_CLK_c), .D(n5930));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5723_5724 (.Q(\REG.mem_59_7 ), .C(FIFO_CLK_c), .D(n5929));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5720_5721 (.Q(\REG.mem_59_6 ), .C(FIFO_CLK_c), .D(n5928));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5717_5718 (.Q(\REG.mem_59_5 ), .C(FIFO_CLK_c), .D(n5927));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5714_5715 (.Q(\REG.mem_59_4 ), .C(FIFO_CLK_c), .D(n5926));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5711_5712 (.Q(\REG.mem_59_3 ), .C(FIFO_CLK_c), .D(n5925));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5708_5709 (.Q(\REG.mem_59_2 ), .C(FIFO_CLK_c), .D(n5924));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5705_5706 (.Q(\REG.mem_59_1 ), .C(FIFO_CLK_c), .D(n5923));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5702_5703 (.Q(\REG.mem_59_0 ), .C(FIFO_CLK_c), .D(n5922));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync2_r__i4 (.Q(rp_sync2_r[4]), .C(FIFO_CLK_c), .D(n5921));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i5 (.Q(rp_sync2_r[5]), .C(FIFO_CLK_c), .D(n5920));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i6 (.Q(rp_sync2_r[6]), .C(FIFO_CLK_c), .D(n5919));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(n5918));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF i74_75 (.Q(\REG.mem_0_12 ), .C(FIFO_CLK_c), .D(n4927));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9392_3_lut (.I0(n12720), .I1(n12564), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11242));
    defparam i9392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9401_3_lut (.I0(n12150), .I1(n13728), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11251));
    defparam i9401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12291_bdd_4_lut (.I0(n12291), .I1(\REG.mem_41_0 ), .I2(\REG.mem_40_0 ), 
            .I3(rd_addr_r[1]), .O(n12294));
    defparam n12291_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9400_3_lut (.I0(n12312), .I1(n12234), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11250));
    defparam i9400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11477 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_26_1 ), 
            .I2(\REG.mem_27_1 ), .I3(rd_addr_r[1]), .O(n13563));
    defparam rd_addr_r_0__bdd_4_lut_11477.LUT_INIT = 16'he4aa;
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .D(n5917));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i3 (.Q(rd_addr_r[3]), .C(SLM_CLK_c), .D(n5916));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_LUT4 i9020_3_lut (.I0(n13620), .I1(n13614), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10870));
    defparam i9020_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF rd_addr_r__i4 (.Q(rd_addr_r[4]), .C(SLM_CLK_c), .D(n5915));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i5 (.Q(rd_addr_r[5]), .C(SLM_CLK_c), .D(n5914));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i6 (.Q(\rd_addr_r[6] ), .C(SLM_CLK_c), .D(n5913));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF i5651_5652 (.Q(\REG.mem_58_15 ), .C(FIFO_CLK_c), .D(n5912));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5648_5649 (.Q(\REG.mem_58_14 ), .C(FIFO_CLK_c), .D(n5911));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5645_5646 (.Q(\REG.mem_58_13 ), .C(FIFO_CLK_c), .D(n5910));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5642_5643 (.Q(\REG.mem_58_12 ), .C(FIFO_CLK_c), .D(n5909));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5639_5640 (.Q(\REG.mem_58_11 ), .C(FIFO_CLK_c), .D(n5908));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5636_5637 (.Q(\REG.mem_58_10 ), .C(FIFO_CLK_c), .D(n5907));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5633_5634 (.Q(\REG.mem_58_9 ), .C(FIFO_CLK_c), .D(n5906));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5630_5631 (.Q(\REG.mem_58_8 ), .C(FIFO_CLK_c), .D(n5905));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5627_5628 (.Q(\REG.mem_58_7 ), .C(FIFO_CLK_c), .D(n5904));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5624_5625 (.Q(\REG.mem_58_6 ), .C(FIFO_CLK_c), .D(n5903));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5621_5622 (.Q(\REG.mem_58_5 ), .C(FIFO_CLK_c), .D(n5902));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10962 (.I0(rd_addr_r[3]), .I1(n11322), 
            .I2(n11323), .I3(rd_addr_r[4]), .O(n12909));
    defparam rd_addr_r_3__bdd_4_lut_10962.LUT_INIT = 16'he4aa;
    SB_LUT4 i9023_3_lut (.I0(n13548), .I1(n13524), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10873));
    defparam i9023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3941_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_24_11 ), .O(n5324));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3941_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4354_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_49_3 ), .O(n5737));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4354_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10415 (.I0(rd_addr_r[2]), .I1(n11444), 
            .I2(n11465), .I3(rd_addr_r[3]), .O(n12285));
    defparam rd_addr_r_2__bdd_4_lut_10415.LUT_INIT = 16'he4aa;
    SB_LUT4 i9856_3_lut (.I0(\REG.mem_8_14 ), .I1(\REG.mem_9_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11706));
    defparam i9856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13563_bdd_4_lut (.I0(n13563), .I1(\REG.mem_25_1 ), .I2(\REG.mem_24_1 ), 
            .I3(rd_addr_r[1]), .O(n13566));
    defparam n13563_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3940_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_24_10 ), .O(n5323));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3940_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9857_3_lut (.I0(\REG.mem_10_14 ), .I1(\REG.mem_11_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11707));
    defparam i9857_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5618_5619 (.Q(\REG.mem_58_4 ), .C(FIFO_CLK_c), .D(n5901));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5615_5616 (.Q(\REG.mem_58_3 ), .C(FIFO_CLK_c), .D(n5900));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5612_5613 (.Q(\REG.mem_58_2 ), .C(FIFO_CLK_c), .D(n5899));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5609_5610 (.Q(\REG.mem_58_1 ), .C(FIFO_CLK_c), .D(n5898));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5606_5607 (.Q(\REG.mem_58_0 ), .C(FIFO_CLK_c), .D(n5897));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5555_5556 (.Q(\REG.mem_57_15 ), .C(FIFO_CLK_c), .D(n5894));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5552_5553 (.Q(\REG.mem_57_14 ), .C(FIFO_CLK_c), .D(n5893));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5549_5550 (.Q(\REG.mem_57_13 ), .C(FIFO_CLK_c), .D(n5892));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5546_5547 (.Q(\REG.mem_57_12 ), .C(FIFO_CLK_c), .D(n5891));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5543_5544 (.Q(\REG.mem_57_11 ), .C(FIFO_CLK_c), .D(n5890));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5540_5541 (.Q(\REG.mem_57_10 ), .C(FIFO_CLK_c), .D(n5889));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5537_5538 (.Q(\REG.mem_57_9 ), .C(FIFO_CLK_c), .D(n5888));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5534_5535 (.Q(\REG.mem_57_8 ), .C(FIFO_CLK_c), .D(n5887));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5531_5532 (.Q(\REG.mem_57_7 ), .C(FIFO_CLK_c), .D(n5886));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3939_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_24_9 ), .O(n5322));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3939_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3938_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_24_8 ), .O(n5321));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3938_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12909_bdd_4_lut (.I0(n12909), .I1(n11311), .I2(n12888), .I3(rd_addr_r[4]), 
            .O(n12912));
    defparam n12909_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12285_bdd_4_lut (.I0(n12285), .I1(n11396), .I2(n11381), .I3(rd_addr_r[3]), 
            .O(n11633));
    defparam n12285_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11467 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_6_8 ), 
            .I2(\REG.mem_7_8 ), .I3(rd_addr_r[1]), .O(n13557));
    defparam rd_addr_r_0__bdd_4_lut_11467.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10410 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_38_15 ), 
            .I2(\REG.mem_39_15 ), .I3(rd_addr_r[1]), .O(n12279));
    defparam rd_addr_r_0__bdd_4_lut_10410.LUT_INIT = 16'he4aa;
    SB_DFF i5528_5529 (.Q(\REG.mem_57_6 ), .C(FIFO_CLK_c), .D(n5885));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13557_bdd_4_lut (.I0(n13557), .I1(\REG.mem_5_8 ), .I2(\REG.mem_4_8 ), 
            .I3(rd_addr_r[1]), .O(n13560));
    defparam n13557_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3937_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_24_7 ), .O(n5320));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3937_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9860_3_lut (.I0(\REG.mem_14_14 ), .I1(\REG.mem_15_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11710));
    defparam i9860_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5525_5526 (.Q(\REG.mem_57_5 ), .C(FIFO_CLK_c), .D(n5884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5522_5523 (.Q(\REG.mem_57_4 ), .C(FIFO_CLK_c), .D(n5883));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5519_5520 (.Q(\REG.mem_57_3 ), .C(FIFO_CLK_c), .D(n5882));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5516_5517 (.Q(\REG.mem_57_2 ), .C(FIFO_CLK_c), .D(n5881));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5513_5514 (.Q(\REG.mem_57_1 ), .C(FIFO_CLK_c), .D(n5880));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5510_5511 (.Q(\REG.mem_57_0 ), .C(FIFO_CLK_c), .D(n5879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5459_5460 (.Q(\REG.mem_56_15 ), .C(FIFO_CLK_c), .D(n5878));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5456_5457 (.Q(\REG.mem_56_14 ), .C(FIFO_CLK_c), .D(n5877));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5453_5454 (.Q(\REG.mem_56_13 ), .C(FIFO_CLK_c), .D(n5876));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5450_5451 (.Q(\REG.mem_56_12 ), .C(FIFO_CLK_c), .D(n5875));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5447_5448 (.Q(\REG.mem_56_11 ), .C(FIFO_CLK_c), .D(n5874));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5444_5445 (.Q(\REG.mem_56_10 ), .C(FIFO_CLK_c), .D(n5873));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5441_5442 (.Q(\REG.mem_56_9 ), .C(FIFO_CLK_c), .D(n5872));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5438_5439 (.Q(\REG.mem_56_8 ), .C(FIFO_CLK_c), .D(n5871));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5435_5436 (.Q(\REG.mem_56_7 ), .C(FIFO_CLK_c), .D(n5870));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5432_5433 (.Q(\REG.mem_56_6 ), .C(FIFO_CLK_c), .D(n5869));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9859_3_lut (.I0(\REG.mem_12_14 ), .I1(\REG.mem_13_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11709));
    defparam i9859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9238_3_lut (.I0(\REG.mem_56_4 ), .I1(\REG.mem_57_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11088));
    defparam i9238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10927 (.I0(rd_addr_r[1]), .I1(n11253), 
            .I2(n11254), .I3(rd_addr_r[2]), .O(n12903));
    defparam rd_addr_r_1__bdd_4_lut_10927.LUT_INIT = 16'he4aa;
    SB_LUT4 i9239_3_lut (.I0(\REG.mem_58_4 ), .I1(\REG.mem_59_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11089));
    defparam i9239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12279_bdd_4_lut (.I0(n12279), .I1(\REG.mem_37_15 ), .I2(\REG.mem_36_15 ), 
            .I3(rd_addr_r[1]), .O(n12282));
    defparam n12279_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9242_3_lut (.I0(\REG.mem_62_4 ), .I1(\REG.mem_63_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11092));
    defparam i9242_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5429_5430 (.Q(\REG.mem_56_5 ), .C(FIFO_CLK_c), .D(n5868));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5426_5427 (.Q(\REG.mem_56_4 ), .C(FIFO_CLK_c), .D(n5867));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5423_5424 (.Q(\REG.mem_56_3 ), .C(FIFO_CLK_c), .D(n5866));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5420_5421 (.Q(\REG.mem_56_2 ), .C(FIFO_CLK_c), .D(n5865));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5417_5418 (.Q(\REG.mem_56_1 ), .C(FIFO_CLK_c), .D(n5864));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5414_5415 (.Q(\REG.mem_56_0 ), .C(FIFO_CLK_c), .D(n5862));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wp_sync1_r__i1 (.Q(wp_sync1_r[1]), .C(SLM_CLK_c), .D(n5861));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i2 (.Q(wp_sync1_r[2]), .C(SLM_CLK_c), .D(n5860));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i3 (.Q(wp_sync1_r[3]), .C(SLM_CLK_c), .D(n5859));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i4 (.Q(wp_sync1_r[4]), .C(SLM_CLK_c), .D(n5858));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i5 (.Q(wp_sync1_r[5]), .C(SLM_CLK_c), .D(n5857));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i6 (.Q(wp_sync1_r[6]), .C(SLM_CLK_c), .D(n5856));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i5363_5364 (.Q(\REG.mem_55_15 ), .C(FIFO_CLK_c), .D(n5855));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5360_5361 (.Q(\REG.mem_55_14 ), .C(FIFO_CLK_c), .D(n5854));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5357_5358 (.Q(\REG.mem_55_13 ), .C(FIFO_CLK_c), .D(n5853));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_6__I_0_141_7 (.CI(n10009), .I0(wr_addr_r[5]), .I1(GND_net), 
            .CO(n10010));
    SB_LUT4 i9241_3_lut (.I0(\REG.mem_60_4 ), .I1(\REG.mem_61_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11091));
    defparam i9241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_141_6_lut (.I0(GND_net), .I1(wr_addr_r[4]), 
            .I2(GND_net), .I3(n10008), .O(wr_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_6 (.CI(n10008), .I0(wr_addr_r[4]), .I1(GND_net), 
            .CO(n10009));
    SB_LUT4 wr_addr_r_6__I_0_141_5_lut (.I0(GND_net), .I1(wr_addr_r[3]), 
            .I2(GND_net), .I3(n10007), .O(wr_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_5 (.CI(n10007), .I0(wr_addr_r[3]), .I1(GND_net), 
            .CO(n10008));
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_3 (.CI(n9962), .I0(wp_sync_w[1]), 
            .I1(n1[1]), .CO(n9963));
    SB_LUT4 wr_addr_r_6__I_0_141_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(GND_net), .I3(n10006), .O(wr_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_2_lut (.I0(GND_net), .I1(wp_sync_w[0]), 
            .I2(n1[0]), .I3(VCC_net), .O(\rd_sig_diff0_w[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_4 (.CI(n10006), .I0(wr_addr_r[2]), .I1(GND_net), 
            .CO(n10007));
    SB_DFF i5354_5355 (.Q(\REG.mem_55_12 ), .C(FIFO_CLK_c), .D(n5852));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5351_5352 (.Q(\REG.mem_55_11 ), .C(FIFO_CLK_c), .D(n5851));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5348_5349 (.Q(\REG.mem_55_10 ), .C(FIFO_CLK_c), .D(n5850));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5345_5346 (.Q(\REG.mem_55_9 ), .C(FIFO_CLK_c), .D(n5849));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5342_5343 (.Q(\REG.mem_55_8 ), .C(FIFO_CLK_c), .D(n5848));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5339_5340 (.Q(\REG.mem_55_7 ), .C(FIFO_CLK_c), .D(n5847));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5336_5337 (.Q(\REG.mem_55_6 ), .C(FIFO_CLK_c), .D(n5846));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5333_5334 (.Q(\REG.mem_55_5 ), .C(FIFO_CLK_c), .D(n5845));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5330_5331 (.Q(\REG.mem_55_4 ), .C(FIFO_CLK_c), .D(n5844));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5327_5328 (.Q(\REG.mem_55_3 ), .C(FIFO_CLK_c), .D(n5843));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5324_5325 (.Q(\REG.mem_55_2 ), .C(FIFO_CLK_c), .D(n5842));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5321_5322 (.Q(\REG.mem_55_1 ), .C(FIFO_CLK_c), .D(n5841));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5318_5319 (.Q(\REG.mem_55_0 ), .C(FIFO_CLK_c), .D(n5840));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wp_sync2_r__i1 (.Q(wp_sync2_r[1]), .C(SLM_CLK_c), .D(n5839));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i2 (.Q(wp_sync2_r[2]), .C(SLM_CLK_c), .D(n5838));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 wr_addr_r_6__I_0_141_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), 
            .I2(GND_net), .I3(n10005), .O(wr_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_6__I_0_151_8_lut (.I0(GND_net), .I1(\rd_addr_r[6] ), 
            .I2(GND_net), .I3(n10016), .O(rd_addr_p1_w[6])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_3 (.CI(n10005), .I0(wr_addr_r[1]), .I1(GND_net), 
            .CO(n10006));
    SB_LUT4 wr_addr_r_6__I_0_141_2_lut (.I0(GND_net), .I1(wr_addr_r[0]), 
            .I2(GND_net), .I3(VCC_net), .O(wr_addr_p1_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_6__I_0_151_7_lut (.I0(GND_net), .I1(rd_addr_r[5]), 
            .I2(GND_net), .I3(n10015), .O(rd_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_141_2 (.CI(VCC_net), .I0(wr_addr_r[0]), .I1(GND_net), 
            .CO(n10005));
    SB_CARRY rd_addr_r_6__I_0_151_7 (.CI(n10015), .I0(rd_addr_r[5]), .I1(GND_net), 
            .CO(n10016));
    SB_LUT4 i9217_3_lut (.I0(\REG.mem_40_4 ), .I1(\REG.mem_41_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11067));
    defparam i9217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_8_lut (.I0(n10828), .I1(wr_grey_sync_r[6]), 
            .I2(n1_adj_1212[6]), .I3(n9973), .O(\afull_flag_impl.af_flag_nxt_w )) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i9218_3_lut (.I0(\REG.mem_42_4 ), .I1(\REG.mem_43_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11068));
    defparam i9218_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF wp_sync2_r__i3 (.Q(wp_sync2_r[3]), .C(SLM_CLK_c), .D(n5836));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i4 (.Q(wp_sync2_r[4]), .C(SLM_CLK_c), .D(n5835));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i5 (.Q(wp_sync2_r[5]), .C(SLM_CLK_c), .D(n5834));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i6 (.Q(wp_sync2_r[6]), .C(SLM_CLK_c), .D(n5833));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i5267_5268 (.Q(\REG.mem_54_15 ), .C(FIFO_CLK_c), .D(n5832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5264_5265 (.Q(\REG.mem_54_14 ), .C(FIFO_CLK_c), .D(n5831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5261_5262 (.Q(\REG.mem_54_13 ), .C(FIFO_CLK_c), .D(n5830));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5258_5259 (.Q(\REG.mem_54_12 ), .C(FIFO_CLK_c), .D(n5829));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5255_5256 (.Q(\REG.mem_54_11 ), .C(FIFO_CLK_c), .D(n5828));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5252_5253 (.Q(\REG.mem_54_10 ), .C(FIFO_CLK_c), .D(n5827));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5249_5250 (.Q(\REG.mem_54_9 ), .C(FIFO_CLK_c), .D(n5826));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5246_5247 (.Q(\REG.mem_54_8 ), .C(FIFO_CLK_c), .D(n5825));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5243_5244 (.Q(\REG.mem_54_7 ), .C(FIFO_CLK_c), .D(n5824));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5240_5241 (.Q(\REG.mem_54_6 ), .C(FIFO_CLK_c), .D(n5823));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5237_5238 (.Q(\REG.mem_54_5 ), .C(FIFO_CLK_c), .D(n5822));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5234_5235 (.Q(\REG.mem_54_4 ), .C(FIFO_CLK_c), .D(n5821));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_r_6__I_0_add_2_7_lut (.I0(n10798), .I1(wr_addr_r[5]), 
            .I2(rp_sync_w[5]), .I3(n9972), .O(n10828)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY wr_addr_r_6__I_0_add_2_7 (.CI(n9972), .I0(wr_addr_r[5]), .I1(rp_sync_w[5]), 
            .CO(n9973));
    SB_LUT4 rd_addr_r_6__I_0_151_6_lut (.I0(GND_net), .I1(rd_addr_r[4]), 
            .I2(GND_net), .I3(n10014), .O(rd_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wr_addr_r_6__I_0_add_2_6_lut (.I0(n2_adj_1188), .I1(wr_addr_r[4]), 
            .I2(rp_sync_w[4]), .I3(n9971), .O(n10778)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_6_lut.LUT_INIT = 16'hebbe;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_2 (.CI(VCC_net), .I0(wp_sync_w[0]), 
            .I1(n1[0]), .CO(n9962));
    SB_CARRY wr_addr_r_6__I_0_add_2_6 (.CI(n9971), .I0(wr_addr_r[4]), .I1(rp_sync_w[4]), 
            .CO(n9972));
    SB_LUT4 i9221_3_lut (.I0(\REG.mem_46_4 ), .I1(\REG.mem_47_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11071));
    defparam i9221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_5_lut (.I0(GND_net), .I1(wr_addr_r[3]), 
            .I2(rp_sync_w[3]), .I3(n9970), .O(wr_sig_diff0_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_add_2_5 (.CI(n9970), .I0(wr_addr_r[3]), .I1(rp_sync_w[3]), 
            .CO(n9971));
    SB_LUT4 n12903_bdd_4_lut (.I0(n12903), .I1(n11236), .I2(n11235), .I3(rd_addr_r[2]), 
            .O(n12906));
    defparam n12903_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9220_3_lut (.I0(\REG.mem_44_4 ), .I1(\REG.mem_45_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11070));
    defparam i9220_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_6__I_0_151_6 (.CI(n10014), .I0(rd_addr_r[4]), .I1(GND_net), 
            .CO(n10015));
    SB_DFF i5231_5232 (.Q(\REG.mem_54_3 ), .C(FIFO_CLK_c), .D(n5820));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5228_5229 (.Q(\REG.mem_54_2 ), .C(FIFO_CLK_c), .D(n5819));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5225_5226 (.Q(\REG.mem_54_1 ), .C(FIFO_CLK_c), .D(n5818));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5222_5223 (.Q(\REG.mem_54_0 ), .C(FIFO_CLK_c), .D(n5817));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5171_5172 (.Q(\REG.mem_53_15 ), .C(FIFO_CLK_c), .D(n5816));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5168_5169 (.Q(\REG.mem_53_14 ), .C(FIFO_CLK_c), .D(n5815));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5165_5166 (.Q(\REG.mem_53_13 ), .C(FIFO_CLK_c), .D(n5814));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5162_5163 (.Q(\REG.mem_53_12 ), .C(FIFO_CLK_c), .D(n5813));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5159_5160 (.Q(\REG.mem_53_11 ), .C(FIFO_CLK_c), .D(n5812));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5156_5157 (.Q(\REG.mem_53_10 ), .C(FIFO_CLK_c), .D(n5811));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5153_5154 (.Q(\REG.mem_53_9 ), .C(FIFO_CLK_c), .D(n5810));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5150_5151 (.Q(\REG.mem_53_8 ), .C(FIFO_CLK_c), .D(n5809));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5147_5148 (.Q(\REG.mem_53_7 ), .C(FIFO_CLK_c), .D(n5808));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5144_5145 (.Q(\REG.mem_53_6 ), .C(FIFO_CLK_c), .D(n5807));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5141_5142 (.Q(\REG.mem_53_5 ), .C(FIFO_CLK_c), .D(n5806));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5138_5139 (.Q(\REG.mem_53_4 ), .C(FIFO_CLK_c), .D(n5805));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4089_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_33_15 ), .O(n5472));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4089_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9193_3_lut (.I0(\REG.mem_24_4 ), .I1(\REG.mem_25_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11043));
    defparam i9193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_6__I_0_151_5_lut (.I0(GND_net), .I1(rd_addr_r[3]), 
            .I2(GND_net), .I3(n10013), .O(rd_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9194_3_lut (.I0(\REG.mem_26_4 ), .I1(\REG.mem_27_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11044));
    defparam i9194_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rd_addr_r_6__I_0_151_5 (.CI(n10013), .I0(rd_addr_r[3]), .I1(GND_net), 
            .CO(n10014));
    SB_DFF i5135_5136 (.Q(\REG.mem_53_3 ), .C(FIFO_CLK_c), .D(n5804));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5132_5133 (.Q(\REG.mem_53_2 ), .C(FIFO_CLK_c), .D(n5803));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5129_5130 (.Q(\REG.mem_53_1 ), .C(FIFO_CLK_c), .D(n5802));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5126_5127 (.Q(\REG.mem_53_0 ), .C(FIFO_CLK_c), .D(n5801));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5075_5076 (.Q(\REG.mem_52_15 ), .C(FIFO_CLK_c), .D(n5800));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5072_5073 (.Q(\REG.mem_52_14 ), .C(FIFO_CLK_c), .D(n5799));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5069_5070 (.Q(\REG.mem_52_13 ), .C(FIFO_CLK_c), .D(n5798));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5066_5067 (.Q(\REG.mem_52_12 ), .C(FIFO_CLK_c), .D(n5797));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5063_5064 (.Q(\REG.mem_52_11 ), .C(FIFO_CLK_c), .D(n5796));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5060_5061 (.Q(\REG.mem_52_10 ), .C(FIFO_CLK_c), .D(n5795));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5057_5058 (.Q(\REG.mem_52_9 ), .C(FIFO_CLK_c), .D(n5794));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5054_5055 (.Q(\REG.mem_52_8 ), .C(FIFO_CLK_c), .D(n5793));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5051_5052 (.Q(\REG.mem_52_7 ), .C(FIFO_CLK_c), .D(n5792));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5048_5049 (.Q(\REG.mem_52_6 ), .C(FIFO_CLK_c), .D(n5791));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5045_5046 (.Q(\REG.mem_52_5 ), .C(FIFO_CLK_c), .D(n5790));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5042_5043 (.Q(\REG.mem_52_4 ), .C(FIFO_CLK_c), .D(n5789));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9200_3_lut (.I0(\REG.mem_30_4 ), .I1(\REG.mem_31_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11050));
    defparam i9200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3936_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_24_6 ), .O(n5319));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3936_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9199_3_lut (.I0(\REG.mem_28_4 ), .I1(\REG.mem_29_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11049));
    defparam i9199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9169_3_lut (.I0(\REG.mem_8_4 ), .I1(\REG.mem_9_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11019));
    defparam i9169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(rp_sync_w[2]), .I3(n9969), .O(wr_sig_diff0_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF i5039_5040 (.Q(\REG.mem_52_3 ), .C(FIFO_CLK_c), .D(n5788));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_6__I_0_add_2_4 (.CI(n9969), .I0(wr_addr_r[2]), .I1(rp_sync_w[2]), 
            .CO(n9970));
    SB_DFF i5036_5037 (.Q(\REG.mem_52_2 ), .C(FIFO_CLK_c), .D(n5787));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5033_5034 (.Q(\REG.mem_52_1 ), .C(FIFO_CLK_c), .D(n5786));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5030_5031 (.Q(\REG.mem_52_0 ), .C(FIFO_CLK_c), .D(n5785));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4979_4980 (.Q(\REG.mem_51_15 ), .C(FIFO_CLK_c), .D(n5784));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4976_4977 (.Q(\REG.mem_51_14 ), .C(FIFO_CLK_c), .D(n5783));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4973_4974 (.Q(\REG.mem_51_13 ), .C(FIFO_CLK_c), .D(n5782));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4970_4971 (.Q(\REG.mem_51_12 ), .C(FIFO_CLK_c), .D(n5781));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4967_4968 (.Q(\REG.mem_51_11 ), .C(FIFO_CLK_c), .D(n5780));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4964_4965 (.Q(\REG.mem_51_10 ), .C(FIFO_CLK_c), .D(n5779));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4961_4962 (.Q(\REG.mem_51_9 ), .C(FIFO_CLK_c), .D(n5778));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4958_4959 (.Q(\REG.mem_51_8 ), .C(FIFO_CLK_c), .D(n5777));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4955_4956 (.Q(\REG.mem_51_7 ), .C(FIFO_CLK_c), .D(n5776));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4952_4953 (.Q(\REG.mem_51_6 ), .C(FIFO_CLK_c), .D(n5775));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4949_4950 (.Q(\REG.mem_51_5 ), .C(FIFO_CLK_c), .D(n5774));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4946_4947 (.Q(\REG.mem_51_4 ), .C(FIFO_CLK_c), .D(n5773));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9170_3_lut (.I0(\REG.mem_10_4 ), .I1(\REG.mem_11_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11020));
    defparam i9170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), 
            .I2(rp_sync_w[1]), .I3(n9968), .O(wr_sig_diff0_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_add_2_3 (.CI(n9968), .I0(wr_addr_r[1]), .I1(rp_sync_w[1]), 
            .CO(n9969));
    SB_LUT4 i9173_3_lut (.I0(\REG.mem_14_4 ), .I1(\REG.mem_15_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11023));
    defparam i9173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9172_3_lut (.I0(\REG.mem_12_4 ), .I1(\REG.mem_13_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11022));
    defparam i9172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_6__I_0_151_4_lut (.I0(GND_net), .I1(rd_addr_r[2]), 
            .I2(GND_net), .I3(n10012), .O(rd_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wr_addr_r_6__I_0_add_2_2_lut (.I0(GND_net), .I1(wr_addr_r[0]), 
            .I2(rp_sync_w[0]), .I3(VCC_net), .O(wr_sig_diff0_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF i4943_4944 (.Q(\REG.mem_51_3 ), .C(FIFO_CLK_c), .D(n5772));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4940_4941 (.Q(\REG.mem_51_2 ), .C(FIFO_CLK_c), .D(n5771));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4937_4938 (.Q(\REG.mem_51_1 ), .C(FIFO_CLK_c), .D(n5770));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4934_4935 (.Q(\REG.mem_51_0 ), .C(FIFO_CLK_c), .D(n5769));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4883_4884 (.Q(\REG.mem_50_15 ), .C(FIFO_CLK_c), .D(n5768));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4880_4881 (.Q(\REG.mem_50_14 ), .C(FIFO_CLK_c), .D(n5767));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4877_4878 (.Q(\REG.mem_50_13 ), .C(FIFO_CLK_c), .D(n5766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4874_4875 (.Q(\REG.mem_50_12 ), .C(FIFO_CLK_c), .D(n5765));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4871_4872 (.Q(\REG.mem_50_11 ), .C(FIFO_CLK_c), .D(n5764));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4868_4869 (.Q(\REG.mem_50_10 ), .C(FIFO_CLK_c), .D(n5763));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4865_4866 (.Q(\REG.mem_50_9 ), .C(FIFO_CLK_c), .D(n5762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4862_4863 (.Q(\REG.mem_50_8 ), .C(FIFO_CLK_c), .D(n5761));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4859_4860 (.Q(\REG.mem_50_7 ), .C(FIFO_CLK_c), .D(n5760));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4856_4857 (.Q(\REG.mem_50_6 ), .C(FIFO_CLK_c), .D(n5759));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4853_4854 (.Q(\REG.mem_50_5 ), .C(FIFO_CLK_c), .D(n5758));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4850_4851 (.Q(\REG.mem_50_4 ), .C(FIFO_CLK_c), .D(n5757));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_6__I_0_add_2_2 (.CI(VCC_net), .I0(wr_addr_r[0]), 
            .I1(rp_sync_w[0]), .CO(n9968));
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_8_lut (.I0(rd_sig_diff0_w[5]), .I1(wp_sync2_r[6]), 
            .I2(n1[6]), .I3(n9967), .O(n10700)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_7_lut (.I0(GND_net), .I1(wp_sync_w[5]), 
            .I2(n1[5]), .I3(n9966), .O(rd_sig_diff0_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3935_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_24_5 ), .O(n5318));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3935_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4847_4848 (.Q(\REG.mem_50_3 ), .C(FIFO_CLK_c), .D(n5756));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY rd_addr_r_6__I_0_151_4 (.CI(n10012), .I0(rd_addr_r[2]), .I1(GND_net), 
            .CO(n10013));
    SB_DFF i4844_4845 (.Q(\REG.mem_50_2 ), .C(FIFO_CLK_c), .D(n5755));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4841_4842 (.Q(\REG.mem_50_1 ), .C(FIFO_CLK_c), .D(n5754));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF \REG.out_buffer__i14  (.Q(\fifo_data_out[14] ), .C(SLM_CLK_c), 
           .D(n4893));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i15  (.Q(\fifo_data_out[15] ), .C(SLM_CLK_c), 
           .D(n4896));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF i4838_4839 (.Q(\REG.mem_50_0 ), .C(FIFO_CLK_c), .D(n5750));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4787_4788 (.Q(\REG.mem_49_15 ), .C(FIFO_CLK_c), .D(n5749));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4784_4785 (.Q(\REG.mem_49_14 ), .C(FIFO_CLK_c), .D(n5748));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4781_4782 (.Q(\REG.mem_49_13 ), .C(FIFO_CLK_c), .D(n5747));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4778_4779 (.Q(\REG.mem_49_12 ), .C(FIFO_CLK_c), .D(n5746));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4775_4776 (.Q(\REG.mem_49_11 ), .C(FIFO_CLK_c), .D(n5745));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4772_4773 (.Q(\REG.mem_49_10 ), .C(FIFO_CLK_c), .D(n5744));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4769_4770 (.Q(\REG.mem_49_9 ), .C(FIFO_CLK_c), .D(n5743));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4766_4767 (.Q(\REG.mem_49_8 ), .C(FIFO_CLK_c), .D(n5742));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4763_4764 (.Q(\REG.mem_49_7 ), .C(FIFO_CLK_c), .D(n5741));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_6__I_0_151_3_lut (.I0(GND_net), .I1(rd_addr_r[1]), 
            .I2(GND_net), .I3(n10011), .O(rd_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3934_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_24_4 ), .O(n5317));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3934_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY rd_addr_r_6__I_0_151_3 (.CI(n10011), .I0(rd_addr_r[1]), .I1(GND_net), 
            .CO(n10012));
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_7 (.CI(n9966), .I0(wp_sync_w[5]), 
            .I1(n1[5]), .CO(n9967));
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10400 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_38_5 ), 
            .I2(\REG.mem_39_5 ), .I3(rd_addr_r[1]), .O(n12273));
    defparam rd_addr_r_0__bdd_4_lut_10400.LUT_INIT = 16'he4aa;
    SB_DFF i4760_4761 (.Q(\REG.mem_49_6 ), .C(FIFO_CLK_c), .D(n5740));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4757_4758 (.Q(\REG.mem_49_5 ), .C(FIFO_CLK_c), .D(n5739));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4754_4755 (.Q(\REG.mem_49_4 ), .C(FIFO_CLK_c), .D(n5738));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4751_4752 (.Q(\REG.mem_49_3 ), .C(FIFO_CLK_c), .D(n5737));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4748_4749 (.Q(\REG.mem_49_2 ), .C(FIFO_CLK_c), .D(n5736));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4745_4746 (.Q(\REG.mem_49_1 ), .C(FIFO_CLK_c), .D(n5735));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4742_4743 (.Q(\REG.mem_49_0 ), .C(FIFO_CLK_c), .D(n5734));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4691_4692 (.Q(\REG.mem_48_15 ), .C(FIFO_CLK_c), .D(n5733));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4688_4689 (.Q(\REG.mem_48_14 ), .C(FIFO_CLK_c), .D(n5732));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4685_4686 (.Q(\REG.mem_48_13 ), .C(FIFO_CLK_c), .D(n5731));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4682_4683 (.Q(\REG.mem_48_12 ), .C(FIFO_CLK_c), .D(n5730));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4679_4680 (.Q(\REG.mem_48_11 ), .C(FIFO_CLK_c), .D(n5729));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4676_4677 (.Q(\REG.mem_48_10 ), .C(FIFO_CLK_c), .D(n5728));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4673_4674 (.Q(\REG.mem_48_9 ), .C(FIFO_CLK_c), .D(n5727));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4670_4671 (.Q(\REG.mem_48_8 ), .C(FIFO_CLK_c), .D(n5726));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3933_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_24_3 ), .O(n5316));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3933_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4667_4668 (.Q(\REG.mem_48_7 ), .C(FIFO_CLK_c), .D(n5725));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4664_4665 (.Q(\REG.mem_48_6 ), .C(FIFO_CLK_c), .D(n5724));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_6_lut (.I0(rd_sig_diff0_w[3]), .I1(wp_sync_w[4]), 
            .I2(n1[4]), .I3(n9965), .O(n10748)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_6_lut.LUT_INIT = 16'hebbe;
    SB_DFF i4661_4662 (.Q(\REG.mem_48_5 ), .C(FIFO_CLK_c), .D(n5723));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4658_4659 (.Q(\REG.mem_48_4 ), .C(FIFO_CLK_c), .D(n5722));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4655_4656 (.Q(\REG.mem_48_3 ), .C(FIFO_CLK_c), .D(n5721));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4652_4653 (.Q(\REG.mem_48_2 ), .C(FIFO_CLK_c), .D(n5720));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4649_4650 (.Q(\REG.mem_48_1 ), .C(FIFO_CLK_c), .D(n5719));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i77_78 (.Q(\REG.mem_0_13 ), .C(FIFO_CLK_c), .D(n4926));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i80_81 (.Q(\REG.mem_0_14 ), .C(FIFO_CLK_c), .D(n4925));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11462 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_42_6 ), 
            .I2(\REG.mem_43_6 ), .I3(rd_addr_r[1]), .O(n13551));
    defparam rd_addr_r_0__bdd_4_lut_11462.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10972 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_26_12 ), 
            .I2(\REG.mem_27_12 ), .I3(rd_addr_r[1]), .O(n12897));
    defparam rd_addr_r_0__bdd_4_lut_10972.LUT_INIT = 16'he4aa;
    SB_DFF i4646_4647 (.Q(\REG.mem_48_0 ), .C(FIFO_CLK_c), .D(n5718));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4595_4596 (.Q(\REG.mem_47_15 ), .C(FIFO_CLK_c), .D(n5717));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13551_bdd_4_lut (.I0(n13551), .I1(\REG.mem_41_6 ), .I2(\REG.mem_40_6 ), 
            .I3(rd_addr_r[1]), .O(n11315));
    defparam n13551_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4592_4593 (.Q(\REG.mem_47_14 ), .C(FIFO_CLK_c), .D(n5716));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4589_4590 (.Q(\REG.mem_47_13 ), .C(FIFO_CLK_c), .D(n5715));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4586_4587 (.Q(\REG.mem_47_12 ), .C(FIFO_CLK_c), .D(n5714));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4583_4584 (.Q(\REG.mem_47_11 ), .C(FIFO_CLK_c), .D(n5713));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4580_4581 (.Q(\REG.mem_47_10 ), .C(FIFO_CLK_c), .D(n5712));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4577_4578 (.Q(\REG.mem_47_9 ), .C(FIFO_CLK_c), .D(n5711));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4574_4575 (.Q(\REG.mem_47_8 ), .C(FIFO_CLK_c), .D(n5710));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4571_4572 (.Q(\REG.mem_47_7 ), .C(FIFO_CLK_c), .D(n5709));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4568_4569 (.Q(\REG.mem_47_6 ), .C(FIFO_CLK_c), .D(n5708));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4565_4566 (.Q(\REG.mem_47_5 ), .C(FIFO_CLK_c), .D(n5707));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4562_4563 (.Q(\REG.mem_47_4 ), .C(FIFO_CLK_c), .D(n5706));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4559_4560 (.Q(\REG.mem_47_3 ), .C(FIFO_CLK_c), .D(n5705));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4556_4557 (.Q(\REG.mem_47_2 ), .C(FIFO_CLK_c), .D(n5704));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4553_4554 (.Q(\REG.mem_47_1 ), .C(FIFO_CLK_c), .D(n5703));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12897_bdd_4_lut (.I0(n12897), .I1(\REG.mem_25_12 ), .I2(\REG.mem_24_12 ), 
            .I3(rd_addr_r[1]), .O(n12900));
    defparam n12897_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i83_84 (.Q(\REG.mem_0_15 ), .C(FIFO_CLK_c), .D(n4924));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12273_bdd_4_lut (.I0(n12273), .I1(\REG.mem_37_5 ), .I2(\REG.mem_36_5 ), 
            .I3(rd_addr_r[1]), .O(n12276));
    defparam n12273_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4550_4551 (.Q(\REG.mem_47_0 ), .C(FIFO_CLK_c), .D(n5702));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11457 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_58_2 ), 
            .I2(\REG.mem_59_2 ), .I3(rd_addr_r[1]), .O(n13545));
    defparam rd_addr_r_0__bdd_4_lut_11457.LUT_INIT = 16'he4aa;
    SB_DFF i4499_4500 (.Q(\REG.mem_46_15 ), .C(FIFO_CLK_c), .D(n5701));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4496_4497 (.Q(\REG.mem_46_14 ), .C(FIFO_CLK_c), .D(n5700));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4493_4494 (.Q(\REG.mem_46_13 ), .C(FIFO_CLK_c), .D(n5699));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3932_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_24_2 ), .O(n5315));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3932_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4490_4491 (.Q(\REG.mem_46_12 ), .C(FIFO_CLK_c), .D(n5698));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4487_4488 (.Q(\REG.mem_46_11 ), .C(FIFO_CLK_c), .D(n5697));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4484_4485 (.Q(\REG.mem_46_10 ), .C(FIFO_CLK_c), .D(n5696));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3931_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_24_1 ), .O(n5314));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3931_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4481_4482 (.Q(\REG.mem_46_9 ), .C(FIFO_CLK_c), .D(n5695));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4478_4479 (.Q(\REG.mem_46_8 ), .C(FIFO_CLK_c), .D(n5694));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4475_4476 (.Q(\REG.mem_46_7 ), .C(FIFO_CLK_c), .D(n5693));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4472_4473 (.Q(\REG.mem_46_6 ), .C(FIFO_CLK_c), .D(n5692));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4469_4470 (.Q(\REG.mem_46_5 ), .C(FIFO_CLK_c), .D(n5691));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4466_4467 (.Q(\REG.mem_46_4 ), .C(FIFO_CLK_c), .D(n5690));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4463_4464 (.Q(\REG.mem_46_3 ), .C(FIFO_CLK_c), .D(n5689));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4460_4461 (.Q(\REG.mem_46_2 ), .C(FIFO_CLK_c), .D(n5688));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4457_4458 (.Q(\REG.mem_46_1 ), .C(FIFO_CLK_c), .D(n5687));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4454_4455 (.Q(\REG.mem_46_0 ), .C(FIFO_CLK_c), .D(n5686));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4403_4404 (.Q(\REG.mem_45_15 ), .C(FIFO_CLK_c), .D(n5685));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4400_4401 (.Q(\REG.mem_45_14 ), .C(FIFO_CLK_c), .D(n5684));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4397_4398 (.Q(\REG.mem_45_13 ), .C(FIFO_CLK_c), .D(n5683));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4394_4395 (.Q(\REG.mem_45_12 ), .C(FIFO_CLK_c), .D(n5682));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4391_4392 (.Q(\REG.mem_45_11 ), .C(FIFO_CLK_c), .D(n5681));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4388_4389 (.Q(\REG.mem_45_10 ), .C(FIFO_CLK_c), .D(n5680));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4385_4386 (.Q(\REG.mem_45_9 ), .C(FIFO_CLK_c), .D(n5679));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3924_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_24_0 ), .O(n5307));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3924_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10395 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_58_12 ), 
            .I2(\REG.mem_59_12 ), .I3(rd_addr_r[1]), .O(n12267));
    defparam rd_addr_r_0__bdd_4_lut_10395.LUT_INIT = 16'he4aa;
    SB_DFF i4382_4383 (.Q(\REG.mem_45_8 ), .C(FIFO_CLK_c), .D(n5678));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13545_bdd_4_lut (.I0(n13545), .I1(\REG.mem_57_2 ), .I2(\REG.mem_56_2 ), 
            .I3(rd_addr_r[1]), .O(n13548));
    defparam n13545_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3977_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_26_15 ), .O(n5360));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3977_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12267_bdd_4_lut (.I0(n12267), .I1(\REG.mem_57_12 ), .I2(\REG.mem_56_12 ), 
            .I3(rd_addr_r[1]), .O(n12270));
    defparam n12267_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10912 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_6_15 ), 
            .I2(\REG.mem_7_15 ), .I3(rd_addr_r[1]), .O(n12891));
    defparam rd_addr_r_0__bdd_4_lut_10912.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10390 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_2_1 ), 
            .I2(\REG.mem_3_1 ), .I3(rd_addr_r[1]), .O(n12261));
    defparam rd_addr_r_0__bdd_4_lut_10390.LUT_INIT = 16'he4aa;
    SB_DFF i4379_4380 (.Q(\REG.mem_45_7 ), .C(FIFO_CLK_c), .D(n5677));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12891_bdd_4_lut (.I0(n12891), .I1(\REG.mem_5_15 ), .I2(\REG.mem_4_15 ), 
            .I3(rd_addr_r[1]), .O(n12894));
    defparam n12891_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4376_4377 (.Q(\REG.mem_45_6 ), .C(FIFO_CLK_c), .D(n5676));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4373_4374 (.Q(\REG.mem_45_5 ), .C(FIFO_CLK_c), .D(n5675));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4370_4371 (.Q(\REG.mem_45_4 ), .C(FIFO_CLK_c), .D(n5674));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4367_4368 (.Q(\REG.mem_45_3 ), .C(FIFO_CLK_c), .D(n5673));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4364_4365 (.Q(\REG.mem_45_2 ), .C(FIFO_CLK_c), .D(n5672));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4361_4362 (.Q(\REG.mem_45_1 ), .C(FIFO_CLK_c), .D(n5671));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4358_4359 (.Q(\REG.mem_45_0 ), .C(FIFO_CLK_c), .D(n5670));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wr_grey_sync_r__i6 (.Q(wr_grey_sync_r[6]), .C(FIFO_CLK_c), .D(n5669));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF i4307_4308 (.Q(\REG.mem_44_15 ), .C(FIFO_CLK_c), .D(n5668));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4304_4305 (.Q(\REG.mem_44_14 ), .C(FIFO_CLK_c), .D(n5667));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4301_4302 (.Q(\REG.mem_44_13 ), .C(FIFO_CLK_c), .D(n5665));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4298_4299 (.Q(\REG.mem_44_12 ), .C(FIFO_CLK_c), .D(n5664));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4295_4296 (.Q(\REG.mem_44_11 ), .C(FIFO_CLK_c), .D(n5663));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4292_4293 (.Q(\REG.mem_44_10 ), .C(FIFO_CLK_c), .D(n5661));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12261_bdd_4_lut (.I0(n12261), .I1(\REG.mem_1_1 ), .I2(\REG.mem_0_1 ), 
            .I3(rd_addr_r[1]), .O(n11006));
    defparam n12261_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3976_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_26_14 ), .O(n5359));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3976_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3975_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_26_13 ), .O(n5358));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3975_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4289_4290 (.Q(\REG.mem_44_9 ), .C(FIFO_CLK_c), .D(n5660));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4286_4287 (.Q(\REG.mem_44_8 ), .C(FIFO_CLK_c), .D(n5659));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4283_4284 (.Q(\REG.mem_44_7 ), .C(FIFO_CLK_c), .D(n5658));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4280_4281 (.Q(\REG.mem_44_6 ), .C(FIFO_CLK_c), .D(n5657));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4277_4278 (.Q(\REG.mem_44_5 ), .C(FIFO_CLK_c), .D(n5656));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4274_4275 (.Q(\REG.mem_44_4 ), .C(FIFO_CLK_c), .D(n5655));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4271_4272 (.Q(\REG.mem_44_3 ), .C(FIFO_CLK_c), .D(n5654));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4268_4269 (.Q(\REG.mem_44_2 ), .C(FIFO_CLK_c), .D(n5653));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4265_4266 (.Q(\REG.mem_44_1 ), .C(FIFO_CLK_c), .D(n5652));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4262_4263 (.Q(\REG.mem_44_0 ), .C(FIFO_CLK_c), .D(n5651));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4211_4212 (.Q(\REG.mem_43_15 ), .C(FIFO_CLK_c), .D(n5650));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4208_4209 (.Q(\REG.mem_43_14 ), .C(FIFO_CLK_c), .D(n5649));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4205_4206 (.Q(\REG.mem_43_13 ), .C(FIFO_CLK_c), .D(n5648));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4202_4203 (.Q(\REG.mem_43_12 ), .C(FIFO_CLK_c), .D(n5647));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4199_4200 (.Q(\REG.mem_43_11 ), .C(FIFO_CLK_c), .D(n5646));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4196_4197 (.Q(\REG.mem_43_10 ), .C(FIFO_CLK_c), .D(n5645));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3974_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_26_12 ), .O(n5357));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3974_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_6 (.CI(n9965), .I0(wp_sync_w[4]), 
            .I1(n1[4]), .CO(n9966));
    SB_DFF i4193_4194 (.Q(\REG.mem_43_9 ), .C(FIFO_CLK_c), .D(n5644));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11557 (.I0(rd_addr_r[1]), .I1(n11784), 
            .I2(n11785), .I3(rd_addr_r[2]), .O(n13539));
    defparam rd_addr_r_1__bdd_4_lut_11557.LUT_INIT = 16'he4aa;
    SB_LUT4 i3973_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_26_11 ), .O(n5356));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3973_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13539_bdd_4_lut (.I0(n13539), .I1(n11722), .I2(n11721), .I3(rd_addr_r[2]), 
            .O(n10900));
    defparam n13539_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_5_lut (.I0(GND_net), .I1(wp_sync_w[3]), 
            .I2(n1[3]), .I3(n9964), .O(rd_sig_diff0_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3972_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_26_10 ), .O(n5355));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3972_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3971_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_26_9 ), .O(n5354));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3971_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3970_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_26_8 ), .O(n5353));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3970_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_6__I_0_151_2_lut (.I0(GND_net), .I1(\rd_addr_r[0] ), 
            .I2(GND_net), .I3(VCC_net), .O(\rd_addr_p1_w[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10385 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_18_7 ), 
            .I2(\REG.mem_19_7 ), .I3(rd_addr_r[1]), .O(n12255));
    defparam rd_addr_r_0__bdd_4_lut_10385.LUT_INIT = 16'he4aa;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_5 (.CI(n9964), .I0(wp_sync_w[3]), 
            .I1(n1[3]), .CO(n9965));
    SB_LUT4 i3969_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_26_7 ), .O(n5352));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3969_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4190_4191 (.Q(\REG.mem_43_8 ), .C(FIFO_CLK_c), .D(n5643));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4187_4188 (.Q(\REG.mem_43_7 ), .C(FIFO_CLK_c), .D(n5642));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4184_4185 (.Q(\REG.mem_43_6 ), .C(FIFO_CLK_c), .D(n5641));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4181_4182 (.Q(\REG.mem_43_5 ), .C(FIFO_CLK_c), .D(n5640));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4178_4179 (.Q(\REG.mem_43_4 ), .C(FIFO_CLK_c), .D(n5639));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4175_4176 (.Q(\REG.mem_43_3 ), .C(FIFO_CLK_c), .D(n5638));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4172_4173 (.Q(\REG.mem_43_2 ), .C(FIFO_CLK_c), .D(n5637));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4169_4170 (.Q(\REG.mem_43_1 ), .C(FIFO_CLK_c), .D(n5636));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4166_4167 (.Q(\REG.mem_43_0 ), .C(FIFO_CLK_c), .D(n5635));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4115_4116 (.Q(\REG.mem_42_15 ), .C(FIFO_CLK_c), .D(n5634));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4112_4113 (.Q(\REG.mem_42_14 ), .C(FIFO_CLK_c), .D(n5633));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4109_4110 (.Q(\REG.mem_42_13 ), .C(FIFO_CLK_c), .D(n5632));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4106_4107 (.Q(\REG.mem_42_12 ), .C(FIFO_CLK_c), .D(n5631));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4103_4104 (.Q(\REG.mem_42_11 ), .C(FIFO_CLK_c), .D(n5630));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4100_4101 (.Q(\REG.mem_42_10 ), .C(FIFO_CLK_c), .D(n5629));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF \genblk16.rd_prev_r_132  (.Q(\genblk16.rd_prev_r ), .C(SLM_CLK_c), 
           .D(n4916));   // src/fifo_dc_32_lut_gen.v(751[29] 761[32])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10405 (.I0(rd_addr_r[2]), .I1(n11153), 
            .I2(n12174), .I3(rd_addr_r[3]), .O(n12219));
    defparam rd_addr_r_2__bdd_4_lut_10405.LUT_INIT = 16'he4aa;
    SB_LUT4 i3968_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_26_6 ), .O(n5351));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3968_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11452 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_46_0 ), 
            .I2(\REG.mem_47_0 ), .I3(rd_addr_r[1]), .O(n13533));
    defparam rd_addr_r_0__bdd_4_lut_11452.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10917 (.I0(rd_addr_r[1]), .I1(n10923), 
            .I2(n10924), .I3(rd_addr_r[2]), .O(n12885));
    defparam rd_addr_r_1__bdd_4_lut_10917.LUT_INIT = 16'he4aa;
    SB_LUT4 n13533_bdd_4_lut (.I0(n13533), .I1(\REG.mem_45_0 ), .I2(\REG.mem_44_0 ), 
            .I3(rd_addr_r[1]), .O(n11807));
    defparam n13533_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3967_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_26_5 ), .O(n5350));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3967_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12885_bdd_4_lut (.I0(n12885), .I1(n10888), .I2(n10887), .I3(rd_addr_r[2]), 
            .O(n12888));
    defparam n12885_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10907 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_22_11 ), 
            .I2(\REG.mem_23_11 ), .I3(rd_addr_r[1]), .O(n12879));
    defparam rd_addr_r_0__bdd_4_lut_10907.LUT_INIT = 16'he4aa;
    SB_LUT4 n12879_bdd_4_lut (.I0(n12879), .I1(\REG.mem_21_11 ), .I2(\REG.mem_20_11 ), 
            .I3(rd_addr_r[1]), .O(n11504));
    defparam n12879_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i167_168 (.Q(\REG.mem_1_11 ), .C(FIFO_CLK_c), .D(n4915));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i152_153 (.Q(\REG.mem_1_6 ), .C(FIFO_CLK_c), .D(n4914));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4097_4098 (.Q(\REG.mem_42_9 ), .C(FIFO_CLK_c), .D(n5628));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4094_4095 (.Q(\REG.mem_42_8 ), .C(FIFO_CLK_c), .D(n5627));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4091_4092 (.Q(\REG.mem_42_7 ), .C(FIFO_CLK_c), .D(n5626));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4088_4089 (.Q(\REG.mem_42_6 ), .C(FIFO_CLK_c), .D(n5625));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4085_4086 (.Q(\REG.mem_42_5 ), .C(FIFO_CLK_c), .D(n5624));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4082_4083 (.Q(\REG.mem_42_4 ), .C(FIFO_CLK_c), .D(n5623));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4079_4080 (.Q(\REG.mem_42_3 ), .C(FIFO_CLK_c), .D(n5622));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4076_4077 (.Q(\REG.mem_42_2 ), .C(FIFO_CLK_c), .D(n5621));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4073_4074 (.Q(\REG.mem_42_1 ), .C(FIFO_CLK_c), .D(n5620));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4070_4071 (.Q(\REG.mem_42_0 ), .C(FIFO_CLK_c), .D(n5619));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4019_4020 (.Q(\REG.mem_41_15 ), .C(FIFO_CLK_c), .D(n5618));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4016_4017 (.Q(\REG.mem_41_14 ), .C(FIFO_CLK_c), .D(n5617));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4013_4014 (.Q(\REG.mem_41_13 ), .C(FIFO_CLK_c), .D(n5616));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4010_4011 (.Q(\REG.mem_41_12 ), .C(FIFO_CLK_c), .D(n5615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4007_4008 (.Q(\REG.mem_41_11 ), .C(FIFO_CLK_c), .D(n5614));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4004_4005 (.Q(\REG.mem_41_10 ), .C(FIFO_CLK_c), .D(n5613));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3966_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_26_4 ), .O(n5349));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3966_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10897 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_26_6 ), 
            .I2(\REG.mem_27_6 ), .I3(rd_addr_r[1]), .O(n12873));
    defparam rd_addr_r_0__bdd_4_lut_10897.LUT_INIT = 16'he4aa;
    SB_LUT4 i4353_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_49_2 ), .O(n5736));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4353_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12873_bdd_4_lut (.I0(n12873), .I1(\REG.mem_25_6 ), .I2(\REG.mem_24_6 ), 
            .I3(rd_addr_r[1]), .O(n11123));
    defparam n12873_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4352_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_49_1 ), .O(n5735));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4352_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11447 (.I0(rd_addr_r[1]), .I1(n11775), 
            .I2(n11776), .I3(rd_addr_r[2]), .O(n13527));
    defparam rd_addr_r_1__bdd_4_lut_11447.LUT_INIT = 16'he4aa;
    SB_LUT4 n13527_bdd_4_lut (.I0(n13527), .I1(n11767), .I2(n11766), .I3(rd_addr_r[2]), 
            .O(n10903));
    defparam n13527_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3965_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_26_3 ), .O(n5348));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3965_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i170_171 (.Q(\REG.mem_1_12 ), .C(FIFO_CLK_c), .D(n4912));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4001_4002 (.Q(\REG.mem_41_9 ), .C(FIFO_CLK_c), .D(n5612));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3998_3999 (.Q(\REG.mem_41_8 ), .C(FIFO_CLK_c), .D(n5611));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3995_3996 (.Q(\REG.mem_41_7 ), .C(FIFO_CLK_c), .D(n5610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3992_3993 (.Q(\REG.mem_41_6 ), .C(FIFO_CLK_c), .D(n5609));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3989_3990 (.Q(\REG.mem_41_5 ), .C(FIFO_CLK_c), .D(n5608));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3986_3987 (.Q(\REG.mem_41_4 ), .C(FIFO_CLK_c), .D(n5607));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3983_3984 (.Q(\REG.mem_41_3 ), .C(FIFO_CLK_c), .D(n5606));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3980_3981 (.Q(\REG.mem_41_2 ), .C(FIFO_CLK_c), .D(n5605));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3977_3978 (.Q(\REG.mem_41_1 ), .C(FIFO_CLK_c), .D(n5604));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3974_3975 (.Q(\REG.mem_41_0 ), .C(FIFO_CLK_c), .D(n5603));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3923_3924 (.Q(\REG.mem_40_15 ), .C(FIFO_CLK_c), .D(n5602));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3920_3921 (.Q(\REG.mem_40_14 ), .C(FIFO_CLK_c), .D(n5601));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3917_3918 (.Q(\REG.mem_40_13 ), .C(FIFO_CLK_c), .D(n5600));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3914_3915 (.Q(\REG.mem_40_12 ), .C(FIFO_CLK_c), .D(n5599));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3911_3912 (.Q(\REG.mem_40_11 ), .C(FIFO_CLK_c), .D(n5598));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3908_3909 (.Q(\REG.mem_40_10 ), .C(FIFO_CLK_c), .D(n5597));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4088_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_33_14 ), .O(n5471));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4088_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3964_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_26_2 ), .O(n5347));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3964_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY rd_addr_r_6__I_0_151_2 (.CI(VCC_net), .I0(\rd_addr_r[0] ), 
            .I1(GND_net), .CO(n10011));
    SB_DFF i155_156 (.Q(\REG.mem_1_7 ), .C(FIFO_CLK_c), .D(n4905));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3963_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_26_1 ), .O(n5346));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3963_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9385_3_lut (.I0(\REG.mem_48_5 ), .I1(\REG.mem_49_5 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11235));
    defparam i9385_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF wp_sync2_r__i0 (.Q(wp_sync2_r[0]), .C(SLM_CLK_c), .D(n4904));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i0 (.Q(wp_sync1_r[0]), .C(SLM_CLK_c), .D(n4903));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i173_174 (.Q(\REG.mem_1_13 ), .C(FIFO_CLK_c), .D(n4902));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rd_addr_r__i0 (.Q(\rd_addr_r[0] ), .C(SLM_CLK_c), .D(n4901));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF i158_159 (.Q(\REG.mem_1_8 ), .C(FIFO_CLK_c), .D(n4900));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync2_r__i0 (.Q(rp_sync2_r[0]), .C(FIFO_CLK_c), .D(n4899));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i3905_3906 (.Q(\REG.mem_40_9 ), .C(FIFO_CLK_c), .D(n5596));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3962_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_26_0 ), .O(n5345));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3962_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3902_3903 (.Q(\REG.mem_40_8 ), .C(FIFO_CLK_c), .D(n5595));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9386_3_lut (.I0(\REG.mem_50_5 ), .I1(\REG.mem_51_5 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11236));
    defparam i9386_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3899_3900 (.Q(\REG.mem_40_7 ), .C(FIFO_CLK_c), .D(n5594));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3896_3897 (.Q(\REG.mem_40_6 ), .C(FIFO_CLK_c), .D(n5593));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3893_3894 (.Q(\REG.mem_40_5 ), .C(FIFO_CLK_c), .D(n5592));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3890_3891 (.Q(\REG.mem_40_4 ), .C(FIFO_CLK_c), .D(n5591));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3887_3888 (.Q(\REG.mem_40_3 ), .C(FIFO_CLK_c), .D(n5590));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3884_3885 (.Q(\REG.mem_40_2 ), .C(FIFO_CLK_c), .D(n5589));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3881_3882 (.Q(\REG.mem_40_1 ), .C(FIFO_CLK_c), .D(n5588));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3878_3879 (.Q(\REG.mem_40_0 ), .C(FIFO_CLK_c), .D(n5587));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3827_3828 (.Q(\REG.mem_39_15 ), .C(FIFO_CLK_c), .D(n5586));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3824_3825 (.Q(\REG.mem_39_14 ), .C(FIFO_CLK_c), .D(n5585));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3821_3822 (.Q(\REG.mem_39_13 ), .C(FIFO_CLK_c), .D(n5584));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3818_3819 (.Q(\REG.mem_39_12 ), .C(FIFO_CLK_c), .D(n5583));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3815_3816 (.Q(\REG.mem_39_11 ), .C(FIFO_CLK_c), .D(n5582));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3812_3813 (.Q(\REG.mem_39_10 ), .C(FIFO_CLK_c), .D(n5581));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync1_r__i0 (.Q(rp_sync1_r[0]), .C(FIFO_CLK_c), .D(n4898));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_LUT4 i4087_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_33_13 ), .O(n5470));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4087_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12219_bdd_4_lut (.I0(n12219), .I1(n11081), .I2(n11006), .I3(rd_addr_r[3]), 
            .O(n12222));
    defparam n12219_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3993_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_27_15 ), .O(n5376));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3993_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_2_lut (.I0(wr_sig_diff0_w[0]), .I1(wr_sig_diff0_w[1]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_1189));   // src/fifo_dc_32_lut_gen.v(403[38:87])
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(DEBUG_5_c), .I1(wr_sig_diff0_w[3]), .I2(n6_adj_1189), 
            .I3(wr_sig_diff0_w[2]), .O(n2_adj_1188));   // src/fifo_dc_32_lut_gen.v(403[38:87])
    defparam i1_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i3992_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_27_14 ), .O(n5375));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3992_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11442 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_62_2 ), 
            .I2(\REG.mem_63_2 ), .I3(rd_addr_r[1]), .O(n13521));
    defparam rd_addr_r_0__bdd_4_lut_11442.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut (.I0(wr_sig_diff0_w[2]), .I1(wr_sig_diff0_w[1]), .I2(wr_sig_diff0_w[0]), 
            .I3(GND_net), .O(n10126));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10922 (.I0(rd_addr_r[3]), .I1(n12750), 
            .I2(n11113), .I3(rd_addr_r[4]), .O(n12867));
    defparam rd_addr_r_3__bdd_4_lut_10922.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10312 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_2_4 ), 
            .I2(\REG.mem_3_4 ), .I3(rd_addr_r[1]), .O(n12165));
    defparam rd_addr_r_0__bdd_4_lut_10312.LUT_INIT = 16'he4aa;
    SB_LUT4 i8949_4_lut (.I0(dc32_fifo_almost_full), .I1(n10778), .I2(n10126), 
            .I3(wr_sig_diff0_w[3]), .O(n10798));
    defparam i8949_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i3991_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_27_13 ), .O(n5374));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3991_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12867_bdd_4_lut (.I0(n12867), .I1(n11110), .I2(n12744), .I3(rd_addr_r[4]), 
            .O(n12870));
    defparam n12867_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3990_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_27_12 ), .O(n5373));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3990_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13521_bdd_4_lut (.I0(n13521), .I1(\REG.mem_61_2 ), .I2(\REG.mem_60_2 ), 
            .I3(rd_addr_r[1]), .O(n13524));
    defparam n13521_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3989_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_27_11 ), .O(n5372));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3989_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11432 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_6_4 ), 
            .I2(\REG.mem_7_4 ), .I3(rd_addr_r[1]), .O(n13515));
    defparam rd_addr_r_0__bdd_4_lut_11432.LUT_INIT = 16'he4aa;
    SB_DFF i3809_3810 (.Q(\REG.mem_39_9 ), .C(FIFO_CLK_c), .D(n5580));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3806_3807 (.Q(\REG.mem_39_8 ), .C(FIFO_CLK_c), .D(n5579));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10892 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_26_11 ), 
            .I2(\REG.mem_27_11 ), .I3(rd_addr_r[1]), .O(n12861));
    defparam rd_addr_r_0__bdd_4_lut_10892.LUT_INIT = 16'he4aa;
    SB_DFF i3803_3804 (.Q(\REG.mem_39_7 ), .C(FIFO_CLK_c), .D(n5578));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3800_3801 (.Q(\REG.mem_39_6 ), .C(FIFO_CLK_c), .D(n5577));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3797_3798 (.Q(\REG.mem_39_5 ), .C(FIFO_CLK_c), .D(n5576));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3794_3795 (.Q(\REG.mem_39_4 ), .C(FIFO_CLK_c), .D(n5575));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3791_3792 (.Q(\REG.mem_39_3 ), .C(FIFO_CLK_c), .D(n5574));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3788_3789 (.Q(\REG.mem_39_2 ), .C(FIFO_CLK_c), .D(n5573));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3785_3786 (.Q(\REG.mem_39_1 ), .C(FIFO_CLK_c), .D(n5572));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3782_3783 (.Q(\REG.mem_39_0 ), .C(FIFO_CLK_c), .D(n5570));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3731_3732 (.Q(\REG.mem_38_15 ), .C(FIFO_CLK_c), .D(n5569));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3728_3729 (.Q(\REG.mem_38_14 ), .C(FIFO_CLK_c), .D(n5568));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3725_3726 (.Q(\REG.mem_38_13 ), .C(FIFO_CLK_c), .D(n5567));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3722_3723 (.Q(\REG.mem_38_12 ), .C(FIFO_CLK_c), .D(n5566));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3719_3720 (.Q(\REG.mem_38_11 ), .C(FIFO_CLK_c), .D(n5565));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3716_3717 (.Q(\REG.mem_38_10 ), .C(FIFO_CLK_c), .D(n5564));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3988_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_27_10 ), .O(n5371));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3988_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3987_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_27_9 ), .O(n5370));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3987_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13515_bdd_4_lut (.I0(n13515), .I1(\REG.mem_5_4 ), .I2(\REG.mem_4_4 ), 
            .I3(rd_addr_r[1]), .O(n13518));
    defparam n13515_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3986_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_27_8 ), .O(n5369));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3986_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3985_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_27_7 ), .O(n5368));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3985_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3984_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_27_6 ), .O(n5367));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3984_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3983_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_27_5 ), .O(n5366));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3983_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3982_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_27_4 ), .O(n5365));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3982_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3981_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_27_3 ), .O(n5364));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3981_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12165_bdd_4_lut (.I0(n12165), .I1(\REG.mem_1_4 ), .I2(\REG.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(n12168));
    defparam n12165_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3980_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_27_2 ), .O(n5363));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3980_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3979_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_27_1 ), .O(n5362));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3979_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3713_3714 (.Q(\REG.mem_38_9 ), .C(FIFO_CLK_c), .D(n5563));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3710_3711 (.Q(\REG.mem_38_8 ), .C(FIFO_CLK_c), .D(n5562));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3707_3708 (.Q(\REG.mem_38_7 ), .C(FIFO_CLK_c), .D(n5561));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3704_3705 (.Q(\REG.mem_38_6 ), .C(FIFO_CLK_c), .D(n5560));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3701_3702 (.Q(\REG.mem_38_5 ), .C(FIFO_CLK_c), .D(n5559));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3698_3699 (.Q(\REG.mem_38_4 ), .C(FIFO_CLK_c), .D(n5558));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3695_3696 (.Q(\REG.mem_38_3 ), .C(FIFO_CLK_c), .D(n5557));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3692_3693 (.Q(\REG.mem_38_2 ), .C(FIFO_CLK_c), .D(n5556));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3689_3690 (.Q(\REG.mem_38_1 ), .C(FIFO_CLK_c), .D(n5555));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3686_3687 (.Q(\REG.mem_38_0 ), .C(FIFO_CLK_c), .D(n5554));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3635_3636 (.Q(\REG.mem_37_15 ), .C(FIFO_CLK_c), .D(n5553));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3632_3633 (.Q(\REG.mem_37_14 ), .C(FIFO_CLK_c), .D(n5552));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3629_3630 (.Q(\REG.mem_37_13 ), .C(FIFO_CLK_c), .D(n5551));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3626_3627 (.Q(\REG.mem_37_12 ), .C(FIFO_CLK_c), .D(n5550));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3623_3624 (.Q(\REG.mem_37_11 ), .C(FIFO_CLK_c), .D(n5549));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFE \REG.out_raw__i16  (.Q(\REG.out_raw[15] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [15]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i15  (.Q(\REG.out_raw[14] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [14]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i14  (.Q(\REG.out_raw[13] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [13]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i13  (.Q(\REG.out_raw[12] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [12]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i12  (.Q(\REG.out_raw[11] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [11]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFF i3620_3621 (.Q(\REG.mem_37_10 ), .C(FIFO_CLK_c), .D(n5548));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3617_3618 (.Q(\REG.mem_37_9 ), .C(FIFO_CLK_c), .D(n5547));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3614_3615 (.Q(\REG.mem_37_8 ), .C(FIFO_CLK_c), .D(n5546));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3611_3612 (.Q(\REG.mem_37_7 ), .C(FIFO_CLK_c), .D(n5545));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3608_3609 (.Q(\REG.mem_37_6 ), .C(FIFO_CLK_c), .D(n5544));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3605_3606 (.Q(\REG.mem_37_5 ), .C(FIFO_CLK_c), .D(n5543));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3602_3603 (.Q(\REG.mem_37_4 ), .C(FIFO_CLK_c), .D(n5542));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3599_3600 (.Q(\REG.mem_37_3 ), .C(FIFO_CLK_c), .D(n5541));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3596_3597 (.Q(\REG.mem_37_2 ), .C(FIFO_CLK_c), .D(n5540));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3593_3594 (.Q(\REG.mem_37_1 ), .C(FIFO_CLK_c), .D(n5539));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3590_3591 (.Q(\REG.mem_37_0 ), .C(FIFO_CLK_c), .D(n5538));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFE \REG.out_raw__i11  (.Q(\REG.out_raw[10] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [10]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 i4086_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_33_12 ), .O(n5469));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4086_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3978_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_27_0 ), .O(n5361));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3978_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_raw__i10  (.Q(\REG.out_raw[9] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [9]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i9  (.Q(\REG.out_raw[8] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [8]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i5 (.Q(wr_grey_sync_r[5]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[5]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i8  (.Q(\REG.out_raw[7] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [7]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i4 (.Q(wr_grey_sync_r[4]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[4]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i7  (.Q(\REG.out_raw[6] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [6]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i3 (.Q(wr_grey_sync_r[3]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[3]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i6  (.Q(\REG.out_raw[5] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [5]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i2 (.Q(wr_grey_sync_r[2]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[2]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i5  (.Q(\REG.out_raw[4] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [4]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFSR wr_grey_sync_r__i1 (.Q(wr_grey_sync_r[1]), .C(FIFO_CLK_c), 
            .D(wr_grey_w[1]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFE \REG.out_raw__i4  (.Q(\REG.out_raw[3] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [3]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i3  (.Q(\REG.out_raw[2] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [2]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i2  (.Q(\REG.out_raw[1] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_559 [1]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 i4009_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_28_15 ), .O(n5392));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4009_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4008_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_28_14 ), .O(n5391));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4008_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4007_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_28_13 ), .O(n5390));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4007_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4006_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_28_12 ), .O(n5389));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4006_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4351_3_lut_4_lut (.I0(n39), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_49_0 ), .O(n5734));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4351_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i3539_3540 (.Q(\REG.mem_36_15 ), .C(FIFO_CLK_c), .D(n5524));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3536_3537 (.Q(\REG.mem_36_14 ), .C(FIFO_CLK_c), .D(n5523));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3533_3534 (.Q(\REG.mem_36_13 ), .C(FIFO_CLK_c), .D(n5522));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3530_3531 (.Q(\REG.mem_36_12 ), .C(FIFO_CLK_c), .D(n5521));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3527_3528 (.Q(\REG.mem_36_11 ), .C(FIFO_CLK_c), .D(n5520));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3524_3525 (.Q(\REG.mem_36_10 ), .C(FIFO_CLK_c), .D(n5519));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3521_3522 (.Q(\REG.mem_36_9 ), .C(FIFO_CLK_c), .D(n5518));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3518_3519 (.Q(\REG.mem_36_8 ), .C(FIFO_CLK_c), .D(n5517));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3515_3516 (.Q(\REG.mem_36_7 ), .C(FIFO_CLK_c), .D(n5516));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4005_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_28_11 ), .O(n5388));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4005_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4004_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_28_10 ), .O(n5387));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4004_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4003_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_28_9 ), .O(n5386));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4003_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_r_6__I_0_141_8_lut (.I0(GND_net), .I1(wr_grey_sync_r[6]), 
            .I2(GND_net), .I3(n10010), .O(wr_addr_p1_w[6])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_4_lut (.I0(GND_net), .I1(wp_sync_w[2]), 
            .I2(n1[2]), .I3(n9963), .O(\rd_sig_diff0_w[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4002_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_28_8 ), .O(n5385));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4002_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3512_3513 (.Q(\REG.mem_36_6 ), .C(FIFO_CLK_c), .D(n5515));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3509_3510 (.Q(\REG.mem_36_5 ), .C(FIFO_CLK_c), .D(n5514));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3506_3507 (.Q(\REG.mem_36_4 ), .C(FIFO_CLK_c), .D(n5513));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3503_3504 (.Q(\REG.mem_36_3 ), .C(FIFO_CLK_c), .D(n5512));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3500_3501 (.Q(\REG.mem_36_2 ), .C(FIFO_CLK_c), .D(n5511));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3497_3498 (.Q(\REG.mem_36_1 ), .C(FIFO_CLK_c), .D(n5510));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3494_3495 (.Q(\REG.mem_36_0 ), .C(FIFO_CLK_c), .D(n5509));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3443_3444 (.Q(\REG.mem_35_15 ), .C(FIFO_CLK_c), .D(n5505));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3440_3441 (.Q(\REG.mem_35_14 ), .C(FIFO_CLK_c), .D(n5504));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3437_3438 (.Q(\REG.mem_35_13 ), .C(FIFO_CLK_c), .D(n5503));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3434_3435 (.Q(\REG.mem_35_12 ), .C(FIFO_CLK_c), .D(n5502));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3431_3432 (.Q(\REG.mem_35_11 ), .C(FIFO_CLK_c), .D(n5501));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3428_3429 (.Q(\REG.mem_35_10 ), .C(FIFO_CLK_c), .D(n5500));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4001_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_28_7 ), .O(n5384));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4001_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4000_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_28_6 ), .O(n5383));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4000_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_4 (.CI(n9963), .I0(wp_sync_w[2]), 
            .I1(n1[2]), .CO(n9964));
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_3_lut (.I0(GND_net), .I1(wp_sync_w[1]), 
            .I2(n1[1]), .I3(n9962), .O(\rd_sig_diff0_w[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3999_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_28_5 ), .O(n5382));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3999_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3425_3426 (.Q(\REG.mem_35_9 ), .C(FIFO_CLK_c), .D(n5499));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3422_3423 (.Q(\REG.mem_35_8 ), .C(FIFO_CLK_c), .D(n5498));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3419_3420 (.Q(\REG.mem_35_7 ), .C(FIFO_CLK_c), .D(n5497));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3416_3417 (.Q(\REG.mem_35_6 ), .C(FIFO_CLK_c), .D(n5496));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3413_3414 (.Q(\REG.mem_35_5 ), .C(FIFO_CLK_c), .D(n5495));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3410_3411 (.Q(\REG.mem_35_4 ), .C(FIFO_CLK_c), .D(n5494));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3407_3408 (.Q(\REG.mem_35_3 ), .C(FIFO_CLK_c), .D(n5493));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3404_3405 (.Q(\REG.mem_35_2 ), .C(FIFO_CLK_c), .D(n5492));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3401_3402 (.Q(\REG.mem_35_1 ), .C(FIFO_CLK_c), .D(n5491));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3398_3399 (.Q(\REG.mem_35_0 ), .C(FIFO_CLK_c), .D(n5490));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3347_3348 (.Q(\REG.mem_34_15 ), .C(FIFO_CLK_c), .D(n5488));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3344_3345 (.Q(\REG.mem_34_14 ), .C(FIFO_CLK_c), .D(n5487));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3341_3342 (.Q(\REG.mem_34_13 ), .C(FIFO_CLK_c), .D(n5486));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3338_3339 (.Q(\REG.mem_34_12 ), .C(FIFO_CLK_c), .D(n5485));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3335_3336 (.Q(\REG.mem_34_11 ), .C(FIFO_CLK_c), .D(n5484));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3998_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_28_4 ), .O(n5381));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3998_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12861_bdd_4_lut (.I0(n12861), .I1(\REG.mem_25_11 ), .I2(\REG.mem_24_11 ), 
            .I3(rd_addr_r[1]), .O(n11507));
    defparam n12861_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11427 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_13 ), 
            .I2(\REG.mem_11_13 ), .I3(rd_addr_r[1]), .O(n13509));
    defparam rd_addr_r_0__bdd_4_lut_11427.LUT_INIT = 16'he4aa;
    SB_LUT4 n13509_bdd_4_lut (.I0(n13509), .I1(\REG.mem_9_13 ), .I2(\REG.mem_8_13 ), 
            .I3(rd_addr_r[1]), .O(n13512));
    defparam n13509_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i3332_3333 (.Q(\REG.mem_34_10 ), .C(FIFO_CLK_c), .D(n5483));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3329_3330 (.Q(\REG.mem_34_9 ), .C(FIFO_CLK_c), .D(n5482));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3326_3327 (.Q(\REG.mem_34_8 ), .C(FIFO_CLK_c), .D(n5481));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3323_3324 (.Q(\REG.mem_34_7 ), .C(FIFO_CLK_c), .D(n5480));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3320_3321 (.Q(\REG.mem_34_6 ), .C(FIFO_CLK_c), .D(n5479));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3317_3318 (.Q(\REG.mem_34_5 ), .C(FIFO_CLK_c), .D(n5478));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3314_3315 (.Q(\REG.mem_34_4 ), .C(FIFO_CLK_c), .D(n5477));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3311_3312 (.Q(\REG.mem_34_3 ), .C(FIFO_CLK_c), .D(n5476));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3308_3309 (.Q(\REG.mem_34_2 ), .C(FIFO_CLK_c), .D(n5475));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3305_3306 (.Q(\REG.mem_34_1 ), .C(FIFO_CLK_c), .D(n5474));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3302_3303 (.Q(\REG.mem_34_0 ), .C(FIFO_CLK_c), .D(n5473));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3251_3252 (.Q(\REG.mem_33_15 ), .C(FIFO_CLK_c), .D(n5472));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3248_3249 (.Q(\REG.mem_33_14 ), .C(FIFO_CLK_c), .D(n5471));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3245_3246 (.Q(\REG.mem_33_13 ), .C(FIFO_CLK_c), .D(n5470));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3242_3243 (.Q(\REG.mem_33_12 ), .C(FIFO_CLK_c), .D(n5469));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3239_3240 (.Q(\REG.mem_33_11 ), .C(FIFO_CLK_c), .D(n5468));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10887 (.I0(rd_addr_r[3]), .I1(n12840), 
            .I2(n11233), .I3(rd_addr_r[4]), .O(n12855));
    defparam rd_addr_r_3__bdd_4_lut_10887.LUT_INIT = 16'he4aa;
    SB_LUT4 n12855_bdd_4_lut (.I0(n12855), .I1(n11230), .I2(n11229), .I3(rd_addr_r[4]), 
            .O(n12858));
    defparam n12855_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3997_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_28_3 ), .O(n5380));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3997_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11422 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_50_0 ), 
            .I2(\REG.mem_51_0 ), .I3(rd_addr_r[1]), .O(n13503));
    defparam rd_addr_r_0__bdd_4_lut_11422.LUT_INIT = 16'he4aa;
    SB_DFF i3236_3237 (.Q(\REG.mem_33_10 ), .C(FIFO_CLK_c), .D(n5467));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3233_3234 (.Q(\REG.mem_33_9 ), .C(FIFO_CLK_c), .D(n5466));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3230_3231 (.Q(\REG.mem_33_8 ), .C(FIFO_CLK_c), .D(n5465));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3227_3228 (.Q(\REG.mem_33_7 ), .C(FIFO_CLK_c), .D(n5464));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3224_3225 (.Q(\REG.mem_33_6 ), .C(FIFO_CLK_c), .D(n5463));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3221_3222 (.Q(\REG.mem_33_5 ), .C(FIFO_CLK_c), .D(n5462));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3218_3219 (.Q(\REG.mem_33_4 ), .C(FIFO_CLK_c), .D(n5461));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3215_3216 (.Q(\REG.mem_33_3 ), .C(FIFO_CLK_c), .D(n5460));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3212_3213 (.Q(\REG.mem_33_2 ), .C(FIFO_CLK_c), .D(n5459));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3209_3210 (.Q(\REG.mem_33_1 ), .C(FIFO_CLK_c), .D(n5458));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3206_3207 (.Q(\REG.mem_33_0 ), .C(FIFO_CLK_c), .D(n5457));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3155_3156 (.Q(\REG.mem_32_15 ), .C(FIFO_CLK_c), .D(n5456));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3152_3153 (.Q(\REG.mem_32_14 ), .C(FIFO_CLK_c), .D(n5455));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3149_3150 (.Q(\REG.mem_32_13 ), .C(FIFO_CLK_c), .D(n5454));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3146_3147 (.Q(\REG.mem_32_12 ), .C(FIFO_CLK_c), .D(n5453));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3996_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_28_2 ), .O(n5379));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3996_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3995_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_28_1 ), .O(n5378));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3995_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3994_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_28_0 ), .O(n5377));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3994_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3143_3144 (.Q(\REG.mem_32_11 ), .C(FIFO_CLK_c), .D(n5452));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4025_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_29_15 ), .O(n5408));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4025_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3140_3141 (.Q(\REG.mem_32_10 ), .C(FIFO_CLK_c), .D(n5451));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3137_3138 (.Q(\REG.mem_32_9 ), .C(FIFO_CLK_c), .D(n5450));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3134_3135 (.Q(\REG.mem_32_8 ), .C(FIFO_CLK_c), .D(n5449));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3131_3132 (.Q(\REG.mem_32_7 ), .C(FIFO_CLK_c), .D(n5448));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3128_3129 (.Q(\REG.mem_32_6 ), .C(FIFO_CLK_c), .D(n5447));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3125_3126 (.Q(\REG.mem_32_5 ), .C(FIFO_CLK_c), .D(n5446));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3122_3123 (.Q(\REG.mem_32_4 ), .C(FIFO_CLK_c), .D(n5445));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3119_3120 (.Q(\REG.mem_32_3 ), .C(FIFO_CLK_c), .D(n5444));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3116_3117 (.Q(\REG.mem_32_2 ), .C(FIFO_CLK_c), .D(n5443));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3113_3114 (.Q(\REG.mem_32_1 ), .C(FIFO_CLK_c), .D(n5442));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3110_3111 (.Q(\REG.mem_32_0 ), .C(FIFO_CLK_c), .D(n5441));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3059_3060 (.Q(\REG.mem_31_15 ), .C(FIFO_CLK_c), .D(n5440));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3056_3057 (.Q(\REG.mem_31_14 ), .C(FIFO_CLK_c), .D(n5439));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3053_3054 (.Q(\REG.mem_31_13 ), .C(FIFO_CLK_c), .D(n5438));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3050_3051 (.Q(\REG.mem_31_12 ), .C(FIFO_CLK_c), .D(n5437));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11152 (.I0(rd_addr_r[2]), .I1(n10853), 
            .I2(n10946), .I3(rd_addr_r[3]), .O(n12849));
    defparam rd_addr_r_2__bdd_4_lut_11152.LUT_INIT = 16'he4aa;
    SB_LUT4 n12849_bdd_4_lut (.I0(n12849), .I1(n11876), .I2(n11864), .I3(rd_addr_r[3]), 
            .O(n11510));
    defparam n12849_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13503_bdd_4_lut (.I0(n13503), .I1(\REG.mem_49_0 ), .I2(\REG.mem_48_0 ), 
            .I3(rd_addr_r[1]), .O(n11819));
    defparam n13503_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i3047_3048 (.Q(\REG.mem_31_11 ), .C(FIFO_CLK_c), .D(n5436));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_r_6__I_0_141_7_lut (.I0(GND_net), .I1(wr_addr_r[5]), 
            .I2(GND_net), .I3(n10009), .O(wr_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4024_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_29_14 ), .O(n5407));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4024_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3044_3045 (.Q(\REG.mem_31_10 ), .C(FIFO_CLK_c), .D(n5435));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3041_3042 (.Q(\REG.mem_31_9 ), .C(FIFO_CLK_c), .D(n5434));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3038_3039 (.Q(\REG.mem_31_8 ), .C(FIFO_CLK_c), .D(n5433));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3035_3036 (.Q(\REG.mem_31_7 ), .C(FIFO_CLK_c), .D(n5432));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3032_3033 (.Q(\REG.mem_31_6 ), .C(FIFO_CLK_c), .D(n5431));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3029_3030 (.Q(\REG.mem_31_5 ), .C(FIFO_CLK_c), .D(n5430));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3026_3027 (.Q(\REG.mem_31_4 ), .C(FIFO_CLK_c), .D(n5429));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3023_3024 (.Q(\REG.mem_31_3 ), .C(FIFO_CLK_c), .D(n5428));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3020_3021 (.Q(\REG.mem_31_2 ), .C(FIFO_CLK_c), .D(n5427));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3017_3018 (.Q(\REG.mem_31_1 ), .C(FIFO_CLK_c), .D(n5426));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3014_3015 (.Q(\REG.mem_31_0 ), .C(FIFO_CLK_c), .D(n5425));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2963_2964 (.Q(\REG.mem_30_15 ), .C(FIFO_CLK_c), .D(n5424));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2960_2961 (.Q(\REG.mem_30_14 ), .C(FIFO_CLK_c), .D(n5423));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2957_2958 (.Q(\REG.mem_30_13 ), .C(FIFO_CLK_c), .D(n5422));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2954_2955 (.Q(\REG.mem_30_12 ), .C(FIFO_CLK_c), .D(n5421));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2951_2952 (.Q(\REG.mem_30_11 ), .C(FIFO_CLK_c), .D(n5420));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4023_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_29_13 ), .O(n5406));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4023_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4022_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_29_12 ), .O(n5405));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4022_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4021_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_29_11 ), .O(n5404));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4021_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut (.I0(dc32_fifo_almost_full), .I1(DEBUG_1_c_c), .I2(GND_net), 
            .I3(GND_net), .O(write_to_dc32_fifo_latched_N_425));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4020_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_29_10 ), .O(n5403));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4020_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11417 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_46_13 ), 
            .I2(\REG.mem_47_13 ), .I3(rd_addr_r[1]), .O(n13497));
    defparam rd_addr_r_0__bdd_4_lut_11417.LUT_INIT = 16'he4aa;
    SB_LUT4 n13497_bdd_4_lut (.I0(n13497), .I1(\REG.mem_45_13 ), .I2(\REG.mem_44_13 ), 
            .I3(rd_addr_r[1]), .O(n11333));
    defparam n13497_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4019_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_29_9 ), .O(n5402));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4019_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10882 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_18_6 ), 
            .I2(\REG.mem_19_6 ), .I3(rd_addr_r[1]), .O(n12843));
    defparam rd_addr_r_0__bdd_4_lut_10882.LUT_INIT = 16'he4aa;
    SB_DFF i2948_2949 (.Q(\REG.mem_30_10 ), .C(FIFO_CLK_c), .D(n5419));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2945_2946 (.Q(\REG.mem_30_9 ), .C(FIFO_CLK_c), .D(n5418));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2942_2943 (.Q(\REG.mem_30_8 ), .C(FIFO_CLK_c), .D(n5417));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2939_2940 (.Q(\REG.mem_30_7 ), .C(FIFO_CLK_c), .D(n5416));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2936_2937 (.Q(\REG.mem_30_6 ), .C(FIFO_CLK_c), .D(n5415));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2933_2934 (.Q(\REG.mem_30_5 ), .C(FIFO_CLK_c), .D(n5414));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2930_2931 (.Q(\REG.mem_30_4 ), .C(FIFO_CLK_c), .D(n5413));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2927_2928 (.Q(\REG.mem_30_3 ), .C(FIFO_CLK_c), .D(n5412));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2924_2925 (.Q(\REG.mem_30_2 ), .C(FIFO_CLK_c), .D(n5411));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2921_2922 (.Q(\REG.mem_30_1 ), .C(FIFO_CLK_c), .D(n5410));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2918_2919 (.Q(\REG.mem_30_0 ), .C(FIFO_CLK_c), .D(n5409));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2867_2868 (.Q(\REG.mem_29_15 ), .C(FIFO_CLK_c), .D(n5408));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2864_2865 (.Q(\REG.mem_29_14 ), .C(FIFO_CLK_c), .D(n5407));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2861_2862 (.Q(\REG.mem_29_13 ), .C(FIFO_CLK_c), .D(n5406));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2858_2859 (.Q(\REG.mem_29_12 ), .C(FIFO_CLK_c), .D(n5405));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2855_2856 (.Q(\REG.mem_29_11 ), .C(FIFO_CLK_c), .D(n5404));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10268 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_46_15 ), 
            .I2(\REG.mem_47_15 ), .I3(rd_addr_r[1]), .O(n12111));
    defparam rd_addr_r_0__bdd_4_lut_10268.LUT_INIT = 16'he4aa;
    SB_LUT4 n12843_bdd_4_lut (.I0(n12843), .I1(\REG.mem_17_6 ), .I2(\REG.mem_16_6 ), 
            .I3(rd_addr_r[1]), .O(n10961));
    defparam n12843_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4018_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_29_8 ), .O(n5401));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4018_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4017_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_29_7 ), .O(n5400));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4017_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4016_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_29_6 ), .O(n5399));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4016_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i2_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[1] ), .O(wr_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4015_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_29_5 ), .O(n5398));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4015_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4014_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_29_4 ), .O(n5397));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4014_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4013_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_29_3 ), .O(n5396));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4013_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4012_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_29_2 ), .O(n5395));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4012_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4011_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_29_1 ), .O(n5394));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4011_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i3_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[3] ), .O(wr_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i3_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10360 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_9 ), 
            .I2(\REG.mem_11_9 ), .I3(rd_addr_r[1]), .O(n12213));
    defparam rd_addr_r_0__bdd_4_lut_10360.LUT_INIT = 16'he4aa;
    SB_LUT4 i4010_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_29_0 ), .O(n5393));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4010_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11412 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_46_6 ), 
            .I2(\REG.mem_47_6 ), .I3(rd_addr_r[1]), .O(n13491));
    defparam rd_addr_r_0__bdd_4_lut_11412.LUT_INIT = 16'he4aa;
    SB_LUT4 i4073_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_32_15 ), .O(n5456));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4073_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4072_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_32_14 ), .O(n5455));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4072_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12213_bdd_4_lut (.I0(n12213), .I1(\REG.mem_9_9 ), .I2(\REG.mem_8_9 ), 
            .I3(rd_addr_r[1]), .O(n12216));
    defparam n12213_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13491_bdd_4_lut (.I0(n13491), .I1(\REG.mem_45_6 ), .I2(\REG.mem_44_6 ), 
            .I3(rd_addr_r[1]), .O(n11336));
    defparam n13491_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2852_2853 (.Q(\REG.mem_29_10 ), .C(FIFO_CLK_c), .D(n5403));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4071_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_32_13 ), .O(n5454));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4071_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2849_2850 (.Q(\REG.mem_29_9 ), .C(FIFO_CLK_c), .D(n5402));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2846_2847 (.Q(\REG.mem_29_8 ), .C(FIFO_CLK_c), .D(n5401));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2843_2844 (.Q(\REG.mem_29_7 ), .C(FIFO_CLK_c), .D(n5400));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2840_2841 (.Q(\REG.mem_29_6 ), .C(FIFO_CLK_c), .D(n5399));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2837_2838 (.Q(\REG.mem_29_5 ), .C(FIFO_CLK_c), .D(n5398));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2834_2835 (.Q(\REG.mem_29_4 ), .C(FIFO_CLK_c), .D(n5397));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2831_2832 (.Q(\REG.mem_29_3 ), .C(FIFO_CLK_c), .D(n5396));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2828_2829 (.Q(\REG.mem_29_2 ), .C(FIFO_CLK_c), .D(n5395));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2825_2826 (.Q(\REG.mem_29_1 ), .C(FIFO_CLK_c), .D(n5394));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2822_2823 (.Q(\REG.mem_29_0 ), .C(FIFO_CLK_c), .D(n5393));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2771_2772 (.Q(\REG.mem_28_15 ), .C(FIFO_CLK_c), .D(n5392));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2768_2769 (.Q(\REG.mem_28_14 ), .C(FIFO_CLK_c), .D(n5391));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2765_2766 (.Q(\REG.mem_28_13 ), .C(FIFO_CLK_c), .D(n5390));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2762_2763 (.Q(\REG.mem_28_12 ), .C(FIFO_CLK_c), .D(n5389));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2759_2760 (.Q(\REG.mem_28_11 ), .C(FIFO_CLK_c), .D(n5388));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2756_2757 (.Q(\REG.mem_28_10 ), .C(FIFO_CLK_c), .D(n5387));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4070_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_32_12 ), .O(n5453));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4070_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10902 (.I0(rd_addr_r[1]), .I1(n11061), 
            .I2(n11062), .I3(rd_addr_r[2]), .O(n12837));
    defparam rd_addr_r_1__bdd_4_lut_10902.LUT_INIT = 16'he4aa;
    SB_LUT4 i4069_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_32_11 ), .O(n5452));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4069_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4068_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_32_10 ), .O(n5451));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4068_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4067_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_32_9 ), .O(n5450));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4067_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4066_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_32_8 ), .O(n5449));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4066_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2753_2754 (.Q(\REG.mem_28_9 ), .C(FIFO_CLK_c), .D(n5386));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4065_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_32_7 ), .O(n5448));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4065_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4650_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(wr_sig_mv_w), .I3(reset_per_frame), .O(n6033));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i4650_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i4064_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_32_6 ), .O(n5447));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4064_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4063_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_32_5 ), .O(n5446));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4063_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4062_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_32_4 ), .O(n5445));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4062_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4061_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_32_3 ), .O(n5444));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4061_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11407 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_13 ), 
            .I2(\REG.mem_15_13 ), .I3(rd_addr_r[1]), .O(n13485));
    defparam rd_addr_r_0__bdd_4_lut_11407.LUT_INIT = 16'he4aa;
    SB_LUT4 i4060_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_32_2 ), .O(n5443));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4060_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4059_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_32_1 ), .O(n5442));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4059_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13485_bdd_4_lut (.I0(n13485), .I1(\REG.mem_13_13 ), .I2(\REG.mem_12_13 ), 
            .I3(rd_addr_r[1]), .O(n13488));
    defparam n13485_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2750_2751 (.Q(\REG.mem_28_8 ), .C(FIFO_CLK_c), .D(n5385));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2747_2748 (.Q(\REG.mem_28_7 ), .C(FIFO_CLK_c), .D(n5384));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2744_2745 (.Q(\REG.mem_28_6 ), .C(FIFO_CLK_c), .D(n5383));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2741_2742 (.Q(\REG.mem_28_5 ), .C(FIFO_CLK_c), .D(n5382));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2738_2739 (.Q(\REG.mem_28_4 ), .C(FIFO_CLK_c), .D(n5381));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2735_2736 (.Q(\REG.mem_28_3 ), .C(FIFO_CLK_c), .D(n5380));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2732_2733 (.Q(\REG.mem_28_2 ), .C(FIFO_CLK_c), .D(n5379));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2729_2730 (.Q(\REG.mem_28_1 ), .C(FIFO_CLK_c), .D(n5378));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2726_2727 (.Q(\REG.mem_28_0 ), .C(FIFO_CLK_c), .D(n5377));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2675_2676 (.Q(\REG.mem_27_15 ), .C(FIFO_CLK_c), .D(n5376));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2672_2673 (.Q(\REG.mem_27_14 ), .C(FIFO_CLK_c), .D(n5375));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2669_2670 (.Q(\REG.mem_27_13 ), .C(FIFO_CLK_c), .D(n5374));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2666_2667 (.Q(\REG.mem_27_12 ), .C(FIFO_CLK_c), .D(n5373));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2663_2664 (.Q(\REG.mem_27_11 ), .C(FIFO_CLK_c), .D(n5372));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2660_2661 (.Q(\REG.mem_27_10 ), .C(FIFO_CLK_c), .D(n5371));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2657_2658 (.Q(\REG.mem_27_9 ), .C(FIFO_CLK_c), .D(n5370));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i134_135 (.Q(\REG.mem_1_0 ), .C(FIFO_CLK_c), .D(n4884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4058_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_32_0 ), .O(n5441));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4058_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4596_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_61_15 ), .O(n5979));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4596_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12837_bdd_4_lut (.I0(n12837), .I1(n11038), .I2(n11037), .I3(rd_addr_r[2]), 
            .O(n12840));
    defparam n12837_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4595_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_61_14 ), .O(n5978));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4595_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_r_6__I_0_inv_0_i7_1_lut (.I0(rp_sync2_r[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1212[6]));   // src/fifo_dc_32_lut_gen.v(212[47:78])
    defparam wr_addr_r_6__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4594_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_61_13 ), .O(n5977));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4594_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i4_2_lut_4_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[3] ), .O(wr_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i4_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11402 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_30_1 ), 
            .I2(\REG.mem_31_1 ), .I3(rd_addr_r[1]), .O(n13479));
    defparam rd_addr_r_0__bdd_4_lut_11402.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i88_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n56));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i88_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 n13479_bdd_4_lut (.I0(n13479), .I1(\REG.mem_29_1 ), .I2(\REG.mem_28_1 ), 
            .I3(rd_addr_r[1]), .O(n13482));
    defparam n13479_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4593_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_61_12 ), .O(n5976));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4593_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4592_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_61_11 ), .O(n5975));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4592_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11397 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_9 ), 
            .I2(\REG.mem_15_9 ), .I3(rd_addr_r[1]), .O(n13473));
    defparam rd_addr_r_0__bdd_4_lut_11397.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10867 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_15 ), 
            .I2(\REG.mem_11_15 ), .I3(rd_addr_r[1]), .O(n12831));
    defparam rd_addr_r_0__bdd_4_lut_10867.LUT_INIT = 16'he4aa;
    SB_DFF i2654_2655 (.Q(\REG.mem_27_8 ), .C(FIFO_CLK_c), .D(n5369));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12831_bdd_4_lut (.I0(n12831), .I1(\REG.mem_9_15 ), .I2(\REG.mem_8_15 ), 
            .I3(rd_addr_r[1]), .O(n12834));
    defparam n12831_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4591_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_61_10 ), .O(n5974));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4591_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2651_2652 (.Q(\REG.mem_27_7 ), .C(FIFO_CLK_c), .D(n5368));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2648_2649 (.Q(\REG.mem_27_6 ), .C(FIFO_CLK_c), .D(n5367));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2645_2646 (.Q(\REG.mem_27_5 ), .C(FIFO_CLK_c), .D(n5366));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2642_2643 (.Q(\REG.mem_27_4 ), .C(FIFO_CLK_c), .D(n5365));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2639_2640 (.Q(\REG.mem_27_3 ), .C(FIFO_CLK_c), .D(n5364));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2636_2637 (.Q(\REG.mem_27_2 ), .C(FIFO_CLK_c), .D(n5363));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2633_2634 (.Q(\REG.mem_27_1 ), .C(FIFO_CLK_c), .D(n5362));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2630_2631 (.Q(\REG.mem_27_0 ), .C(FIFO_CLK_c), .D(n5361));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2579_2580 (.Q(\REG.mem_26_15 ), .C(FIFO_CLK_c), .D(n5360));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2576_2577 (.Q(\REG.mem_26_14 ), .C(FIFO_CLK_c), .D(n5359));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2573_2574 (.Q(\REG.mem_26_13 ), .C(FIFO_CLK_c), .D(n5358));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2570_2571 (.Q(\REG.mem_26_12 ), .C(FIFO_CLK_c), .D(n5357));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2567_2568 (.Q(\REG.mem_26_11 ), .C(FIFO_CLK_c), .D(n5356));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2564_2565 (.Q(\REG.mem_26_10 ), .C(FIFO_CLK_c), .D(n5355));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2561_2562 (.Q(\REG.mem_26_9 ), .C(FIFO_CLK_c), .D(n5354));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2558_2559 (.Q(\REG.mem_26_8 ), .C(FIFO_CLK_c), .D(n5353));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4590_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_61_9 ), .O(n5973));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4590_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10857 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_7 ), 
            .I2(\REG.mem_11_7 ), .I3(rd_addr_r[1]), .O(n12825));
    defparam rd_addr_r_0__bdd_4_lut_10857.LUT_INIT = 16'he4aa;
    SB_LUT4 i4589_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_61_8 ), .O(n5972));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4589_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2555_2556 (.Q(\REG.mem_26_7 ), .C(FIFO_CLK_c), .D(n5352));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13473_bdd_4_lut (.I0(n13473), .I1(\REG.mem_13_9 ), .I2(\REG.mem_12_9 ), 
            .I3(rd_addr_r[1]), .O(n13476));
    defparam n13473_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4588_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_61_7 ), .O(n5971));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4588_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4587_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_61_6 ), .O(n5970));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4587_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4586_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_61_5 ), .O(n5969));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4586_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2552_2553 (.Q(\REG.mem_26_6 ), .C(FIFO_CLK_c), .D(n5351));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i5_2_lut_4_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[5] ), .O(wr_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_DFF i2549_2550 (.Q(\REG.mem_26_5 ), .C(FIFO_CLK_c), .D(n5350));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2546_2547 (.Q(\REG.mem_26_4 ), .C(FIFO_CLK_c), .D(n5349));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2543_2544 (.Q(\REG.mem_26_3 ), .C(FIFO_CLK_c), .D(n5348));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2540_2541 (.Q(\REG.mem_26_2 ), .C(FIFO_CLK_c), .D(n5347));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2537_2538 (.Q(\REG.mem_26_1 ), .C(FIFO_CLK_c), .D(n5346));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2534_2535 (.Q(\REG.mem_26_0 ), .C(FIFO_CLK_c), .D(n5345));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2483_2484 (.Q(\REG.mem_25_15 ), .C(FIFO_CLK_c), .D(n5344));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2480_2481 (.Q(\REG.mem_25_14 ), .C(FIFO_CLK_c), .D(n5343));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2477_2478 (.Q(\REG.mem_25_13 ), .C(FIFO_CLK_c), .D(n5342));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2474_2475 (.Q(\REG.mem_25_12 ), .C(FIFO_CLK_c), .D(n5341));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2471_2472 (.Q(\REG.mem_25_11 ), .C(FIFO_CLK_c), .D(n5340));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2468_2469 (.Q(\REG.mem_25_10 ), .C(FIFO_CLK_c), .D(n5339));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2465_2466 (.Q(\REG.mem_25_9 ), .C(FIFO_CLK_c), .D(n5338));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2462_2463 (.Q(\REG.mem_25_8 ), .C(FIFO_CLK_c), .D(n5337));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2459_2460 (.Q(\REG.mem_25_7 ), .C(FIFO_CLK_c), .D(n5336));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_r_6__I_0_135_i2_3_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(wr_sig_mv_w), .I3(GND_net), .O(\wr_addr_nxt_c[1] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11392 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_18_13 ), 
            .I2(\REG.mem_19_13 ), .I3(rd_addr_r[1]), .O(n13467));
    defparam rd_addr_r_0__bdd_4_lut_11392.LUT_INIT = 16'he4aa;
    SB_LUT4 n12825_bdd_4_lut (.I0(n12825), .I1(\REG.mem_9_7 ), .I2(\REG.mem_8_7 ), 
            .I3(rd_addr_r[1]), .O(n12828));
    defparam n12825_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4585_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_61_4 ), .O(n5968));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4585_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4584_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_61_3 ), .O(n5967));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4584_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13467_bdd_4_lut (.I0(n13467), .I1(\REG.mem_17_13 ), .I2(\REG.mem_16_13 ), 
            .I3(rd_addr_r[1]), .O(n13470));
    defparam n13467_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2456_2457 (.Q(\REG.mem_25_6 ), .C(FIFO_CLK_c), .D(n5335));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2453_2454 (.Q(\REG.mem_25_5 ), .C(FIFO_CLK_c), .D(n5334));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2450_2451 (.Q(\REG.mem_25_4 ), .C(FIFO_CLK_c), .D(n5333));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4583_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_61_2 ), .O(n5966));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4583_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9511_3_lut (.I0(\REG.mem_56_7 ), .I1(\REG.mem_57_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11361));
    defparam i9511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4582_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_61_1 ), .O(n5965));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4582_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2447_2448 (.Q(\REG.mem_25_3 ), .C(FIFO_CLK_c), .D(n5332));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2444_2445 (.Q(\REG.mem_25_2 ), .C(FIFO_CLK_c), .D(n5331));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4581_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_61_0 ), .O(n5964));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4581_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9512_3_lut (.I0(\REG.mem_58_7 ), .I1(\REG.mem_59_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11362));
    defparam i9512_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2441_2442 (.Q(\REG.mem_25_1 ), .C(FIFO_CLK_c), .D(n5330));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2438_2439 (.Q(\REG.mem_25_0 ), .C(FIFO_CLK_c), .D(n5329));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2387_2388 (.Q(\REG.mem_24_15 ), .C(FIFO_CLK_c), .D(n5328));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2384_2385 (.Q(\REG.mem_24_14 ), .C(FIFO_CLK_c), .D(n5327));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2381_2382 (.Q(\REG.mem_24_13 ), .C(FIFO_CLK_c), .D(n5326));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2378_2379 (.Q(\REG.mem_24_12 ), .C(FIFO_CLK_c), .D(n5325));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2375_2376 (.Q(\REG.mem_24_11 ), .C(FIFO_CLK_c), .D(n5324));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2372_2373 (.Q(\REG.mem_24_10 ), .C(FIFO_CLK_c), .D(n5323));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2369_2370 (.Q(\REG.mem_24_9 ), .C(FIFO_CLK_c), .D(n5322));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2366_2367 (.Q(\REG.mem_24_8 ), .C(FIFO_CLK_c), .D(n5321));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2363_2364 (.Q(\REG.mem_24_7 ), .C(FIFO_CLK_c), .D(n5320));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2360_2361 (.Q(\REG.mem_24_6 ), .C(FIFO_CLK_c), .D(n5319));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2357_2358 (.Q(\REG.mem_24_5 ), .C(FIFO_CLK_c), .D(n5318));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2354_2355 (.Q(\REG.mem_24_4 ), .C(FIFO_CLK_c), .D(n5317));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2351_2352 (.Q(\REG.mem_24_3 ), .C(FIFO_CLK_c), .D(n5316));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2348_2349 (.Q(\REG.mem_24_2 ), .C(FIFO_CLK_c), .D(n5315));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2345_2346 (.Q(\REG.mem_24_1 ), .C(FIFO_CLK_c), .D(n5314));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4648_2_lut_4_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(wr_sig_mv_w), .I3(reset_per_frame), .O(n6031));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i4648_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 EnabledDecoder_2_i96_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n52));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i96_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10852 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_30_12 ), 
            .I2(\REG.mem_31_12 ), .I3(rd_addr_r[1]), .O(n12819));
    defparam rd_addr_r_0__bdd_4_lut_10852.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11387 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_54_0 ), 
            .I2(\REG.mem_55_0 ), .I3(rd_addr_r[1]), .O(n13461));
    defparam rd_addr_r_0__bdd_4_lut_11387.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i95_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n20));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i95_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 n13461_bdd_4_lut (.I0(n13461), .I1(\REG.mem_53_0 ), .I2(\REG.mem_52_0 ), 
            .I3(rd_addr_r[1]), .O(n11828));
    defparam n13461_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2342_2343 (.Q(\REG.mem_24_0 ), .C(FIFO_CLK_c), .D(n5307));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9533_3_lut (.I0(\REG.mem_62_7 ), .I1(\REG.mem_63_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11383));
    defparam i9533_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2291_2292 (.Q(\REG.mem_23_15 ), .C(FIFO_CLK_c), .D(n5306));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2288_2289 (.Q(\REG.mem_23_14 ), .C(FIFO_CLK_c), .D(n5305));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2285_2286 (.Q(\REG.mem_23_13 ), .C(FIFO_CLK_c), .D(n5304));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2282_2283 (.Q(\REG.mem_23_12 ), .C(FIFO_CLK_c), .D(n5303));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3567_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_2_2 ), .O(n4950));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3567_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i2279_2280 (.Q(\REG.mem_23_11 ), .C(FIFO_CLK_c), .D(n5302));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2276_2277 (.Q(\REG.mem_23_10 ), .C(FIFO_CLK_c), .D(n5301));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2273_2274 (.Q(\REG.mem_23_9 ), .C(FIFO_CLK_c), .D(n5300));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2270_2271 (.Q(\REG.mem_23_8 ), .C(FIFO_CLK_c), .D(n5299));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2267_2268 (.Q(\REG.mem_23_7 ), .C(FIFO_CLK_c), .D(n5298));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2264_2265 (.Q(\REG.mem_23_6 ), .C(FIFO_CLK_c), .D(n5297));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2261_2262 (.Q(\REG.mem_23_5 ), .C(FIFO_CLK_c), .D(n5296));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2258_2259 (.Q(\REG.mem_23_4 ), .C(FIFO_CLK_c), .D(n5295));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2255_2256 (.Q(\REG.mem_23_3 ), .C(FIFO_CLK_c), .D(n5294));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2252_2253 (.Q(\REG.mem_23_2 ), .C(FIFO_CLK_c), .D(n5293));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2249_2250 (.Q(\REG.mem_23_1 ), .C(FIFO_CLK_c), .D(n5292));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2246_2247 (.Q(\REG.mem_23_0 ), .C(FIFO_CLK_c), .D(n5291));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2195_2196 (.Q(\REG.mem_22_15 ), .C(FIFO_CLK_c), .D(n5290));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2192_2193 (.Q(\REG.mem_22_14 ), .C(FIFO_CLK_c), .D(n5289));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2189_2190 (.Q(\REG.mem_22_13 ), .C(FIFO_CLK_c), .D(n5288));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2186_2187 (.Q(\REG.mem_22_12 ), .C(FIFO_CLK_c), .D(n5287));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2183_2184 (.Q(\REG.mem_22_11 ), .C(FIFO_CLK_c), .D(n5286));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2180_2181 (.Q(\REG.mem_22_10 ), .C(FIFO_CLK_c), .D(n5285));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12819_bdd_4_lut (.I0(n12819), .I1(\REG.mem_29_12 ), .I2(\REG.mem_28_12 ), 
            .I3(rd_addr_r[1]), .O(n12822));
    defparam n12819_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9532_3_lut (.I0(\REG.mem_60_7 ), .I1(\REG.mem_61_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11382));
    defparam i9532_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR rd_grey_sync_r__i5 (.Q(\rd_grey_sync_r[5] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[5]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i4 (.Q(\rd_grey_sync_r[4] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[4]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i3 (.Q(\rd_grey_sync_r[3] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[3]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i2 (.Q(\rd_grey_sync_r[2] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[2]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i1 (.Q(\rd_grey_sync_r[1] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[1]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFF i2177_2178 (.Q(\REG.mem_22_9 ), .C(FIFO_CLK_c), .D(n5284));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9637_3_lut (.I0(\REG.mem_32_8 ), .I1(\REG.mem_33_8 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11487));
    defparam i9637_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2174_2175 (.Q(\REG.mem_22_8 ), .C(FIFO_CLK_c), .D(n5283));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2171_2172 (.Q(\REG.mem_22_7 ), .C(FIFO_CLK_c), .D(n5282));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2168_2169 (.Q(\REG.mem_22_6 ), .C(FIFO_CLK_c), .D(n5281));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2165_2166 (.Q(\REG.mem_22_5 ), .C(FIFO_CLK_c), .D(n5280));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2162_2163 (.Q(\REG.mem_22_4 ), .C(FIFO_CLK_c), .D(n5279));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2159_2160 (.Q(\REG.mem_22_3 ), .C(FIFO_CLK_c), .D(n5278));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2156_2157 (.Q(\REG.mem_22_2 ), .C(FIFO_CLK_c), .D(n5277));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2153_2154 (.Q(\REG.mem_22_1 ), .C(FIFO_CLK_c), .D(n5276));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2150_2151 (.Q(\REG.mem_22_0 ), .C(FIFO_CLK_c), .D(n5275));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2099_2100 (.Q(\REG.mem_21_15 ), .C(FIFO_CLK_c), .D(n5274));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2096_2097 (.Q(\REG.mem_21_14 ), .C(FIFO_CLK_c), .D(n5273));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2093_2094 (.Q(\REG.mem_21_13 ), .C(FIFO_CLK_c), .D(n5272));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2090_2091 (.Q(\REG.mem_21_12 ), .C(FIFO_CLK_c), .D(n5271));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2087_2088 (.Q(\REG.mem_21_11 ), .C(FIFO_CLK_c), .D(n5270));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2084_2085 (.Q(\REG.mem_21_10 ), .C(FIFO_CLK_c), .D(n5269));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11382 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_3 ), 
            .I2(\REG.mem_15_3 ), .I3(rd_addr_r[1]), .O(n13455));
    defparam rd_addr_r_0__bdd_4_lut_11382.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10847 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_38_9 ), 
            .I2(\REG.mem_39_9 ), .I3(rd_addr_r[1]), .O(n12813));
    defparam rd_addr_r_0__bdd_4_lut_10847.LUT_INIT = 16'he4aa;
    SB_LUT4 i3566_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_2_1 ), .O(n4949));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3566_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9638_3_lut (.I0(\REG.mem_34_8 ), .I1(\REG.mem_35_8 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11488));
    defparam i9638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_40 (.I0(wp_sync2_r[1]), .I1(wp_sync_w[2]), .I2(GND_net), 
            .I3(GND_net), .O(wp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_40.LUT_INIT = 16'h6666;
    SB_DFF i2081_2082 (.Q(\REG.mem_21_9 ), .C(FIFO_CLK_c), .D(n5268));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2078_2079 (.Q(\REG.mem_21_8 ), .C(FIFO_CLK_c), .D(n5267));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2075_2076 (.Q(\REG.mem_21_7 ), .C(FIFO_CLK_c), .D(n5266));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2072_2073 (.Q(\REG.mem_21_6 ), .C(FIFO_CLK_c), .D(n5265));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2069_2070 (.Q(\REG.mem_21_5 ), .C(FIFO_CLK_c), .D(n5264));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2066_2067 (.Q(\REG.mem_21_4 ), .C(FIFO_CLK_c), .D(n5263));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2063_2064 (.Q(\REG.mem_21_3 ), .C(FIFO_CLK_c), .D(n5262));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2060_2061 (.Q(\REG.mem_21_2 ), .C(FIFO_CLK_c), .D(n5261));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2057_2058 (.Q(\REG.mem_21_1 ), .C(FIFO_CLK_c), .D(n5260));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2054_2055 (.Q(\REG.mem_21_0 ), .C(FIFO_CLK_c), .D(n5259));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2003_2004 (.Q(\REG.mem_20_15 ), .C(FIFO_CLK_c), .D(n5258));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2000_2001 (.Q(\REG.mem_20_14 ), .C(FIFO_CLK_c), .D(n5257));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1997_1998 (.Q(\REG.mem_20_13 ), .C(FIFO_CLK_c), .D(n5256));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1994_1995 (.Q(\REG.mem_20_12 ), .C(FIFO_CLK_c), .D(n5255));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1991_1992 (.Q(\REG.mem_20_11 ), .C(FIFO_CLK_c), .D(n5254));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1988_1989 (.Q(\REG.mem_20_10 ), .C(FIFO_CLK_c), .D(n5253));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i1_2_lut_adj_41 (.I0(wp_sync2_r[3]), .I1(wp_sync_w[4]), .I2(GND_net), 
            .I3(GND_net), .O(wp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_41.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_42 (.I0(wp_sync2_r[6]), .I1(wp_sync2_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n4274));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_42.LUT_INIT = 16'h6666;
    SB_LUT4 i8923_4_lut (.I0(\rd_addr_r[0] ), .I1(rd_addr_r[4]), .I2(wp_sync_w[0]), 
            .I3(wp_sync_w[4]), .O(n10772));
    defparam i8923_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i1_1_lut (.I0(\rd_addr_r[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n13455_bdd_4_lut (.I0(n13455), .I1(\REG.mem_13_3 ), .I2(\REG.mem_12_3 ), 
            .I3(rd_addr_r[1]), .O(n10907));
    defparam n13455_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1985_1986 (.Q(\REG.mem_20_9 ), .C(FIFO_CLK_c), .D(n5252));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i2_1_lut (.I0(rd_addr_r[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n12813_bdd_4_lut (.I0(n12813), .I1(\REG.mem_37_9 ), .I2(\REG.mem_36_9 ), 
            .I3(rd_addr_r[1]), .O(n12816));
    defparam n12813_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10842 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_30_11 ), 
            .I2(\REG.mem_31_11 ), .I3(rd_addr_r[1]), .O(n12807));
    defparam rd_addr_r_0__bdd_4_lut_10842.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11377 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_8 ), 
            .I2(\REG.mem_11_8 ), .I3(rd_addr_r[1]), .O(n13449));
    defparam rd_addr_r_0__bdd_4_lut_11377.LUT_INIT = 16'he4aa;
    SB_LUT4 n13449_bdd_4_lut (.I0(n13449), .I1(\REG.mem_9_8 ), .I2(\REG.mem_8_8 ), 
            .I3(rd_addr_r[1]), .O(n13452));
    defparam n13449_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4085_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_33_11 ), .O(n5468));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4085_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8873_4_lut (.I0(rd_addr_r[5]), .I1(rd_addr_r[3]), .I2(n4274), 
            .I3(wp_sync_w[3]), .O(n10722));
    defparam i8873_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_2_lut_adj_43 (.I0(rd_addr_p1_w[4]), .I1(wp_sync_w[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4298));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_43.LUT_INIT = 16'h6666;
    SB_LUT4 n12807_bdd_4_lut (.I0(n12807), .I1(\REG.mem_29_11 ), .I2(\REG.mem_28_11 ), 
            .I3(rd_addr_r[1]), .O(n11519));
    defparam n12807_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut (.I0(rd_addr_p1_w[5]), .I1(rd_addr_p1_w[3]), .I2(n4274), 
            .I3(wp_sync_w[3]), .O(n10_c));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_44 (.I0(wp_sync2_r[6]), .I1(rd_addr_p1_w[1]), .I2(rd_addr_p1_w[6]), 
            .I3(wp_sync_w[1]), .O(n8_adj_1191));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i1_4_lut_adj_44.LUT_INIT = 16'h7bde;
    SB_DFF i1982_1983 (.Q(\REG.mem_20_8 ), .C(FIFO_CLK_c), .D(n5251));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5_4_lut (.I0(\rd_addr_p1_w[0] ), .I1(n10_c), .I2(n4298), 
            .I3(wp_sync_w[0]), .O(n12));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i5_4_lut.LUT_INIT = 16'hfdfe;
    SB_DFF i1979_1980 (.Q(\REG.mem_20_7 ), .C(FIFO_CLK_c), .D(n5250));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1976_1977 (.Q(\REG.mem_20_6 ), .C(FIFO_CLK_c), .D(n5249));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1973_1974 (.Q(\REG.mem_20_5 ), .C(FIFO_CLK_c), .D(n5248));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1970_1971 (.Q(\REG.mem_20_4 ), .C(FIFO_CLK_c), .D(n5247));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1967_1968 (.Q(\REG.mem_20_3 ), .C(FIFO_CLK_c), .D(n5246));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1964_1965 (.Q(\REG.mem_20_2 ), .C(FIFO_CLK_c), .D(n5245));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1961_1962 (.Q(\REG.mem_20_1 ), .C(FIFO_CLK_c), .D(n5244));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1958_1959 (.Q(\REG.mem_20_0 ), .C(FIFO_CLK_c), .D(n5243));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1907_1908 (.Q(\REG.mem_19_15 ), .C(FIFO_CLK_c), .D(n5242));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1904_1905 (.Q(\REG.mem_19_14 ), .C(FIFO_CLK_c), .D(n5241));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1901_1902 (.Q(\REG.mem_19_13 ), .C(FIFO_CLK_c), .D(n5240));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1898_1899 (.Q(\REG.mem_19_12 ), .C(FIFO_CLK_c), .D(n5239));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1895_1896 (.Q(\REG.mem_19_11 ), .C(FIFO_CLK_c), .D(n5238));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1892_1893 (.Q(\REG.mem_19_10 ), .C(FIFO_CLK_c), .D(n5237));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10837 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_54_1 ), 
            .I2(\REG.mem_55_1 ), .I3(rd_addr_r[1]), .O(n12801));
    defparam rd_addr_r_0__bdd_4_lut_10837.LUT_INIT = 16'he4aa;
    SB_LUT4 i8988_3_lut (.I0(n10766), .I1(n10722), .I2(n10772), .I3(GND_net), 
            .O(n10838));
    defparam i8988_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut (.I0(rd_addr_p1_w[2]), .I1(n12), .I2(n8_adj_1191), 
            .I3(wp_sync_w[2]), .O(n10130));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i6_4_lut.LUT_INIT = 16'hfdfe;
    SB_LUT4 empty_nxt_c_I_7_4_lut (.I0(n10130), .I1(n10838), .I2(DEBUG_3_c), 
            .I3(get_next_word), .O(empty_nxt_c_N_629));   // src/fifo_dc_32_lut_gen.v(555[46:103])
    defparam empty_nxt_c_I_7_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i9683_3_lut (.I0(\REG.mem_38_8 ), .I1(\REG.mem_39_8 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11533));
    defparam i9683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9682_3_lut (.I0(\REG.mem_36_8 ), .I1(\REG.mem_37_8 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11532));
    defparam i9682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9835_3_lut (.I0(\REG.mem_16_2 ), .I1(\REG.mem_17_2 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11685));
    defparam i9835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3565_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_2_0 ), .O(n4948));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3565_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3580_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_2_15 ), .O(n4963));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3580_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11372 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_50_13 ), 
            .I2(\REG.mem_51_13 ), .I3(rd_addr_r[1]), .O(n13443));
    defparam rd_addr_r_0__bdd_4_lut_11372.LUT_INIT = 16'he4aa;
    SB_LUT4 n12801_bdd_4_lut (.I0(n12801), .I1(\REG.mem_53_1 ), .I2(\REG.mem_52_1 ), 
            .I3(rd_addr_r[1]), .O(n12804));
    defparam n12801_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9836_3_lut (.I0(\REG.mem_18_2 ), .I1(\REG.mem_19_2 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11686));
    defparam i9836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13443_bdd_4_lut (.I0(n13443), .I1(\REG.mem_49_13 ), .I2(\REG.mem_48_13 ), 
            .I3(rd_addr_r[1]), .O(n11351));
    defparam n13443_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1889_1890 (.Q(\REG.mem_19_9 ), .C(FIFO_CLK_c), .D(n5236));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9878_3_lut (.I0(\REG.mem_22_2 ), .I1(\REG.mem_23_2 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11728));
    defparam i9878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9877_3_lut (.I0(\REG.mem_20_2 ), .I1(\REG.mem_21_2 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11727));
    defparam i9877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10832 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_34_11 ), 
            .I2(\REG.mem_35_11 ), .I3(rd_addr_r[1]), .O(n12795));
    defparam rd_addr_r_0__bdd_4_lut_10832.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11367 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_18_3 ), 
            .I2(\REG.mem_19_3 ), .I3(rd_addr_r[1]), .O(n13437));
    defparam rd_addr_r_0__bdd_4_lut_11367.LUT_INIT = 16'he4aa;
    SB_LUT4 n12795_bdd_4_lut (.I0(n12795), .I1(\REG.mem_33_11 ), .I2(\REG.mem_32_11 ), 
            .I3(rd_addr_r[1]), .O(n11525));
    defparam n12795_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1886_1887 (.Q(\REG.mem_19_8 ), .C(FIFO_CLK_c), .D(n5235));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1883_1884 (.Q(\REG.mem_19_7 ), .C(FIFO_CLK_c), .D(n5234));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1880_1881 (.Q(\REG.mem_19_6 ), .C(FIFO_CLK_c), .D(n5233));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1877_1878 (.Q(\REG.mem_19_5 ), .C(FIFO_CLK_c), .D(n5232));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1874_1875 (.Q(\REG.mem_19_4 ), .C(FIFO_CLK_c), .D(n5231));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1871_1872 (.Q(\REG.mem_19_3 ), .C(FIFO_CLK_c), .D(n5230));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1868_1869 (.Q(\REG.mem_19_2 ), .C(FIFO_CLK_c), .D(n5229));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1865_1866 (.Q(\REG.mem_19_1 ), .C(FIFO_CLK_c), .D(n5228));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1862_1863 (.Q(\REG.mem_19_0 ), .C(FIFO_CLK_c), .D(n5227));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1811_1812 (.Q(\REG.mem_18_15 ), .C(FIFO_CLK_c), .D(n5226));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1808_1809 (.Q(\REG.mem_18_14 ), .C(FIFO_CLK_c), .D(n5225));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1805_1806 (.Q(\REG.mem_18_13 ), .C(FIFO_CLK_c), .D(n5224));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1802_1803 (.Q(\REG.mem_18_12 ), .C(FIFO_CLK_c), .D(n5223));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1799_1800 (.Q(\REG.mem_18_11 ), .C(FIFO_CLK_c), .D(n5222));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1796_1797 (.Q(\REG.mem_18_10 ), .C(FIFO_CLK_c), .D(n5221));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1793_1794 (.Q(\REG.mem_18_9 ), .C(FIFO_CLK_c), .D(n5220));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_6__I_0_i1_3_lut (.I0(\rd_addr_r[0] ), .I1(\rd_addr_p1_w[0] ), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(rd_addr_nxt_c_6__N_498[0]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13437_bdd_4_lut (.I0(n13437), .I1(\REG.mem_17_3 ), .I2(\REG.mem_16_3 ), 
            .I3(rd_addr_r[1]), .O(n10910));
    defparam n13437_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9694_3_lut (.I0(\REG.mem_16_15 ), .I1(\REG.mem_17_15 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11544));
    defparam i9694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9695_3_lut (.I0(\REG.mem_18_15 ), .I1(\REG.mem_19_15 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11545));
    defparam i9695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9716_3_lut (.I0(\REG.mem_22_15 ), .I1(\REG.mem_23_15 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11566));
    defparam i9716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3579_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_2_14 ), .O(n4962));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3579_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9715_3_lut (.I0(\REG.mem_20_15 ), .I1(\REG.mem_21_15 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11565));
    defparam i9715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3578_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_2_13 ), .O(n4961));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3578_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4084_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_33_10 ), .O(n5467));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4084_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3577_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_2_12 ), .O(n4960));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3577_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1790_1791 (.Q(\REG.mem_18_8 ), .C(FIFO_CLK_c), .D(n5219));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1787_1788 (.Q(\REG.mem_18_7 ), .C(FIFO_CLK_c), .D(n5218));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1784_1785 (.Q(\REG.mem_18_6 ), .C(FIFO_CLK_c), .D(n5217));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1781_1782 (.Q(\REG.mem_18_5 ), .C(FIFO_CLK_c), .D(n5216));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1778_1779 (.Q(\REG.mem_18_4 ), .C(FIFO_CLK_c), .D(n5215));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1775_1776 (.Q(\REG.mem_18_3 ), .C(FIFO_CLK_c), .D(n5214));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1772_1773 (.Q(\REG.mem_18_2 ), .C(FIFO_CLK_c), .D(n5213));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1769_1770 (.Q(\REG.mem_18_1 ), .C(FIFO_CLK_c), .D(n5212));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1766_1767 (.Q(\REG.mem_18_0 ), .C(FIFO_CLK_c), .D(n5211));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1715_1716 (.Q(\REG.mem_17_15 ), .C(FIFO_CLK_c), .D(n5210));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1712_1713 (.Q(\REG.mem_17_14 ), .C(FIFO_CLK_c), .D(n5209));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1709_1710 (.Q(\REG.mem_17_13 ), .C(FIFO_CLK_c), .D(n5208));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1706_1707 (.Q(\REG.mem_17_12 ), .C(FIFO_CLK_c), .D(n5207));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1703_1704 (.Q(\REG.mem_17_11 ), .C(FIFO_CLK_c), .D(n5206));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1700_1701 (.Q(\REG.mem_17_10 ), .C(FIFO_CLK_c), .D(n5205));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1697_1698 (.Q(\REG.mem_17_9 ), .C(FIFO_CLK_c), .D(n5204));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3576_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_2_11 ), .O(n4959));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3576_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3575_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_2_10 ), .O(n4958));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3575_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3574_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_2_9 ), .O(n4957));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3574_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1694_1695 (.Q(\REG.mem_17_8 ), .C(FIFO_CLK_c), .D(n5203));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11502 (.I0(rd_addr_r[3]), .I1(n12600), 
            .I2(n10903), .I3(rd_addr_r[4]), .O(n13431));
    defparam rd_addr_r_3__bdd_4_lut_11502.LUT_INIT = 16'he4aa;
    SB_LUT4 i3573_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_2_8 ), .O(n4956));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3573_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3572_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_2_7 ), .O(n4955));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3572_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1691_1692 (.Q(\REG.mem_17_7 ), .C(FIFO_CLK_c), .D(n5202));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3571_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_2_6 ), .O(n4954));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3571_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4083_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_33_9 ), .O(n5466));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4083_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1688_1689 (.Q(\REG.mem_17_6 ), .C(FIFO_CLK_c), .D(n5201));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10827 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_50_3 ), 
            .I2(\REG.mem_51_3 ), .I3(rd_addr_r[1]), .O(n12789));
    defparam rd_addr_r_0__bdd_4_lut_10827.LUT_INIT = 16'he4aa;
    SB_LUT4 n13431_bdd_4_lut (.I0(n13431), .I1(n10879), .I2(n10878), .I3(rd_addr_r[4]), 
            .O(n13434));
    defparam n13431_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3570_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_2_5 ), .O(n4953));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3570_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12789_bdd_4_lut (.I0(n12789), .I1(\REG.mem_49_3 ), .I2(\REG.mem_48_3 ), 
            .I3(rd_addr_r[1]), .O(n10964));
    defparam n12789_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1685_1686 (.Q(\REG.mem_17_5 ), .C(FIFO_CLK_c), .D(n5200));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1682_1683 (.Q(\REG.mem_17_4 ), .C(FIFO_CLK_c), .D(n5199));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1679_1680 (.Q(\REG.mem_17_3 ), .C(FIFO_CLK_c), .D(n5198));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1676_1677 (.Q(\REG.mem_17_2 ), .C(FIFO_CLK_c), .D(n5197));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1673_1674 (.Q(\REG.mem_17_1 ), .C(FIFO_CLK_c), .D(n5196));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1670_1671 (.Q(\REG.mem_17_0 ), .C(FIFO_CLK_c), .D(n5195));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1619_1620 (.Q(\REG.mem_16_15 ), .C(FIFO_CLK_c), .D(n5190));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1616_1617 (.Q(\REG.mem_16_14 ), .C(FIFO_CLK_c), .D(n5188));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1613_1614 (.Q(\REG.mem_16_13 ), .C(FIFO_CLK_c), .D(n5187));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1610_1611 (.Q(\REG.mem_16_12 ), .C(FIFO_CLK_c), .D(n5186));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12111_bdd_4_lut (.I0(n12111), .I1(\REG.mem_45_15 ), .I2(\REG.mem_44_15 ), 
            .I3(rd_addr_r[1]), .O(n12114));
    defparam n12111_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1607_1608 (.Q(\REG.mem_16_11 ), .C(FIFO_CLK_c), .D(n5185));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10822 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_38_11 ), 
            .I2(\REG.mem_39_11 ), .I3(rd_addr_r[1]), .O(n12783));
    defparam rd_addr_r_0__bdd_4_lut_10822.LUT_INIT = 16'he4aa;
    SB_DFF i1604_1605 (.Q(\REG.mem_16_10 ), .C(FIFO_CLK_c), .D(n5184));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11362 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_26_8 ), 
            .I2(\REG.mem_27_8 ), .I3(rd_addr_r[1]), .O(n13425));
    defparam rd_addr_r_0__bdd_4_lut_11362.LUT_INIT = 16'he4aa;
    SB_LUT4 n12783_bdd_4_lut (.I0(n12783), .I1(\REG.mem_37_11 ), .I2(\REG.mem_36_11 ), 
            .I3(rd_addr_r[1]), .O(n11528));
    defparam n12783_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13425_bdd_4_lut (.I0(n13425), .I1(\REG.mem_25_8 ), .I2(\REG.mem_24_8 ), 
            .I3(rd_addr_r[1]), .O(n13428));
    defparam n13425_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9404_3_lut (.I0(\REG.mem_54_5 ), .I1(\REG.mem_55_5 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11254));
    defparam i9404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9403_3_lut (.I0(\REG.mem_52_5 ), .I1(\REG.mem_53_5 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11253));
    defparam i9403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11472 (.I0(rd_addr_r[2]), .I1(n13242), 
            .I2(n12210), .I3(rd_addr_r[3]), .O(n13419));
    defparam rd_addr_r_2__bdd_4_lut_11472.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10862 (.I0(rd_addr_r[1]), .I1(n11847), 
            .I2(n11848), .I3(rd_addr_r[2]), .O(n12777));
    defparam rd_addr_r_1__bdd_4_lut_10862.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10346 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_62_0 ), 
            .I2(\REG.mem_63_0 ), .I3(rd_addr_r[1]), .O(n12207));
    defparam rd_addr_r_0__bdd_4_lut_10346.LUT_INIT = 16'he4aa;
    SB_LUT4 n13419_bdd_4_lut (.I0(n13419), .I1(n11828), .I2(n11819), .I3(rd_addr_r[3]), 
            .O(n11834));
    defparam n13419_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12207_bdd_4_lut (.I0(n12207), .I1(\REG.mem_61_0 ), .I2(\REG.mem_60_0 ), 
            .I3(rd_addr_r[1]), .O(n12210));
    defparam n12207_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10341 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_2_2 ), 
            .I2(\REG.mem_3_2 ), .I3(rd_addr_r[1]), .O(n12201));
    defparam rd_addr_r_0__bdd_4_lut_10341.LUT_INIT = 16'he4aa;
    SB_LUT4 n12777_bdd_4_lut (.I0(n12777), .I1(n11842), .I2(n11841), .I3(rd_addr_r[2]), 
            .O(n12780));
    defparam n12777_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11352 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_22_3 ), 
            .I2(\REG.mem_23_3 ), .I3(rd_addr_r[1]), .O(n13413));
    defparam rd_addr_r_0__bdd_4_lut_11352.LUT_INIT = 16'he4aa;
    SB_LUT4 i3569_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_2_4 ), .O(n4952));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3569_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13413_bdd_4_lut (.I0(n13413), .I1(\REG.mem_21_3 ), .I2(\REG.mem_20_3 ), 
            .I3(rd_addr_r[1]), .O(n10916));
    defparam n13413_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10817 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_2_0 ), 
            .I2(\REG.mem_3_0 ), .I3(rd_addr_r[1]), .O(n12771));
    defparam rd_addr_r_0__bdd_4_lut_10817.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11437 (.I0(rd_addr_r[1]), .I1(n11283), 
            .I2(n11284), .I3(rd_addr_r[2]), .O(n13407));
    defparam rd_addr_r_1__bdd_4_lut_11437.LUT_INIT = 16'he4aa;
    SB_DFF i1601_1602 (.Q(\REG.mem_16_9 ), .C(FIFO_CLK_c), .D(n5183));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1598_1599 (.Q(\REG.mem_16_8 ), .C(FIFO_CLK_c), .D(n5182));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1595_1596 (.Q(\REG.mem_16_7 ), .C(FIFO_CLK_c), .D(n5181));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1592_1593 (.Q(\REG.mem_16_6 ), .C(FIFO_CLK_c), .D(n5180));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1589_1590 (.Q(\REG.mem_16_5 ), .C(FIFO_CLK_c), .D(n5179));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1586_1587 (.Q(\REG.mem_16_4 ), .C(FIFO_CLK_c), .D(n5178));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1583_1584 (.Q(\REG.mem_16_3 ), .C(FIFO_CLK_c), .D(n5177));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12771_bdd_4_lut (.I0(n12771), .I1(\REG.mem_1_0 ), .I2(\REG.mem_0_0 ), 
            .I3(rd_addr_r[1]), .O(n12774));
    defparam n12771_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9904_3_lut (.I0(\REG.mem_32_2 ), .I1(\REG.mem_33_2 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11754));
    defparam i9904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13407_bdd_4_lut (.I0(n13407), .I1(n11272), .I2(n11271), .I3(rd_addr_r[2]), 
            .O(n11365));
    defparam n13407_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9905_3_lut (.I0(\REG.mem_34_2 ), .I1(\REG.mem_35_2 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11755));
    defparam i9905_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1580_1581 (.Q(\REG.mem_16_2 ), .C(FIFO_CLK_c), .D(n5176));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9908_3_lut (.I0(\REG.mem_38_2 ), .I1(\REG.mem_39_2 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11758));
    defparam i9908_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i137_138 (.Q(\REG.mem_1_1 ), .C(FIFO_CLK_c), .D(n4879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9907_3_lut (.I0(\REG.mem_36_2 ), .I1(\REG.mem_37_2 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11757));
    defparam i9907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3568_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_2_3 ), .O(n4951));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3568_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11347 (.I0(rd_addr_r[2]), .I1(n11291), 
            .I2(n11333), .I3(rd_addr_r[3]), .O(n13401));
    defparam rd_addr_r_2__bdd_4_lut_11347.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10807 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_6_0 ), 
            .I2(\REG.mem_7_0 ), .I3(rd_addr_r[1]), .O(n12765));
    defparam rd_addr_r_0__bdd_4_lut_10807.LUT_INIT = 16'he4aa;
    SB_LUT4 n13401_bdd_4_lut (.I0(n13401), .I1(n12126), .I2(n12984), .I3(rd_addr_r[3]), 
            .O(n11840));
    defparam n13401_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1577_1578 (.Q(\REG.mem_16_1 ), .C(FIFO_CLK_c), .D(n5175));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1574_1575 (.Q(\REG.mem_16_0 ), .C(FIFO_CLK_c), .D(n5174));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1523_1524 (.Q(\REG.mem_15_15 ), .C(FIFO_CLK_c), .D(n5171));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1520_1521 (.Q(\REG.mem_15_14 ), .C(FIFO_CLK_c), .D(n5170));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1517_1518 (.Q(\REG.mem_15_13 ), .C(FIFO_CLK_c), .D(n5169));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1514_1515 (.Q(\REG.mem_15_12 ), .C(FIFO_CLK_c), .D(n5168));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1511_1512 (.Q(\REG.mem_15_11 ), .C(FIFO_CLK_c), .D(n5167));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11357 (.I0(rd_addr_r[3]), .I1(n11736), 
            .I2(n11737), .I3(rd_addr_r[4]), .O(n13395));
    defparam rd_addr_r_3__bdd_4_lut_11357.LUT_INIT = 16'he4aa;
    SB_LUT4 n13395_bdd_4_lut (.I0(n13395), .I1(n11725), .I2(n11724), .I3(rd_addr_r[4]), 
            .O(n13398));
    defparam n13395_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1508_1509 (.Q(\REG.mem_15_10 ), .C(FIFO_CLK_c), .D(n5166));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1505_1506 (.Q(\REG.mem_15_9 ), .C(FIFO_CLK_c), .D(n5165));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1502_1503 (.Q(\REG.mem_15_8 ), .C(FIFO_CLK_c), .D(n5164));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1499_1500 (.Q(\REG.mem_15_7 ), .C(FIFO_CLK_c), .D(n5163));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1496_1497 (.Q(\REG.mem_15_6 ), .C(FIFO_CLK_c), .D(n5162));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12765_bdd_4_lut (.I0(n12765), .I1(\REG.mem_5_0 ), .I2(\REG.mem_4_0 ), 
            .I3(rd_addr_r[1]), .O(n12768));
    defparam n12765_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1493_1494 (.Q(\REG.mem_15_5 ), .C(FIFO_CLK_c), .D(n5161));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9461_3_lut (.I0(n13206), .I1(n12462), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11311));
    defparam i9461_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1490_1491 (.Q(\REG.mem_15_4 ), .C(FIFO_CLK_c), .D(n5160));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1487_1488 (.Q(\REG.mem_15_3 ), .C(FIFO_CLK_c), .D(n5159));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1484_1485 (.Q(\REG.mem_15_2 ), .C(FIFO_CLK_c), .D(n5158));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1481_1482 (.Q(\REG.mem_15_1 ), .C(FIFO_CLK_c), .D(n5157));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1478_1479 (.Q(\REG.mem_15_0 ), .C(FIFO_CLK_c), .D(n5156));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1427_1428 (.Q(\REG.mem_14_15 ), .C(FIFO_CLK_c), .D(n5155));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1424_1425 (.Q(\REG.mem_14_14 ), .C(FIFO_CLK_c), .D(n5154));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1421_1422 (.Q(\REG.mem_14_13 ), .C(FIFO_CLK_c), .D(n5153));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1418_1419 (.Q(\REG.mem_14_12 ), .C(FIFO_CLK_c), .D(n5152));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1415_1416 (.Q(\REG.mem_14_11 ), .C(FIFO_CLK_c), .D(n5151));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1412_1413 (.Q(\REG.mem_14_10 ), .C(FIFO_CLK_c), .D(n5150));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1409_1410 (.Q(\REG.mem_14_9 ), .C(FIFO_CLK_c), .D(n5149));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1406_1407 (.Q(\REG.mem_14_8 ), .C(FIFO_CLK_c), .D(n5148));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1403_1404 (.Q(\REG.mem_14_7 ), .C(FIFO_CLK_c), .D(n5147));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1400_1401 (.Q(\REG.mem_14_6 ), .C(FIFO_CLK_c), .D(n5146));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1397_1398 (.Q(\REG.mem_14_5 ), .C(FIFO_CLK_c), .D(n5145));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1394_1395 (.Q(\REG.mem_14_4 ), .C(FIFO_CLK_c), .D(n5144));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1391_1392 (.Q(\REG.mem_14_3 ), .C(FIFO_CLK_c), .D(n5143));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1388_1389 (.Q(\REG.mem_14_2 ), .C(FIFO_CLK_c), .D(n5142));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1385_1386 (.Q(\REG.mem_14_1 ), .C(FIFO_CLK_c), .D(n5141));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1382_1383 (.Q(\REG.mem_14_0 ), .C(FIFO_CLK_c), .D(n5140));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1331_1332 (.Q(\REG.mem_13_15 ), .C(FIFO_CLK_c), .D(n5139));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1328_1329 (.Q(\REG.mem_13_14 ), .C(FIFO_CLK_c), .D(n5138));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1325_1326 (.Q(\REG.mem_13_13 ), .C(FIFO_CLK_c), .D(n5137));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1322_1323 (.Q(\REG.mem_13_12 ), .C(FIFO_CLK_c), .D(n5136));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1319_1320 (.Q(\REG.mem_13_11 ), .C(FIFO_CLK_c), .D(n5135));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1316_1317 (.Q(\REG.mem_13_10 ), .C(FIFO_CLK_c), .D(n5134));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1313_1314 (.Q(\REG.mem_13_9 ), .C(FIFO_CLK_c), .D(n5133));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1310_1311 (.Q(\REG.mem_13_8 ), .C(FIFO_CLK_c), .D(n5132));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9940_3_lut (.I0(\REG.mem_48_2 ), .I1(\REG.mem_49_2 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11790));
    defparam i9940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9941_3_lut (.I0(\REG.mem_50_2 ), .I1(\REG.mem_51_2 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11791));
    defparam i9941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11342 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_34_1 ), 
            .I2(\REG.mem_35_1 ), .I3(rd_addr_r[1]), .O(n13389));
    defparam rd_addr_r_0__bdd_4_lut_11342.LUT_INIT = 16'he4aa;
    SB_LUT4 n13389_bdd_4_lut (.I0(n13389), .I1(\REG.mem_33_1 ), .I2(\REG.mem_32_1 ), 
            .I3(rd_addr_r[1]), .O(n13392));
    defparam n13389_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1307_1308 (.Q(\REG.mem_13_7 ), .C(FIFO_CLK_c), .D(n5131));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10872 (.I0(rd_addr_r[2]), .I1(n12576), 
            .I2(n12492), .I3(rd_addr_r[3]), .O(n12759));
    defparam rd_addr_r_2__bdd_4_lut_10872.LUT_INIT = 16'he4aa;
    SB_LUT4 n12759_bdd_4_lut (.I0(n12759), .I1(n12588), .I2(n12654), .I3(rd_addr_r[3]), 
            .O(n12762));
    defparam n12759_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i106_2_lut_3_lut_4_lut (.I0(n18_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n47));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i106_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11327 (.I0(rd_addr_r[3]), .I1(n12906), 
            .I2(n11365), .I3(rd_addr_r[4]), .O(n13383));
    defparam rd_addr_r_3__bdd_4_lut_11327.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i105_2_lut_3_lut_4_lut (.I0(n18_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n15));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i105_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i4579_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_60_15 ), .O(n5962));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4579_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13383_bdd_4_lut (.I0(n13383), .I1(n11344), .I2(n11343), .I3(rd_addr_r[4]), 
            .O(n13386));
    defparam n13383_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4578_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_60_14 ), .O(n5961));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4578_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i100_2_lut_3_lut (.I0(n35_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n50));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i100_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i4577_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_60_13 ), .O(n5960));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4577_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1304_1305 (.Q(\REG.mem_13_6 ), .C(FIFO_CLK_c), .D(n5130));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4576_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_60_12 ), .O(n5959));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4576_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4575_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_60_11 ), .O(n5958));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4575_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i99_2_lut_3_lut (.I0(n35_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n18));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i99_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10877 (.I0(rd_addr_r[3]), .I1(n12738), 
            .I2(n11107), .I3(rd_addr_r[4]), .O(n12753));
    defparam rd_addr_r_3__bdd_4_lut_10877.LUT_INIT = 16'he4aa;
    SB_DFF i1301_1302 (.Q(\REG.mem_13_5 ), .C(FIFO_CLK_c), .D(n5129));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1298_1299 (.Q(\REG.mem_13_4 ), .C(FIFO_CLK_c), .D(n5128));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1295_1296 (.Q(\REG.mem_13_3 ), .C(FIFO_CLK_c), .D(n5127));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11322 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_22_6 ), 
            .I2(\REG.mem_23_6 ), .I3(rd_addr_r[1]), .O(n13377));
    defparam rd_addr_r_0__bdd_4_lut_11322.LUT_INIT = 16'he4aa;
    SB_DFF i1292_1293 (.Q(\REG.mem_13_2 ), .C(FIFO_CLK_c), .D(n5126));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4574_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_60_10 ), .O(n5957));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4574_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13377_bdd_4_lut (.I0(n13377), .I1(\REG.mem_21_6 ), .I2(\REG.mem_20_6 ), 
            .I3(rd_addr_r[1]), .O(n11048));
    defparam n13377_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4573_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_60_9 ), .O(n5956));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4573_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1289_1290 (.Q(\REG.mem_13_1 ), .C(FIFO_CLK_c), .D(n5125));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12753_bdd_4_lut (.I0(n12753), .I1(n11101), .I2(n11100), .I3(rd_addr_r[4]), 
            .O(n12756));
    defparam n12753_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4572_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_60_8 ), .O(n5955));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4572_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1286_1287 (.Q(\REG.mem_13_0 ), .C(FIFO_CLK_c), .D(n5124));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1235_1236 (.Q(\REG.mem_12_15 ), .C(FIFO_CLK_c), .D(n5123));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1232_1233 (.Q(\REG.mem_12_14 ), .C(FIFO_CLK_c), .D(n5122));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10812 (.I0(rd_addr_r[1]), .I1(n11085), 
            .I2(n11086), .I3(rd_addr_r[2]), .O(n12747));
    defparam rd_addr_r_1__bdd_4_lut_10812.LUT_INIT = 16'he4aa;
    SB_LUT4 i4571_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_60_7 ), .O(n5954));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4571_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11312 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_50_6 ), 
            .I2(\REG.mem_51_6 ), .I3(rd_addr_r[1]), .O(n13371));
    defparam rd_addr_r_0__bdd_4_lut_11312.LUT_INIT = 16'he4aa;
    SB_LUT4 n12747_bdd_4_lut (.I0(n12747), .I1(n11077), .I2(n11076), .I3(rd_addr_r[2]), 
            .O(n12750));
    defparam n12747_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13371_bdd_4_lut (.I0(n13371), .I1(\REG.mem_49_6 ), .I2(\REG.mem_48_6 ), 
            .I3(rd_addr_r[1]), .O(n11381));
    defparam n13371_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1229_1230 (.Q(\REG.mem_12_13 ), .C(FIFO_CLK_c), .D(n5121));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1226_1227 (.Q(\REG.mem_12_12 ), .C(FIFO_CLK_c), .D(n5120));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4570_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_60_6 ), .O(n5953));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4570_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1223_1224 (.Q(\REG.mem_12_11 ), .C(FIFO_CLK_c), .D(n5119));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1220_1221 (.Q(\REG.mem_12_10 ), .C(FIFO_CLK_c), .D(n5118));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4569_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_60_5 ), .O(n5952));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4569_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12201_bdd_4_lut (.I0(n12201), .I1(\REG.mem_1_2 ), .I2(\REG.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(n12204));
    defparam n12201_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10787 (.I0(rd_addr_r[1]), .I1(n11064), 
            .I2(n11065), .I3(rd_addr_r[2]), .O(n12741));
    defparam rd_addr_r_1__bdd_4_lut_10787.LUT_INIT = 16'he4aa;
    SB_DFF i1217_1218 (.Q(\REG.mem_12_9 ), .C(FIFO_CLK_c), .D(n5117));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9947_3_lut (.I0(\REG.mem_54_2 ), .I1(\REG.mem_55_2 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11797));
    defparam i9947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12741_bdd_4_lut (.I0(n12741), .I1(n11059), .I2(n11058), .I3(rd_addr_r[2]), 
            .O(n12744));
    defparam n12741_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1214_1215 (.Q(\REG.mem_12_8 ), .C(FIFO_CLK_c), .D(n5116));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11332 (.I0(rd_addr_r[2]), .I1(n13002), 
            .I2(n12480), .I3(rd_addr_r[3]), .O(n13365));
    defparam rd_addr_r_2__bdd_4_lut_11332.LUT_INIT = 16'he4aa;
    SB_LUT4 n13365_bdd_4_lut (.I0(n13365), .I1(n13128), .I2(n11351), .I3(rd_addr_r[3]), 
            .O(n11846));
    defparam n13365_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4568_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_60_4 ), .O(n5951));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4568_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4567_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_60_3 ), .O(n5950));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4567_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9946_3_lut (.I0(\REG.mem_52_2 ), .I1(\REG.mem_53_2 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11796));
    defparam i9946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9473_3_lut (.I0(n13158), .I1(n12990), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11323));
    defparam i9473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9847_3_lut (.I0(\REG.mem_0_14 ), .I1(\REG.mem_1_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11697));
    defparam i9847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11307 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_2_12 ), 
            .I2(\REG.mem_3_12 ), .I3(rd_addr_r[1]), .O(n13359));
    defparam rd_addr_r_0__bdd_4_lut_11307.LUT_INIT = 16'he4aa;
    SB_LUT4 i9848_3_lut (.I0(\REG.mem_2_14 ), .I1(\REG.mem_3_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11698));
    defparam i9848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9472_3_lut (.I0(n12138), .I1(n13344), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11322));
    defparam i9472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4566_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_60_2 ), .O(n5949));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4566_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4565_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_60_1 ), .O(n5948));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4565_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13359_bdd_4_lut (.I0(n13359), .I1(\REG.mem_1_12 ), .I2(\REG.mem_0_12 ), 
            .I3(rd_addr_r[1]), .O(n13362));
    defparam n13359_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10336 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_42_5 ), 
            .I2(\REG.mem_43_5 ), .I3(rd_addr_r[1]), .O(n12195));
    defparam rd_addr_r_0__bdd_4_lut_10336.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10782 (.I0(rd_addr_r[1]), .I1(n11040), 
            .I2(n11041), .I3(rd_addr_r[2]), .O(n12735));
    defparam rd_addr_r_1__bdd_4_lut_10782.LUT_INIT = 16'he4aa;
    SB_LUT4 i4564_3_lut_4_lut (.I0(n61_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_60_0 ), .O(n5947));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4564_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1211_1212 (.Q(\REG.mem_12_7 ), .C(FIFO_CLK_c), .D(n5115));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1208_1209 (.Q(\REG.mem_12_6 ), .C(FIFO_CLK_c), .D(n5114));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1205_1206 (.Q(\REG.mem_12_5 ), .C(FIFO_CLK_c), .D(n5113));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i61_2_lut_3_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n61_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i61_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n12735_bdd_4_lut (.I0(n12735), .I1(n11029), .I2(n11028), .I3(rd_addr_r[2]), 
            .O(n12738));
    defparam n12735_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4082_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_33_8 ), .O(n5465));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4082_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12195_bdd_4_lut (.I0(n12195), .I1(\REG.mem_41_5 ), .I2(\REG.mem_40_5 ), 
            .I3(rd_addr_r[1]), .O(n12198));
    defparam n12195_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1202_1203 (.Q(\REG.mem_12_4 ), .C(FIFO_CLK_c), .D(n5112));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_4__bdd_4_lut (.I0(rd_addr_r[4]), .I1(n12300), .I2(n11834), 
            .I3(rd_addr_r[5]), .O(n13353));
    defparam rd_addr_r_4__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i94_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n53));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i94_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i4081_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_33_7 ), .O(n5464));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4081_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i93_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n21));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i93_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10802 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_0 ), 
            .I2(\REG.mem_11_0 ), .I3(rd_addr_r[1]), .O(n12729));
    defparam rd_addr_r_0__bdd_4_lut_10802.LUT_INIT = 16'he4aa;
    SB_LUT4 n13353_bdd_4_lut (.I0(n13353), .I1(n12762), .I2(n13188), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_559 [0]));
    defparam n13353_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i13_2_lut_3_lut_4_lut (.I0(wr_sig_mv_w), .I1(wr_addr_r[0]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[1]), .O(n13));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i13_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 n12729_bdd_4_lut (.I0(n12729), .I1(\REG.mem_9_0 ), .I2(\REG.mem_8_0 ), 
            .I3(rd_addr_r[1]), .O(n12732));
    defparam n12729_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1199_1200 (.Q(\REG.mem_12_3 ), .C(FIFO_CLK_c), .D(n5111));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i14_2_lut_3_lut_4_lut (.I0(wr_sig_mv_w), .I1(wr_addr_r[0]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[1]), .O(n14));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i14_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i4554_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_59_15 ), .O(n5937));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4554_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4553_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_59_14 ), .O(n5936));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4553_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4552_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_59_13 ), .O(n5935));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4552_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4551_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_59_12 ), .O(n5934));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4551_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4550_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_59_11 ), .O(n5933));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4550_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1196_1197 (.Q(\REG.mem_12_2 ), .C(FIFO_CLK_c), .D(n5110));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1193_1194 (.Q(\REG.mem_12_1 ), .C(FIFO_CLK_c), .D(n5109));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10792 (.I0(rd_addr_r[3]), .I1(n12636), 
            .I2(n10921), .I3(rd_addr_r[4]), .O(n12723));
    defparam rd_addr_r_3__bdd_4_lut_10792.LUT_INIT = 16'he4aa;
    SB_LUT4 i4549_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_59_10 ), .O(n5932));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4549_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4548_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_59_9 ), .O(n5931));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4548_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4547_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_59_8 ), .O(n5930));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4547_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12723_bdd_4_lut (.I0(n12723), .I1(n10876), .I2(n12546), .I3(rd_addr_r[4]), 
            .O(n12726));
    defparam n12723_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1190_1191 (.Q(\REG.mem_12_0 ), .C(FIFO_CLK_c), .D(n5108));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4546_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_59_7 ), .O(n5929));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4546_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10772 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_42_9 ), 
            .I2(\REG.mem_43_9 ), .I3(rd_addr_r[1]), .O(n12717));
    defparam rd_addr_r_0__bdd_4_lut_10772.LUT_INIT = 16'he4aa;
    SB_LUT4 i4545_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_59_6 ), .O(n5928));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4545_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10331 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_30_6 ), 
            .I2(\REG.mem_31_6 ), .I3(rd_addr_r[1]), .O(n12189));
    defparam rd_addr_r_0__bdd_4_lut_10331.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i98_2_lut_3_lut (.I0(n33), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n51));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i98_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 n12717_bdd_4_lut (.I0(n12717), .I1(\REG.mem_41_9 ), .I2(\REG.mem_40_9 ), 
            .I3(rd_addr_r[1]), .O(n12720));
    defparam n12717_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4544_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_59_5 ), .O(n5927));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4544_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4080_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_33_6 ), .O(n5463));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4080_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i97_2_lut_3_lut (.I0(n33), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n19));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i97_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i4543_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_59_4 ), .O(n5926));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4543_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4542_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_59_3 ), .O(n5925));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4542_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4541_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_59_2 ), .O(n5924));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4541_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1139_1140 (.Q(\REG.mem_11_15 ), .C(FIFO_CLK_c), .D(n5107));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4540_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_59_1 ), .O(n5923));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4540_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11297 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_26_3 ), 
            .I2(\REG.mem_27_3 ), .I3(rd_addr_r[1]), .O(n13347));
    defparam rd_addr_r_0__bdd_4_lut_11297.LUT_INIT = 16'he4aa;
    SB_LUT4 i4539_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_59_0 ), .O(n5922));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4539_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13347_bdd_4_lut (.I0(n13347), .I1(\REG.mem_25_3 ), .I2(\REG.mem_24_3 ), 
            .I3(rd_addr_r[1]), .O(n10919));
    defparam n13347_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i92_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n54));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i92_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i91_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n22));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i91_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i4079_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_33_5 ), .O(n5462));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4079_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10762 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_15 ), 
            .I2(\REG.mem_15_15 ), .I3(rd_addr_r[1]), .O(n12711));
    defparam rd_addr_r_0__bdd_4_lut_10762.LUT_INIT = 16'he4aa;
    SB_DFF i1136_1137 (.Q(\REG.mem_11_14 ), .C(FIFO_CLK_c), .D(n5106));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12189_bdd_4_lut (.I0(n12189), .I1(\REG.mem_29_6 ), .I2(\REG.mem_28_6 ), 
            .I3(rd_addr_r[1]), .O(n12192));
    defparam n12189_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12711_bdd_4_lut (.I0(n12711), .I1(\REG.mem_13_15 ), .I2(\REG.mem_12_15 ), 
            .I3(rd_addr_r[1]), .O(n12714));
    defparam n12711_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11287 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_22_5 ), 
            .I2(\REG.mem_23_5 ), .I3(rd_addr_r[1]), .O(n13341));
    defparam rd_addr_r_0__bdd_4_lut_11287.LUT_INIT = 16'he4aa;
    SB_DFF i1133_1134 (.Q(\REG.mem_11_13 ), .C(FIFO_CLK_c), .D(n5105));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1130_1131 (.Q(\REG.mem_11_12 ), .C(FIFO_CLK_c), .D(n5104));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1127_1128 (.Q(\REG.mem_11_11 ), .C(FIFO_CLK_c), .D(n5103));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1124_1125 (.Q(\REG.mem_11_10 ), .C(FIFO_CLK_c), .D(n5102));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1121_1122 (.Q(\REG.mem_11_9 ), .C(FIFO_CLK_c), .D(n5101));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1118_1119 (.Q(\REG.mem_11_8 ), .C(FIFO_CLK_c), .D(n5100));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1115_1116 (.Q(\REG.mem_11_7 ), .C(FIFO_CLK_c), .D(n5099));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1112_1113 (.Q(\REG.mem_11_6 ), .C(FIFO_CLK_c), .D(n5098));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i140_141 (.Q(\REG.mem_1_2 ), .C(FIFO_CLK_c), .D(n4868));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i176_177 (.Q(\REG.mem_1_14 ), .C(FIFO_CLK_c), .D(n4867));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(FIFO_CLK_c), .D(n4866));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i143_144 (.Q(\REG.mem_1_3 ), .C(FIFO_CLK_c), .D(n4861));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3564_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_0_0 ), .O(n4947));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3564_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1109_1110 (.Q(\REG.mem_11_5 ), .C(FIFO_CLK_c), .D(n5097));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3541_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_0_15 ), .O(n4924));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3541_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3542_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_0_14 ), .O(n4925));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3542_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13341_bdd_4_lut (.I0(n13341), .I1(\REG.mem_21_5 ), .I2(\REG.mem_20_5 ), 
            .I3(rd_addr_r[1]), .O(n13344));
    defparam n13341_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3543_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_0_13 ), .O(n4926));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3543_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_6__I_0_i6_3_lut (.I0(rd_addr_r[5]), .I1(rd_addr_p1_w[5]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_498[5] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1106_1107 (.Q(\REG.mem_11_4 ), .C(FIFO_CLK_c), .D(n5096));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1103_1104 (.Q(\REG.mem_11_3 ), .C(FIFO_CLK_c), .D(n5095));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1100_1101 (.Q(\REG.mem_11_2 ), .C(FIFO_CLK_c), .D(n5094));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1097_1098 (.Q(\REG.mem_11_1 ), .C(FIFO_CLK_c), .D(n5093));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1094_1095 (.Q(\REG.mem_11_0 ), .C(FIFO_CLK_c), .D(n5092));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1043_1044 (.Q(\REG.mem_10_15 ), .C(FIFO_CLK_c), .D(n5091));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1040_1041 (.Q(\REG.mem_10_14 ), .C(FIFO_CLK_c), .D(n5090));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1037_1038 (.Q(\REG.mem_10_13 ), .C(FIFO_CLK_c), .D(n5089));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11282 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_54_6 ), 
            .I2(\REG.mem_55_6 ), .I3(rd_addr_r[1]), .O(n13335));
    defparam rd_addr_r_0__bdd_4_lut_11282.LUT_INIT = 16'he4aa;
    SB_DFF i1034_1035 (.Q(\REG.mem_10_12 ), .C(FIFO_CLK_c), .D(n5088));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10757 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_34_12 ), 
            .I2(\REG.mem_35_12 ), .I3(rd_addr_r[1]), .O(n12705));
    defparam rd_addr_r_0__bdd_4_lut_10757.LUT_INIT = 16'he4aa;
    SB_LUT4 i3544_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_0_12 ), .O(n4927));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3544_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12705_bdd_4_lut (.I0(n12705), .I1(\REG.mem_33_12 ), .I2(\REG.mem_32_12 ), 
            .I3(rd_addr_r[1]), .O(n12708));
    defparam n12705_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3545_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_0_11 ), .O(n4928));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3545_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13335_bdd_4_lut (.I0(n13335), .I1(\REG.mem_53_6 ), .I2(\REG.mem_52_6 ), 
            .I3(rd_addr_r[1]), .O(n11396));
    defparam n13335_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3546_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_0_10 ), .O(n4929));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3546_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1031_1032 (.Q(\REG.mem_10_11 ), .C(FIFO_CLK_c), .D(n5087));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1028_1029 (.Q(\REG.mem_10_10 ), .C(FIFO_CLK_c), .D(n5086));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1025_1026 (.Q(\REG.mem_10_9 ), .C(FIFO_CLK_c), .D(n5085));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1022_1023 (.Q(\REG.mem_10_8 ), .C(FIFO_CLK_c), .D(n5084));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1019_1020 (.Q(\REG.mem_10_7 ), .C(FIFO_CLK_c), .D(n5083));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1016_1017 (.Q(\REG.mem_10_6 ), .C(FIFO_CLK_c), .D(n5082));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1013_1014 (.Q(\REG.mem_10_5 ), .C(FIFO_CLK_c), .D(n5081));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1010_1011 (.Q(\REG.mem_10_4 ), .C(FIFO_CLK_c), .D(n5080));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3547_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_0_9 ), .O(n4930));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3547_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_6__I_0_i4_3_lut (.I0(rd_addr_r[3]), .I1(rd_addr_p1_w[3]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_498[3] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1007_1008 (.Q(\REG.mem_10_3 ), .C(FIFO_CLK_c), .D(n5079));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3548_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_0_8 ), .O(n4931));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3548_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3549_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_0_7 ), .O(n4932));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3549_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3550_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_0_6 ), .O(n4933));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3550_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3551_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_0_5 ), .O(n4934));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3551_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3552_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_0_4 ), .O(n4935));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3552_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3560_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_0_3 ), .O(n4943));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3560_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3561_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_0_2 ), .O(n4944));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3561_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3563_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_0_1 ), .O(n4946));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3563_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11292 (.I0(rd_addr_r[4]), .I1(n11840), 
            .I2(n11846), .I3(rd_addr_r[5]), .O(n13329));
    defparam rd_addr_r_4__bdd_4_lut_11292.LUT_INIT = 16'he4aa;
    SB_LUT4 n13329_bdd_4_lut (.I0(n13329), .I1(n11762), .I2(n11690), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_559 [13]));
    defparam n13329_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_6__I_0_i3_3_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_498[2] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i38_2_lut_3_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n38));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i38_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i102_2_lut_3_lut_4_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n49));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i102_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 EnabledDecoder_2_i101_2_lut_3_lut_4_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n17));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i101_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i4_2_lut_4_lut (.I0(rd_addr_r[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_498[3] ), .O(rd_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i4_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11277 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_38_1 ), 
            .I2(\REG.mem_39_1 ), .I3(rd_addr_r[1]), .O(n13323));
    defparam rd_addr_r_0__bdd_4_lut_11277.LUT_INIT = 16'he4aa;
    SB_LUT4 n13323_bdd_4_lut (.I0(n13323), .I1(\REG.mem_37_1 ), .I2(\REG.mem_36_1 ), 
            .I3(rd_addr_r[1]), .O(n13326));
    defparam n13323_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10752 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_42_11 ), 
            .I2(\REG.mem_43_11 ), .I3(rd_addr_r[1]), .O(n12699));
    defparam rd_addr_r_0__bdd_4_lut_10752.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i5_2_lut_4_lut (.I0(rd_addr_r[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_498[5] ), .O(rd_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4532_2_lut_4_lut (.I0(rd_addr_r[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5915));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4532_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11267 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_50_14 ), 
            .I2(\REG.mem_51_14 ), .I3(rd_addr_r[1]), .O(n13317));
    defparam rd_addr_r_0__bdd_4_lut_11267.LUT_INIT = 16'he4aa;
    SB_LUT4 n13317_bdd_4_lut (.I0(n13317), .I1(\REG.mem_49_14 ), .I2(\REG.mem_48_14 ), 
            .I3(rd_addr_r[1]), .O(n11861));
    defparam n13317_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12699_bdd_4_lut (.I0(n12699), .I1(\REG.mem_41_11 ), .I2(\REG.mem_40_11 ), 
            .I3(rd_addr_r[1]), .O(n11543));
    defparam n12699_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i6_2_lut_4_lut (.I0(\rd_addr_r[6] ), 
            .I1(rd_addr_p1_w[6]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_498[5] ), 
            .O(rd_grey_w[5]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i6_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11337 (.I0(rd_addr_r[1]), .I1(n11286), 
            .I2(n11287), .I3(rd_addr_r[2]), .O(n13311));
    defparam rd_addr_r_1__bdd_4_lut_11337.LUT_INIT = 16'he4aa;
    SB_LUT4 n13311_bdd_4_lut (.I0(n13311), .I1(n11278), .I2(n11277), .I3(rd_addr_r[2]), 
            .O(n11401));
    defparam n13311_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4530_2_lut_4_lut (.I0(\rd_addr_r[6] ), .I1(rd_addr_p1_w[6]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5913));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4530_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i9851_3_lut (.I0(\REG.mem_6_14 ), .I1(\REG.mem_7_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11701));
    defparam i9851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9850_3_lut (.I0(\REG.mem_4_14 ), .I1(\REG.mem_5_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11700));
    defparam i9850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10747 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_54_3 ), 
            .I2(\REG.mem_55_3 ), .I3(rd_addr_r[1]), .O(n12693));
    defparam rd_addr_r_0__bdd_4_lut_10747.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i87_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n24));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i87_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i1004_1005 (.Q(\REG.mem_10_2 ), .C(FIFO_CLK_c), .D(n5078));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12693_bdd_4_lut (.I0(n12693), .I1(\REG.mem_53_3 ), .I2(\REG.mem_52_3 ), 
            .I3(rd_addr_r[1]), .O(n10970));
    defparam n12693_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4529_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_58_15 ), .O(n5912));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4529_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4528_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_58_14 ), .O(n5911));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4528_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4527_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_58_13 ), .O(n5910));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4527_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11262 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_2_6 ), 
            .I2(\REG.mem_3_6 ), .I3(rd_addr_r[1]), .O(n13305));
    defparam rd_addr_r_0__bdd_4_lut_11262.LUT_INIT = 16'he4aa;
    SB_LUT4 i4526_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_58_12 ), .O(n5909));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4526_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9010_3_lut (.I0(n12204), .I1(n12132), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10860));
    defparam i9010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4525_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_58_11 ), .O(n5908));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4525_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1001_1002 (.Q(\REG.mem_10_1 ), .C(FIFO_CLK_c), .D(n5077));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10302 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_58_9 ), 
            .I2(\REG.mem_59_9 ), .I3(rd_addr_r[1]), .O(n12147));
    defparam rd_addr_r_0__bdd_4_lut_10302.LUT_INIT = 16'he4aa;
    SB_LUT4 i4524_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_58_10 ), .O(n5907));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4524_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13305_bdd_4_lut (.I0(n13305), .I1(\REG.mem_1_6 ), .I2(\REG.mem_0_6 ), 
            .I3(rd_addr_r[1]), .O(n11864));
    defparam n13305_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4523_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_58_9 ), .O(n5906));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4523_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4522_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_58_8 ), .O(n5905));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4522_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4521_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_58_7 ), .O(n5904));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4521_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10777 (.I0(rd_addr_r[1]), .I1(n11835), 
            .I2(n11836), .I3(rd_addr_r[2]), .O(n12681));
    defparam rd_addr_r_1__bdd_4_lut_10777.LUT_INIT = 16'he4aa;
    SB_LUT4 i9011_3_lut (.I0(n12120), .I1(n13734), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10861));
    defparam i9011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4520_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_58_6 ), .O(n5903));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4520_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4519_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_58_5 ), .O(n5902));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4519_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4518_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_58_4 ), .O(n5901));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4518_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i998_999 (.Q(\REG.mem_10_0 ), .C(FIFO_CLK_c), .D(n5076));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9014_3_lut (.I0(n13686), .I1(n13680), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10864));
    defparam i9014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12681_bdd_4_lut (.I0(n12681), .I1(n11830), .I2(n11829), .I3(rd_addr_r[2]), 
            .O(n12684));
    defparam n12681_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4517_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_58_3 ), .O(n5900));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4517_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11257 (.I0(rd_addr_r[1]), .I1(n11268), 
            .I2(n11269), .I3(rd_addr_r[2]), .O(n13299));
    defparam rd_addr_r_1__bdd_4_lut_11257.LUT_INIT = 16'he4aa;
    SB_DFF i947_948 (.Q(\REG.mem_9_15 ), .C(FIFO_CLK_c), .D(n5075));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13299_bdd_4_lut (.I0(n13299), .I1(n11239), .I2(n11238), .I3(rd_addr_r[2]), 
            .O(n13302));
    defparam n13299_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10742 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_2_9 ), 
            .I2(\REG.mem_3_9 ), .I3(rd_addr_r[1]), .O(n12675));
    defparam rd_addr_r_0__bdd_4_lut_10742.LUT_INIT = 16'he4aa;
    SB_LUT4 i4516_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_58_2 ), .O(n5899));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4516_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4515_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_58_1 ), .O(n5898));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4515_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11247 (.I0(rd_addr_r[1]), .I1(n11763), 
            .I2(n11764), .I3(rd_addr_r[2]), .O(n13293));
    defparam rd_addr_r_1__bdd_4_lut_11247.LUT_INIT = 16'he4aa;
    SB_LUT4 n13293_bdd_4_lut (.I0(n13293), .I1(n11740), .I2(n11739), .I3(rd_addr_r[2]), 
            .O(n10921));
    defparam n13293_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4514_3_lut_4_lut (.I0(n57_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_58_0 ), .O(n5897));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4514_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12675_bdd_4_lut (.I0(n12675), .I1(\REG.mem_1_9 ), .I2(\REG.mem_0_9 ), 
            .I3(rd_addr_r[1]), .O(n12678));
    defparam n12675_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i944_945 (.Q(\REG.mem_9_14 ), .C(FIFO_CLK_c), .D(n5074));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4078_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_33_4 ), .O(n5461));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4078_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i941_942 (.Q(\REG.mem_9_13 ), .C(FIFO_CLK_c), .D(n5073));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i20_2_lut (.I0(n11_c), .I1(wr_addr_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n20_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i20_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 EnabledDecoder_2_i90_2_lut_3_lut_4_lut (.I0(n18_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n55));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i90_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i89_2_lut_3_lut_4_lut (.I0(n18_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n23));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i89_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 EnabledDecoder_2_i120_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n40));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i120_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10767 (.I0(rd_addr_r[3]), .I1(n11871), 
            .I2(n11872), .I3(rd_addr_r[4]), .O(n12669));
    defparam rd_addr_r_3__bdd_4_lut_10767.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i119_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n8));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i119_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n12669_bdd_4_lut (.I0(n12669), .I1(n11854), .I2(n11853), .I3(rd_addr_r[4]), 
            .O(n12672));
    defparam n12669_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i23_2_lut_3_lut (.I0(n12_adj_1199), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n23_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i23_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i938_939 (.Q(\REG.mem_9_12 ), .C(FIFO_CLK_c), .D(n5072));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i132_2_lut_3_lut (.I0(n35_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n34));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i132_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11252 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_54_14 ), 
            .I2(\REG.mem_55_14 ), .I3(rd_addr_r[1]), .O(n13287));
    defparam rd_addr_r_0__bdd_4_lut_11252.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i40_2_lut_3_lut_4_lut (.I0(n12_adj_1199), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n40_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i40_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_DFF i146_147 (.Q(\REG.mem_1_4 ), .C(FIFO_CLK_c), .D(n4837));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i39_2_lut_3_lut_4_lut (.I0(n12_adj_1199), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n39));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i39_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_DFF i935_936 (.Q(\REG.mem_9_11 ), .C(FIFO_CLK_c), .D(n5071));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10728 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_58_3 ), 
            .I2(\REG.mem_59_3 ), .I3(rd_addr_r[1]), .O(n12663));
    defparam rd_addr_r_0__bdd_4_lut_10728.LUT_INIT = 16'he4aa;
    SB_DFF i932_933 (.Q(\REG.mem_9_10 ), .C(FIFO_CLK_c), .D(n5070));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13287_bdd_4_lut (.I0(n13287), .I1(\REG.mem_53_14 ), .I2(\REG.mem_52_14 ), 
            .I3(rd_addr_r[1]), .O(n11867));
    defparam n13287_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12663_bdd_4_lut (.I0(n12663), .I1(\REG.mem_57_3 ), .I2(\REG.mem_56_3 ), 
            .I3(rd_addr_r[1]), .O(n10976));
    defparam n12663_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4495_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_56_15 ), .O(n5878));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4495_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4077_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_33_3 ), .O(n5460));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4077_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4494_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_56_14 ), .O(n5877));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4494_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i929_930 (.Q(\REG.mem_9_9 ), .C(FIFO_CLK_c), .D(n5069));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i131_2_lut_3_lut (.I0(n35_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n2));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i131_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11242 (.I0(rd_addr_r[1]), .I1(n11811), 
            .I2(n11812), .I3(rd_addr_r[2]), .O(n13281));
    defparam rd_addr_r_1__bdd_4_lut_11242.LUT_INIT = 16'he4aa;
    SB_LUT4 i4493_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_56_13 ), .O(n5876));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4493_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4492_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_56_12 ), .O(n5875));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4492_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i149_150 (.Q(\REG.mem_1_5 ), .C(FIFO_CLK_c), .D(n4835));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i926_927 (.Q(\REG.mem_9_8 ), .C(FIFO_CLK_c), .D(n5068));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i923_924 (.Q(\REG.mem_9_7 ), .C(FIFO_CLK_c), .D(n5067));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4076_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_33_2 ), .O(n5459));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4076_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4491_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_56_11 ), .O(n5874));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4491_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4490_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_56_10 ), .O(n5873));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4490_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i36_2_lut_3_lut (.I0(n11_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n36));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i36_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i4489_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_56_9 ), .O(n5872));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4489_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10718 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_0 ), 
            .I2(\REG.mem_15_0 ), .I3(rd_addr_r[1]), .O(n12657));
    defparam rd_addr_r_0__bdd_4_lut_10718.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i35_2_lut_3_lut (.I0(n11_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n35_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i35_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF i920_921 (.Q(\REG.mem_9_6 ), .C(FIFO_CLK_c), .D(n5066));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i917_918 (.Q(\REG.mem_9_5 ), .C(FIFO_CLK_c), .D(n5065));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12657_bdd_4_lut (.I0(n12657), .I1(\REG.mem_13_0 ), .I2(\REG.mem_12_0 ), 
            .I3(rd_addr_r[1]), .O(n12660));
    defparam n12657_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13281_bdd_4_lut (.I0(n13281), .I1(n11794), .I2(n11793), .I3(rd_addr_r[2]), 
            .O(n13284));
    defparam n13281_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12141_bdd_4_lut (.I0(n12141), .I1(\REG.mem_41_15 ), .I2(\REG.mem_40_15 ), 
            .I3(rd_addr_r[1]), .O(n12144));
    defparam n12141_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9535_3_lut (.I0(\REG.mem_56_10 ), .I1(\REG.mem_57_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11385));
    defparam i9535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4488_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_56_8 ), .O(n5871));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4488_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i914_915 (.Q(\REG.mem_9_4 ), .C(FIFO_CLK_c), .D(n5064));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4487_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_56_7 ), .O(n5870));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4487_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11237 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_30_3 ), 
            .I2(\REG.mem_31_3 ), .I3(rd_addr_r[1]), .O(n13275));
    defparam rd_addr_r_0__bdd_4_lut_11237.LUT_INIT = 16'he4aa;
    SB_LUT4 i4486_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_56_6 ), .O(n5869));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4486_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9536_3_lut (.I0(\REG.mem_58_10 ), .I1(\REG.mem_59_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11386));
    defparam i9536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9539_3_lut (.I0(\REG.mem_62_10 ), .I1(\REG.mem_63_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11389));
    defparam i9539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9538_3_lut (.I0(\REG.mem_60_10 ), .I1(\REG.mem_61_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11388));
    defparam i9538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4485_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_56_5 ), .O(n5868));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4485_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i911_912 (.Q(\REG.mem_9_3 ), .C(FIFO_CLK_c), .D(n5063));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10713 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_18_0 ), 
            .I2(\REG.mem_19_0 ), .I3(rd_addr_r[1]), .O(n12651));
    defparam rd_addr_r_0__bdd_4_lut_10713.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_45 (.I0(DEBUG_3_c), .I1(get_next_word), .I2(GND_net), 
            .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i1_2_lut_adj_45.LUT_INIT = 16'h4444;
    SB_LUT4 i4484_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_56_4 ), .O(n5867));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4484_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13275_bdd_4_lut (.I0(n13275), .I1(\REG.mem_29_3 ), .I2(\REG.mem_28_3 ), 
            .I3(rd_addr_r[1]), .O(n10928));
    defparam n13275_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4483_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_56_3 ), .O(n5866));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4483_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i908_909 (.Q(\REG.mem_9_2 ), .C(FIFO_CLK_c), .D(n5062));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rp_sync2_r_6__I_0_136_i1_2_lut (.I0(rp_sync2_r[5]), .I1(rp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(rp_sync_w[5]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam rp_sync2_r_6__I_0_136_i1_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 n12651_bdd_4_lut (.I0(n12651), .I1(\REG.mem_17_0 ), .I2(\REG.mem_16_0 ), 
            .I3(rd_addr_r[1]), .O(n12654));
    defparam n12651_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_46 (.I0(rp_sync2_r[3]), .I1(rp_sync_w[4]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_adj_46.LUT_INIT = 16'h6666;
    SB_DFF i905_906 (.Q(\REG.mem_9_1 ), .C(FIFO_CLK_c), .D(n5061));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11227 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_34_3 ), 
            .I2(\REG.mem_35_3 ), .I3(rd_addr_r[1]), .O(n13269));
    defparam rd_addr_r_0__bdd_4_lut_11227.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i6_2_lut_4_lut (.I0(wr_grey_sync_r[6]), 
            .I1(wr_addr_p1_w[6]), .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[5] ), 
            .O(wr_grey_w[5]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i6_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4286_2_lut_4_lut (.I0(wr_grey_sync_r[6]), .I1(wr_addr_p1_w[6]), 
            .I2(wr_sig_mv_w), .I3(reset_per_frame), .O(n5669));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i4286_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i4482_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_56_2 ), .O(n5865));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4482_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13269_bdd_4_lut (.I0(n13269), .I1(\REG.mem_33_3 ), .I2(\REG.mem_32_3 ), 
            .I3(rd_addr_r[1]), .O(n10931));
    defparam n13269_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4481_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_56_1 ), .O(n5864));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4481_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9415_3_lut (.I0(\REG.mem_0_10 ), .I1(\REG.mem_1_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11265));
    defparam i9415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_47 (.I0(rp_sync2_r[1]), .I1(rp_sync_w[2]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_adj_47.LUT_INIT = 16'h6666;
    SB_DFF i902_903 (.Q(\REG.mem_9_0 ), .C(FIFO_CLK_c), .D(n5060));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i851_852 (.Q(\REG.mem_8_15 ), .C(FIFO_CLK_c), .D(n5059));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i848_849 (.Q(\REG.mem_8_14 ), .C(FIFO_CLK_c), .D(n5058));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i845_846 (.Q(\REG.mem_8_13 ), .C(FIFO_CLK_c), .D(n5057));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i842_843 (.Q(\REG.mem_8_12 ), .C(FIFO_CLK_c), .D(n5056));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i839_840 (.Q(\REG.mem_8_11 ), .C(FIFO_CLK_c), .D(n5055));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i836_837 (.Q(\REG.mem_8_10 ), .C(FIFO_CLK_c), .D(n5054));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i833_834 (.Q(\REG.mem_8_9 ), .C(FIFO_CLK_c), .D(n5053));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i830_831 (.Q(\REG.mem_8_8 ), .C(FIFO_CLK_c), .D(n5052));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i827_828 (.Q(\REG.mem_8_7 ), .C(FIFO_CLK_c), .D(n5051));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i824_825 (.Q(\REG.mem_8_6 ), .C(FIFO_CLK_c), .D(n5050));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i821_822 (.Q(\REG.mem_8_5 ), .C(FIFO_CLK_c), .D(n5049));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i818_819 (.Q(\REG.mem_8_4 ), .C(FIFO_CLK_c), .D(n5048));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i815_816 (.Q(\REG.mem_8_3 ), .C(FIFO_CLK_c), .D(n5047));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i812_813 (.Q(\REG.mem_8_2 ), .C(FIFO_CLK_c), .D(n5046));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i809_810 (.Q(\REG.mem_8_1 ), .C(FIFO_CLK_c), .D(n5045));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i806_807 (.Q(\REG.mem_8_0 ), .C(FIFO_CLK_c), .D(n5044));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i755_756 (.Q(\REG.mem_7_15 ), .C(FIFO_CLK_c), .D(n5043));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i752_753 (.Q(\REG.mem_7_14 ), .C(FIFO_CLK_c), .D(n5042));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i749_750 (.Q(\REG.mem_7_13 ), .C(FIFO_CLK_c), .D(n5041));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i746_747 (.Q(\REG.mem_7_12 ), .C(FIFO_CLK_c), .D(n5040));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i743_744 (.Q(\REG.mem_7_11 ), .C(FIFO_CLK_c), .D(n5039));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i740_741 (.Q(\REG.mem_7_10 ), .C(FIFO_CLK_c), .D(n5038));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i737_738 (.Q(\REG.mem_7_9 ), .C(FIFO_CLK_c), .D(n5037));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i734_735 (.Q(\REG.mem_7_8 ), .C(FIFO_CLK_c), .D(n5036));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i731_732 (.Q(\REG.mem_7_7 ), .C(FIFO_CLK_c), .D(n5035));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i728_729 (.Q(\REG.mem_7_6 ), .C(FIFO_CLK_c), .D(n5034));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i725_726 (.Q(\REG.mem_7_5 ), .C(FIFO_CLK_c), .D(n5033));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i722_723 (.Q(\REG.mem_7_4 ), .C(FIFO_CLK_c), .D(n5032));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i719_720 (.Q(\REG.mem_7_3 ), .C(FIFO_CLK_c), .D(n5031));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i716_717 (.Q(\REG.mem_7_2 ), .C(FIFO_CLK_c), .D(n5030));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i713_714 (.Q(\REG.mem_7_1 ), .C(FIFO_CLK_c), .D(n5029));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i710_711 (.Q(\REG.mem_7_0 ), .C(FIFO_CLK_c), .D(n5028));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i659_660 (.Q(\REG.mem_6_15 ), .C(FIFO_CLK_c), .D(n5027));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i656_657 (.Q(\REG.mem_6_14 ), .C(FIFO_CLK_c), .D(n5026));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i653_654 (.Q(\REG.mem_6_13 ), .C(FIFO_CLK_c), .D(n5025));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i650_651 (.Q(\REG.mem_6_12 ), .C(FIFO_CLK_c), .D(n5024));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i647_648 (.Q(\REG.mem_6_11 ), .C(FIFO_CLK_c), .D(n5023));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i644_645 (.Q(\REG.mem_6_10 ), .C(FIFO_CLK_c), .D(n5022));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i641_642 (.Q(\REG.mem_6_9 ), .C(FIFO_CLK_c), .D(n5021));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i638_639 (.Q(\REG.mem_6_8 ), .C(FIFO_CLK_c), .D(n5020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i635_636 (.Q(\REG.mem_6_7 ), .C(FIFO_CLK_c), .D(n5019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i632_633 (.Q(\REG.mem_6_6 ), .C(FIFO_CLK_c), .D(n5018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i629_630 (.Q(\REG.mem_6_5 ), .C(FIFO_CLK_c), .D(n5017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i626_627 (.Q(\REG.mem_6_4 ), .C(FIFO_CLK_c), .D(n5016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i623_624 (.Q(\REG.mem_6_3 ), .C(FIFO_CLK_c), .D(n5015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i620_621 (.Q(\REG.mem_6_2 ), .C(FIFO_CLK_c), .D(n5014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i617_618 (.Q(\REG.mem_6_1 ), .C(FIFO_CLK_c), .D(n5013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i614_615 (.Q(\REG.mem_6_0 ), .C(FIFO_CLK_c), .D(n5012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i563_564 (.Q(\REG.mem_5_15 ), .C(FIFO_CLK_c), .D(n5011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i560_561 (.Q(\REG.mem_5_14 ), .C(FIFO_CLK_c), .D(n5010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i557_558 (.Q(\REG.mem_5_13 ), .C(FIFO_CLK_c), .D(n5009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i554_555 (.Q(\REG.mem_5_12 ), .C(FIFO_CLK_c), .D(n5008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i551_552 (.Q(\REG.mem_5_11 ), .C(FIFO_CLK_c), .D(n5007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i548_549 (.Q(\REG.mem_5_10 ), .C(FIFO_CLK_c), .D(n5006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i545_546 (.Q(\REG.mem_5_9 ), .C(FIFO_CLK_c), .D(n5005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i542_543 (.Q(\REG.mem_5_8 ), .C(FIFO_CLK_c), .D(n5004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i539_540 (.Q(\REG.mem_5_7 ), .C(FIFO_CLK_c), .D(n5003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i536_537 (.Q(\REG.mem_5_6 ), .C(FIFO_CLK_c), .D(n5002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i533_534 (.Q(\REG.mem_5_5 ), .C(FIFO_CLK_c), .D(n5001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i530_531 (.Q(\REG.mem_5_4 ), .C(FIFO_CLK_c), .D(n5000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i527_528 (.Q(\REG.mem_5_3 ), .C(FIFO_CLK_c), .D(n4999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i524_525 (.Q(\REG.mem_5_2 ), .C(FIFO_CLK_c), .D(n4998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i521_522 (.Q(\REG.mem_5_1 ), .C(FIFO_CLK_c), .D(n4997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i518_519 (.Q(\REG.mem_5_0 ), .C(FIFO_CLK_c), .D(n4996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i467_468 (.Q(\REG.mem_4_15 ), .C(FIFO_CLK_c), .D(n4995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i464_465 (.Q(\REG.mem_4_14 ), .C(FIFO_CLK_c), .D(n4994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i461_462 (.Q(\REG.mem_4_13 ), .C(FIFO_CLK_c), .D(n4993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i458_459 (.Q(\REG.mem_4_12 ), .C(FIFO_CLK_c), .D(n4992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i455_456 (.Q(\REG.mem_4_11 ), .C(FIFO_CLK_c), .D(n4991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i452_453 (.Q(\REG.mem_4_10 ), .C(FIFO_CLK_c), .D(n4990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i449_450 (.Q(\REG.mem_4_9 ), .C(FIFO_CLK_c), .D(n4989));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i446_447 (.Q(\REG.mem_4_8 ), .C(FIFO_CLK_c), .D(n4988));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i443_444 (.Q(\REG.mem_4_7 ), .C(FIFO_CLK_c), .D(n4987));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i440_441 (.Q(\REG.mem_4_6 ), .C(FIFO_CLK_c), .D(n4986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i437_438 (.Q(\REG.mem_4_5 ), .C(FIFO_CLK_c), .D(n4985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i434_435 (.Q(\REG.mem_4_4 ), .C(FIFO_CLK_c), .D(n4984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i431_432 (.Q(\REG.mem_4_3 ), .C(FIFO_CLK_c), .D(n4983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i428_429 (.Q(\REG.mem_4_2 ), .C(FIFO_CLK_c), .D(n4982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i425_426 (.Q(\REG.mem_4_1 ), .C(FIFO_CLK_c), .D(n4981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i422_423 (.Q(\REG.mem_4_0 ), .C(FIFO_CLK_c), .D(n4980));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i371_372 (.Q(\REG.mem_3_15 ), .C(FIFO_CLK_c), .D(n4979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i368_369 (.Q(\REG.mem_3_14 ), .C(FIFO_CLK_c), .D(n4978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i365_366 (.Q(\REG.mem_3_13 ), .C(FIFO_CLK_c), .D(n4977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i362_363 (.Q(\REG.mem_3_12 ), .C(FIFO_CLK_c), .D(n4976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i359_360 (.Q(\REG.mem_3_11 ), .C(FIFO_CLK_c), .D(n4975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i356_357 (.Q(\REG.mem_3_10 ), .C(FIFO_CLK_c), .D(n4974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i353_354 (.Q(\REG.mem_3_9 ), .C(FIFO_CLK_c), .D(n4973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i350_351 (.Q(\REG.mem_3_8 ), .C(FIFO_CLK_c), .D(n4972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i347_348 (.Q(\REG.mem_3_7 ), .C(FIFO_CLK_c), .D(n4971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i344_345 (.Q(\REG.mem_3_6 ), .C(FIFO_CLK_c), .D(n4970));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i341_342 (.Q(\REG.mem_3_5 ), .C(FIFO_CLK_c), .D(n4969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4479_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_56_0 ), .O(n5862));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4479_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9416_3_lut (.I0(\REG.mem_2_10 ), .I1(\REG.mem_3_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11266));
    defparam i9416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_48 (.I0(rp_sync2_r[5]), .I1(rp_sync2_r[4]), .I2(rp_sync2_r[6]), 
            .I3(GND_net), .O(rp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i2_3_lut_adj_48.LUT_INIT = 16'h6969;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11222 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_6_12 ), 
            .I2(\REG.mem_7_12 ), .I3(rd_addr_r[1]), .O(n13263));
    defparam rd_addr_r_0__bdd_4_lut_11222.LUT_INIT = 16'he4aa;
    SB_LUT4 i4075_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_33_1 ), .O(n5458));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4075_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_p1_w_6__I_0_2_lut (.I0(wr_addr_p1_w[6]), .I1(rp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(full_max_w));   // src/fifo_dc_32_lut_gen.v(296[27:88])
    defparam wr_addr_p1_w_6__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8911_4_lut (.I0(wr_addr_p1_w[4]), .I1(wr_addr_p1_w[1]), .I2(rp_sync_w[4]), 
            .I3(rp_sync_w[1]), .O(n10760));
    defparam i8911_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i8875_4_lut (.I0(wr_addr_p1_w[5]), .I1(wr_addr_p1_w[3]), .I2(rp_sync_w[5]), 
            .I3(rp_sync_w[3]), .O(n10724));
    defparam i8875_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i5_4_lut_adj_49 (.I0(wr_addr_p1_w[0]), .I1(n10760), .I2(full_max_w), 
            .I3(rp_sync_w[0]), .O(n12_adj_1201));
    defparam i5_4_lut_adj_49.LUT_INIT = 16'h1020;
    SB_LUT4 i8897_4_lut (.I0(wr_addr_r[5]), .I1(wr_addr_r[1]), .I2(rp_sync_w[5]), 
            .I3(rp_sync_w[1]), .O(n10746));
    defparam i8897_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i8887_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_r[0]), .I2(rp_sync_w[2]), 
            .I3(rp_sync_w[0]), .O(n10736));
    defparam i8887_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i10135_4_lut (.I0(wr_addr_p1_w[2]), .I1(n12_adj_1201), .I2(n10724), 
            .I3(rp_sync_w[2]), .O(n11883));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam i10135_4_lut.LUT_INIT = 16'h0408;
    SB_LUT4 i8986_3_lut (.I0(n10744), .I1(n10736), .I2(n10746), .I3(GND_net), 
            .O(n10836));
    defparam i8986_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 full_nxt_c_I_6_4_lut (.I0(n10836), .I1(n11883), .I2(wr_sig_mv_w), 
            .I3(full_o), .O(full_nxt_c_N_626));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam full_nxt_c_I_6_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i1_2_lut_adj_50 (.I0(dc32_fifo_almost_full), .I1(DEBUG_1_c_c), 
            .I2(GND_net), .I3(GND_net), .O(FT_OE_N_420));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    defparam i1_2_lut_adj_50.LUT_INIT = 16'heeee;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10708 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_62_3 ), 
            .I2(\REG.mem_63_3 ), .I3(rd_addr_r[1]), .O(n12645));
    defparam rd_addr_r_0__bdd_4_lut_10708.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i53_2_lut_3_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n53_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i53_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n12645_bdd_4_lut (.I0(n12645), .I1(\REG.mem_61_3 ), .I2(\REG.mem_60_3 ), 
            .I3(rd_addr_r[1]), .O(n10979));
    defparam n12645_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4074_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_33_0 ), .O(n5457));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4074_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13263_bdd_4_lut (.I0(n13263), .I1(\REG.mem_5_12 ), .I2(\REG.mem_4_12 ), 
            .I3(rd_addr_r[1]), .O(n13266));
    defparam n13263_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i86_2_lut_3_lut_4_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n57));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i86_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_DFF i161_162 (.Q(\REG.mem_1_9 ), .C(FIFO_CLK_c), .D(n4833));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10797 (.I0(rd_addr_r[2]), .I1(n10895), 
            .I2(n10907), .I3(rd_addr_r[3]), .O(n12639));
    defparam rd_addr_r_2__bdd_4_lut_10797.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i85_2_lut_3_lut_4_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n25));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i85_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11217 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_38_3 ), 
            .I2(\REG.mem_39_3 ), .I3(rd_addr_r[1]), .O(n13257));
    defparam rd_addr_r_0__bdd_4_lut_11217.LUT_INIT = 16'he4aa;
    SB_DFF i179_180 (.Q(\REG.mem_1_15 ), .C(FIFO_CLK_c), .D(n4832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13257_bdd_4_lut (.I0(n13257), .I1(\REG.mem_37_3 ), .I2(\REG.mem_36_3 ), 
            .I3(rd_addr_r[1]), .O(n10937));
    defparam n13257_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11232 (.I0(rd_addr_r[1]), .I1(n11319), 
            .I2(n11320), .I3(rd_addr_r[2]), .O(n13251));
    defparam rd_addr_r_1__bdd_4_lut_11232.LUT_INIT = 16'he4aa;
    SB_LUT4 n13251_bdd_4_lut (.I0(n13251), .I1(n11308), .I2(n11307), .I3(rd_addr_r[2]), 
            .O(n11410));
    defparam n13251_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_en_i_I_0_2_lut (.I0(DEBUG_5_c), .I1(full_o), .I2(GND_net), 
            .I3(GND_net), .O(wr_sig_mv_w));   // src/fifo_dc_32_lut_gen.v(293[28:49])
    defparam wr_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_DFF i164_165 (.Q(\REG.mem_1_10 ), .C(FIFO_CLK_c), .D(n4831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12639_bdd_4_lut (.I0(n12639), .I1(n10892), .I2(n10886), .I3(rd_addr_r[3]), 
            .O(n10982));
    defparam n12639_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11212 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_42_3 ), 
            .I2(\REG.mem_43_3 ), .I3(rd_addr_r[1]), .O(n13245));
    defparam rd_addr_r_0__bdd_4_lut_11212.LUT_INIT = 16'he4aa;
    SB_LUT4 n13245_bdd_4_lut (.I0(n13245), .I1(\REG.mem_41_3 ), .I2(\REG.mem_40_3 ), 
            .I3(rd_addr_r[1]), .O(n10940));
    defparam n13245_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10733 (.I0(rd_addr_r[1]), .I1(n11718), 
            .I2(n11719), .I3(rd_addr_r[2]), .O(n12633));
    defparam rd_addr_r_1__bdd_4_lut_10733.LUT_INIT = 16'he4aa;
    SB_LUT4 n12633_bdd_4_lut (.I0(n12633), .I1(n11716), .I2(n11715), .I3(rd_addr_r[2]), 
            .O(n12636));
    defparam n12633_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11202 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_58_0 ), 
            .I2(\REG.mem_59_0 ), .I3(rd_addr_r[1]), .O(n13239));
    defparam rd_addr_r_0__bdd_4_lut_11202.LUT_INIT = 16'he4aa;
    SB_LUT4 n13239_bdd_4_lut (.I0(n13239), .I1(\REG.mem_57_0 ), .I2(\REG.mem_56_0 ), 
            .I3(rd_addr_r[1]), .O(n13242));
    defparam n13239_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i2_2_lut_4_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1_w[1]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_498[2] ), .O(rd_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4535_2_lut_4_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1_w[1]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5918));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4535_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i1_2_lut_4_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1_w[1]), 
            .I2(rd_fifo_en_w), .I3(rd_addr_nxt_c_6__N_498[0]), .O(rd_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10703 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_38_12 ), 
            .I2(\REG.mem_39_12 ), .I3(rd_addr_r[1]), .O(n12627));
    defparam rd_addr_r_0__bdd_4_lut_10703.LUT_INIT = 16'he4aa;
    SB_LUT4 n12627_bdd_4_lut (.I0(n12627), .I1(\REG.mem_37_12 ), .I2(\REG.mem_36_12 ), 
            .I3(rd_addr_r[1]), .O(n12630));
    defparam n12627_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4105_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_34_15 ), .O(n5488));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4105_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i116_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n42));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i116_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i18_2_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n18_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i18_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 EnabledDecoder_2_i115_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n10));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i115_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3483_2_lut_4_lut (.I0(wr_addr_r[0]), .I1(wr_addr_p1_w[0]), 
            .I2(wr_sig_mv_w), .I3(reset_per_frame), .O(n4866));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i3483_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i4104_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_34_14 ), .O(n5487));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4104_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i1_2_lut_4_lut (.I0(wr_addr_r[0]), .I1(wr_addr_p1_w[0]), 
            .I2(wr_sig_mv_w), .I3(\wr_addr_nxt_c[1] ), .O(wr_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4103_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_34_13 ), .O(n5486));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4103_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i84_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n58));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i84_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11197 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_6 ), 
            .I2(\REG.mem_15_6 ), .I3(rd_addr_r[1]), .O(n13233));
    defparam rd_addr_r_0__bdd_4_lut_11197.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10688 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_1 ), 
            .I2(\REG.mem_11_1 ), .I3(rd_addr_r[1]), .O(n12621));
    defparam rd_addr_r_0__bdd_4_lut_10688.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i83_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n26));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i83_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i114_2_lut_3_lut (.I0(n34_adj_1205), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n43));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i114_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 n13233_bdd_4_lut (.I0(n13233), .I1(\REG.mem_13_6 ), .I2(\REG.mem_12_6 ), 
            .I3(rd_addr_r[1]), .O(n10946));
    defparam n13233_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i130_2_lut_3_lut (.I0(n33), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n35));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i130_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i113_2_lut_3_lut (.I0(n34_adj_1205), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n11));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i113_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i129_2_lut_3_lut (.I0(n33), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n3));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i129_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n12621_bdd_4_lut (.I0(n12621), .I1(\REG.mem_9_1 ), .I2(\REG.mem_8_1 ), 
            .I3(rd_addr_r[1]), .O(n11153));
    defparam n12621_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9425_3_lut (.I0(\REG.mem_6_10 ), .I1(\REG.mem_7_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11275));
    defparam i9425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9424_3_lut (.I0(\REG.mem_4_10 ), .I1(\REG.mem_5_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11274));
    defparam i9424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9202_3_lut (.I0(\REG.mem_0_7 ), .I1(\REG.mem_1_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11052));
    defparam i9202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11192 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_2_8 ), 
            .I2(\REG.mem_3_8 ), .I3(rd_addr_r[1]), .O(n13227));
    defparam rd_addr_r_0__bdd_4_lut_11192.LUT_INIT = 16'he4aa;
    SB_LUT4 n13227_bdd_4_lut (.I0(n13227), .I1(\REG.mem_1_8 ), .I2(\REG.mem_0_8 ), 
            .I3(rd_addr_r[1]), .O(n13230));
    defparam n13227_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9203_3_lut (.I0(\REG.mem_2_7 ), .I1(\REG.mem_3_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11053));
    defparam i9203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10683 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_34_5 ), 
            .I2(\REG.mem_35_5 ), .I3(rd_addr_r[1]), .O(n12615));
    defparam rd_addr_r_0__bdd_4_lut_10683.LUT_INIT = 16'he4aa;
    SB_LUT4 i4102_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_34_12 ), .O(n5485));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4102_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4101_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_34_11 ), .O(n5484));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4101_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11317 (.I0(rd_addr_r[3]), .I1(n12594), 
            .I2(n10900), .I3(rd_addr_r[4]), .O(n13221));
    defparam rd_addr_r_3__bdd_4_lut_11317.LUT_INIT = 16'he4aa;
    SB_LUT4 i9245_3_lut (.I0(\REG.mem_6_7 ), .I1(\REG.mem_7_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11095));
    defparam i9245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12615_bdd_4_lut (.I0(n12615), .I1(\REG.mem_33_5 ), .I2(\REG.mem_32_5 ), 
            .I3(rd_addr_r[1]), .O(n12618));
    defparam n12615_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9244_3_lut (.I0(\REG.mem_4_7 ), .I1(\REG.mem_5_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11094));
    defparam i9244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4433_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_53_15 ), .O(n5816));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4433_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4100_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_34_10 ), .O(n5483));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4100_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i34_2_lut_3_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n34_adj_1205));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i34_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 n13221_bdd_4_lut (.I0(n13221), .I1(n10855), .I2(n12504), .I3(rd_addr_r[4]), 
            .O(n13224));
    defparam n13221_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9448_3_lut (.I0(\REG.mem_16_10 ), .I1(\REG.mem_17_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11298));
    defparam i9448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i33_2_lut_3_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n33));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i33_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i9449_3_lut (.I0(\REG.mem_18_10 ), .I1(\REG.mem_19_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11299));
    defparam i9449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4432_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_53_14 ), .O(n5815));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4432_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i338_339 (.Q(\REG.mem_3_4 ), .C(FIFO_CLK_c), .D(n4968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9445_3_lut (.I0(\REG.mem_40_7 ), .I1(\REG.mem_41_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11295));
    defparam i9445_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i335_336 (.Q(\REG.mem_3_3 ), .C(FIFO_CLK_c), .D(n4967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9446_3_lut (.I0(\REG.mem_42_7 ), .I1(\REG.mem_43_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11296));
    defparam i9446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11272 (.I0(rd_addr_r[4]), .I1(n11753), 
            .I2(n11789), .I3(rd_addr_r[5]), .O(n12609));
    defparam rd_addr_r_4__bdd_4_lut_11272.LUT_INIT = 16'he4aa;
    SB_LUT4 i4431_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_53_13 ), .O(n5814));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4431_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11207 (.I0(rd_addr_r[1]), .I1(n11358), 
            .I2(n11359), .I3(rd_addr_r[2]), .O(n13215));
    defparam rd_addr_r_1__bdd_4_lut_11207.LUT_INIT = 16'he4aa;
    SB_LUT4 n12609_bdd_4_lut (.I0(n12609), .I1(n11696), .I2(n12222), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_559 [1]));
    defparam n12609_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13215_bdd_4_lut (.I0(n13215), .I1(n11347), .I2(n11346), .I3(rd_addr_r[2]), 
            .O(n11413));
    defparam n13215_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i332_333 (.Q(\REG.mem_3_2 ), .C(FIFO_CLK_c), .D(n4966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4430_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_53_12 ), .O(n5813));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4430_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i329_330 (.Q(\REG.mem_3_1 ), .C(FIFO_CLK_c), .D(n4965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10723 (.I0(rd_addr_r[3]), .I1(n12516), 
            .I2(n10867), .I3(rd_addr_r[4]), .O(n12603));
    defparam rd_addr_r_3__bdd_4_lut_10723.LUT_INIT = 16'he4aa;
    SB_DFF i326_327 (.Q(\REG.mem_3_0 ), .C(FIFO_CLK_c), .D(n4964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4429_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_53_11 ), .O(n5812));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4429_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12603_bdd_4_lut (.I0(n12603), .I1(n11800), .I2(n11799), .I3(rd_addr_r[4]), 
            .O(n12606));
    defparam n12603_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11187 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_6_6 ), 
            .I2(\REG.mem_7_6 ), .I3(rd_addr_r[1]), .O(n13209));
    defparam rd_addr_r_0__bdd_4_lut_11187.LUT_INIT = 16'he4aa;
    SB_LUT4 i4099_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_34_9 ), .O(n5482));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4099_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4428_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_53_10 ), .O(n5811));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4428_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13209_bdd_4_lut (.I0(n13209), .I1(\REG.mem_5_6 ), .I2(\REG.mem_4_6 ), 
            .I3(rd_addr_r[1]), .O(n11876));
    defparam n13209_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4427_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_53_9 ), .O(n5810));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4427_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4098_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_34_8 ), .O(n5481));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4098_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4426_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_53_8 ), .O(n5809));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4426_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11172 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_5 ), 
            .I2(\REG.mem_11_5 ), .I3(rd_addr_r[1]), .O(n13203));
    defparam rd_addr_r_0__bdd_4_lut_11172.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10693 (.I0(rd_addr_r[1]), .I1(n11742), 
            .I2(n11743), .I3(rd_addr_r[2]), .O(n12597));
    defparam rd_addr_r_1__bdd_4_lut_10693.LUT_INIT = 16'he4aa;
    SB_LUT4 n13203_bdd_4_lut (.I0(n13203), .I1(\REG.mem_9_5 ), .I2(\REG.mem_8_5 ), 
            .I3(rd_addr_r[1]), .O(n13206));
    defparam n13203_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i15_2_lut (.I0(n12_adj_1199), .I1(wr_addr_r[2]), 
            .I2(GND_net), .I3(GND_net), .O(n15_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i15_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n12597_bdd_4_lut (.I0(n12597), .I1(n11731), .I2(n11730), .I3(rd_addr_r[2]), 
            .O(n12600));
    defparam n12597_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11177 (.I0(rd_addr_r[1]), .I1(n11247), 
            .I2(n11248), .I3(rd_addr_r[2]), .O(n13197));
    defparam rd_addr_r_1__bdd_4_lut_11177.LUT_INIT = 16'he4aa;
    SB_DFF i275_276 (.Q(\REG.mem_2_15 ), .C(FIFO_CLK_c), .D(n4963));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4425_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_53_7 ), .O(n5808));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4425_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13197_bdd_4_lut (.I0(n13197), .I1(n11227), .I2(n11226), .I3(rd_addr_r[2]), 
            .O(n11419));
    defparam n13197_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4424_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_53_6 ), .O(n5807));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4424_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4423_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_53_5 ), .O(n5806));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4423_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4422_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_53_4 ), .O(n5805));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4422_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10663 (.I0(rd_addr_r[1]), .I1(n11712), 
            .I2(n11713), .I3(rd_addr_r[2]), .O(n12591));
    defparam rd_addr_r_1__bdd_4_lut_10663.LUT_INIT = 16'he4aa;
    SB_LUT4 n12591_bdd_4_lut (.I0(n12591), .I1(n11704), .I2(n11703), .I3(rd_addr_r[2]), 
            .O(n12594));
    defparam n12591_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4421_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_53_3 ), .O(n5804));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4421_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i272_273 (.Q(\REG.mem_2_14 ), .C(FIFO_CLK_c), .D(n4962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4420_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_53_2 ), .O(n5803));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4420_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i269_270 (.Q(\REG.mem_2_13 ), .C(FIFO_CLK_c), .D(n4961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10326 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_14_1 ), 
            .I2(\REG.mem_15_1 ), .I3(rd_addr_r[1]), .O(n12171));
    defparam rd_addr_r_0__bdd_4_lut_10326.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10678 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_22_0 ), 
            .I2(\REG.mem_23_0 ), .I3(rd_addr_r[1]), .O(n12585));
    defparam rd_addr_r_0__bdd_4_lut_10678.LUT_INIT = 16'he4aa;
    SB_LUT4 n12585_bdd_4_lut (.I0(n12585), .I1(\REG.mem_21_0 ), .I2(\REG.mem_20_0 ), 
            .I3(rd_addr_r[1]), .O(n12588));
    defparam n12585_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4097_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_34_7 ), .O(n5480));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4097_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4096_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_34_6 ), .O(n5479));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4096_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11167 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_10_12 ), 
            .I2(\REG.mem_11_12 ), .I3(rd_addr_r[1]), .O(n13191));
    defparam rd_addr_r_0__bdd_4_lut_11167.LUT_INIT = 16'he4aa;
    SB_LUT4 n13191_bdd_4_lut (.I0(n13191), .I1(\REG.mem_9_12 ), .I2(\REG.mem_8_12 ), 
            .I3(rd_addr_r[1]), .O(n13194));
    defparam n13191_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4419_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_53_1 ), .O(n5802));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4419_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10653 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_46_11 ), 
            .I2(\REG.mem_47_11 ), .I3(rd_addr_r[1]), .O(n12579));
    defparam rd_addr_r_0__bdd_4_lut_10653.LUT_INIT = 16'he4aa;
    SB_DFF i266_267 (.Q(\REG.mem_2_12 ), .C(FIFO_CLK_c), .D(n4960));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i263_264 (.Q(\REG.mem_2_11 ), .C(FIFO_CLK_c), .D(n4959));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11302 (.I0(rd_addr_r[2]), .I1(n12732), 
            .I2(n12660), .I3(rd_addr_r[3]), .O(n13185));
    defparam rd_addr_r_2__bdd_4_lut_11302.LUT_INIT = 16'he4aa;
    SB_LUT4 i9452_3_lut (.I0(\REG.mem_22_10 ), .I1(\REG.mem_23_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11302));
    defparam i9452_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i260_261 (.Q(\REG.mem_2_10 ), .C(FIFO_CLK_c), .D(n4958));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13185_bdd_4_lut (.I0(n13185), .I1(n12768), .I2(n12774), .I3(rd_addr_r[3]), 
            .O(n13188));
    defparam n13185_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4418_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_53_0 ), .O(n5801));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4418_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9451_3_lut (.I0(\REG.mem_20_10 ), .I1(\REG.mem_21_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11301));
    defparam i9451_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i257_258 (.Q(\REG.mem_2_9 ), .C(FIFO_CLK_c), .D(n4957));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i254_255 (.Q(\REG.mem_2_8 ), .C(FIFO_CLK_c), .D(n4956));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4095_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_34_5 ), .O(n5478));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4095_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i251_252 (.Q(\REG.mem_2_7 ), .C(FIFO_CLK_c), .D(n4955));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9478_3_lut (.I0(\REG.mem_32_10 ), .I1(\REG.mem_33_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11328));
    defparam i9478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12579_bdd_4_lut (.I0(n12579), .I1(\REG.mem_45_11 ), .I2(\REG.mem_44_11 ), 
            .I3(rd_addr_r[1]), .O(n11552));
    defparam n12579_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i80_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n60));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i80_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i4094_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_34_4 ), .O(n5477));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4094_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9479_3_lut (.I0(\REG.mem_34_10 ), .I1(\REG.mem_35_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11329));
    defparam i9479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i79_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n28));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i79_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 n12171_bdd_4_lut (.I0(n12171), .I1(\REG.mem_13_1 ), .I2(\REG.mem_12_1 ), 
            .I3(rd_addr_r[1]), .O(n12174));
    defparam n12171_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11157 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_22_13 ), 
            .I2(\REG.mem_23_13 ), .I3(rd_addr_r[1]), .O(n13179));
    defparam rd_addr_r_0__bdd_4_lut_11157.LUT_INIT = 16'he4aa;
    SB_LUT4 n13179_bdd_4_lut (.I0(n13179), .I1(\REG.mem_21_13 ), .I2(\REG.mem_20_13 ), 
            .I3(rd_addr_r[1]), .O(n13182));
    defparam n13179_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9491_3_lut (.I0(\REG.mem_38_10 ), .I1(\REG.mem_39_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11341));
    defparam i9491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9490_3_lut (.I0(\REG.mem_36_10 ), .I1(\REG.mem_37_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11340));
    defparam i9490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i82_2_lut_3_lut (.I0(n34_adj_1205), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n59));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i82_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i81_2_lut_3_lut (.I0(n34_adj_1205), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n27));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i81_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11147 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_30_8 ), 
            .I2(\REG.mem_31_8 ), .I3(rd_addr_r[1]), .O(n13173));
    defparam rd_addr_r_0__bdd_4_lut_11147.LUT_INIT = 16'he4aa;
    SB_LUT4 i4093_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_34_3 ), .O(n5476));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4093_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4092_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_34_2 ), .O(n5475));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4092_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4091_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_34_1 ), .O(n5474));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4091_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9467_3_lut (.I0(\REG.mem_46_7 ), .I1(\REG.mem_47_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11317));
    defparam i9467_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i248_249 (.Q(\REG.mem_2_6 ), .C(FIFO_CLK_c), .D(n4954));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10648 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_26_0 ), 
            .I2(\REG.mem_27_0 ), .I3(rd_addr_r[1]), .O(n12573));
    defparam rd_addr_r_0__bdd_4_lut_10648.LUT_INIT = 16'he4aa;
    SB_DFF i245_246 (.Q(\REG.mem_2_5 ), .C(FIFO_CLK_c), .D(n4953));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4090_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_34_0 ), .O(n5473));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4090_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i242_243 (.Q(\REG.mem_2_4 ), .C(FIFO_CLK_c), .D(n4952));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13173_bdd_4_lut (.I0(n13173), .I1(\REG.mem_29_8 ), .I2(\REG.mem_28_8 ), 
            .I3(rd_addr_r[1]), .O(n13176));
    defparam n13173_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i239_240 (.Q(\REG.mem_2_3 ), .C(FIFO_CLK_c), .D(n4951));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3532_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_1_11 ), .O(n4915));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3532_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11142 (.I0(\rd_addr_r[0] ), .I1(\REG.mem_42_1 ), 
            .I2(\REG.mem_43_1 ), .I3(rd_addr_r[1]), .O(n13167));
    defparam rd_addr_r_0__bdd_4_lut_11142.LUT_INIT = 16'he4aa;
    SB_LUT4 i9466_3_lut (.I0(\REG.mem_44_7 ), .I1(\REG.mem_45_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11316));
    defparam i9466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12573_bdd_4_lut (.I0(n12573), .I1(\REG.mem_25_0 ), .I2(\REG.mem_24_0 ), 
            .I3(rd_addr_r[1]), .O(n12576));
    defparam n12573_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13167_bdd_4_lut (.I0(n13167), .I1(\REG.mem_41_1 ), .I2(\REG.mem_40_1 ), 
            .I3(rd_addr_r[1]), .O(n13170));
    defparam n13167_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3519_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_1_13 ), .O(n4902));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3519_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4417_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_52_15 ), .O(n5800));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4417_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9211_3_lut (.I0(\REG.mem_20_9 ), .I1(\REG.mem_21_9 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11061));
    defparam i9211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9212_3_lut (.I0(\REG.mem_22_9 ), .I1(\REG.mem_23_9 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11062));
    defparam i9212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4416_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_52_14 ), .O(n5799));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4416_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9188_3_lut (.I0(\REG.mem_18_9 ), .I1(\REG.mem_19_9 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11038));
    defparam i9188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9187_3_lut (.I0(\REG.mem_16_9 ), .I1(\REG.mem_17_9 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11037));
    defparam i9187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4415_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_52_13 ), .O(n5798));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4415_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4414_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_52_12 ), .O(n5797));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4414_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4413_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_52_11 ), .O(n5796));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4413_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4412_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_52_10 ), .O(n5795));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4412_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4411_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_52_9 ), .O(n5794));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4411_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i3_2_lut (.I0(\rd_addr_nxt_c_6__N_498[2] ), 
            .I1(\rd_addr_nxt_c_6__N_498[3] ), .I2(GND_net), .I3(GND_net), 
            .O(rd_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(504[28:66])
    defparam rd_addr_nxt_c_6__I_0_152_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4410_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_52_8 ), .O(n5793));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4410_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4409_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_52_7 ), .O(n5792));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4409_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4408_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_52_6 ), .O(n5791));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4408_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4407_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_52_5 ), .O(n5790));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4407_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4406_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_52_4 ), .O(n5789));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4406_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9029_3_lut (.I0(n12144), .I1(n12114), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10879));
    defparam i9029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9028_3_lut (.I0(n12360), .I1(n12282), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10878));
    defparam i9028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4405_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_52_3 ), .O(n5788));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4405_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4404_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_52_2 ), .O(n5787));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4404_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9997_3_lut (.I0(\REG.mem_44_14 ), .I1(\REG.mem_45_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11847));
    defparam i9997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9998_3_lut (.I0(\REG.mem_46_14 ), .I1(\REG.mem_47_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11848));
    defparam i9998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9992_3_lut (.I0(\REG.mem_42_14 ), .I1(\REG.mem_43_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11842));
    defparam i9992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9991_3_lut (.I0(\REG.mem_40_14 ), .I1(\REG.mem_41_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11841));
    defparam i9991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9433_3_lut (.I0(\REG.mem_60_5 ), .I1(\REG.mem_61_5 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11283));
    defparam i9433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9434_3_lut (.I0(\REG.mem_62_5 ), .I1(\REG.mem_63_5 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11284));
    defparam i9434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9422_3_lut (.I0(\REG.mem_58_5 ), .I1(\REG.mem_59_5 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11272));
    defparam i9422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9421_3_lut (.I0(\REG.mem_56_5 ), .I1(\REG.mem_57_5 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11271));
    defparam i9421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4403_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_52_1 ), .O(n5786));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4403_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3529_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_1_12 ), .O(n4912));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3529_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9886_3_lut (.I0(n13044), .I1(n13014), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11736));
    defparam i9886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9887_3_lut (.I0(n12900), .I1(n12822), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11737));
    defparam i9887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9875_3_lut (.I0(n13194), .I1(n13110), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11725));
    defparam i9875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9874_3_lut (.I0(n13362), .I1(n13266), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11724));
    defparam i9874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3448_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_1_10 ), .O(n4831));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3448_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3450_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_1_9 ), .O(n4833));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3450_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4402_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_52_0 ), .O(n5785));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4402_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i45_2_lut_3_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n45));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i45_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i78_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n61));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i78_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i47_2_lut_3_lut_4_lut (.I0(n12_adj_1199), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n47_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i47_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i3484_3_lut_4_lut (.I0(n40_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_1_14 ), .O(n4867));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3484_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i77_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n29));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i77_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i9494_3_lut (.I0(n12198), .I1(n13704), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11344));
    defparam i9494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9493_3_lut (.I0(n12618), .I1(n12276), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11343));
    defparam i9493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9250_3_lut (.I0(n12168), .I1(n13518), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11100));
    defparam i9250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4401_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_51_15 ), .O(n5784));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4401_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8895_4_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_r[4]), .I2(rp_sync2_r[3]), 
            .I3(rp_sync_w[4]), .O(n10744));
    defparam i8895_4_lut_4_lut.LUT_INIT = 16'hdeb7;
    SB_LUT4 i9235_3_lut (.I0(\REG.mem_52_4 ), .I1(\REG.mem_53_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11085));
    defparam i9235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9236_3_lut (.I0(\REG.mem_54_4 ), .I1(\REG.mem_55_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11086));
    defparam i9236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9227_3_lut (.I0(\REG.mem_50_4 ), .I1(\REG.mem_51_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11077));
    defparam i9227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9226_3_lut (.I0(\REG.mem_48_4 ), .I1(\REG.mem_49_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11076));
    defparam i9226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9214_3_lut (.I0(\REG.mem_36_4 ), .I1(\REG.mem_37_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11064));
    defparam i9214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9215_3_lut (.I0(\REG.mem_38_4 ), .I1(\REG.mem_39_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11065));
    defparam i9215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9209_3_lut (.I0(\REG.mem_34_4 ), .I1(\REG.mem_35_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11059));
    defparam i9209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9208_3_lut (.I0(\REG.mem_32_4 ), .I1(\REG.mem_33_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11058));
    defparam i9208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9190_3_lut (.I0(\REG.mem_20_4 ), .I1(\REG.mem_21_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11040));
    defparam i9190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9191_3_lut (.I0(\REG.mem_22_4 ), .I1(\REG.mem_23_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11041));
    defparam i9191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9179_3_lut (.I0(\REG.mem_18_4 ), .I1(\REG.mem_19_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11029));
    defparam i9179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9178_3_lut (.I0(\REG.mem_16_4 ), .I1(\REG.mem_17_4 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11028));
    defparam i9178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4400_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_51_14 ), .O(n5783));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4400_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut (.I0(rp_sync2_r[2]), .I1(rp_sync2_r[3]), .I2(rp_sync_w[4]), 
            .I3(GND_net), .O(rp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_51 (.I0(rp_sync2_r[0]), .I1(rp_sync2_r[1]), 
            .I2(rp_sync_w[2]), .I3(GND_net), .O(rp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_3_lut_adj_51.LUT_INIT = 16'h9696;
    SB_LUT4 rd_fifo_en_w_I_0_158_2_lut_3_lut (.I0(DEBUG_3_c), .I1(get_next_word), 
            .I2(\genblk16.rd_prev_r ), .I3(GND_net), .O(t_rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(747[41:67])
    defparam rd_fifo_en_w_I_0_158_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_LUT4 EnabledDecoder_2_i11_2_lut_3_lut_4_lut (.I0(DEBUG_5_c), .I1(full_o), 
            .I2(wr_addr_r[0]), .I3(wr_addr_r[1]), .O(n11_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i12_2_lut_3_lut_4_lut (.I0(DEBUG_5_c), .I1(full_o), 
            .I2(wr_addr_r[0]), .I3(wr_addr_r[1]), .O(n12_adj_1199));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i12_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i4399_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_51_13 ), .O(n5782));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4399_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i57_2_lut_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n57_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i57_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i9840_3_lut (.I0(n13284), .I1(n11689), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n11690));
    defparam i9840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9839_3_lut (.I0(n13512), .I1(n13488), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11689));
    defparam i9839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9436_3_lut (.I0(\REG.mem_12_10 ), .I1(\REG.mem_13_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11286));
    defparam i9436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9437_3_lut (.I0(\REG.mem_14_10 ), .I1(\REG.mem_15_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11287));
    defparam i9437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9428_3_lut (.I0(\REG.mem_10_10 ), .I1(\REG.mem_11_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11278));
    defparam i9428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9427_3_lut (.I0(\REG.mem_8_10 ), .I1(\REG.mem_9_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11277));
    defparam i9427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3289_1_lut (.I0(\fifo_data_out[10] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4672));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3289_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9985_3_lut (.I0(\REG.mem_36_14 ), .I1(\REG.mem_37_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11835));
    defparam i9985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9986_3_lut (.I0(\REG.mem_38_14 ), .I1(\REG.mem_39_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11836));
    defparam i9986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3288_1_lut (.I0(\fifo_data_out[9] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4671));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3288_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9980_3_lut (.I0(\REG.mem_34_14 ), .I1(\REG.mem_35_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11830));
    defparam i9980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9979_3_lut (.I0(\REG.mem_32_14 ), .I1(\REG.mem_33_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11829));
    defparam i9979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9418_3_lut (.I0(\REG.mem_20_1 ), .I1(\REG.mem_21_1 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11268));
    defparam i9418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9419_3_lut (.I0(\REG.mem_22_1 ), .I1(\REG.mem_23_1 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11269));
    defparam i9419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4398_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_51_12 ), .O(n5781));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4398_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i59_2_lut_3_lut_4_lut (.I0(n11_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n59_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i59_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i9389_3_lut (.I0(\REG.mem_18_1 ), .I1(\REG.mem_19_1 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11239));
    defparam i9389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9388_3_lut (.I0(\REG.mem_16_1 ), .I1(\REG.mem_17_1 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11238));
    defparam i9388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9913_3_lut (.I0(\REG.mem_28_14 ), .I1(\REG.mem_29_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11763));
    defparam i9913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9914_3_lut (.I0(\REG.mem_30_14 ), .I1(\REG.mem_31_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11764));
    defparam i9914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3287_1_lut (.I0(\fifo_data_out[11] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4670));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3287_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9890_3_lut (.I0(\REG.mem_26_14 ), .I1(\REG.mem_27_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11740));
    defparam i9890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9889_3_lut (.I0(\REG.mem_24_14 ), .I1(\REG.mem_25_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11739));
    defparam i9889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3286_1_lut (.I0(\fifo_data_out[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4669));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3286_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3285_1_lut (.I0(\fifo_data_out[13] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4668));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3285_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10021_3_lut (.I0(n13692), .I1(n13578), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11871));
    defparam i10021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10022_3_lut (.I0(n13428), .I1(n13176), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11872));
    defparam i10022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10004_3_lut (.I0(n13452), .I1(n12414), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11854));
    defparam i10004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10003_3_lut (.I0(n13230), .I1(n13560), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11853));
    defparam i10003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i9_2_lut_3_lut_4_lut (.I0(DEBUG_5_c), .I1(full_o), 
            .I2(wr_addr_r[0]), .I3(wr_addr_r[1]), .O(n9));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i9_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i3284_1_lut (.I0(\fifo_data_out[14] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4667));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3284_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9961_3_lut (.I0(\REG.mem_4_13 ), .I1(\REG.mem_5_13 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11811));
    defparam i9961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9962_3_lut (.I0(\REG.mem_6_13 ), .I1(\REG.mem_7_13 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11812));
    defparam i9962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i42_2_lut_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n42_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i42_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i9944_3_lut (.I0(\REG.mem_2_13 ), .I1(\REG.mem_3_13 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11794));
    defparam i9944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9943_3_lut (.I0(\REG.mem_0_13 ), .I1(\REG.mem_1_13 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11793));
    defparam i9943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4397_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_51_11 ), .O(n5780));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4397_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8917_4_lut_4_lut (.I0(rd_addr_r[1]), .I1(rd_addr_r[2]), .I2(wp_sync2_r[1]), 
            .I3(wp_sync_w[2]), .O(n10766));
    defparam i8917_4_lut_4_lut.LUT_INIT = 16'hb7de;
    SB_LUT4 i4396_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_51_10 ), .O(n5779));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4396_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_52 (.I0(wp_sync2_r[4]), .I1(wp_sync2_r[6]), 
            .I2(wp_sync2_r[5]), .I3(GND_net), .O(wp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_52.LUT_INIT = 16'h9696;
    SB_LUT4 i4395_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_51_9 ), .O(n5778));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4395_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_53 (.I0(wp_sync2_r[0]), .I1(wp_sync2_r[1]), 
            .I2(wp_sync_w[2]), .I3(GND_net), .O(wp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_53.LUT_INIT = 16'h9696;
    SB_LUT4 i4394_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_51_8 ), .O(n5777));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4394_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_54 (.I0(wp_sync2_r[2]), .I1(wp_sync2_r[3]), 
            .I2(wp_sync_w[4]), .I3(GND_net), .O(wp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_54.LUT_INIT = 16'h9696;
    SB_LUT4 i4393_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_51_7 ), .O(n5776));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4393_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i63_2_lut_3_lut_4_lut (.I0(n12_adj_1199), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n63));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i63_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4392_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_51_6 ), .O(n5775));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4392_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4391_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_51_5 ), .O(n5774));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4391_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4390_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_51_4 ), .O(n5773));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4390_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4389_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_51_3 ), .O(n5772));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4389_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4388_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_51_2 ), .O(n5771));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4388_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4387_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_51_1 ), .O(n5770));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4387_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4386_3_lut_4_lut (.I0(n43_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_51_0 ), .O(n5769));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4386_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9469_3_lut (.I0(\REG.mem_28_10 ), .I1(\REG.mem_29_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11319));
    defparam i9469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9470_3_lut (.I0(\REG.mem_30_10 ), .I1(\REG.mem_31_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11320));
    defparam i9470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9458_3_lut (.I0(\REG.mem_26_10 ), .I1(\REG.mem_27_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11308));
    defparam i9458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9457_3_lut (.I0(\REG.mem_24_10 ), .I1(\REG.mem_25_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11307));
    defparam i9457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3283_1_lut (.I0(\fifo_data_out[8] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4666));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9868_3_lut (.I0(\REG.mem_20_14 ), .I1(\REG.mem_21_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11718));
    defparam i9868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9869_3_lut (.I0(\REG.mem_22_14 ), .I1(\REG.mem_23_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11719));
    defparam i9869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9866_3_lut (.I0(\REG.mem_18_14 ), .I1(\REG.mem_19_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11716));
    defparam i9866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9865_3_lut (.I0(\REG.mem_16_14 ), .I1(\REG.mem_17_14 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11715));
    defparam i9865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3282_1_lut (.I0(\fifo_data_out[15] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4665));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3282_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3281_1_lut (.I0(\fifo_data_out[7] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4664));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3281_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3280_1_lut (.I0(\fifo_data_out[6] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4663));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3280_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3279_1_lut (.I0(\fifo_data_out[5] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4662));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3279_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3278_1_lut (.I0(\fifo_data_out[4] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4661));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3278_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9005_3_lut (.I0(n12396), .I1(n13710), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10855));
    defparam i9005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3277_1_lut (.I0(\fifo_data_out[3] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4660));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3277_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9508_3_lut (.I0(\REG.mem_44_10 ), .I1(\REG.mem_45_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11358));
    defparam i9508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9509_3_lut (.I0(\REG.mem_46_10 ), .I1(\REG.mem_47_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11359));
    defparam i9509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9846_3_lut (.I0(n13302), .I1(n11695), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n11696));
    defparam i9846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9845_3_lut (.I0(n13566), .I1(n13482), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11695));
    defparam i9845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9497_3_lut (.I0(\REG.mem_42_10 ), .I1(\REG.mem_43_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11347));
    defparam i9497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9496_3_lut (.I0(\REG.mem_40_10 ), .I1(\REG.mem_41_10 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11346));
    defparam i9496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9017_3_lut (.I0(n12438), .I1(n12384), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10867));
    defparam i9017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9950_3_lut (.I0(n12834), .I1(n12714), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11800));
    defparam i9950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9949_3_lut (.I0(n13026), .I1(n12894), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11799));
    defparam i9949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9892_3_lut (.I0(\REG.mem_52_15 ), .I1(\REG.mem_53_15 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11742));
    defparam i9892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9893_3_lut (.I0(\REG.mem_54_15 ), .I1(\REG.mem_55_15 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11743));
    defparam i9893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3276_1_lut (.I0(\fifo_data_out[2] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4659));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3276_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9881_3_lut (.I0(\REG.mem_50_15 ), .I1(\REG.mem_51_15 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11731));
    defparam i9881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9880_3_lut (.I0(\REG.mem_48_15 ), .I1(\REG.mem_49_15 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11730));
    defparam i9880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9397_3_lut (.I0(\REG.mem_28_7 ), .I1(\REG.mem_29_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11247));
    defparam i9397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9398_3_lut (.I0(\REG.mem_30_7 ), .I1(\REG.mem_31_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11248));
    defparam i9398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9377_3_lut (.I0(\REG.mem_26_7 ), .I1(\REG.mem_27_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11227));
    defparam i9377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9376_3_lut (.I0(\REG.mem_24_7 ), .I1(\REG.mem_25_7 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11226));
    defparam i9376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3275_1_lut (.I0(\fifo_data_out[1] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4658));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    defparam i3275_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9862_3_lut (.I0(\REG.mem_52_8 ), .I1(\REG.mem_53_8 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11712));
    defparam i9862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9863_3_lut (.I0(\REG.mem_54_8 ), .I1(\REG.mem_55_8 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11713));
    defparam i9863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9854_3_lut (.I0(\REG.mem_50_8 ), .I1(\REG.mem_51_8 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11704));
    defparam i9854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9853_3_lut (.I0(\REG.mem_48_8 ), .I1(\REG.mem_49_8 ), .I2(\rd_addr_r[0] ), 
            .I3(GND_net), .O(n11703));
    defparam i9853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i43_2_lut_3_lut_4_lut (.I0(n11_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n43_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i43_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=20) 
//

module \uart_rx(CLKS_PER_BIT=20)  (SLM_CLK_c, r_Rx_Data, GND_net, debug_led3, 
            n4248, n4253, n4, n4_adj_1, n7347, n6083, pc_data_rx, 
            VCC_net, n6067, n6066, n6064, n6063, n6062, n6060, 
            n4_adj_2, n10211, UART_RX_c, n6030) /* synthesis syn_module_defined=1 */ ;
    input SLM_CLK_c;
    output r_Rx_Data;
    input GND_net;
    output debug_led3;
    output n4248;
    output n4253;
    output n4;
    output n4_adj_1;
    output n7347;
    input n6083;
    output [7:0]pc_data_rx;
    input VCC_net;
    input n6067;
    input n6066;
    input n6064;
    input n6063;
    input n6062;
    input n6060;
    output n4_adj_2;
    output n10211;
    input UART_RX_c;
    input n6030;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n3;
    wire [2:0]r_SM_Main;   // src/uart_rx.v(36[17:26])
    
    wire r_Rx_Data_R;
    wire [2:0]r_SM_Main_2__N_765;
    
    wire n55, n145, n3_adj_1182;
    wire [9:0]n45;
    
    wire n6689;
    wire [9:0]r_Clock_Count;   // src/uart_rx.v(32[17:30])
    
    wire n6680, n4335, n10278, n151;
    wire [2:0]r_Bit_Index;   // src/uart_rx.v(33[17:28])
    
    wire n10320, n4367, n5863, n10085, n10084, n10083, n13, n125, 
        n10082, n10081, n10080, n10079;
    wire [2:0]n340;
    
    wire n4691, n149, n6, n140, n8, n4_adj_1186, n10078, n6714, 
        n6699, n10077;
    
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n3), .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(SLM_CLK_c), .D(r_Rx_Data_R));   // src/uart_rx.v(41[10] 45[8])
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_765[2]), .I2(GND_net), 
            .I3(GND_net), .O(n55));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5340_4_lut (.I0(r_Rx_Data), .I1(n55), .I2(r_SM_Main[1]), 
            .I3(n145), .O(n3_adj_1182));   // src/uart_rx.v(36[17:26])
    defparam i5340_4_lut.LUT_INIT = 16'h3530;
    SB_DFFESR r_Clock_Count_1191__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n6689), .D(n45[0]), .R(n6680));   // src/uart_rx.v(120[34:51])
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_765[2]), 
            .I3(r_SM_Main[0]), .O(n4335));
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n4335), 
            .I3(debug_led3), .O(n10278));
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i1_2_lut_3_lut (.I0(r_SM_Main[0]), .I1(n151), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n4248));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_33 (.I0(r_SM_Main[0]), .I1(n151), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n4253));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_adj_33.LUT_INIT = 16'hbfbf;
    SB_LUT4 equal_140_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // src/uart_rx.v(97[17:39])
    defparam equal_140_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_137_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // src/uart_rx.v(97[17:39])
    defparam equal_137_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i5971_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n7347));
    defparam i5971_2_lut.LUT_INIT = 16'h8888;
    SB_DFF r_Rx_Byte_i0 (.Q(pc_data_rx[0]), .C(SLM_CLK_c), .D(n6083));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Rx_DV_52 (.Q(debug_led3), .C(SLM_CLK_c), .E(VCC_net), .D(n10278));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n10320));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_4_lut (.I0(r_SM_Main_2__N_765[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main[2]), .O(n4367));
    defparam i2_4_lut.LUT_INIT = 16'h0023;
    SB_DFF r_Rx_Byte_i7 (.Q(pc_data_rx[7]), .C(SLM_CLK_c), .D(n6067));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(pc_data_rx[6]), .C(SLM_CLK_c), .D(n6066));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(pc_data_rx[5]), .C(SLM_CLK_c), .D(n6064));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(pc_data_rx[4]), .C(SLM_CLK_c), .D(n6063));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(pc_data_rx[3]), .C(SLM_CLK_c), .D(n6062));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(pc_data_rx[2]), .C(SLM_CLK_c), .D(n6060));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i12_3_lut (.I0(n4367), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n10320));   // src/uart_rx.v(36[17:26])
    defparam i12_3_lut.LUT_INIT = 16'h6464;
    SB_LUT4 equal_141_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // src/uart_rx.v(97[17:39])
    defparam equal_141_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[0]), .I1(n151), .I2(n4_adj_2), .I3(r_Bit_Index[0]), 
            .O(n10211));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(SLM_CLK_c), .D(UART_RX_c));   // src/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Byte_i1 (.Q(pc_data_rx[1]), .C(SLM_CLK_c), .D(n6030));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(n5863));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n3_adj_1182), 
            .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_1191_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n10085), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1191_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n10084), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Clock_Count_1191__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n6689), .D(n45[9]), .R(n6680));   // src/uart_rx.v(120[34:51])
    SB_CARRY r_Clock_Count_1191_add_4_10 (.CI(n10084), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n10085));
    SB_LUT4 r_Clock_Count_1191_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n10083), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Clock_Count_1191__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n6689), .D(n45[8]), .R(n6680));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1191__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n6689), .D(n45[7]), .R(n6680));   // src/uart_rx.v(120[34:51])
    SB_CARRY r_Clock_Count_1191_add_4_9 (.CI(n10083), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n10084));
    SB_LUT4 i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main[0]), .I2(n13), .I3(GND_net), 
            .O(n125));   // src/uart_rx.v(30[17:26])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i10207_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[2]), .I2(n145), 
            .I3(r_SM_Main[1]), .O(n6689));
    defparam i10207_4_lut.LUT_INIT = 16'h3313;
    SB_DFFESR r_Clock_Count_1191__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n6689), .D(n45[6]), .R(n6680));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1191__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n6689), .D(n45[5]), .R(n6680));   // src/uart_rx.v(120[34:51])
    SB_LUT4 r_Clock_Count_1191_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n10082), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1191_add_4_8 (.CI(n10082), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n10083));
    SB_DFFESR r_Clock_Count_1191__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n6689), .D(n45[4]), .R(n6680));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1191__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n6689), .D(n45[3]), .R(n6680));   // src/uart_rx.v(120[34:51])
    SB_LUT4 r_Clock_Count_1191_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n10081), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_34 (.I0(r_SM_Main[0]), .I1(n151), .I2(GND_net), 
            .I3(GND_net), .O(n5863));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_34.LUT_INIT = 16'h8888;
    SB_DFFESR r_Clock_Count_1191__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n6689), .D(n45[2]), .R(n6680));   // src/uart_rx.v(120[34:51])
    SB_CARRY r_Clock_Count_1191_add_4_7 (.CI(n10081), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n10082));
    SB_DFFESR r_Clock_Count_1191__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n6689), .D(n45[1]), .R(n6680));   // src/uart_rx.v(120[34:51])
    SB_LUT4 r_Clock_Count_1191_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n10080), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1191_add_4_6 (.CI(n10080), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n10081));
    SB_LUT4 r_Clock_Count_1191_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n10079), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(SLM_CLK_c), .E(n4367), 
            .D(n340[1]), .R(n4691));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(SLM_CLK_c), .E(n4367), 
            .D(n340[2]), .R(n4691));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1350_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n340[2]));   // src/uart_rx.v(49[10] 144[8])
    defparam i1350_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n149));   // src/uart_rx.v(49[10] 144[8])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY r_Clock_Count_1191_add_4_5 (.CI(n10079), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n10080));
    SB_LUT4 i1_2_lut_adj_35 (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // src/uart_rx.v(32[17:30])
    defparam i1_2_lut_adj_35.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[9]), 
            .I3(n6), .O(n140));   // src/uart_rx.v(32[17:30])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_36 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), 
            .I2(r_Clock_Count[3]), .I3(r_Clock_Count[4]), .O(n8));
    defparam i3_4_lut_adj_36.LUT_INIT = 16'hffdf;
    SB_LUT4 i4_3_lut (.I0(n140), .I1(n8), .I2(r_Clock_Count[2]), .I3(GND_net), 
            .O(n13));
    defparam i4_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_37 (.I0(r_SM_Main[0]), .I1(n13), .I2(GND_net), 
            .I3(GND_net), .O(n145));   // src/uart_rx.v(36[17:26])
    defparam i1_2_lut_adj_37.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_adj_38 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), 
            .I2(r_Clock_Count[1]), .I3(GND_net), .O(n4_adj_1186));   // src/uart_rx.v(118[17:47])
    defparam i1_3_lut_adj_38.LUT_INIT = 16'hecec;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[4]), .I1(n140), .I2(r_Clock_Count[3]), 
            .I3(n4_adj_1186), .O(r_SM_Main_2__N_765[2]));   // src/uart_rx.v(32[17:30])
    defparam i1_4_lut.LUT_INIT = 16'heeec;
    SB_LUT4 r_Clock_Count_1191_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n10078), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5332_3_lut (.I0(n149), .I1(r_SM_Main[0]), .I2(r_SM_Main_2__N_765[2]), 
            .I3(GND_net), .O(n6714));   // src/uart_rx.v(36[17:26])
    defparam i5332_3_lut.LUT_INIT = 16'h2c2c;
    SB_CARRY r_Clock_Count_1191_add_4_4 (.CI(n10078), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n10079));
    SB_LUT4 i5333_3_lut (.I0(n6699), .I1(n6714), .I2(r_SM_Main[1]), .I3(GND_net), 
            .O(n3));   // src/uart_rx.v(36[17:26])
    defparam i5333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_1191_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n10077), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1191_add_4_3 (.CI(n10077), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n10078));
    SB_LUT4 i5298_4_lut_4_lut (.I0(r_SM_Main_2__N_765[2]), .I1(r_SM_Main[2]), 
            .I2(n125), .I3(r_SM_Main[1]), .O(n6680));   // src/uart_rx.v(49[10] 144[8])
    defparam i5298_4_lut_4_lut.LUT_INIT = 16'h2203;
    SB_LUT4 r_Clock_Count_1191_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1191_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_39 (.I0(r_SM_Main_2__N_765[2]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n151));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_adj_39.LUT_INIT = 16'h2020;
    SB_CARRY r_Clock_Count_1191_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n10077));
    SB_LUT4 i1343_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n340[1]));   // src/uart_rx.v(102[36:51])
    defparam i1343_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3308_3_lut (.I0(n4367), .I1(r_SM_Main[1]), .I2(n149), .I3(GND_net), 
            .O(n4691));   // src/uart_rx.v(49[10] 144[8])
    defparam i3308_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i5317_4_lut_3_lut (.I0(r_SM_Main[0]), .I1(n13), .I2(r_Rx_Data), 
            .I3(GND_net), .O(n6699));   // src/uart_rx.v(30[17:26])
    defparam i5317_4_lut_3_lut.LUT_INIT = 16'h8d8d;
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word
//

module FIFO_Quad_Word (rd_fifo_en_w, \mem_LUT.data_raw_r[7] , SLM_CLK_c, 
            \mem_LUT.data_raw_r[6] , rd_addr_r, \rd_addr_p1_w[2] , GND_net, 
            \mem_LUT.data_raw_r[5] , n13895, \mem_LUT.data_raw_r[0] , 
            \mem_LUT.data_raw_r[4] , \mem_LUT.data_raw_r[3] , reset_all_w, 
            n8, wr_addr_r, \mem_LUT.data_raw_r[2] , \mem_LUT.data_raw_r[1] , 
            n4941, VCC_net, n4938, rx_buf_byte, n6112, \fifo_temp_output[1] , 
            n10302, is_tx_fifo_full_flag, n6073, \fifo_temp_output[0] , 
            n1, \wr_addr_p1_w[2] , n10098, n5310, \fifo_temp_output[4] , 
            n5313, \fifo_temp_output[5] , n4882, \fifo_temp_output[2] , 
            n4887, \fifo_temp_output[3] , n5534, \fifo_temp_output[6] , 
            n5537, \fifo_temp_output[7] , n10632, is_fifo_empty_flag, 
            n4919, n4922, fifo_write_cmd, wr_fifo_en_w, n4878, rd_fifo_en_prev_r, 
            fifo_read_cmd) /* synthesis syn_module_defined=1 */ ;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[7] ;
    input SLM_CLK_c;
    output \mem_LUT.data_raw_r[6] ;
    output [2:0]rd_addr_r;
    output \rd_addr_p1_w[2] ;
    input GND_net;
    output \mem_LUT.data_raw_r[5] ;
    output n13895;
    output \mem_LUT.data_raw_r[0] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[3] ;
    input reset_all_w;
    input n8;
    output [2:0]wr_addr_r;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[1] ;
    input n4941;
    input VCC_net;
    input n4938;
    input [7:0]rx_buf_byte;
    input n6112;
    output \fifo_temp_output[1] ;
    input n10302;
    output is_tx_fifo_full_flag;
    input n6073;
    output \fifo_temp_output[0] ;
    output n1;
    output \wr_addr_p1_w[2] ;
    output n10098;
    input n5310;
    output \fifo_temp_output[4] ;
    input n5313;
    output \fifo_temp_output[5] ;
    input n4882;
    output \fifo_temp_output[2] ;
    input n4887;
    output \fifo_temp_output[3] ;
    input n5534;
    output \fifo_temp_output[6] ;
    input n5537;
    output \fifo_temp_output[7] ;
    input n10632;
    output is_fifo_empty_flag;
    input n4919;
    input n4922;
    input fifo_write_cmd;
    output wr_fifo_en_w;
    input n4878;
    output rd_fifo_en_prev_r;
    input fifo_read_cmd;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2 lscc_fifo_inst (.rd_fifo_en_w(rd_fifo_en_w), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r[7] ), .SLM_CLK_c(SLM_CLK_c), 
            .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r[6] ), .rd_addr_r({rd_addr_r}), 
            .\rd_addr_p1_w[2] (\rd_addr_p1_w[2] ), .GND_net(GND_net), .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r[5] ), 
            .n13895(n13895), .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r[0] ), 
            .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r[4] ), .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r[3] ), 
            .reset_all_w(reset_all_w), .n8(n8), .wr_addr_r({wr_addr_r}), 
            .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r[2] ), .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r[1] ), 
            .n4941(n4941), .VCC_net(VCC_net), .n4938(n4938), .rx_buf_byte({rx_buf_byte}), 
            .n6112(n6112), .\fifo_temp_output[1] (\fifo_temp_output[1] ), 
            .n10302(n10302), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .n6073(n6073), .\fifo_temp_output[0] (\fifo_temp_output[0] ), 
            .n1(n1), .\wr_addr_p1_w[2] (\wr_addr_p1_w[2] ), .n10098(n10098), 
            .n5310(n5310), .\fifo_temp_output[4] (\fifo_temp_output[4] ), 
            .n5313(n5313), .\fifo_temp_output[5] (\fifo_temp_output[5] ), 
            .n4882(n4882), .\fifo_temp_output[2] (\fifo_temp_output[2] ), 
            .n4887(n4887), .\fifo_temp_output[3] (\fifo_temp_output[3] ), 
            .n5534(n5534), .\fifo_temp_output[6] (\fifo_temp_output[6] ), 
            .n5537(n5537), .\fifo_temp_output[7] (\fifo_temp_output[7] ), 
            .n10632(n10632), .is_fifo_empty_flag(is_fifo_empty_flag), .n4919(n4919), 
            .n4922(n4922), .fifo_write_cmd(fifo_write_cmd), .wr_fifo_en_w(wr_fifo_en_w), 
            .n4878(n4878), .rd_fifo_en_prev_r(rd_fifo_en_prev_r), .fifo_read_cmd(fifo_read_cmd)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_quad_word_mod.v(20[37:380])
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2
//

module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2 (rd_fifo_en_w, 
            \mem_LUT.data_raw_r[7] , SLM_CLK_c, \mem_LUT.data_raw_r[6] , 
            rd_addr_r, \rd_addr_p1_w[2] , GND_net, \mem_LUT.data_raw_r[5] , 
            n13895, \mem_LUT.data_raw_r[0] , \mem_LUT.data_raw_r[4] , 
            \mem_LUT.data_raw_r[3] , reset_all_w, n8, wr_addr_r, \mem_LUT.data_raw_r[2] , 
            \mem_LUT.data_raw_r[1] , n4941, VCC_net, n4938, rx_buf_byte, 
            n6112, \fifo_temp_output[1] , n10302, is_tx_fifo_full_flag, 
            n6073, \fifo_temp_output[0] , n1, \wr_addr_p1_w[2] , n10098, 
            n5310, \fifo_temp_output[4] , n5313, \fifo_temp_output[5] , 
            n4882, \fifo_temp_output[2] , n4887, \fifo_temp_output[3] , 
            n5534, \fifo_temp_output[6] , n5537, \fifo_temp_output[7] , 
            n10632, is_fifo_empty_flag, n4919, n4922, fifo_write_cmd, 
            wr_fifo_en_w, n4878, rd_fifo_en_prev_r, fifo_read_cmd) /* synthesis syn_module_defined=1 */ ;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[7] ;
    input SLM_CLK_c;
    output \mem_LUT.data_raw_r[6] ;
    output [2:0]rd_addr_r;
    output \rd_addr_p1_w[2] ;
    input GND_net;
    output \mem_LUT.data_raw_r[5] ;
    output n13895;
    output \mem_LUT.data_raw_r[0] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[3] ;
    input reset_all_w;
    input n8;
    output [2:0]wr_addr_r;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[1] ;
    input n4941;
    input VCC_net;
    input n4938;
    input [7:0]rx_buf_byte;
    input n6112;
    output \fifo_temp_output[1] ;
    input n10302;
    output is_tx_fifo_full_flag;
    input n6073;
    output \fifo_temp_output[0] ;
    output n1;
    output \wr_addr_p1_w[2] ;
    output n10098;
    input n5310;
    output \fifo_temp_output[4] ;
    input n5313;
    output \fifo_temp_output[5] ;
    input n4882;
    output \fifo_temp_output[2] ;
    input n4887;
    output \fifo_temp_output[3] ;
    input n5534;
    output \fifo_temp_output[6] ;
    input n5537;
    output \fifo_temp_output[7] ;
    input n10632;
    output is_fifo_empty_flag;
    input n4919;
    input n4922;
    input fifo_write_cmd;
    output wr_fifo_en_w;
    input n4878;
    output rd_fifo_en_prev_r;
    input fifo_read_cmd;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [31:0]\mem_LUT.data_raw_r_31__N_1084 ;
    wire [2:0]n12;
    
    wire \mem_LUT.mem_2_4 , \mem_LUT.mem_3_4 , n12243, \mem_LUT.mem_1_4 , 
        \mem_LUT.mem_0_4 , \mem_LUT.mem_2_3 , \mem_LUT.mem_3_3 , n12237, 
        \mem_LUT.mem_1_3 , \mem_LUT.mem_0_3 , n3, \mem_LUT.mem_3_7 , 
        n6057, \mem_LUT.mem_3_6 , n6056, \mem_LUT.mem_3_5 , n6055, 
        n6054, n6053, \mem_LUT.mem_3_2 , n6052, \mem_LUT.mem_3_1 , 
        n6051, \mem_LUT.mem_3_0 , n6050, \mem_LUT.mem_2_2 , n12225, 
        \mem_LUT.mem_2_7 , n12333, \mem_LUT.mem_1_7 , \mem_LUT.mem_0_7 , 
        n2, n6042, n6041, \mem_LUT.mem_2_6 , n6040, \mem_LUT.mem_2_5 , 
        n6039, n6038, n6037, n6036, \mem_LUT.mem_2_1 , n6035, \mem_LUT.mem_2_0 , 
        n12321, \mem_LUT.mem_1_6 , \mem_LUT.mem_0_6 , n6029, n6028, 
        n6027, \mem_LUT.mem_1_5 , n6026, n6025, n6024, \mem_LUT.mem_1_2 , 
        n6023, \mem_LUT.mem_1_1 , n6022, \mem_LUT.mem_1_0 , n6021, 
        n6020, n6019, \mem_LUT.mem_0_5 , n6018, n12315, n6017, n6016, 
        \mem_LUT.mem_0_2 , n6015, \mem_LUT.mem_0_1 , n6014, \mem_LUT.mem_0_0 , 
        n4, n12183, n12177;
    
    SB_DFFE \mem_LUT.data_raw_r__i8  (.Q(\mem_LUT.data_raw_r[7] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [7]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i7  (.Q(\mem_LUT.data_raw_r[6] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [6]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 i1416_3_lut (.I0(rd_addr_r[2]), .I1(rd_addr_r[1]), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(\rd_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1416_3_lut.LUT_INIT = 16'h6a6a;
    SB_DFFE \mem_LUT.data_raw_r__i6  (.Q(\mem_LUT.data_raw_r[5] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [5]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 i1409_rep_148_2_lut (.I0(rd_addr_r[1]), .I1(rd_addr_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n13895));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1409_rep_148_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE \mem_LUT.data_raw_r__i1  (.Q(\mem_LUT.data_raw_r[0] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [0]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i5  (.Q(\mem_LUT.data_raw_r[4] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [4]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i4  (.Q(\mem_LUT.data_raw_r[3] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [3]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFSR rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n12[0]), 
            .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFSR wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(SLM_CLK_c), .D(n8), .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFE \mem_LUT.data_raw_r__i3  (.Q(\mem_LUT.data_raw_r[2] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [2]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i2  (.Q(\mem_LUT.data_raw_r[1] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1084 [1]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10430 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_4 ), 
            .I2(\mem_LUT.mem_3_4 ), .I3(rd_addr_r[1]), .O(n12243));
    defparam rd_addr_r_0__bdd_4_lut_10430.LUT_INIT = 16'he4aa;
    SB_LUT4 n12243_bdd_4_lut (.I0(n12243), .I1(\mem_LUT.mem_1_4 ), .I2(\mem_LUT.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [4]));
    defparam n12243_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n4941));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFE wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n4938));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10370 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_3 ), 
            .I2(\mem_LUT.mem_3_3 ), .I3(rd_addr_r[1]), .O(n12237));
    defparam rd_addr_r_0__bdd_4_lut_10370.LUT_INIT = 16'he4aa;
    SB_LUT4 n12237_bdd_4_lut (.I0(n12237), .I1(\mem_LUT.mem_1_3 ), .I2(\mem_LUT.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [3]));
    defparam n12237_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4674_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_3_7 ), .O(n6057));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4674_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4673_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_3_6 ), .O(n6056));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4673_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4672_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_3_5 ), .O(n6055));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4672_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4671_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_3_4 ), .O(n6054));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4671_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4670_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_3_3 ), .O(n6053));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4670_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE \mem_LUT.data_buff_r__i1  (.Q(\fifo_temp_output[1] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6112));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 i4669_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_3_2 ), .O(n6052));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4669_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4668_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_3_1 ), .O(n6051));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4668_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4667_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_3_0 ), .O(n6050));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4667_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10365 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_2 ), 
            .I2(\mem_LUT.mem_3_2 ), .I3(rd_addr_r[1]), .O(n12225));
    defparam rd_addr_r_0__bdd_4_lut_10365.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_7 ), 
            .I2(\mem_LUT.mem_3_7 ), .I3(rd_addr_r[1]), .O(n12333));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n12333_bdd_4_lut (.I0(n12333), .I1(\mem_LUT.mem_1_7 ), .I2(\mem_LUT.mem_0_7 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [7]));
    defparam n12333_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE full_r_84 (.Q(is_tx_fifo_full_flag), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n10302));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFE \mem_LUT.data_buff_r__i0  (.Q(\fifo_temp_output[0] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6073));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF i347_348 (.Q(\mem_LUT.mem_3_7 ), .C(SLM_CLK_c), .D(n6057));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i344_345 (.Q(\mem_LUT.mem_3_6 ), .C(SLM_CLK_c), .D(n6056));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 wr_addr_r_1__I_0_i1_2_lut (.I0(wr_addr_r[0]), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(GND_net), .O(n1));   // src/fifo_quad_word_mod.v(115[26:58])
    defparam wr_addr_r_1__I_0_i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF i341_342 (.Q(\mem_LUT.mem_3_5 ), .C(SLM_CLK_c), .D(n6055));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 i1_4_lut (.I0(n1), .I1(\wr_addr_p1_w[2] ), .I2(n2), .I3(rd_addr_r[2]), 
            .O(n10098));
    defparam i1_4_lut.LUT_INIT = 16'h0208;
    SB_DFF i338_339 (.Q(\mem_LUT.mem_3_4 ), .C(SLM_CLK_c), .D(n6054));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i335_336 (.Q(\mem_LUT.mem_3_3 ), .C(SLM_CLK_c), .D(n6053));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i332_333 (.Q(\mem_LUT.mem_3_2 ), .C(SLM_CLK_c), .D(n6052));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i329_330 (.Q(\mem_LUT.mem_3_1 ), .C(SLM_CLK_c), .D(n6051));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i326_327 (.Q(\mem_LUT.mem_3_0 ), .C(SLM_CLK_c), .D(n6050));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i251_252 (.Q(\mem_LUT.mem_2_7 ), .C(SLM_CLK_c), .D(n6042));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i248_249 (.Q(\mem_LUT.mem_2_6 ), .C(SLM_CLK_c), .D(n6041));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i245_246 (.Q(\mem_LUT.mem_2_5 ), .C(SLM_CLK_c), .D(n6040));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i242_243 (.Q(\mem_LUT.mem_2_4 ), .C(SLM_CLK_c), .D(n6039));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i239_240 (.Q(\mem_LUT.mem_2_3 ), .C(SLM_CLK_c), .D(n6038));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i236_237 (.Q(\mem_LUT.mem_2_2 ), .C(SLM_CLK_c), .D(n6037));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i233_234 (.Q(\mem_LUT.mem_2_1 ), .C(SLM_CLK_c), .D(n6036));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i230_231 (.Q(\mem_LUT.mem_2_0 ), .C(SLM_CLK_c), .D(n6035));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10445 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_6 ), 
            .I2(\mem_LUT.mem_3_6 ), .I3(rd_addr_r[1]), .O(n12321));
    defparam rd_addr_r_0__bdd_4_lut_10445.LUT_INIT = 16'he4aa;
    SB_LUT4 n12321_bdd_4_lut (.I0(n12321), .I1(\mem_LUT.mem_1_6 ), .I2(\mem_LUT.mem_0_6 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [6]));
    defparam n12321_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i155_156 (.Q(\mem_LUT.mem_1_7 ), .C(SLM_CLK_c), .D(n6029));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i152_153 (.Q(\mem_LUT.mem_1_6 ), .C(SLM_CLK_c), .D(n6028));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i149_150 (.Q(\mem_LUT.mem_1_5 ), .C(SLM_CLK_c), .D(n6027));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i146_147 (.Q(\mem_LUT.mem_1_4 ), .C(SLM_CLK_c), .D(n6026));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i143_144 (.Q(\mem_LUT.mem_1_3 ), .C(SLM_CLK_c), .D(n6025));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i140_141 (.Q(\mem_LUT.mem_1_2 ), .C(SLM_CLK_c), .D(n6024));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i137_138 (.Q(\mem_LUT.mem_1_1 ), .C(SLM_CLK_c), .D(n6023));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i134_135 (.Q(\mem_LUT.mem_1_0 ), .C(SLM_CLK_c), .D(n6022));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i59_60 (.Q(\mem_LUT.mem_0_7 ), .C(SLM_CLK_c), .D(n6021));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i56_57 (.Q(\mem_LUT.mem_0_6 ), .C(SLM_CLK_c), .D(n6020));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i53_54 (.Q(\mem_LUT.mem_0_5 ), .C(SLM_CLK_c), .D(n6019));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i50_51 (.Q(\mem_LUT.mem_0_4 ), .C(SLM_CLK_c), .D(n6018));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10435 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_5 ), 
            .I2(\mem_LUT.mem_3_5 ), .I3(rd_addr_r[1]), .O(n12315));
    defparam rd_addr_r_0__bdd_4_lut_10435.LUT_INIT = 16'he4aa;
    SB_LUT4 n12315_bdd_4_lut (.I0(n12315), .I1(\mem_LUT.mem_1_5 ), .I2(\mem_LUT.mem_0_5 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [5]));
    defparam n12315_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i47_48 (.Q(\mem_LUT.mem_0_3 ), .C(SLM_CLK_c), .D(n6017));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i44_45 (.Q(\mem_LUT.mem_0_2 ), .C(SLM_CLK_c), .D(n6016));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i41_42 (.Q(\mem_LUT.mem_0_1 ), .C(SLM_CLK_c), .D(n6015));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i38_39 (.Q(\mem_LUT.mem_0_0 ), .C(SLM_CLK_c), .D(n6014));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 n12225_bdd_4_lut (.I0(n12225), .I1(\mem_LUT.mem_1_2 ), .I2(\mem_LUT.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [2]));
    defparam n12225_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF \mem_LUT.data_buff_r__i4  (.Q(\fifo_temp_output[4] ), .C(SLM_CLK_c), 
           .D(n5310));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i5  (.Q(\fifo_temp_output[5] ), .C(SLM_CLK_c), 
           .D(n5313));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i2  (.Q(\fifo_temp_output[2] ), .C(SLM_CLK_c), 
           .D(n4882));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i3  (.Q(\fifo_temp_output[3] ), .C(SLM_CLK_c), 
           .D(n4887));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i6  (.Q(\fifo_temp_output[6] ), .C(SLM_CLK_c), 
           .D(n5534));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i7  (.Q(\fifo_temp_output[7] ), .C(SLM_CLK_c), 
           .D(n5537));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF empty_r_85 (.Q(is_fifo_empty_flag), .C(SLM_CLK_c), .D(n10632));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i1394_3_lut (.I0(wr_addr_r[2]), .I1(wr_addr_r[1]), .I2(wr_addr_r[0]), 
            .I3(GND_net), .O(\wr_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam i1394_3_lut.LUT_INIT = 16'h6a6a;
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(n4919));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .D(n4922));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i4659_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_2_7 ), .O(n6042));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4659_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4658_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_2_6 ), .O(n6041));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4658_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4657_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_2_5 ), .O(n6040));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4657_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4656_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_2_4 ), .O(n6039));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4656_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4655_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_2_3 ), .O(n6038));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4655_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4654_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_2_2 ), .O(n6037));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4654_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4653_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_2_1 ), .O(n6036));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4653_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4652_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_2_0 ), .O(n6035));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4652_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_en_i_I_0_2_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(GND_net), .I3(GND_net), .O(wr_fifo_en_w));   // src/fifo_quad_word_mod.v(103[21:60])
    defparam wr_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4646_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_1_7 ), .O(n6029));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4646_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4645_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_1_6 ), .O(n6028));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4645_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4644_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_1_5 ), .O(n6027));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4644_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4643_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_1_4 ), .O(n6026));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4643_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4642_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_1_3 ), .O(n6025));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4642_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4641_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_1_2 ), .O(n6024));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4641_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF rd_fifo_en_prev_r_86 (.Q(rd_fifo_en_prev_r), .C(SLM_CLK_c), .D(n4878));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    SB_LUT4 i4640_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_1_1 ), .O(n6023));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4640_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_en_i_I_0_2_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(GND_net), .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_quad_word_mod.v(62[29:51])
    defparam rd_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4639_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_1_0 ), .O(n6022));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4639_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4638_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_0_7 ), .O(n6021));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4638_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4637_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_0_6 ), .O(n6020));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4637_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4636_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_0_5 ), .O(n6019));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4636_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4635_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_0_4 ), .O(n6018));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4635_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4634_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_0_3 ), .O(n6017));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4634_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4633_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_0_2 ), .O(n6016));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4633_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4632_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_0_1 ), .O(n6015));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4632_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4631_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_0_0 ), .O(n6014));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4631_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10355 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_1 ), 
            .I2(\mem_LUT.mem_3_1 ), .I3(rd_addr_r[1]), .O(n12183));
    defparam rd_addr_r_0__bdd_4_lut_10355.LUT_INIT = 16'he4aa;
    SB_LUT4 n12183_bdd_4_lut (.I0(n12183), .I1(\mem_LUT.mem_1_1 ), .I2(\mem_LUT.mem_0_1 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [1]));
    defparam n12183_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10321 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_0 ), 
            .I2(\mem_LUT.mem_3_0 ), .I3(rd_addr_r[1]), .O(n12177));
    defparam rd_addr_r_0__bdd_4_lut_10321.LUT_INIT = 16'he4aa;
    SB_LUT4 n12177_bdd_4_lut (.I0(n12177), .I1(\mem_LUT.mem_1_0 ), .I2(\mem_LUT.mem_0_0 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1084 [0]));
    defparam n12177_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_p1_w_1__I_0_i2_2_lut_3_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[0]), 
            .I2(rd_addr_r[1]), .I3(GND_net), .O(n2));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam wr_addr_p1_w_1__I_0_i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1603_2_lut_4_lut (.I0(rd_addr_r[0]), .I1(fifo_read_cmd), .I2(is_fifo_empty_flag), 
            .I3(reset_all_w), .O(n12[0]));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1603_2_lut_4_lut.LUT_INIT = 16'h55a6;
    SB_LUT4 EnabledDecoder_2_i3_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n3));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i3_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i4_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n4));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i4_2_lut_3_lut.LUT_INIT = 16'h0202;
    
endmodule
//
// Verilog Description of module clock
//

module clock (GND_net, VCC_net, ICE_SYSCLK_c, pll_clk_unbuf) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    input ICE_SYSCLK_c;
    output pll_clk_unbuf;
    
    
    SB_PLL40_CORE pll_config (.REFERENCECLK(ICE_SYSCLK_c), .PLLOUTGLOBAL(pll_clk_unbuf), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=14, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/top.v(222[7] 228[3])
    defparam pll_config.FEEDBACK_PATH = "SIMPLE";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll_config.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll_config.FDA_FEEDBACK = 0;
    defparam pll_config.FDA_RELATIVE = 0;
    defparam pll_config.PLLOUT_SELECT = "GENCLK";
    defparam pll_config.DIVR = 4'b0001;
    defparam pll_config.DIVF = 7'b1010010;
    defparam pll_config.DIVQ = 3'b100;
    defparam pll_config.FILTER_RANGE = 3'b001;
    defparam pll_config.ENABLE_ICEGATE = 1'b0;
    defparam pll_config.TEST_MODE = 1'b0;
    defparam pll_config.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module usb3_if
//

module usb3_if (reset_per_frame, reset_per_frame_latched, SLM_CLK_c, write_to_dc32_fifo_latched_N_425, 
            n2352, DEBUG_3_c, DEBUG_2_c, FIFO_CLK_c, \dc32_fifo_data_in[0] , 
            DEBUG_5_c, buffer_switch_done, buffer_switch_done_latched, 
            n571, n575, GND_net, VCC_net, FT_OE_N_420, n4911, n4910, 
            n4907, dc32_fifo_almost_full, FT_OE_c, FIFO_D15_c_15, FIFO_D14_c_14, 
            FIFO_D13_c_13, FIFO_D12_c_12, FIFO_D11_c_11, FIFO_D10_c_10, 
            FIFO_D9_c_9, FIFO_D8_c_8, FIFO_D7_c_7, FIFO_D6_c_6, FIFO_D5_c_5, 
            FIFO_D4_c_4, FIFO_D3_c_3, FIFO_D2_c_2, FIFO_D1_c_1, \dc32_fifo_data_in[15] , 
            \dc32_fifo_data_in[14] , \dc32_fifo_data_in[13] , \dc32_fifo_data_in[12] , 
            \dc32_fifo_data_in[11] , \dc32_fifo_data_in[10] , \dc32_fifo_data_in[9] , 
            \dc32_fifo_data_in[8] , \dc32_fifo_data_in[7] , \dc32_fifo_data_in[6] , 
            \dc32_fifo_data_in[5] , \dc32_fifo_data_in[4] , \dc32_fifo_data_in[3] , 
            \dc32_fifo_data_in[2] , \dc32_fifo_data_in[1] , DEBUG_1_c_c) /* synthesis syn_module_defined=1 */ ;
    input reset_per_frame;
    output reset_per_frame_latched;
    input SLM_CLK_c;
    input write_to_dc32_fifo_latched_N_425;
    output n2352;
    input DEBUG_3_c;
    output DEBUG_2_c;
    input FIFO_CLK_c;
    output \dc32_fifo_data_in[0] ;
    output DEBUG_5_c;
    input buffer_switch_done;
    output buffer_switch_done_latched;
    output n571;
    output n575;
    input GND_net;
    input VCC_net;
    input FT_OE_N_420;
    input n4911;
    input n4910;
    input n4907;
    input dc32_fifo_almost_full;
    output FT_OE_c;
    input FIFO_D15_c_15;
    input FIFO_D14_c_14;
    input FIFO_D13_c_13;
    input FIFO_D12_c_12;
    input FIFO_D11_c_11;
    input FIFO_D10_c_10;
    input FIFO_D9_c_9;
    input FIFO_D8_c_8;
    input FIFO_D7_c_7;
    input FIFO_D6_c_6;
    input FIFO_D5_c_5;
    input FIFO_D4_c_4;
    input FIFO_D3_c_3;
    input FIFO_D2_c_2;
    input FIFO_D1_c_1;
    output \dc32_fifo_data_in[15] ;
    output \dc32_fifo_data_in[14] ;
    output \dc32_fifo_data_in[13] ;
    output \dc32_fifo_data_in[12] ;
    output \dc32_fifo_data_in[11] ;
    output \dc32_fifo_data_in[10] ;
    output \dc32_fifo_data_in[9] ;
    output \dc32_fifo_data_in[8] ;
    output \dc32_fifo_data_in[7] ;
    output \dc32_fifo_data_in[6] ;
    output \dc32_fifo_data_in[5] ;
    output \dc32_fifo_data_in[4] ;
    output \dc32_fifo_data_in[3] ;
    output \dc32_fifo_data_in[2] ;
    output \dc32_fifo_data_in[1] ;
    input DEBUG_1_c_c;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    
    wire n613;
    wire [15:0]n562;
    
    wire dc32_fifo_empty_latched, FT_RD_N_422;
    wire [31:0]dc32_fifo_data_in_latched;   // src/usb3_if.v(68[12:37])
    
    wire write_to_dc32_fifo_latched, n3004, n618, n3002, n3014, n608, 
        n2992, n10154;
    wire [3:0]state_timeout_counter;   // src/usb3_if.v(66[11:32])
    
    wire n3942, n3938, n524, n606, n2415, n2408;
    wire [10:0]num_lines_clocked_out_10__N_371;
    wire [10:0]num_lines_clocked_out;   // src/usb3_if.v(65[12:33])
    
    wire n10027, n4181, FT_OE_N_419, n10028;
    wire [10:0]n1;
    
    wire n10036, n10035, n10034, n10033, n10032, n10031, n10030, 
        n10029, n520, n551, n4, n21, n4224, n18, n16, n20, 
        n522, n2400, n4310, n4703, n2401, n2402, n2983, n4486, 
        n2399, n2390, n3940, n10629, n2266, n11921, n11881;
    
    SB_DFF reset_per_frame_latched_89 (.Q(reset_per_frame_latched), .C(SLM_CLK_c), 
           .D(reset_per_frame));   // src/usb3_if.v(72[8] 85[4])
    SB_LUT4 i1116_4_lut (.I0(n613), .I1(reset_per_frame_latched), .I2(write_to_dc32_fifo_latched_N_425), 
            .I3(n562[5]), .O(n2352));   // src/usb3_if.v(97[10] 190[8])
    defparam i1116_4_lut.LUT_INIT = 16'hcfdd;
    SB_DFF dc32_fifo_empty_latched_90 (.Q(dc32_fifo_empty_latched), .C(SLM_CLK_c), 
           .D(DEBUG_3_c));   // src/usb3_if.v(72[8] 85[4])
    SB_DFFSS FT_RD_92 (.Q(DEBUG_2_c), .C(FIFO_CLK_c), .D(FT_RD_N_422), 
            .S(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFN dc32_fifo_data_in_i1 (.Q(\dc32_fifo_data_in[0] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[0]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN write_to_dc32_fifo_99 (.Q(DEBUG_5_c), .C(FIFO_CLK_c), .D(write_to_dc32_fifo_latched));   // src/usb3_if.v(194[8] 197[4])
    SB_DFF buffer_switch_done_latched_88 (.Q(buffer_switch_done_latched), 
           .C(SLM_CLK_c), .D(buffer_switch_done));   // src/usb3_if.v(72[8] 85[4])
    SB_DFFSS state_FSM_i1 (.Q(n562[0]), .C(FIFO_CLK_c), .D(n3004), .S(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_DFFSR state_FSM_i8 (.Q(n571), .C(FIFO_CLK_c), .D(n618), .R(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_DFFSR state_FSM_i7 (.Q(n562[6]), .C(FIFO_CLK_c), .D(n3002), .R(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_DFFSR state_FSM_i6 (.Q(n562[5]), .C(FIFO_CLK_c), .D(n3014), .R(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_DFFSR state_FSM_i4 (.Q(n575), .C(FIFO_CLK_c), .D(n608), .R(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_DFFSR state_FSM_i3 (.Q(n562[2]), .C(FIFO_CLK_c), .D(n2992), .R(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_DFFSR state_FSM_i2 (.Q(n562[1]), .C(FIFO_CLK_c), .D(n10154), .R(reset_per_frame_latched));   // src/usb3_if.v(98[9] 189[16])
    SB_LUT4 i1_3_lut_4_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(state_timeout_counter[2]), .I3(state_timeout_counter[3]), 
            .O(n3942));   // src/usb3_if.v(150[42:69])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h01fe;
    SB_LUT4 i1_2_lut_3_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(state_timeout_counter[2]), .I3(GND_net), .O(n3938));   // src/usb3_if.v(150[42:69])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1e1e;
    SB_LUT4 i1600_3_lut_4_lut (.I0(n562[2]), .I1(n562[0]), .I2(n524), 
            .I3(n606), .O(n2415));   // src/usb3_if.v(98[9] 189[16])
    defparam i1600_3_lut_4_lut.LUT_INIT = 16'h20fd;
    SB_LUT4 i1166_2_lut_3_lut (.I0(n562[2]), .I1(n562[0]), .I2(n524), 
            .I3(GND_net), .O(n2408));   // src/usb3_if.v(98[9] 189[16])
    defparam i1166_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 sub_113_add_2_3_lut (.I0(GND_net), .I1(num_lines_clocked_out[1]), 
            .I2(VCC_net), .I3(n10027), .O(num_lines_clocked_out_10__N_371[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i234_3_lut (.I0(n4181), .I1(FT_OE_N_420), .I2(n562[5]), .I3(GND_net), 
            .O(FT_OE_N_419));   // src/usb3_if.v(98[9] 189[16])
    defparam i234_3_lut.LUT_INIT = 16'hc5c5;
    SB_CARRY sub_113_add_2_3 (.CI(n10027), .I0(num_lines_clocked_out[1]), 
            .I1(VCC_net), .CO(n10028));
    SB_LUT4 sub_113_add_2_2_lut (.I0(GND_net), .I1(num_lines_clocked_out[0]), 
            .I2(n1[0]), .I3(VCC_net), .O(num_lines_clocked_out_10__N_371[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_2 (.CI(VCC_net), .I0(num_lines_clocked_out[0]), 
            .I1(n1[0]), .CO(n10027));
    SB_LUT4 sub_113_add_2_12_lut (.I0(GND_net), .I1(num_lines_clocked_out[10]), 
            .I2(VCC_net), .I3(n10036), .O(num_lines_clocked_out_10__N_371[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_113_add_2_11_lut (.I0(GND_net), .I1(num_lines_clocked_out[9]), 
            .I2(VCC_net), .I3(n10035), .O(num_lines_clocked_out_10__N_371[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_11 (.CI(n10035), .I0(num_lines_clocked_out[9]), 
            .I1(VCC_net), .CO(n10036));
    SB_LUT4 sub_113_add_2_10_lut (.I0(GND_net), .I1(num_lines_clocked_out[8]), 
            .I2(VCC_net), .I3(n10034), .O(num_lines_clocked_out_10__N_371[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_10 (.CI(n10034), .I0(num_lines_clocked_out[8]), 
            .I1(VCC_net), .CO(n10035));
    SB_LUT4 sub_113_add_2_9_lut (.I0(GND_net), .I1(num_lines_clocked_out[7]), 
            .I2(VCC_net), .I3(n10033), .O(num_lines_clocked_out_10__N_371[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_9 (.CI(n10033), .I0(num_lines_clocked_out[7]), 
            .I1(VCC_net), .CO(n10034));
    SB_LUT4 sub_113_add_2_8_lut (.I0(GND_net), .I1(num_lines_clocked_out[6]), 
            .I2(VCC_net), .I3(n10032), .O(num_lines_clocked_out_10__N_371[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_8 (.CI(n10032), .I0(num_lines_clocked_out[6]), 
            .I1(VCC_net), .CO(n10033));
    SB_LUT4 sub_113_add_2_7_lut (.I0(GND_net), .I1(num_lines_clocked_out[5]), 
            .I2(VCC_net), .I3(n10031), .O(num_lines_clocked_out_10__N_371[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_7 (.CI(n10031), .I0(num_lines_clocked_out[5]), 
            .I1(VCC_net), .CO(n10032));
    SB_LUT4 sub_113_add_2_6_lut (.I0(GND_net), .I1(num_lines_clocked_out[4]), 
            .I2(VCC_net), .I3(n10030), .O(num_lines_clocked_out_10__N_371[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_6 (.CI(n10030), .I0(num_lines_clocked_out[4]), 
            .I1(VCC_net), .CO(n10031));
    SB_LUT4 sub_113_add_2_5_lut (.I0(GND_net), .I1(num_lines_clocked_out[3]), 
            .I2(VCC_net), .I3(n10029), .O(num_lines_clocked_out_10__N_371[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_5 (.CI(n10029), .I0(num_lines_clocked_out[3]), 
            .I1(VCC_net), .CO(n10030));
    SB_DFF state_FSM_i5 (.Q(n562[4]), .C(FIFO_CLK_c), .D(n4911));   // src/usb3_if.v(98[9] 189[16])
    SB_DFF state_FSM_i9 (.Q(n562[8]), .C(FIFO_CLK_c), .D(n4910));   // src/usb3_if.v(98[9] 189[16])
    SB_LUT4 sub_113_add_2_4_lut (.I0(GND_net), .I1(num_lines_clocked_out[2]), 
            .I2(VCC_net), .I3(n10028), .O(num_lines_clocked_out_10__N_371[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF dc32_fifo_data_in_latched__i1 (.Q(dc32_fifo_data_in_latched[0]), 
           .C(FIFO_CLK_c), .D(n4907));   // src/usb3_if.v(88[8] 191[4])
    SB_LUT4 i1_4_lut (.I0(n520), .I1(n562[1]), .I2(n562[0]), .I3(n551), 
            .O(n4));   // src/usb3_if.v(98[9] 189[16])
    defparam i1_4_lut.LUT_INIT = 16'heca0;
    SB_LUT4 i2_3_lut (.I0(n21), .I1(n4), .I2(n4224), .I3(GND_net), .O(n10154));   // src/usb3_if.v(98[9] 189[16])
    defparam i2_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i200_2_lut (.I0(dc32_fifo_almost_full), .I1(n562[5]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // src/usb3_if.v(98[9] 189[16])
    defparam i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1626_4_lut (.I0(n562[2]), .I1(n606), .I2(n524), .I3(dc32_fifo_empty_latched), 
            .O(n2992));   // src/usb3_if.v(98[9] 189[16])
    defparam i1626_4_lut.LUT_INIT = 16'hecee;
    SB_DFFESS FT_OE_91 (.Q(FT_OE_c), .C(FIFO_CLK_c), .E(VCC_net), .D(FT_OE_N_419), 
            .S(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i16 (.Q(dc32_fifo_data_in_latched[15]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D15_c_15), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i15 (.Q(dc32_fifo_data_in_latched[14]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D14_c_14), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i14 (.Q(dc32_fifo_data_in_latched[13]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D13_c_13), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i13 (.Q(dc32_fifo_data_in_latched[12]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D12_c_12), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i12 (.Q(dc32_fifo_data_in_latched[11]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D11_c_11), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i11 (.Q(dc32_fifo_data_in_latched[10]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D10_c_10), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i10 (.Q(dc32_fifo_data_in_latched[9]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D9_c_9), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i9 (.Q(dc32_fifo_data_in_latched[8]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D8_c_8), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i8 (.Q(dc32_fifo_data_in_latched[7]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D7_c_7), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i7 (.Q(dc32_fifo_data_in_latched[6]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D6_c_6), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i6 (.Q(dc32_fifo_data_in_latched[5]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D5_c_5), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i5 (.Q(dc32_fifo_data_in_latched[4]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D4_c_4), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i4 (.Q(dc32_fifo_data_in_latched[3]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D3_c_3), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i3 (.Q(dc32_fifo_data_in_latched[2]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D2_c_2), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR dc32_fifo_data_in_latched__i2 (.Q(dc32_fifo_data_in_latched[1]), 
            .C(FIFO_CLK_c), .E(VCC_net), .D(FIFO_D1_c_1), .R(n2352));   // src/usb3_if.v(88[8] 191[4])
    SB_LUT4 i1635_4_lut (.I0(n562[6]), .I1(write_to_dc32_fifo_latched_N_425), 
            .I2(n551), .I3(n562[5]), .O(n3002));   // src/usb3_if.v(98[9] 189[16])
    defparam i1635_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 i212_2_lut (.I0(n551), .I1(n562[6]), .I2(GND_net), .I3(GND_net), 
            .O(n618));   // src/usb3_if.v(98[9] 189[16])
    defparam i212_2_lut.LUT_INIT = 16'h4444;
    SB_DFFN dc32_fifo_data_in_i16 (.Q(\dc32_fifo_data_in[15] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[15]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i15 (.Q(\dc32_fifo_data_in[14] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[14]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i14 (.Q(\dc32_fifo_data_in[13] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[13]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i13 (.Q(\dc32_fifo_data_in[12] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[12]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i12 (.Q(\dc32_fifo_data_in[11] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[11]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i11 (.Q(\dc32_fifo_data_in[10] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[10]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i10 (.Q(\dc32_fifo_data_in[9] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[9]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i9 (.Q(\dc32_fifo_data_in[8] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[8]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i8 (.Q(\dc32_fifo_data_in[7] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[7]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i7 (.Q(\dc32_fifo_data_in[6] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[6]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i6 (.Q(\dc32_fifo_data_in[5] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[5]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i5 (.Q(\dc32_fifo_data_in[4] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[4]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i4 (.Q(\dc32_fifo_data_in[3] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[3]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i3 (.Q(\dc32_fifo_data_in[2] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[2]));   // src/usb3_if.v(194[8] 197[4])
    SB_DFFN dc32_fifo_data_in_i2 (.Q(\dc32_fifo_data_in[1] ), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[1]));   // src/usb3_if.v(194[8] 197[4])
    SB_LUT4 i3_4_lut (.I0(state_timeout_counter[0]), .I1(state_timeout_counter[2]), 
            .I2(state_timeout_counter[1]), .I3(state_timeout_counter[3]), 
            .O(n524));   // src/usb3_if.v(151[21:49])
    defparam i3_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_3_lut_adj_31 (.I0(n524), .I1(n562[2]), .I2(dc32_fifo_empty_latched), 
            .I3(GND_net), .O(n4224));   // src/usb3_if.v(98[9] 189[16])
    defparam i2_3_lut_adj_31.LUT_INIT = 16'h4040;
    SB_LUT4 i7_4_lut (.I0(num_lines_clocked_out[7]), .I1(num_lines_clocked_out[2]), 
            .I2(num_lines_clocked_out[9]), .I3(num_lines_clocked_out[0]), 
            .O(n18));   // src/usb3_if.v(175[29:57])
    defparam i7_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i5_2_lut (.I0(num_lines_clocked_out[1]), .I1(num_lines_clocked_out[5]), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // src/usb3_if.v(175[29:57])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut (.I0(num_lines_clocked_out[6]), .I1(n18), .I2(num_lines_clocked_out[3]), 
            .I3(num_lines_clocked_out[10]), .O(n20));   // src/usb3_if.v(175[29:57])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(num_lines_clocked_out[4]), .I1(n20), .I2(n16), 
            .I3(num_lines_clocked_out[8]), .O(n21));   // src/usb3_if.v(175[29:57])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1637_4_lut (.I0(n562[0]), .I1(n21), .I2(n522), .I3(n4224), 
            .O(n3004));   // src/usb3_if.v(98[9] 189[16])
    defparam i1637_4_lut.LUT_INIT = 16'hb3a0;
    SB_DFFESR state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(FIFO_CLK_c), 
            .E(n4310), .D(n2400), .R(n4703));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESS state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(FIFO_CLK_c), 
            .E(n4310), .D(n2401), .S(n4703));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(FIFO_CLK_c), 
            .E(n4310), .D(n2402), .R(n4703));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFSR write_to_dc32_fifo_latched_94 (.Q(write_to_dc32_fifo_latched), 
            .C(FIFO_CLK_c), .D(write_to_dc32_fifo_latched_N_425), .R(n2983));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i0 (.Q(num_lines_clocked_out[0]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[0]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(FIFO_CLK_c), 
            .E(n4310), .D(n2399), .R(n4703));   // src/usb3_if.v(88[8] 191[4])
    SB_LUT4 i150_2_lut_3_lut (.I0(buffer_switch_done_latched), .I1(dc32_fifo_empty_latched), 
            .I2(DEBUG_1_c_c), .I3(GND_net), .O(n522));   // src/usb3_if.v(100[21:96])
    defparam i150_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i148_2_lut_3_lut (.I0(buffer_switch_done_latched), .I1(dc32_fifo_empty_latched), 
            .I2(DEBUG_1_c_c), .I3(GND_net), .O(n520));   // src/usb3_if.v(100[21:96])
    defparam i148_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFFESR num_lines_clocked_out_i1 (.Q(num_lines_clocked_out[1]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[1]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_LUT4 reduce_or_206_i1_2_lut (.I0(n562[8]), .I1(n562[4]), .I2(GND_net), 
            .I3(GND_net), .O(n613));   // src/usb3_if.v(98[9] 189[16])
    defparam reduce_or_206_i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i231_3_lut (.I0(n613), .I1(FT_OE_N_420), .I2(n562[5]), .I3(GND_net), 
            .O(FT_RD_N_422));   // src/usb3_if.v(98[9] 189[16])
    defparam i231_3_lut.LUT_INIT = 16'hc5c5;
    SB_DFFESR num_lines_clocked_out_i2 (.Q(num_lines_clocked_out[2]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[2]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i3 (.Q(num_lines_clocked_out[3]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[3]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i4 (.Q(num_lines_clocked_out[4]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[4]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i5 (.Q(num_lines_clocked_out[5]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[5]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i6 (.Q(num_lines_clocked_out[6]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[6]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i7 (.Q(num_lines_clocked_out[7]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[7]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESS num_lines_clocked_out_i8 (.Q(num_lines_clocked_out[8]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[8]), .S(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESR num_lines_clocked_out_i9 (.Q(num_lines_clocked_out[9]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[9]), .R(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_DFFESS num_lines_clocked_out_i10 (.Q(num_lines_clocked_out[10]), .C(FIFO_CLK_c), 
            .E(n4486), .D(num_lines_clocked_out_10__N_371[10]), .S(reset_per_frame_latched));   // src/usb3_if.v(88[8] 191[4])
    SB_CARRY sub_113_add_2_4 (.CI(n10028), .I0(num_lines_clocked_out[2]), 
            .I1(VCC_net), .CO(n10029));
    SB_LUT4 sub_113_inv_0_i1_1_lut (.I0(dc32_fifo_empty_latched), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // src/usb3_if.v(174[50:77])
    defparam sub_113_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i202_2_lut_3_lut_4_lut (.I0(n524), .I1(dc32_fifo_almost_full), 
            .I2(DEBUG_1_c_c), .I3(n562[1]), .O(n608));   // src/usb3_if.v(98[9] 189[16])
    defparam i202_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1151_4_lut_4_lut (.I0(n562[5]), .I1(dc32_fifo_almost_full), 
            .I2(DEBUG_1_c_c), .I3(n524), .O(n2390));   // src/usb3_if.v(98[9] 189[16])
    defparam i1151_4_lut_4_lut.LUT_INIT = 16'h2276;
    SB_LUT4 mux_1159_i2_4_lut (.I0(n2408), .I1(n3940), .I2(n2415), .I3(dc32_fifo_empty_latched), 
            .O(n2400));   // src/usb3_if.v(98[9] 189[16])
    defparam mux_1159_i2_4_lut.LUT_INIT = 16'h3f35;
    SB_LUT4 i1_2_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n3940));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10259_3_lut (.I0(n10629), .I1(reset_per_frame_latched), .I2(n4181), 
            .I3(GND_net), .O(n4310));   // src/usb3_if.v(97[10] 190[8])
    defparam i10259_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_4_lut_adj_32 (.I0(n562[0]), .I1(n2266), .I2(n520), .I3(DEBUG_1_c_c), 
            .O(n10629));   // src/usb3_if.v(97[10] 190[8])
    defparam i1_4_lut_adj_32.LUT_INIT = 16'h0ace;
    SB_LUT4 i3321_4_lut (.I0(n4310), .I1(n562[2]), .I2(n562[0]), .I3(n2390), 
            .O(n4703));   // src/usb3_if.v(88[8] 191[4])
    defparam i3321_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1050_2_lut (.I0(n562[5]), .I1(dc32_fifo_almost_full), .I2(GND_net), 
            .I3(GND_net), .O(n2266));
    defparam i1050_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1159_i3_4_lut (.I0(n2408), .I1(n3938), .I2(n2415), .I3(n1[0]), 
            .O(n2401));   // src/usb3_if.v(98[9] 189[16])
    defparam mux_1159_i3_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 mux_1159_i4_4_lut (.I0(n11921), .I1(n3942), .I2(n2415), .I3(n2408), 
            .O(n2402));   // src/usb3_if.v(98[9] 189[16])
    defparam mux_1159_i4_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i10105_2_lut (.I0(n21), .I1(dc32_fifo_empty_latched), .I2(GND_net), 
            .I3(GND_net), .O(n11921));   // src/usb3_if.v(98[9] 189[16])
    defparam i10105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10200_2_lut (.I0(n562[5]), .I1(reset_per_frame_latched), .I2(GND_net), 
            .I3(GND_net), .O(n2983));   // src/usb3_if.v(88[8] 191[4])
    defparam i10200_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_3_lut (.I0(n524), .I1(reset_per_frame_latched), .I2(n562[2]), 
            .I3(GND_net), .O(n4486));
    defparam i1_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 mux_1159_i1_4_lut (.I0(n11881), .I1(state_timeout_counter[0]), 
            .I2(n2415), .I3(n2408), .O(n2399));   // src/usb3_if.v(98[9] 189[16])
    defparam mux_1159_i1_4_lut.LUT_INIT = 16'h3a3f;
    SB_LUT4 i10109_2_lut (.I0(n21), .I1(dc32_fifo_empty_latched), .I2(GND_net), 
            .I3(GND_net), .O(n11881));   // src/usb3_if.v(98[9] 189[16])
    defparam i10109_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i179_2_lut_3_lut (.I0(n524), .I1(dc32_fifo_almost_full), .I2(DEBUG_1_c_c), 
            .I3(GND_net), .O(n551));   // src/usb3_if.v(155[26] 157[24])
    defparam i179_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1647_3_lut_4_lut (.I0(n562[5]), .I1(n562[8]), .I2(n562[4]), 
            .I3(FT_OE_N_420), .O(n3014));   // src/usb3_if.v(98[9] 189[16])
    defparam i1647_3_lut_4_lut.LUT_INIT = 16'hfcfe;
    SB_LUT4 i2_3_lut_4_lut (.I0(n575), .I1(n571), .I2(n562[8]), .I3(n562[4]), 
            .O(n4181));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module \uart_tx(CLKS_PER_BIT=20) 
//

module \uart_tx(CLKS_PER_BIT=20)  (UART_TX_c, SLM_CLK_c, r_SM_Main, GND_net, 
            \r_SM_Main_2__N_841[1] , \r_SM_Main_2__N_844[0] , n3794, VCC_net, 
            n13737, n4890, r_Tx_Data, n4889, tx_uart_active_flag, 
            n5194, n5193, n5192, n5191, n5189, n5173, n5172, n10653) /* synthesis syn_module_defined=1 */ ;
    output UART_TX_c;
    input SLM_CLK_c;
    output [2:0]r_SM_Main;
    input GND_net;
    output \r_SM_Main_2__N_841[1] ;
    input \r_SM_Main_2__N_844[0] ;
    output n3794;
    input VCC_net;
    input n13737;
    input n4890;
    output [7:0]r_Tx_Data;
    input n4889;
    output tx_uart_active_flag;
    input n5194;
    input n5193;
    input n5192;
    input n5191;
    input n5189;
    input n5173;
    input n5172;
    output n10653;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n3, n1, n3063;
    wire [9:0]n45;
    wire [9:0]r_Clock_Count;   // src/uart_tx.v(32[16:29])
    
    wire n4798, n7448, n10796, n10816;
    wire [2:0]r_Bit_Index;   // src/uart_tx.v(33[16:27])
    
    wire n6076, n3_adj_1180, n10094, n10093, n10092, n10091, n10090, 
        n10089, n10088, n10087, n10086;
    wire [2:0]n312;
    
    wire n4, n8, n7, n3062, o_Tx_Serial_N_873, n10950, n10951, 
        n12687, n10933, n10932;
    
    SB_DFFE o_Tx_Serial_44 (.Q(UART_TX_c), .C(SLM_CLK_c), .E(n1), .D(n3));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n3063), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Clock_Count_1193__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[0]), .R(n4798));   // src/uart_tx.v(116[34:51])
    SB_LUT4 i10210_2_lut_3_lut (.I0(n7448), .I1(r_SM_Main[1]), .I2(n10796), 
            .I3(GND_net), .O(n10816));   // src/uart_tx.v(41[7] 140[14])
    defparam i10210_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i4693_3_lut_4_lut (.I0(n7448), .I1(r_SM_Main[1]), .I2(r_Bit_Index[0]), 
            .I3(n10796), .O(n6076));   // src/uart_tx.v(41[7] 140[14])
    defparam i4693_3_lut_4_lut.LUT_INIT = 16'h04f0;
    SB_LUT4 i10256_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_841[1] ), .O(n10796));
    defparam i10256_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_844[0] ), .O(n3794));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n6076));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n3_adj_1180), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(n13737));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 r_Clock_Count_1193_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n10094), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1193_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n10093), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_10 (.CI(n10093), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n10094));
    SB_LUT4 r_Clock_Count_1193_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n10092), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_9 (.CI(n10092), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n10093));
    SB_LUT4 r_Clock_Count_1193_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n10091), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_8 (.CI(n10091), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n10092));
    SB_LUT4 r_Clock_Count_1193_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n10090), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_7 (.CI(n10090), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n10091));
    SB_LUT4 r_Clock_Count_1193_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n10089), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_6 (.CI(n10089), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n10090));
    SB_LUT4 r_Clock_Count_1193_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n10088), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_5 (.CI(n10088), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n10089));
    SB_LUT4 r_Clock_Count_1193_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n10087), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_4 (.CI(n10087), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n10088));
    SB_LUT4 r_Clock_Count_1193_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n10086), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_3 (.CI(n10086), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n10087));
    SB_LUT4 r_Clock_Count_1193_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1193_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1193_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n10086));
    SB_DFFESR r_Clock_Count_1193__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[9]), .R(n4798));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[8]), .R(n4798));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[7]), .R(n4798));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[6]), .R(n4798));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[5]), .R(n4798));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[4]), .R(n4798));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[3]), .R(n4798));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[2]), .R(n4798));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1193__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[1]), .R(n4798));   // src/uart_tx.v(116[34:51])
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(SLM_CLK_c), .D(n4890));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Active_46 (.Q(tx_uart_active_flag), .C(SLM_CLK_c), .D(n4889));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(SLM_CLK_c), .E(n10796), 
            .D(n312[1]), .R(n10816));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(SLM_CLK_c), .E(n10796), 
            .D(n312[2]), .R(n10816));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i10203_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_841[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n4798));
    defparam i10203_4_lut.LUT_INIT = 16'h4445;
    SB_DFF r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(SLM_CLK_c), .D(n5194));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(SLM_CLK_c), .D(n5193));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(SLM_CLK_c), .D(n5192));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(SLM_CLK_c), .D(n5191));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(SLM_CLK_c), .D(n5189));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(SLM_CLK_c), .D(n5173));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(SLM_CLK_c), .D(n5172));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n4));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[9]), .I2(GND_net), 
            .I3(GND_net), .O(n8));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[4]), 
            .I3(n4), .O(n7));
    defparam i1_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i5_4_lut (.I0(r_Clock_Count[5]), .I1(n7), .I2(r_Clock_Count[8]), 
            .I3(n8), .O(\r_SM_Main_2__N_841[1] ));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1694_4_lut (.I0(\r_SM_Main_2__N_844[0] ), .I1(n7448), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_841[1] ), .O(n3062));   // src/uart_tx.v(41[7] 140[14])
    defparam i1694_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1695_3_lut (.I0(n3062), .I1(\r_SM_Main_2__N_841[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n3063));   // src/uart_tx.v(41[7] 140[14])
    defparam i1695_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10173_4_lut_4_lut (.I0(\r_SM_Main_2__N_841[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_844[0] ), .O(n10653));
    defparam i10173_4_lut_4_lut.LUT_INIT = 16'h8380;
    SB_LUT4 i2385_2_lut_3_lut (.I0(\r_SM_Main_2__N_841[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_1180));
    defparam i2385_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_SM_Main_2__I_0_55_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_873), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // src/uart_tx.v(41[7] 140[14])
    defparam r_SM_Main_2__I_0_55_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n10950), 
            .I2(n10951), .I3(r_Bit_Index[2]), .O(n12687));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n12687_bdd_4_lut (.I0(n12687), .I1(n10933), .I2(n10932), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_873));
    defparam n12687_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1372_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n312[2]));
    defparam i1372_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n7448));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1365_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n312[1]));   // src/uart_tx.v(96[36:51])
    defparam i1365_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9100_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n10950));
    defparam i9100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9101_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n10951));
    defparam i9101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9083_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n10933));
    defparam i9083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9082_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n10932));
    defparam i9082_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module spi
//

module spi (SEN_c_1, SLM_CLK_c, SOUT_c, n4312, \rx_shift_reg[0] , 
            \tx_data_byte[3] , n2086, GND_net, \tx_data_byte[4] , \tx_data_byte[5] , 
            n4319, SDAT_c_15, \tx_data_byte[6] , \tx_data_byte[7] , 
            tx_addr_byte, VCC_net, n10300, \tx_shift_reg[0] , n6049, 
            rx_buf_byte, n6048, n6047, n6046, n6045, n6044, n6043, 
            spi_rx_byte_ready, SCK_c_0, spi_start_transfer_r, n4897, 
            n4888, \rx_shift_reg[1] , n4883, \rx_shift_reg[2] , n4877, 
            \rx_shift_reg[3] , n4869, \rx_shift_reg[4] , n4838, \rx_shift_reg[5] , 
            n4836, \rx_shift_reg[6] , n4834, \rx_shift_reg[7] , multi_byte_spi_trans_flag_r, 
            \tx_data_byte[2] , \tx_data_byte[1] , n3495) /* synthesis syn_module_defined=1 */ ;
    output SEN_c_1;
    input SLM_CLK_c;
    input SOUT_c;
    output n4312;
    output \rx_shift_reg[0] ;
    input \tx_data_byte[3] ;
    output n2086;
    input GND_net;
    input \tx_data_byte[4] ;
    input \tx_data_byte[5] ;
    output n4319;
    output SDAT_c_15;
    input \tx_data_byte[6] ;
    input \tx_data_byte[7] ;
    input [7:0]tx_addr_byte;
    input VCC_net;
    input n10300;
    output \tx_shift_reg[0] ;
    input n6049;
    output [7:0]rx_buf_byte;
    input n6048;
    input n6047;
    input n6046;
    input n6045;
    input n6044;
    input n6043;
    output spi_rx_byte_ready;
    output SCK_c_0;
    input spi_start_transfer_r;
    input n4897;
    input n4888;
    output \rx_shift_reg[1] ;
    input n4883;
    output \rx_shift_reg[2] ;
    input n4877;
    output \rx_shift_reg[3] ;
    input n4869;
    output \rx_shift_reg[4] ;
    input n4838;
    output \rx_shift_reg[5] ;
    input n4836;
    output \rx_shift_reg[6] ;
    input n4834;
    output \rx_shift_reg[7] ;
    input multi_byte_spi_trans_flag_r;
    input \tx_data_byte[2] ;
    input \tx_data_byte[1] ;
    output n3495;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [2:0]n970;
    wire [3:0]state_3__N_938;
    
    wire n10665;
    wire [3:0]state;   // src/spi.v(71[11:16])
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    wire [15:0]n2087;
    
    wire n7098, n11946;
    wire [9:0]counter;   // src/spi.v(69[11:18])
    
    wire n11947;
    wire [9:0]n45;
    
    wire n4380, n4709, n10075, n10076, n24, n11943, n10074, n10073, 
        n10072, n10071, n10070, n10069, n10068;
    wire [7:0]n315;
    wire [7:0]multi_byte_counter;   // src/spi.v(68[11:29])
    wire [7:0]n2142;
    
    wire n10043, n10042, n10041, n10040, n10039, n10038, n10037, 
        n10780, n4, n37, n2, n51_adj_1168, n11916, n3748, n11917, 
        n14, n19, n11915, n11924, n34, n37_adj_1169, n10762, n4236, 
        n10624, n7, n4358, n10664, n4_adj_1170, n4629, n19_adj_1171, 
        n10666, n10638, n34_adj_1172, n4541, n4687, n10, n14_adj_1173, 
        n10_adj_1174, n14_adj_1175, n11933, n7_adj_1176, n3, n3_adj_1177, 
        n21, n22, n10802, n3_adj_1178, n4519, n11949, n7_adj_1179, 
        n11950;
    
    SB_DFF byte_recv_92_i2 (.Q(SEN_c_1), .C(SLM_CLK_c), .D(n970[1]));   // src/spi.v(88[9] 219[16])
    SB_DFFE rx_shift_reg_i0 (.Q(\rx_shift_reg[0] ), .C(SLM_CLK_c), .E(n4312), 
            .D(SOUT_c));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n10665), .D(state_3__N_938[0]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_981_i4_3_lut (.I0(\tx_data_byte[3] ), .I1(tx_shift_reg[2]), 
            .I2(n2086), .I3(GND_net), .O(n2087[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i5_3_lut (.I0(\tx_data_byte[4] ), .I1(tx_shift_reg[3]), 
            .I2(n2086), .I3(GND_net), .O(n2087[4]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10146_4_lut (.I0(n7098), .I1(state[1]), .I2(state[0]), .I3(state[2]), 
            .O(n11946));   // src/spi.v(88[9] 219[16])
    defparam i10146_4_lut.LUT_INIT = 16'hc08c;
    SB_LUT4 i1_4_lut (.I0(counter[4]), .I1(n11946), .I2(n11947), .I3(state[3]), 
            .O(n970[0]));   // src/spi.v(76[8] 221[4])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 mux_981_i6_3_lut (.I0(\tx_data_byte[5] ), .I1(tx_shift_reg[4]), 
            .I2(n2086), .I3(GND_net), .O(n2087[5]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR counter_1189__i0 (.Q(counter[0]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[0]), .R(n4709));   // src/spi.v(183[28:41])
    SB_DFFE tx_shift_reg_i0_i15 (.Q(SDAT_c_15), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[15]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_981_i7_3_lut (.I0(\tx_data_byte[6] ), .I1(tx_shift_reg[5]), 
            .I2(n2086), .I3(GND_net), .O(n2087[6]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i8_3_lut (.I0(\tx_data_byte[7] ), .I1(tx_shift_reg[6]), 
            .I2(n2086), .I3(GND_net), .O(n2087[7]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i9_3_lut (.I0(tx_addr_byte[0]), .I1(tx_shift_reg[7]), 
            .I2(n2086), .I3(GND_net), .O(n2087[8]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i10_3_lut (.I0(tx_addr_byte[1]), .I1(tx_shift_reg[8]), 
            .I2(n2086), .I3(GND_net), .O(n2087[9]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i11_3_lut (.I0(tx_addr_byte[2]), .I1(tx_shift_reg[9]), 
            .I2(n2086), .I3(GND_net), .O(n2087[10]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i12_3_lut (.I0(tx_addr_byte[3]), .I1(tx_shift_reg[10]), 
            .I2(n2086), .I3(GND_net), .O(n2087[11]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i13_3_lut (.I0(tx_addr_byte[4]), .I1(tx_shift_reg[11]), 
            .I2(n2086), .I3(GND_net), .O(n2087[12]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_1189_add_4_10 (.CI(n10075), .I0(VCC_net), .I1(counter[8]), 
            .CO(n10076));
    SB_LUT4 i1_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n24));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i10142_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n11943));
    defparam i10142_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mux_981_i14_3_lut (.I0(tx_addr_byte[5]), .I1(tx_shift_reg[12]), 
            .I2(n2086), .I3(GND_net), .O(n2087[13]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i15_3_lut (.I0(tx_addr_byte[6]), .I1(tx_shift_reg[13]), 
            .I2(n2086), .I3(GND_net), .O(n2087[14]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_1189_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[7]), 
            .I3(n10074), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_9 (.CI(n10074), .I0(VCC_net), .I1(counter[7]), 
            .CO(n10075));
    SB_DFFE tx_shift_reg_i0_i0 (.Q(\tx_shift_reg[0] ), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n10300));   // src/spi.v(76[8] 221[4])
    SB_LUT4 counter_1189_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[6]), 
            .I3(n10073), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF Rx_Recv_Byte_i1 (.Q(rx_buf_byte[1]), .C(SLM_CLK_c), .D(n6049));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i2 (.Q(rx_buf_byte[2]), .C(SLM_CLK_c), .D(n6048));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i3 (.Q(rx_buf_byte[3]), .C(SLM_CLK_c), .D(n6047));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i4 (.Q(rx_buf_byte[4]), .C(SLM_CLK_c), .D(n6046));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i5 (.Q(rx_buf_byte[5]), .C(SLM_CLK_c), .D(n6045));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i6 (.Q(rx_buf_byte[6]), .C(SLM_CLK_c), .D(n6044));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i7 (.Q(rx_buf_byte[7]), .C(SLM_CLK_c), .D(n6043));   // src/spi.v(76[8] 221[4])
    SB_CARRY counter_1189_add_4_8 (.CI(n10073), .I0(VCC_net), .I1(counter[6]), 
            .CO(n10074));
    SB_LUT4 counter_1189_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[5]), 
            .I3(n10072), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_7 (.CI(n10072), .I0(VCC_net), .I1(counter[5]), 
            .CO(n10073));
    SB_LUT4 counter_1189_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[4]), 
            .I3(n10071), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_6 (.CI(n10071), .I0(VCC_net), .I1(counter[4]), 
            .CO(n10072));
    SB_LUT4 counter_1189_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[3]), 
            .I3(n10070), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_5 (.CI(n10070), .I0(VCC_net), .I1(counter[3]), 
            .CO(n10071));
    SB_LUT4 counter_1189_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[2]), 
            .I3(n10069), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_4 (.CI(n10069), .I0(VCC_net), .I1(counter[2]), 
            .CO(n10070));
    SB_LUT4 counter_1189_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[1]), 
            .I3(n10068), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_3 (.CI(n10068), .I0(VCC_net), .I1(counter[1]), 
            .CO(n10069));
    SB_LUT4 counter_1189_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1189_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n10068));
    SB_LUT4 add_995_9_lut (.I0(GND_net), .I1(multi_byte_counter[7]), .I2(n2142[5]), 
            .I3(n10043), .O(n315[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_995_8_lut (.I0(GND_net), .I1(multi_byte_counter[6]), .I2(n2142[5]), 
            .I3(n10042), .O(n315[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_8 (.CI(n10042), .I0(multi_byte_counter[6]), .I1(n2142[5]), 
            .CO(n10043));
    SB_LUT4 add_995_7_lut (.I0(GND_net), .I1(multi_byte_counter[5]), .I2(n2142[5]), 
            .I3(n10041), .O(n315[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_7 (.CI(n10041), .I0(multi_byte_counter[5]), .I1(n2142[5]), 
            .CO(n10042));
    SB_LUT4 add_995_6_lut (.I0(GND_net), .I1(multi_byte_counter[4]), .I2(n2142[5]), 
            .I3(n10040), .O(n315[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_6 (.CI(n10040), .I0(multi_byte_counter[4]), .I1(n2142[5]), 
            .CO(n10041));
    SB_LUT4 add_995_5_lut (.I0(GND_net), .I1(multi_byte_counter[3]), .I2(n2142[5]), 
            .I3(n10039), .O(n315[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_5 (.CI(n10039), .I0(multi_byte_counter[3]), .I1(n2142[5]), 
            .CO(n10040));
    SB_LUT4 add_995_4_lut (.I0(GND_net), .I1(multi_byte_counter[2]), .I2(n2142[5]), 
            .I3(n10038), .O(n315[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_4 (.CI(n10038), .I0(multi_byte_counter[2]), .I1(n2142[5]), 
            .CO(n10039));
    SB_LUT4 add_995_3_lut (.I0(GND_net), .I1(multi_byte_counter[1]), .I2(n2142[5]), 
            .I3(n10037), .O(n315[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_3 (.CI(n10037), .I0(multi_byte_counter[1]), .I1(n2142[5]), 
            .CO(n10038));
    SB_LUT4 add_995_2_lut (.I0(GND_net), .I1(multi_byte_counter[0]), .I2(n2142[5]), 
            .I3(GND_net), .O(n315[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_995_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_995_2 (.CI(GND_net), .I0(multi_byte_counter[0]), .I1(n2142[5]), 
            .CO(n10037));
    SB_LUT4 i8931_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n10780));
    defparam i8931_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(state[3]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n4));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE tx_shift_reg_i0_i14 (.Q(tx_shift_reg[14]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[14]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i13 (.Q(tx_shift_reg[13]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[13]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i12 (.Q(tx_shift_reg[12]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[12]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i11 (.Q(tx_shift_reg[11]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[11]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i10 (.Q(tx_shift_reg[10]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[10]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_4_lut_adj_14 (.I0(n37), .I1(n4), .I2(n2), .I3(n10780), 
            .O(n2086));
    defparam i1_4_lut_adj_14.LUT_INIT = 16'ha0a8;
    SB_DFFE tx_shift_reg_i0_i9 (.Q(tx_shift_reg[9]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[9]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i8 (.Q(tx_shift_reg[8]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[8]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i7 (.Q(tx_shift_reg[7]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[7]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i6 (.Q(tx_shift_reg[6]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[6]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_2_lut_adj_15 (.I0(counter[4]), .I1(n51_adj_1168), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // src/spi.v(183[28:41])
    defparam i1_2_lut_adj_15.LUT_INIT = 16'h4444;
    SB_DFF byte_recv_92_i3 (.Q(spi_rx_byte_ready), .C(SLM_CLK_c), .D(n970[2]));   // src/spi.v(88[9] 219[16])
    SB_DFFE tx_shift_reg_i0_i5 (.Q(tx_shift_reg[5]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[5]));   // src/spi.v(76[8] 221[4])
    SB_DFF byte_recv_92_i1 (.Q(SCK_c_0), .C(SLM_CLK_c), .D(n970[0]));   // src/spi.v(88[9] 219[16])
    SB_DFFE tx_shift_reg_i0_i4 (.Q(tx_shift_reg[4]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[4]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i3 (.Q(tx_shift_reg[3]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[3]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i10133_4_lut (.I0(spi_start_transfer_r), .I1(state[0]), .I2(n37), 
            .I3(state[3]), .O(n11916));   // src/spi.v(71[11:16])
    defparam i10133_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_4_lut_adj_16 (.I0(n3748), .I1(n11916), .I2(n11917), .I3(state[1]), 
            .O(n4319));
    defparam i1_4_lut_adj_16.LUT_INIT = 16'h5044;
    SB_LUT4 mux_981_i16_3_lut (.I0(tx_addr_byte[7]), .I1(tx_shift_reg[14]), 
            .I2(n2086), .I3(GND_net), .O(n2087[15]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), .I3(GND_net), 
            .O(n14));   // src/spi.v(88[9] 219[16])
    defparam i1_3_lut.LUT_INIT = 16'hcdcd;
    SB_LUT4 i10131_3_lut (.I0(state[0]), .I1(state[2]), .I2(n19), .I3(GND_net), 
            .O(n11915));
    defparam i10131_3_lut.LUT_INIT = 16'h4d4d;
    SB_LUT4 i10144_3_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), 
            .I3(GND_net), .O(n11924));
    defparam i10144_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i65_3_lut (.I0(n14), .I1(n11915), .I2(state[1]), .I3(GND_net), 
            .O(n34));
    defparam i65_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i66_4_lut (.I0(n11924), .I1(n2142[5]), .I2(state[1]), .I3(state[3]), 
            .O(n37_adj_1169));
    defparam i66_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut_adj_17 (.I0(state[3]), .I1(n37_adj_1169), .I2(n34), 
            .I3(n10762), .O(n4709));
    defparam i1_4_lut_adj_17.LUT_INIT = 16'h50dc;
    SB_LUT4 i10238_4_lut (.I0(state[3]), .I1(state[1]), .I2(n4236), .I3(n14), 
            .O(n4380));   // src/spi.v(88[9] 219[16])
    defparam i10238_4_lut.LUT_INIT = 16'h4c5f;
    SB_DFF Rx_Recv_Byte_i0 (.Q(rx_buf_byte[0]), .C(SLM_CLK_c), .D(n4897));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i1 (.Q(\rx_shift_reg[1] ), .C(SLM_CLK_c), .D(n4888));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i2 (.Q(tx_shift_reg[2]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i1 (.Q(tx_shift_reg[1]), .C(SLM_CLK_c), .E(n4319), 
            .D(n2087[1]));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i2 (.Q(\rx_shift_reg[2] ), .C(SLM_CLK_c), .D(n4883));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_1189__i1 (.Q(counter[1]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[1]), .R(n4709));   // src/spi.v(183[28:41])
    SB_LUT4 i2_3_lut (.I0(state[3]), .I1(n19), .I2(state[1]), .I3(GND_net), 
            .O(n10624));
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_DFFESR counter_1189__i2 (.Q(counter[2]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[2]), .R(n4709));   // src/spi.v(183[28:41])
    SB_LUT4 i4_4_lut (.I0(n7), .I1(state[3]), .I2(spi_start_transfer_r), 
            .I3(state[0]), .O(n4358));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_18 (.I0(n4358), .I1(n10624), .I2(state[0]), .I3(state[2]), 
            .O(n10664));
    defparam i1_4_lut_adj_18.LUT_INIT = 16'h8aaa;
    SB_LUT4 i2_2_lut (.I0(state[1]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n7));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESR counter_1189__i3 (.Q(counter[3]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[3]), .R(n4709));   // src/spi.v(183[28:41])
    SB_LUT4 i1_2_lut_adj_19 (.I0(n19), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_1170));
    defparam i1_2_lut_adj_19.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut_adj_20 (.I0(n7), .I1(n10664), .I2(state[3]), .I3(n4_adj_1170), 
            .O(n10665));
    defparam i1_4_lut_adj_20.LUT_INIT = 16'h4c0c;
    SB_LUT4 i3_4_lut (.I0(counter[0]), .I1(counter[3]), .I2(counter[2]), 
            .I3(counter[1]), .O(n51_adj_1168));   // src/spi.v(183[28:41])
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_DFFESR counter_1189__i4 (.Q(counter[4]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[4]), .R(n4709));   // src/spi.v(183[28:41])
    SB_LUT4 i8913_2_lut (.I0(state[0]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n10762));
    defparam i8913_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_21 (.I0(state[2]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3748));   // src/spi.v(88[9] 219[16])
    defparam i1_2_lut_adj_21.LUT_INIT = 16'h2222;
    SB_LUT4 i10248_3_lut (.I0(counter[4]), .I1(n4629), .I2(n51_adj_1168), 
            .I3(GND_net), .O(n4312));   // src/spi.v(88[9] 219[16])
    defparam i10248_3_lut.LUT_INIT = 16'h2020;
    SB_DFFESR counter_1189__i5 (.Q(counter[5]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[5]), .R(n4709));   // src/spi.v(183[28:41])
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(n19_adj_1171), .D(state_3__N_938[3]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n10666), .D(state_3__N_938[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n10638), .D(state_3__N_938[1]));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i3 (.Q(\rx_shift_reg[3] ), .C(SLM_CLK_c), .D(n4877));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_1189__i6 (.Q(counter[6]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[6]), .R(n4709));   // src/spi.v(183[28:41])
    SB_DFF rx_shift_reg_i4 (.Q(\rx_shift_reg[4] ), .C(SLM_CLK_c), .D(n4869));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_1189__i9 (.Q(counter[9]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[9]), .R(n4709));   // src/spi.v(183[28:41])
    SB_DFFESS counter_1189__i8 (.Q(counter[8]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[8]), .S(n4709));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1189__i7 (.Q(counter[7]), .C(SLM_CLK_c), .E(n4380), 
            .D(n45[7]), .R(n4709));   // src/spi.v(183[28:41])
    SB_LUT4 i2_3_lut_adj_22 (.I0(counter[2]), .I1(counter[1]), .I2(counter[3]), 
            .I3(GND_net), .O(n34_adj_1172));   // src/spi.v(183[28:41])
    defparam i2_3_lut_adj_22.LUT_INIT = 16'hfefe;
    SB_DFFESR multi_byte_counter_i1 (.Q(multi_byte_counter[1]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[1]), .R(n4687));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i2_2_lut_adj_23 (.I0(counter[6]), .I1(counter[7]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // src/spi.v(141[21:41])
    defparam i2_2_lut_adj_23.LUT_INIT = 16'heeee;
    SB_DFFESR multi_byte_counter_i2 (.Q(multi_byte_counter[2]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[2]), .R(n4687));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i0 (.Q(multi_byte_counter[0]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[0]), .R(n4687));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i6_4_lut (.I0(counter[4]), .I1(counter[5]), .I2(counter[9]), 
            .I3(n34_adj_1172), .O(n14_adj_1173));   // src/spi.v(141[21:41])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR multi_byte_counter_i3 (.Q(multi_byte_counter[3]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[3]), .R(n4687));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i7_4_lut (.I0(counter[0]), .I1(n14_adj_1173), .I2(n10), .I3(counter[8]), 
            .O(n19));   // src/spi.v(141[21:41])
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_2_lut_adj_24 (.I0(multi_byte_counter[2]), .I1(multi_byte_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_1174));   // src/spi.v(208[21:52])
    defparam i2_2_lut_adj_24.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_25 (.I0(multi_byte_counter[3]), .I1(multi_byte_counter[1]), 
            .I2(multi_byte_counter[5]), .I3(multi_byte_counter[7]), .O(n14_adj_1175));   // src/spi.v(208[21:52])
    defparam i6_4_lut_adj_25.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_26 (.I0(multi_byte_counter[0]), .I1(n14_adj_1175), 
            .I2(n10_adj_1174), .I3(multi_byte_counter[6]), .O(n2142[5]));   // src/spi.v(208[21:52])
    defparam i7_4_lut_adj_26.LUT_INIT = 16'hfffd;
    SB_LUT4 i10154_3_lut (.I0(n2142[5]), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n11933));   // src/spi.v(88[9] 219[16])
    defparam i10154_3_lut.LUT_INIT = 16'hc4c4;
    SB_DFFESR multi_byte_counter_i4 (.Q(multi_byte_counter[4]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[4]), .R(n4687));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_344_Mux_1_i7_4_lut (.I0(state[0]), .I1(state[2]), .I2(n19), 
            .I3(state[1]), .O(n7_adj_1176));   // src/spi.v(88[9] 219[16])
    defparam mux_344_Mux_1_i7_4_lut.LUT_INIT = 16'h02dd;
    SB_LUT4 mux_344_Mux_1_i15_4_lut (.I0(n7_adj_1176), .I1(n11933), .I2(state[3]), 
            .I3(state[2]), .O(n970[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_344_Mux_1_i15_4_lut.LUT_INIT = 16'hfaca;
    SB_DFFESS multi_byte_counter_i5 (.Q(multi_byte_counter[5]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[5]), .S(n4687));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i6 (.Q(multi_byte_counter[6]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[6]), .R(n4687));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i5 (.Q(\rx_shift_reg[5] ), .C(SLM_CLK_c), .D(n4838));   // src/spi.v(76[8] 221[4])
    SB_DFFESS multi_byte_counter_i7 (.Q(multi_byte_counter[7]), .C(SLM_CLK_c), 
            .E(n4541), .D(n315[7]), .S(n4687));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i6 (.Q(\rx_shift_reg[6] ), .C(SLM_CLK_c), .D(n4836));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i7 (.Q(\rx_shift_reg[7] ), .C(SLM_CLK_c), .D(n4834));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_56_Mux_1_i3_3_lut_3_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(GND_net), .O(n3));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i3_3_lut_3_lut.LUT_INIT = 16'h3e3e;
    SB_LUT4 mux_56_Mux_0_i3_4_lut_4_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(n19), .O(n3_adj_1177));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_0_i3_4_lut_4_lut.LUT_INIT = 16'hc131;
    SB_LUT4 i43_4_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(state[1]), 
            .I3(state[0]), .O(n21));
    defparam i43_4_lut_4_lut.LUT_INIT = 16'hf01a;
    SB_LUT4 i3273_3_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), 
            .I3(n3_adj_1177), .O(state_3__N_938[0]));
    defparam i3273_3_lut_4_lut.LUT_INIT = 16'h1f0e;
    SB_LUT4 counter_1189_add_4_11_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[9]), 
            .I3(n10076), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1189_add_4_10_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[8]), 
            .I3(n10075), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1189_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(state[1]), 
            .I3(state[3]), .O(n2));   // src/spi.v(88[9] 219[16])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h00b0;
    SB_LUT4 mux_981_i3_3_lut (.I0(\tx_data_byte[2] ), .I1(tx_shift_reg[1]), 
            .I2(n2086), .I3(GND_net), .O(n2087[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_981_i2_3_lut (.I0(\tx_data_byte[1] ), .I1(\tx_shift_reg[0] ), 
            .I2(n2086), .I3(GND_net), .O(n2087[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_981_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_56_Mux_3_i15_4_lut (.I0(n11943), .I1(state[1]), .I2(state[3]), 
            .I3(n2142[5]), .O(state_3__N_938[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_3_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i10235_4_lut (.I0(n22), .I1(n10802), .I2(n24), .I3(state[3]), 
            .O(n19_adj_1171));
    defparam i10235_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i1_2_lut_adj_27 (.I0(n19), .I1(n21), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i1_2_lut_adj_27.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[2]), .I1(n10624), .I2(n4358), .I3(state[0]), 
            .O(n10666));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hc0e0;
    SB_LUT4 mux_56_Mux_2_i15_4_lut (.I0(n3_adj_1178), .I1(state[2]), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_938[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 mux_56_Mux_2_i3_3_lut (.I0(multi_byte_spi_trans_flag_r), .I1(state[0]), 
            .I2(state[1]), .I3(GND_net), .O(n3_adj_1178));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i3_3_lut.LUT_INIT = 16'hc2c2;
    SB_LUT4 i1_2_lut_adj_28 (.I0(state[2]), .I1(n10624), .I2(GND_net), 
            .I3(GND_net), .O(n4519));
    defparam i1_2_lut_adj_28.LUT_INIT = 16'heeee;
    SB_LUT4 i8953_3_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(spi_start_transfer_r), 
            .I3(state[2]), .O(n10802));
    defparam i8953_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_56_Mux_1_i7_4_lut (.I0(n3), .I1(n11949), .I2(state[2]), 
            .I3(state[1]), .O(n7_adj_1179));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i7_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i10165_2_lut (.I0(n19), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n11949));   // src/spi.v(88[9] 219[16])
    defparam i10165_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_4_lut (.I0(state[3]), .I1(n4519), .I2(n24), .I3(n4358), 
            .O(n10638));
    defparam i2_4_lut.LUT_INIT = 16'h4c00;
    SB_LUT4 i10145_2_lut_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(n7098), .O(n11947));   // src/spi.v(88[9] 219[16])
    defparam i10145_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i2050_4_lut_4_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(state[3]), .O(n4629));   // src/spi.v(88[9] 219[16])
    defparam i2050_4_lut_4_lut_4_lut.LUT_INIT = 16'hfe75;
    SB_LUT4 i1_4_lut_adj_29 (.I0(state[1]), .I1(n4), .I2(n11950), .I3(state[0]), 
            .O(n4541));
    defparam i1_4_lut_adj_29.LUT_INIT = 16'ha088;
    SB_LUT4 i10164_3_lut (.I0(state[3]), .I1(state[2]), .I2(n19), .I3(GND_net), 
            .O(n11950));
    defparam i10164_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i3304_2_lut (.I0(n4541), .I1(state[3]), .I2(GND_net), .I3(GND_net), 
            .O(n4687));   // src/spi.v(76[8] 221[4])
    defparam i3304_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_4_lut (.I0(n2142[5]), .I1(state[0]), .I2(state[2]), 
            .I3(state[1]), .O(n4236));   // src/spi.v(88[9] 219[16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i10106_2_lut_3_lut (.I0(counter[4]), .I1(n51_adj_1168), .I2(state[3]), 
            .I3(GND_net), .O(n11917));   // src/spi.v(71[11:16])
    defparam i10106_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i2123_4_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(state[1]), 
            .I3(state[3]), .O(n3495));   // src/spi.v(88[9] 219[16])
    defparam i2123_4_lut_4_lut.LUT_INIT = 16'hfdfb;
    SB_LUT4 mux_344_Mux_2_i15_4_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[2]), .I3(state[3]), .O(n970[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_344_Mux_2_i15_4_lut_4_lut.LUT_INIT = 16'h0420;
    SB_LUT4 mux_56_Mux_1_i15_3_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[3]), .I3(n7_adj_1179), .O(state_3__N_938[1]));
    defparam mux_56_Mux_1_i15_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i1_2_lut_4_lut_adj_30 (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(counter[3]), .O(n7098));   // src/spi.v(183[28:41])
    defparam i1_2_lut_4_lut_adj_30.LUT_INIT = 16'hfffe;
    
endmodule

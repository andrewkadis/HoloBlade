// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue Mar 30 03:01:22 2021
//
// Verilog Description of module top
//

module top (ICE_SYSCLK, DCD, DSR, DTR, CTS, RST, UART_RX, UART_TX, 
            SEN, SCK, SOUT, SDAT, UPDATE, RESET, SLM_CLK, INVERT, 
            SYNC, VALID, DATA31, DATA0, DATA30, DATA29, DATA1, 
            DATA28, DATA27, DATA2, DATA26, DATA25, DATA3, DATA24, 
            DATA23, DATA4, DATA22, DATA21, DATA5, DATA20, DATA19, 
            DATA6, DATA18, DATA17, DATA7, DATA16, DATA15, DATA8, 
            DATA14, DATA13, DATA12, DATA11, DATA9, DATA10, FT_OE, 
            FT_RD, FT_WR, FT_SIWU, FR_RXF, FT_TXE, FIFO_BE3, FIFO_BE2, 
            FIFO_BE1, FIFO_BE0, FIFO_D31, FIFO_D30, FIFO_D29, FIFO_D28, 
            FIFO_D27, FIFO_CLK, FIFO_D26, FIFO_D25, FIFO_D24, FIFO_D23, 
            FIFO_D22, FIFO_D21, FIFO_D20, FIFO_D19, FIFO_D18, FIFO_D17, 
            FIFO_D16, FIFO_D15, FIFO_D14, FIFO_D13, FIFO_D12, FIFO_D11, 
            FIFO_D10, FIFO_D9, FIFO_D8, FIFO_D7, FIFO_D6, FIFO_D5, 
            FIFO_D4, FIFO_D3, FIFO_D2, FIFO_D1, FIFO_D0, DEBUG_0, 
            DEBUG_1, DEBUG_2, DEBUG_3, DEBUG_5, DEBUG_6, DEBUG_8, 
            DEBUG_9, ICE_CLK, ICE_CDONE, ICE_CREST) /* synthesis syn_module_defined=1 */ ;   // src/top.v(5[8:11])
    input ICE_SYSCLK;   // src/top.v(8[11:21])
    output DCD;   // src/top.v(11[12:15])
    output DSR;   // src/top.v(12[12:15])
    output DTR;   // src/top.v(13[12:15])
    output CTS;   // src/top.v(14[12:15])
    output RST;   // src/top.v(15[12:15])
    input UART_RX;   // src/top.v(16[12:19])
    output UART_TX;   // src/top.v(17[12:19])
    output SEN;   // src/top.v(20[12:15])
    output SCK;   // src/top.v(21[12:15])
    input SOUT;   // src/top.v(22[12:16])
    output SDAT;   // src/top.v(23[12:16])
    output UPDATE;   // src/top.v(27[12:18])
    output RESET;   // src/top.v(28[12:17])
    output SLM_CLK;   // src/top.v(29[12:19])
    output INVERT;   // src/top.v(30[12:18])
    output SYNC;   // src/top.v(31[12:16])
    output VALID;   // src/top.v(32[12:17])
    output DATA31;   // src/top.v(34[12:18])
    output DATA0;   // src/top.v(35[12:17])
    output DATA30;   // src/top.v(36[12:18])
    output DATA29;   // src/top.v(37[12:18])
    output DATA1;   // src/top.v(38[12:17])
    output DATA28;   // src/top.v(39[12:18])
    output DATA27;   // src/top.v(40[12:18])
    output DATA2;   // src/top.v(41[12:17])
    output DATA26;   // src/top.v(42[12:18])
    output DATA25;   // src/top.v(43[12:18])
    output DATA3;   // src/top.v(44[12:17])
    output DATA24;   // src/top.v(45[12:18])
    output DATA23;   // src/top.v(46[12:18])
    output DATA4;   // src/top.v(47[12:17])
    output DATA22;   // src/top.v(48[12:18])
    output DATA21;   // src/top.v(49[12:18])
    output DATA5;   // src/top.v(50[12:17])
    output DATA20;   // src/top.v(51[12:18])
    output DATA19;   // src/top.v(52[12:18])
    output DATA6;   // src/top.v(53[12:17])
    output DATA18;   // src/top.v(54[12:18])
    output DATA17;   // src/top.v(55[12:18])
    output DATA7;   // src/top.v(56[12:17])
    output DATA16;   // src/top.v(57[12:18])
    output DATA15;   // src/top.v(58[12:18])
    output DATA8;   // src/top.v(59[12:17])
    output DATA14;   // src/top.v(60[12:18])
    output DATA13;   // src/top.v(61[12:18])
    output DATA12;   // src/top.v(62[12:18])
    output DATA11;   // src/top.v(63[12:18])
    output DATA9;   // src/top.v(64[12:17])
    output DATA10;   // src/top.v(65[12:18])
    output FT_OE;   // src/top.v(69[12:17])
    output FT_RD;   // src/top.v(70[12:17])
    output FT_WR;   // src/top.v(71[12:17])
    output FT_SIWU;   // src/top.v(72[12:19])
    input FR_RXF;   // src/top.v(73[12:18])
    input FT_TXE;   // src/top.v(74[12:18])
    input FIFO_BE3;   // src/top.v(75[12:20])
    input FIFO_BE2;   // src/top.v(76[12:20])
    input FIFO_BE1;   // src/top.v(77[12:20])
    input FIFO_BE0;   // src/top.v(78[12:20])
    input FIFO_D31;   // src/top.v(79[12:20])
    input FIFO_D30;   // src/top.v(80[12:20])
    input FIFO_D29;   // src/top.v(81[12:20])
    input FIFO_D28;   // src/top.v(82[12:20])
    input FIFO_D27;   // src/top.v(83[12:20])
    input FIFO_CLK;   // src/top.v(84[12:20])
    input FIFO_D26;   // src/top.v(85[12:20])
    input FIFO_D25;   // src/top.v(86[12:20])
    input FIFO_D24;   // src/top.v(87[12:20])
    input FIFO_D23;   // src/top.v(88[12:20])
    input FIFO_D22;   // src/top.v(89[12:20])
    input FIFO_D21;   // src/top.v(90[12:20])
    input FIFO_D20;   // src/top.v(91[12:20])
    input FIFO_D19;   // src/top.v(92[12:20])
    input FIFO_D18;   // src/top.v(93[12:20])
    input FIFO_D17;   // src/top.v(94[12:20])
    input FIFO_D16;   // src/top.v(95[12:20])
    input FIFO_D15;   // src/top.v(97[11:19])
    input FIFO_D14;   // src/top.v(98[11:19])
    input FIFO_D13;   // src/top.v(99[11:19])
    input FIFO_D12;   // src/top.v(100[11:19])
    input FIFO_D11;   // src/top.v(101[11:19])
    input FIFO_D10;   // src/top.v(102[11:19])
    input FIFO_D9;   // src/top.v(103[11:18])
    input FIFO_D8;   // src/top.v(104[11:18])
    input FIFO_D7;   // src/top.v(105[11:18])
    input FIFO_D6;   // src/top.v(106[11:18])
    input FIFO_D5;   // src/top.v(107[11:18])
    input FIFO_D4;   // src/top.v(108[11:18])
    input FIFO_D3;   // src/top.v(109[11:18])
    input FIFO_D2;   // src/top.v(110[11:18])
    input FIFO_D1;   // src/top.v(111[11:18])
    input FIFO_D0;   // src/top.v(112[11:18])
    output DEBUG_0;   // src/top.v(115[12:19])
    output DEBUG_1;   // src/top.v(116[12:19])
    output DEBUG_2;   // src/top.v(117[12:19])
    output DEBUG_3;   // src/top.v(118[12:19])
    output DEBUG_5;   // src/top.v(119[12:19])
    output DEBUG_6;   // src/top.v(120[12:19])
    output DEBUG_8;   // src/top.v(121[12:19])
    output DEBUG_9;   // src/top.v(122[12:19])
    output ICE_CLK;   // src/top.v(125[12:19])
    output ICE_CDONE;   // src/top.v(126[12:21])
    output ICE_CREST;   // src/top.v(127[12:21])
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire FIFO_CLK_c /* synthesis SET_AS_NETWORK=FIFO_CLK_c, is_clock=1 */ ;   // src/top.v(84[12:20])
    
    wire GND_net, VCC_net, ICE_SYSCLK_c, DEBUG_2_c_c, DEBUG_1_c, SEN_c_1, 
        SCK_c_0, SOUT_c, SDAT_c_15, UPDATE_c_3, RESET_c, INVERT_c_4, 
        SYNC_c, DEBUG_6_c, DATA31_c_31, DEBUG_8_c, DATA30_c_30, DATA29_c_29, 
        DATA1_c_1, DATA28_c_28, DATA27_c_27, DATA2_c_2, DATA26_c_26, 
        DATA25_c_25, DATA3_c_3, DATA24_c_24, DATA23_c_23, DATA4_c_4, 
        DATA22_c_22, DATA21_c_21, DATA5_c_5, DATA20_c_20, DATA19_c_19, 
        DATA6_c_6, DATA18_c_18, DATA17_c_17, DATA7_c_7, DATA16_c_16, 
        DATA15_c_15, DATA8_c_8, DATA14_c_14, DATA13_c_13, DATA12_c_12, 
        DATA11_c_11, DATA9_c_9, DATA10_c_10, FT_OE_c, FT_RD_c, DEBUG_9_c_c, 
        FIFO_D31_c_0, FIFO_D30_c_1, FIFO_D29_c_2, FIFO_D28_c_3, FIFO_D27_c_4, 
        FIFO_D26_c_5, FIFO_D25_c_6, FIFO_D24_c_7, FIFO_D23_c_8, FIFO_D22_c_9, 
        FIFO_D21_c_10, FIFO_D20_c_11, FIFO_D19_c_12, FIFO_D18_c_13, 
        FIFO_D17_c_14, FIFO_D16_c_15, FIFO_D15_c_16, FIFO_D14_c_17, 
        FIFO_D13_c_18, FIFO_D12_c_19, FIFO_D11_c_20, FIFO_D10_c_21, 
        FIFO_D9_c_22, FIFO_D8_c_23, FIFO_D7_c_24, FIFO_D6_c_25, FIFO_D5_c_26, 
        FIFO_D4_c_27, FIFO_D3_c_28, FIFO_D2_c_29, FIFO_D1_c_30, FIFO_D0_c_31, 
        DEBUG_0_c_24, DEBUG_5_c, debug_led3, reset_all_w;
    wire [3:0]reset_clk_counter;   // src/top.v(242[10:27])
    
    wire reset_all, reset_per_frame, buffer_switch_done, dc32_fifo_full, 
        line_of_data_available;
    wire [31:0]dc32_fifo_data_in;   // src/top.v(574[13:30])
    
    wire dc32_fifo_empty, dc32_fifo_read_enable;
    wire [31:0]dc32_fifo_data_out;   // src/top.v(484[23:41])
    
    wire sc32_fifo_write_enable, sc32_fifo_read_enable;
    wire [3:0]state;   // src/timing_controller.v(78[11:16])
    wire [31:0]sc32_fifo_data_out;   // src/top.v(646[12:30])
    
    wire sc32_fifo_almost_empty;
    wire [7:0]pc_data_rx;   // src/top.v(809[11:21])
    
    wire tx_uart_active_flag, spi_start_transfer_r, multi_byte_spi_trans_flag_r;
    wire [7:0]tx_addr_byte;   // src/top.v(931[11:23])
    wire [7:0]tx_data_byte;   // src/top.v(933[11:23])
    wire [7:0]rx_buf_byte;   // src/top.v(940[11:22])
    
    wire is_tx_fifo_full_flag, fifo_write_cmd, spi_rx_byte_ready, fifo_read_cmd, 
        is_fifo_empty_flag;
    wire [31:0]fifo_temp_output;   // src/top.v(1030[12:28])
    
    wire even_byte_flag, uart_rx_complete_rising_edge, uart_rx_complete_prev, 
        get_next_word, dc32_fifo_almost_full, reset_all_w_N_61, start_tx_N_64, 
        pll_clk_unbuf, multi_byte_spi_trans_flag_r_N_72, \REG.mem_11_19 , 
        \REG.mem_11_18 , \REG.mem_11_17 , \REG.mem_11_16 , \REG.mem_11_15 , 
        \REG.mem_11_14 , \REG.mem_11_13 , \REG.mem_11_12 , \REG.mem_11_11 , 
        \REG.mem_11_10 , \REG.mem_11_9 , \REG.mem_11_8 , \REG.mem_11_7 , 
        \REG.mem_11_6 , \REG.mem_11_5 , \REG.mem_11_4 , \REG.mem_23_17 , 
        \REG.mem_23_16 , \REG.mem_23_15 , \REG.mem_23_14 , \REG.mem_23_13 , 
        \REG.mem_23_12 , \REG.mem_23_11 , \REG.mem_23_10 , \REG.mem_23_9 , 
        \REG.mem_23_8 , \REG.mem_23_7 , \REG.mem_23_6 , \REG.mem_23_5 , 
        \REG.mem_23_4 , \REG.mem_23_3 , \REG.mem_23_2 , \REG.mem_23_1 , 
        \REG.mem_23_0 , \REG.mem_22_31 , \REG.mem_22_30 , \REG.mem_22_29 , 
        \REG.mem_22_28 , \REG.mem_22_27 , \REG.mem_22_26 , \REG.mem_22_25 , 
        \REG.mem_22_24 , \REG.mem_22_23 , \REG.mem_11_3 , \REG.mem_11_2 , 
        \REG.mem_11_1 , \REG.mem_11_0 , \REG.mem_22_22 , \REG.mem_22_21 , 
        \REG.mem_22_20 , \REG.mem_22_19 , \REG.mem_22_18 , \REG.mem_22_17 , 
        \REG.mem_22_16 , \REG.mem_22_15 , \REG.mem_22_14 , \REG.mem_22_13 , 
        \REG.mem_22_12 , \REG.mem_22_11 , \REG.mem_22_10 , \REG.mem_22_9 , 
        \REG.mem_22_8 , \REG.mem_22_7 , \REG.mem_22_6 , \REG.mem_22_5 , 
        \REG.mem_22_4 , \REG.mem_22_3 , \REG.mem_22_2 , \REG.mem_22_1 , 
        \REG.mem_22_0 , \REG.mem_21_31 , \REG.mem_21_30 , \REG.mem_21_29 , 
        \REG.mem_21_28 , \REG.mem_21_27 , \REG.mem_21_26 , \REG.mem_21_25 , 
        \REG.mem_21_24 , \REG.mem_21_23 , \REG.mem_21_22 , \REG.mem_21_21 , 
        \REG.mem_21_20 , \REG.mem_21_19 , \REG.mem_21_18 , \REG.mem_21_17 , 
        \REG.mem_21_16 , \REG.mem_21_15 , \REG.mem_21_14 , \REG.mem_21_13 , 
        \REG.mem_21_12 , \REG.mem_21_11 , \REG.mem_21_10 , \REG.mem_21_9 , 
        \REG.mem_21_8 , \REG.mem_21_7 , \REG.mem_21_6 , \REG.mem_21_5 , 
        \REG.mem_21_4 , \REG.mem_21_3 , \REG.mem_21_2 , \REG.mem_21_1 , 
        \REG.mem_21_0 , buffer_switch_done_latched, n1224, n12, n14076, 
        n2438, FT_OE_N_496, n2555, n15935, n910, n5390, n5391, 
        n5392, n5412, n5411, n5410, n5409, n5408, n5407, n5406, 
        n5405, n5703, bluejay_data_out_31__N_919, bluejay_data_out_31__N_920, 
        bluejay_data_out_31__N_921, bluejay_data_out_31__N_922, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // src/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main_adj_1451;   // src/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_1453;   // src/uart_tx.v(33[16:27])
    wire [7:0]r_Tx_Data;   // src/uart_tx.v(34[16:25])
    wire [2:0]r_SM_Main_2__N_1029;
    wire [2:0]r_SM_Main_2__N_1026;
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    wire [15:0]rx_shift_reg;   // src/spi.v(72[12:24])
    
    wire n2283, \REG.mem_11_31 , \REG.mem_11_30 , \REG.mem_11_29 , \REG.mem_11_28 , 
        \REG.mem_11_27 , \REG.mem_11_26 , \REG.mem_11_25 , \REG.mem_11_24 , 
        \REG.mem_11_23 , n5414, n5664, n5658, \REG.mem_11_22 , n5386, 
        \REG.mem_11_21 , \REG.mem_11_20 ;
    wire [5:0]wr_addr_r;   // src/fifo_dc_32_lut_gen.v(196[29:38])
    wire [5:0]wr_addr_nxt_c;   // src/fifo_dc_32_lut_gen.v(198[29:42])
    wire [5:0]wr_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(200[30:42])
    wire [5:0]rp_sync1_r;   // src/fifo_dc_32_lut_gen.v(201[37:47])
    wire [5:0]wr_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(204[37:51])
    wire [5:0]wp_sync1_r;   // src/fifo_dc_32_lut_gen.v(222[37:47])
    wire [5:0]rd_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(225[37:51])
    
    wire wr_fifo_en_w, rd_fifo_en_w, \aempty_flag_impl.ae_flag_nxt_w ;
    wire [5:0]rd_addr_nxt_c_5__N_573;
    
    wire empty_nxt_c_N_636, \REG.mem_7_31 , \REG.mem_7_30 , \REG.mem_7_29 , 
        \REG.mem_7_28 , \REG.mem_7_27 , \REG.mem_7_26 , \REG.mem_7_25 , 
        \REG.mem_7_24 , \REG.mem_7_23 , \REG.mem_7_22 , \REG.mem_7_21 , 
        \REG.mem_7_20 , \REG.mem_7_19 , \REG.mem_7_18 , \REG.mem_7_17 , 
        \REG.mem_7_16 , \REG.mem_7_15 , \REG.mem_7_14 , \REG.mem_7_13 , 
        \REG.mem_7_12 , \REG.mem_7_11 , \REG.mem_7_10 , \REG.mem_7_9 , 
        \MISC.empty_flag_r , n5413, n5385, n32, \REG.mem_7_8 , \REG.mem_7_7 , 
        \REG.mem_7_6 , \REG.mem_7_5 , \REG.mem_7_4 , \REG.mem_7_3 , 
        \REG.mem_7_2 , \REG.mem_7_1 , \REG.mem_7_0 , \REG.mem_6_31 , 
        \REG.mem_6_30 , \REG.mem_6_29 , \REG.mem_6_28 , \REG.mem_6_27 , 
        \REG.mem_6_26 , \REG.mem_6_25 , \REG.mem_6_24 , \REG.mem_6_23 , 
        \REG.mem_6_22 , \REG.mem_6_21 , \REG.mem_6_20 , \REG.mem_6_19 , 
        \REG.mem_6_18 , \REG.mem_6_17 , \REG.mem_6_16 , \REG.mem_6_15 , 
        \REG.mem_6_14 , \REG.mem_6_13 , \REG.mem_6_12 , \REG.mem_6_11 , 
        \REG.mem_6_10 , \REG.mem_6_9 , n5403, wr_fifo_en_w_adj_1412, 
        rd_fifo_en_w_adj_1413;
    wire [2:0]wr_addr_r_adj_1502;   // src/fifo_quad_word_mod.v(65[31:40])
    wire [2:0]wr_addr_p1_w_adj_1504;   // src/fifo_quad_word_mod.v(67[32:44])
    wire [2:0]rd_addr_r_adj_1505;   // src/fifo_quad_word_mod.v(69[31:40])
    wire [2:0]rd_addr_p1_w_adj_1507;   // src/fifo_quad_word_mod.v(71[32:44])
    
    wire n3414;
    wire [31:0]\mem_LUT.data_raw_r ;   // src/fifo_quad_word_mod.v(449[42:52])
    
    wire \REG.mem_6_8 , \REG.mem_6_7 , \REG.mem_6_6 , \REG.mem_6_5 , 
        \REG.mem_6_4 , \REG.mem_6_3 , \REG.mem_6_2 , \REG.mem_6_1 , 
        \REG.mem_6_0 , \REG.mem_5_31 , \REG.mem_5_30 , \REG.mem_5_29 , 
        \REG.mem_5_28 , \REG.mem_5_27 , \REG.mem_5_26 , \REG.mem_5_25 , 
        \REG.mem_5_24 , \REG.mem_5_23 , \REG.mem_5_22 , \REG.mem_5_21 , 
        \REG.mem_5_20 , \REG.mem_5_19 , \REG.mem_5_18 , \REG.mem_5_17 , 
        \REG.mem_5_16 , \REG.mem_5_15 , \REG.mem_5_14 , \REG.mem_5_13 , 
        \REG.mem_5_12 , \REG.mem_5_11 , \REG.mem_5_10 , \REG.mem_5_9 , 
        \REG.mem_5_8 , \REG.mem_5_7 , \REG.mem_5_6 , \REG.mem_5_5 , 
        \REG.mem_5_4 , \REG.mem_5_3 , \REG.mem_5_2 , \REG.mem_5_1 , 
        \REG.mem_5_0 , n3531, n8, n14096, n5648, n5647, n5207, 
        n989, n1028, n5431, n5642, n2178, \REG.mem_23_31 , \REG.mem_23_30 , 
        \REG.mem_23_29 , \REG.mem_23_28 , \REG.mem_23_27 , \REG.mem_23_26 , 
        \REG.mem_23_25 , \REG.mem_23_24 , \REG.mem_23_23 , \REG.mem_23_22 , 
        \REG.mem_23_21 , \REG.mem_23_20 , \REG.mem_23_19 , \REG.mem_23_18 , 
        n14298, n5639, \REG.mem_27_0 , \REG.mem_27_1 , \REG.mem_27_2 , 
        \REG.mem_27_3 , \REG.mem_27_4 , \REG.mem_27_5 , \REG.mem_27_6 , 
        \REG.mem_27_7 , \REG.mem_27_8 , \REG.mem_27_9 , \REG.mem_27_10 , 
        \REG.mem_27_11 , \REG.mem_27_12 , \REG.mem_27_13 , \REG.mem_27_14 , 
        \REG.mem_27_15 , \REG.mem_27_16 , \REG.mem_27_17 , \REG.mem_27_18 , 
        \REG.mem_27_19 , \REG.mem_27_20 , \REG.mem_27_21 , \REG.mem_27_22 , 
        \REG.mem_27_23 , \REG.mem_27_24 , \REG.mem_27_25 , \REG.mem_27_26 , 
        \REG.mem_27_27 , \REG.mem_27_28 , \REG.mem_27_29 , \REG.mem_27_30 , 
        \REG.mem_27_31 , n6, n10, n11, n12_adj_1415, n22, n26, 
        n27, n28, n10059, n10051, n14706, n14692, n9873, n14690, 
        n14688, n14684, n7067, n7064, n7061, n7058, n7055, n7052, 
        n7049, n7038, n7037, n7036, n7035, n7034, n7033, n7032, 
        n7031, n7030, n7029, n7028, n7027, n7025, n7023, n7022, 
        n7021, n7020, n7019, n7018, n7017, n7016, n7015, n7014, 
        n7013, n7012, n7011, n7010, n7009, n7008, n7007, n7006, 
        n7005, n7004, n7003, n7002, n7001, n7000, n6999, n6998, 
        n6997, n6996, n6995, n6994, n6993, n6992, n6991, n6990, 
        n6989, n6988, n6987, n6986, n14118, n6982, n6981, n6977, 
        n6974, n14710, n6970, n6964, n6963, n6962, n6961, n6960, 
        n6959, n6958, n6957, n6955, n6953, n6532, n6531, n6530, 
        n6529, n6528, n6527, n6526, n6525, n6524, n6523, n6522, 
        n6521, n6520, n6519, n6518, n6517, n6516, n6515, n6514, 
        n6513, n6512, n6511, n6510, n6509, n6508, n6507, n6506, 
        n6505, n6504, n6503, n6502, n6501, n6404, n6403, n6402, 
        n6401, n6400, n6399, n6398, n6397, n6396, n6395, n6394, 
        n6393, n6392, n6391, n6390, n6389, n6388, n6387, n6386, 
        n6385, n6384, n6383, n6382, n6381, n6380, n6379, n6378, 
        n6377, n6376, n6375, n6374, n6373, n6372, n6371, n6370, 
        n6369, n6368, n6367, n6366, n6365, n6364, n6363, n6362, 
        n6361, n6360, n6359, n6358, n6357, n6356, n6355, n6354, 
        n6353, n6352, n6351, n6350, n6349, n6348, n6347, n6346, 
        n6345, n6344, n6343, n6342, n6341, n6340, n6339, n6338, 
        n6337, n6336, n6335, n6334, n6333, n6332, n6331, n6330, 
        n6329, n6328, n6327, n6326, n6325, n6324, n6323, n6322, 
        n6321, n6320, n6319, n6318, n6317, n6316, n6315, n6314, 
        n6313, n6312, n6311, n6310, n6309, n6020, n6019, n6018, 
        n6017, n6016, n6015, n6014, n6013, n6012, n6011, n6010, 
        n6009, n6008, n6007, n6006, n6005, n6004, n6003, n6002, 
        n6001, n6000, n5999, n5998, n5997, n5996, n5995, n5994, 
        n5993, n5992, n5991, n5990, n5989, n5638, n5636, n5384, 
        n5387, n5388, n5398, n5399, n5629, n5628, n63, n5400, 
        n5394, n5395, n5892, n5891, n5890, n5889, n14672, n5888, 
        n5887, n5886, n5624, n5885, n5884, n5883, n5882, n5881, 
        n5880, n5879, n5878, n5877, n5876, n5875, n5874, n5873, 
        n5872, n5871, n5870, n5869, n5868, n5867, n5866, n5865, 
        n5864, n5863, n5862, n5861, n4, n5860, n5859, n5858, 
        n5857, n5856, n5855, n5854, n5853, n5852, n5851, n5850, 
        n5849, n5848, n5847, n5846, n5845, n5844, n5843, n5842, 
        n5841, n5840, n5839, n5838, n5837, n5836, n5835, n5834, 
        n5620, n5618, n5833, n5077, n5832, n5831, n5830, n5829, 
        n5828, n5614, n4_adj_1416, n5827, n5826, n5613, n5825, 
        n5824, n5823, n4_adj_1417, n5822, n5821, n5820, n5819, 
        n5818, n5817, n5816, n5815, n5814, n5813, n5812, n5811, 
        n5810, n5809, n5808, n5807, n5806, n5805, n5804, n5803, 
        n5389, n5043, n5802, n5801, n5800, n14508, n5799, n5798, 
        n5797, n5401, n5612, n5611, n5609, n5608, n5605, n25, 
        n5025, n2, n3, n4_adj_1418, n5, n6_adj_1419, n7, n8_adj_1420, 
        n9, n10_adj_1421, n11_adj_1422, n12_adj_1423, n13, n14, 
        n15, n16, n17, n18, n19, n20, n21, n22_adj_1424, n23, 
        n24, n25_adj_1425, n14567, n14657, n106, n107, n108, n109, 
        n110, n111, n112, n113, n114, n115, n116, n117, n118, 
        n119, n120, n121, n122, n123, n124, n125, n126, n127, 
        n128, n129, n130, n13865, n5397, n5396, n14482, n9752, 
        n5404, n4999, n4086, n5393, n14116, n13776, n13775, n13774, 
        n13773, n13772, n13771, n13770, n13769, n13768, n13767, 
        n13766, n13765, n13764, n13763, n13762, n13761, n13760, 
        n13759, n8_adj_1426, n13758, n13757, n13756, n7_adj_1427, 
        n13755, n13754, n13753, n2_adj_1428, n14603, n4843, n13820, 
        n5529, n15_adj_1429, n5528, n5597, n5418, n25_adj_1430, 
        n4435, n5402, n4942, n4938, n4935, n4566, n4_adj_1431, 
        n14647, n14542, n13902, n13900, n13898, n18034;
    
    VCC i2 (.Y(VCC_net));
    timing_controller timing_controller_inst (.SLM_CLK_c(SLM_CLK_c), .sc32_fifo_write_enable(sc32_fifo_write_enable), 
            .sc32_fifo_read_enable(sc32_fifo_read_enable), .n14567(n14567), 
            .state({state}), .dc32_fifo_read_enable(dc32_fifo_read_enable), 
            .buffer_switch_done(buffer_switch_done), .n5043(n5043), .GND_net(GND_net), 
            .VCC_net(VCC_net), .n2283(n2283), .n14118(n14118), .n1224(n1224), 
            .n63(n63), .n5077(n5077), .line_of_data_available(line_of_data_available), 
            .n2178(n2178), .INVERT_c_4(INVERT_c_4), .n7(n7_adj_1427), 
            .n8(n8_adj_1426), .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .get_next_word(get_next_word), .dc32_fifo_full(dc32_fifo_full), 
            .reset_all(reset_all), .n9752(n9752), .n10059(n10059), .n14542(n14542), 
            .reset_per_frame(reset_per_frame), .n25(n25_adj_1430), .UPDATE_c_3(UPDATE_c_3), 
            .n14692(n14692), .n10051(n10051), .n4843(n4843), .n910(n910), 
            .n989(n989), .n1028(n1028), .buffer_switch_done_latched(buffer_switch_done_latched), 
            .n14482(n14482), .n5529(n5529), .bluejay_data_out_31__N_920(bluejay_data_out_31__N_920), 
            .n5528(n5528), .bluejay_data_out_31__N_919(bluejay_data_out_31__N_919), 
            .n5431(n5431)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(473[19] 494[2])
    SB_DFF uart_rx_complete_prev_83 (.Q(uart_rx_complete_prev), .C(SLM_CLK_c), 
           .D(debug_led3));   // src/top.v(1189[8] 1195[4])
    bluejay_data bluejay_data_inst (.DEBUG_6_c(DEBUG_6_c), .SLM_CLK_c(SLM_CLK_c), 
            .buffer_switch_done(buffer_switch_done), .buffer_switch_done_latched(buffer_switch_done_latched), 
            .GND_net(GND_net), .n910(n910), .line_of_data_available(line_of_data_available), 
            .n989(n989), .bluejay_data_out_31__N_921(bluejay_data_out_31__N_921), 
            .bluejay_data_out_31__N_920(bluejay_data_out_31__N_920), .bluejay_data_out_31__N_922(bluejay_data_out_31__N_922), 
            .n5043(n5043), .n14482(n14482), .n6982(n6982), .DEBUG_8_c(DEBUG_8_c), 
            .n5431(n5431), .VCC_net(VCC_net), .DATA10_c_10(DATA10_c_10), 
            .n5414(n5414), .DATA9_c_9(DATA9_c_9), .n5413(n5413), .DATA11_c_11(DATA11_c_11), 
            .n5412(n5412), .DATA12_c_12(DATA12_c_12), .n5411(n5411), .n14298(n14298), 
            .n1028(n1028), .bluejay_data_out_31__N_919(bluejay_data_out_31__N_919), 
            .SYNC_c(SYNC_c), .DATA13_c_13(DATA13_c_13), .n5410(n5410), 
            .DATA14_c_14(DATA14_c_14), .n5409(n5409), .DATA8_c_8(DATA8_c_8), 
            .n5408(n5408), .DATA15_c_15(DATA15_c_15), .n5407(n5407), .DATA16_c_16(DATA16_c_16), 
            .n5406(n5406), .DATA7_c_7(DATA7_c_7), .n5405(n5405), .DATA17_c_17(DATA17_c_17), 
            .n5404(n5404), .DATA18_c_18(DATA18_c_18), .n5403(n5403), .DATA6_c_6(DATA6_c_6), 
            .n5402(n5402), .DATA19_c_19(DATA19_c_19), .n5401(n5401), .DATA20_c_20(DATA20_c_20), 
            .n5400(n5400), .DATA5_c_5(DATA5_c_5), .n5399(n5399), .DATA21_c_21(DATA21_c_21), 
            .n5398(n5398), .DATA22_c_22(DATA22_c_22), .n5397(n5397), .DATA4_c_4(DATA4_c_4), 
            .n5396(n5396), .DATA23_c_23(DATA23_c_23), .n5395(n5395), .DATA24_c_24(DATA24_c_24), 
            .n5394(n5394), .n5529(n5529), .n5528(n5528), .DATA3_c_3(DATA3_c_3), 
            .n5393(n5393), .get_next_word(get_next_word), .DATA25_c_25(DATA25_c_25), 
            .n5392(n5392), .DATA26_c_26(DATA26_c_26), .n5391(n5391), .DATA2_c_2(DATA2_c_2), 
            .n5390(n5390), .DATA27_c_27(DATA27_c_27), .n5389(n5389), .DATA28_c_28(DATA28_c_28), 
            .n5388(n5388), .DATA1_c_1(DATA1_c_1), .n5387(n5387), .DATA29_c_29(DATA29_c_29), 
            .n5386(n5386), .DATA30_c_30(DATA30_c_30), .n5385(n5385), .DATA31_c_31(DATA31_c_31), 
            .n5384(n5384), .sc32_fifo_almost_empty(sc32_fifo_almost_empty)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(750[14] 763[2])
    SB_GB clk_gb (.GLOBAL_BUFFER_OUTPUT(SLM_CLK_c), .USER_SIGNAL_TO_GLOBAL_BUFFER(pll_clk_unbuf)) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/clock.v(82[7:96])
    SB_IO UART_TX_pad (.PACKAGE_PIN(UART_TX), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_1_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_TX_pad.PIN_TYPE = 6'b011001;
    defparam UART_TX_pad.PULLUP = 1'b0;
    defparam UART_TX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_TX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4815_3_lut (.I0(\REG.mem_21_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6314));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4816_3_lut (.I0(\REG.mem_21_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6315));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4817_3_lut (.I0(\REG.mem_21_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6316));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4818_3_lut (.I0(\REG.mem_21_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6317));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4819_3_lut (.I0(\REG.mem_21_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6318));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4820_3_lut (.I0(\REG.mem_21_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6319));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4821_3_lut (.I0(\REG.mem_21_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6320));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4822_3_lut (.I0(\REG.mem_21_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6321));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4823_3_lut (.I0(\REG.mem_21_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6322));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4824_3_lut (.I0(\REG.mem_21_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6323));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4825_3_lut (.I0(\REG.mem_21_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6324));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4826_3_lut (.I0(\REG.mem_21_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6325));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4827_3_lut (.I0(\REG.mem_21_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6326));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4828_3_lut (.I0(\REG.mem_21_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6327));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4829_3_lut (.I0(\REG.mem_21_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6328));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4830_3_lut (.I0(\REG.mem_21_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6329));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4831_3_lut (.I0(\REG.mem_21_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6330));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4832_3_lut (.I0(\REG.mem_21_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6331));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4833_3_lut (.I0(\REG.mem_21_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6332));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4834_3_lut (.I0(\REG.mem_21_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6333));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4835_3_lut (.I0(\REG.mem_21_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6334));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4836_3_lut (.I0(\REG.mem_21_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6335));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4837_3_lut (.I0(\REG.mem_21_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6336));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4838_3_lut (.I0(\REG.mem_21_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6337));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4839_3_lut (.I0(\REG.mem_21_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6338));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4840_3_lut (.I0(\REG.mem_21_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6339));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4840_3_lut.LUT_INIT = 16'hcaca;
    SB_IO RST_pad (.PACKAGE_PIN(RST), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RST_pad.PIN_TYPE = 6'b011001;
    defparam RST_pad.PULLUP = 1'b0;
    defparam RST_pad.NEG_TRIGGER = 1'b0;
    defparam RST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CTS_pad (.PACKAGE_PIN(CTS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CTS_pad.PIN_TYPE = 6'b011001;
    defparam CTS_pad.PULLUP = 1'b0;
    defparam CTS_pad.NEG_TRIGGER = 1'b0;
    defparam CTS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4841_3_lut (.I0(\REG.mem_21_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6340));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4842_3_lut (.I0(\REG.mem_22_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n11), .I3(GND_net), .O(n6341));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4842_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DTR_pad (.PACKAGE_PIN(DTR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DTR_pad.PIN_TYPE = 6'b011001;
    defparam DTR_pad.PULLUP = 1'b0;
    defparam DTR_pad.NEG_TRIGGER = 1'b0;
    defparam DTR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DSR_pad (.PACKAGE_PIN(DSR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DSR_pad.PIN_TYPE = 6'b011001;
    defparam DSR_pad.PULLUP = 1'b0;
    defparam DSR_pad.NEG_TRIGGER = 1'b0;
    defparam DSR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4843_3_lut (.I0(\REG.mem_22_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n11), .I3(GND_net), .O(n6342));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4844_3_lut (.I0(\REG.mem_22_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n11), .I3(GND_net), .O(n6343));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4844_3_lut.LUT_INIT = 16'hcaca;
    SB_IO SEN_pad (.PACKAGE_PIN(SEN), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SEN_c_1)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SEN_pad.PIN_TYPE = 6'b011001;
    defparam SEN_pad.PULLUP = 1'b0;
    defparam SEN_pad.NEG_TRIGGER = 1'b0;
    defparam SEN_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4845_3_lut (.I0(\REG.mem_22_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n11), .I3(GND_net), .O(n6344));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4846_3_lut (.I0(\REG.mem_22_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n11), .I3(GND_net), .O(n6345));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4847_3_lut (.I0(\REG.mem_22_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n11), .I3(GND_net), .O(n6346));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4848_3_lut (.I0(\REG.mem_22_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n11), .I3(GND_net), .O(n6347));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4849_3_lut (.I0(\REG.mem_22_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n11), .I3(GND_net), .O(n6348));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4850_3_lut (.I0(\REG.mem_22_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n11), .I3(GND_net), .O(n6349));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4851_3_lut (.I0(\REG.mem_22_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n11), .I3(GND_net), .O(n6350));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4852_3_lut (.I0(\REG.mem_22_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n11), .I3(GND_net), .O(n6351));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4852_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_all_r_77 (.Q(reset_all_w), .C(SLM_CLK_c), .D(reset_all_w_N_61));   // src/top.v(246[8] 264[4])
    SB_LUT4 i4853_3_lut (.I0(\REG.mem_22_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n11), .I3(GND_net), .O(n6352));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4854_3_lut (.I0(\REG.mem_22_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n11), .I3(GND_net), .O(n6353));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4855_3_lut (.I0(\REG.mem_22_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n11), .I3(GND_net), .O(n6354));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4856_3_lut (.I0(\REG.mem_22_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n11), .I3(GND_net), .O(n6355));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4857_3_lut (.I0(\REG.mem_22_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n11), .I3(GND_net), .O(n6356));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4858_3_lut (.I0(\REG.mem_22_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n11), .I3(GND_net), .O(n6357));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4859_3_lut (.I0(\REG.mem_22_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n11), .I3(GND_net), .O(n6358));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4860_3_lut (.I0(\REG.mem_22_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n11), .I3(GND_net), .O(n6359));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4861_3_lut (.I0(\REG.mem_22_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n11), .I3(GND_net), .O(n6360));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4862_3_lut (.I0(\REG.mem_22_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n11), .I3(GND_net), .O(n6361));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4863_3_lut (.I0(\REG.mem_22_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n11), .I3(GND_net), .O(n6362));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12535_2_lut (.I0(tx_data_byte[5]), .I1(tx_data_byte[7]), .I2(GND_net), 
            .I3(GND_net), .O(n14657));
    defparam i12535_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12587_4_lut (.I0(tx_data_byte[3]), .I1(tx_data_byte[2]), .I2(tx_data_byte[4]), 
            .I3(n14657), .O(n14710));
    defparam i12587_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i13957_4_lut (.I0(tx_data_byte[0]), .I1(tx_data_byte[1]), .I2(tx_data_byte[6]), 
            .I3(n14710), .O(multi_byte_spi_trans_flag_r_N_72));   // src/top.v(1247[10:31])
    defparam i13957_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i4864_3_lut (.I0(\REG.mem_22_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n11), .I3(GND_net), .O(n6363));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4865_3_lut (.I0(\REG.mem_22_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n11), .I3(GND_net), .O(n6364));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4866_3_lut (.I0(\REG.mem_22_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n11), .I3(GND_net), .O(n6365));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4867_3_lut (.I0(\REG.mem_22_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n11), .I3(GND_net), .O(n6366));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4868_3_lut (.I0(\REG.mem_22_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n11), .I3(GND_net), .O(n6367));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4868_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DCD_pad (.PACKAGE_PIN(DCD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DCD_pad.PIN_TYPE = 6'b011001;
    defparam DCD_pad.PULLUP = 1'b0;
    defparam DCD_pad.NEG_TRIGGER = 1'b0;
    defparam DCD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SCK_pad (.PACKAGE_PIN(SCK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SCK_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SCK_pad.PIN_TYPE = 6'b011001;
    defparam SCK_pad.PULLUP = 1'b0;
    defparam SCK_pad.NEG_TRIGGER = 1'b0;
    defparam SCK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4869_3_lut (.I0(\REG.mem_22_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n11), .I3(GND_net), .O(n6368));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4870_3_lut (.I0(\REG.mem_22_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n11), .I3(GND_net), .O(n6369));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4871_3_lut (.I0(\REG.mem_22_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n11), .I3(GND_net), .O(n6370));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4872_3_lut (.I0(\REG.mem_22_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n11), .I3(GND_net), .O(n6371));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4873_3_lut (.I0(\REG.mem_22_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n11), .I3(GND_net), .O(n6372));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4874_3_lut (.I0(\REG.mem_23_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n10), .I3(GND_net), .O(n6373));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4875_3_lut (.I0(\REG.mem_23_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n10), .I3(GND_net), .O(n6374));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4876_3_lut (.I0(\REG.mem_23_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n10), .I3(GND_net), .O(n6375));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4877_3_lut (.I0(\REG.mem_23_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n10), .I3(GND_net), .O(n6376));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4878_3_lut (.I0(\REG.mem_23_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n10), .I3(GND_net), .O(n6377));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4879_3_lut (.I0(\REG.mem_23_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n10), .I3(GND_net), .O(n6378));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4880_3_lut (.I0(\REG.mem_23_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n10), .I3(GND_net), .O(n6379));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4881_3_lut (.I0(\REG.mem_23_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n10), .I3(GND_net), .O(n6380));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4882_3_lut (.I0(\REG.mem_23_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n10), .I3(GND_net), .O(n6381));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4883_3_lut (.I0(\REG.mem_23_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n10), .I3(GND_net), .O(n6382));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19_4_lut (.I0(n4843), .I1(n15935), .I2(state[3]), .I3(n63), 
            .O(n14118));   // src/timing_controller.v(153[8] 229[4])
    defparam i19_4_lut.LUT_INIT = 16'hfcac;
    SB_LUT4 i4884_3_lut (.I0(\REG.mem_23_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n10), .I3(GND_net), .O(n6383));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4885_3_lut (.I0(\REG.mem_23_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n10), .I3(GND_net), .O(n6384));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4886_3_lut (.I0(\REG.mem_23_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n10), .I3(GND_net), .O(n6385));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4098_3_lut (.I0(tx_data_byte[0]), .I1(pc_data_rx[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5597));   // src/top.v(1198[8] 1265[4])
    defparam i4098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4109_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[7]), .I2(r_Bit_Index[0]), 
            .I3(n4935), .O(n5608));   // src/uart_rx.v(49[10] 144[8])
    defparam i4109_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i4110_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[6]), .I2(r_Bit_Index[0]), 
            .I3(n4935), .O(n5609));   // src/uart_rx.v(49[10] 144[8])
    defparam i4110_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4112_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[5]), .I2(n4), 
            .I3(n4942), .O(n5611));   // src/uart_rx.v(49[10] 144[8])
    defparam i4112_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4113_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[4]), .I2(n4), 
            .I3(n4938), .O(n5612));   // src/uart_rx.v(49[10] 144[8])
    defparam i4113_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4114_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[3]), .I2(n4_adj_1417), 
            .I3(n4942), .O(n5613));   // src/uart_rx.v(49[10] 144[8])
    defparam i4114_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4115_3_lut (.I0(tx_addr_byte[0]), .I1(tx_data_byte[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5614));   // src/top.v(1198[8] 1265[4])
    defparam i4115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4119_2_lut (.I0(uart_rx_complete_prev), .I1(debug_led3), .I2(GND_net), 
            .I3(GND_net), .O(n5618));   // src/top.v(1189[8] 1195[4])
    defparam i4119_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4121_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[2]), .I2(n4_adj_1417), 
            .I3(n4938), .O(n5620));   // src/uart_rx.v(49[10] 144[8])
    defparam i4121_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4298_3_lut (.I0(\REG.mem_5_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n28), .I3(GND_net), .O(n5797));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4125_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[1]), .I2(n4_adj_1416), 
            .I3(n4942), .O(n5624));   // src/uart_rx.v(49[10] 144[8])
    defparam i4125_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4299_3_lut (.I0(\REG.mem_5_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n28), .I3(GND_net), .O(n5798));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4300_3_lut (.I0(\REG.mem_5_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n28), .I3(GND_net), .O(n5799));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4130_3_lut (.I0(r_Tx_Data[0]), .I1(fifo_temp_output[0]), .I2(n4435), 
            .I3(GND_net), .O(n5629));   // src/uart_tx.v(38[10] 141[8])
    defparam i4130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut (.I0(n63), .I1(state[3]), .I2(state[2]), .I3(n9873), 
            .O(n14542));   // src/timing_controller.v(159[5] 228[12])
    defparam i3_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i4137_3_lut (.I0(rx_buf_byte[0]), .I1(rx_shift_reg[0]), .I2(n4086), 
            .I3(GND_net), .O(n5636));   // src/spi.v(76[8] 221[4])
    defparam i4137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4139_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5638));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4139_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4140_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5639));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4140_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4143_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5642));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4143_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4887_3_lut (.I0(\REG.mem_23_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n10), .I3(GND_net), .O(n6386));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5454_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6953));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i5454_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5456_2_lut (.I0(reset_per_frame), .I1(wr_addr_nxt_c[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6955));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i5456_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5458_3_lut (.I0(tx_data_byte[7]), .I1(pc_data_rx[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6957));   // src/top.v(1198[8] 1265[4])
    defparam i5458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5459_3_lut (.I0(tx_data_byte[6]), .I1(pc_data_rx[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6958));   // src/top.v(1198[8] 1265[4])
    defparam i5459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5460_3_lut (.I0(tx_data_byte[5]), .I1(pc_data_rx[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6959));   // src/top.v(1198[8] 1265[4])
    defparam i5460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5461_3_lut (.I0(tx_data_byte[4]), .I1(pc_data_rx[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6960));   // src/top.v(1198[8] 1265[4])
    defparam i5461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5462_3_lut (.I0(tx_data_byte[3]), .I1(pc_data_rx[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6961));   // src/top.v(1198[8] 1265[4])
    defparam i5462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5463_3_lut (.I0(tx_data_byte[2]), .I1(pc_data_rx[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6962));   // src/top.v(1198[8] 1265[4])
    defparam i5463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5464_3_lut (.I0(tx_data_byte[1]), .I1(pc_data_rx[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6963));   // src/top.v(1198[8] 1265[4])
    defparam i5464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13954_2_lut (.I0(is_fifo_empty_flag), .I1(tx_uart_active_flag), 
            .I2(GND_net), .I3(GND_net), .O(start_tx_N_64));
    defparam i13954_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i4888_3_lut (.I0(\REG.mem_23_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n10), .I3(GND_net), .O(n6387));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4889_3_lut (.I0(\REG.mem_23_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n10), .I3(GND_net), .O(n6388));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n25));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4890_3_lut (.I0(\REG.mem_23_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n10), .I3(GND_net), .O(n6389));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4891_3_lut (.I0(\REG.mem_23_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n10), .I3(GND_net), .O(n6390));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4892_3_lut (.I0(\REG.mem_23_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n10), .I3(GND_net), .O(n6391));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4893_3_lut (.I0(\REG.mem_23_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n10), .I3(GND_net), .O(n6392));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4894_3_lut (.I0(\REG.mem_23_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n10), .I3(GND_net), .O(n6393));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12483_4_lut (.I0(n4566), .I1(fifo_read_cmd), .I2(wr_addr_r_adj_1502[1]), 
            .I3(rd_addr_r_adj_1505[1]), .O(n14603));
    defparam i12483_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i4895_3_lut (.I0(\REG.mem_23_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n10), .I3(GND_net), .O(n6394));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4896_3_lut (.I0(\REG.mem_23_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n10), .I3(GND_net), .O(n6395));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(reset_all_w), .I1(n15_adj_1429), .I2(wr_fifo_en_w_adj_1412), 
            .I3(n13820), .O(n14076));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut.LUT_INIT = 16'h5444;
    SB_LUT4 i4897_3_lut (.I0(\REG.mem_23_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n10), .I3(GND_net), .O(n6396));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4898_3_lut (.I0(\REG.mem_23_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n10), .I3(GND_net), .O(n6397));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4301_3_lut (.I0(\REG.mem_5_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n28), .I3(GND_net), .O(n5800));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5471_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[0]), .I2(\mem_LUT.data_raw_r [0]), 
            .I3(n5207), .O(n6970));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i5471_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i2053_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n3531));   // src/top.v(1198[8] 1265[4])
    defparam i2053_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5475_3_lut (.I0(n14690), .I1(r_Bit_Index_adj_1453[0]), .I2(n14684), 
            .I3(GND_net), .O(n6974));   // src/uart_tx.v(38[10] 141[8])
    defparam i5475_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i5478_3_lut (.I0(n14688), .I1(r_Bit_Index[0]), .I2(n14672), 
            .I3(GND_net), .O(n6977));   // src/uart_rx.v(49[10] 144[8])
    defparam i5478_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i4899_3_lut (.I0(\REG.mem_23_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n10), .I3(GND_net), .O(n6398));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4900_3_lut (.I0(\REG.mem_23_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n10), .I3(GND_net), .O(n6399));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4901_3_lut (.I0(\REG.mem_23_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n10), .I3(GND_net), .O(n6400));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4902_3_lut (.I0(\REG.mem_23_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n10), .I3(GND_net), .O(n6401));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5482_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[0]), .I2(n4_adj_1416), 
            .I3(n4938), .O(n6981));   // src/uart_rx.v(49[10] 144[8])
    defparam i5482_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4903_3_lut (.I0(\REG.mem_23_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n10), .I3(GND_net), .O(n6402));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut (.I0(tx_shift_reg[0]), .I1(n2555), .I2(n4999), .I3(tx_data_byte[0]), 
            .O(n14116));   // src/spi.v(76[8] 221[4])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i4904_3_lut (.I0(\REG.mem_23_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n10), .I3(GND_net), .O(n6403));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5487_3_lut (.I0(tx_addr_byte[7]), .I1(tx_data_byte[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6986));   // src/top.v(1198[8] 1265[4])
    defparam i5487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4905_3_lut (.I0(\REG.mem_23_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n10), .I3(GND_net), .O(n6404));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5488_3_lut (.I0(tx_addr_byte[6]), .I1(tx_data_byte[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6987));   // src/top.v(1198[8] 1265[4])
    defparam i5488_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_addr_byte_r_i0_i1 (.Q(tx_addr_byte[1]), .C(SLM_CLK_c), .D(n6992));   // src/top.v(1198[8] 1265[4])
    SB_DFF tx_addr_byte_r_i0_i2 (.Q(tx_addr_byte[2]), .C(SLM_CLK_c), .D(n6991));   // src/top.v(1198[8] 1265[4])
    SB_DFF tx_addr_byte_r_i0_i3 (.Q(tx_addr_byte[3]), .C(SLM_CLK_c), .D(n6990));   // src/top.v(1198[8] 1265[4])
    SB_DFF tx_addr_byte_r_i0_i4 (.Q(tx_addr_byte[4]), .C(SLM_CLK_c), .D(n6989));   // src/top.v(1198[8] 1265[4])
    SB_DFF tx_addr_byte_r_i0_i5 (.Q(tx_addr_byte[5]), .C(SLM_CLK_c), .D(n6988));   // src/top.v(1198[8] 1265[4])
    SB_DFF tx_addr_byte_r_i0_i6 (.Q(tx_addr_byte[6]), .C(SLM_CLK_c), .D(n6987));   // src/top.v(1198[8] 1265[4])
    SB_DFF tx_addr_byte_r_i0_i7 (.Q(tx_addr_byte[7]), .C(SLM_CLK_c), .D(n6986));   // src/top.v(1198[8] 1265[4])
    SB_DFF spi_start_transfer_r_84 (.Q(spi_start_transfer_r), .C(SLM_CLK_c), 
           .D(n3531));   // src/top.v(1198[8] 1265[4])
    SB_DFF start_tx_81 (.Q(r_SM_Main_2__N_1029[0]), .C(SLM_CLK_c), .D(n6964));   // src/top.v(1034[8] 1052[4])
    SB_DFF tx_data_byte_r_i0_i1 (.Q(tx_data_byte[1]), .C(SLM_CLK_c), .D(n6963));   // src/top.v(1198[8] 1265[4])
    SB_DFF tx_data_byte_r_i0_i2 (.Q(tx_data_byte[2]), .C(SLM_CLK_c), .D(n6962));   // src/top.v(1198[8] 1265[4])
    SB_DFF tx_data_byte_r_i0_i3 (.Q(tx_data_byte[3]), .C(SLM_CLK_c), .D(n6961));   // src/top.v(1198[8] 1265[4])
    SB_DFF tx_data_byte_r_i0_i4 (.Q(tx_data_byte[4]), .C(SLM_CLK_c), .D(n6960));   // src/top.v(1198[8] 1265[4])
    SB_DFF tx_data_byte_r_i0_i5 (.Q(tx_data_byte[5]), .C(SLM_CLK_c), .D(n6959));   // src/top.v(1198[8] 1265[4])
    SB_DFF tx_data_byte_r_i0_i6 (.Q(tx_data_byte[6]), .C(SLM_CLK_c), .D(n6958));   // src/top.v(1198[8] 1265[4])
    SB_DFF tx_data_byte_r_i0_i7 (.Q(tx_data_byte[7]), .C(SLM_CLK_c), .D(n6957));   // src/top.v(1198[8] 1265[4])
    SB_LUT4 i5489_3_lut (.I0(tx_addr_byte[5]), .I1(tx_data_byte[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6988));   // src/top.v(1198[8] 1265[4])
    defparam i5489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5490_3_lut (.I0(tx_addr_byte[4]), .I1(tx_data_byte[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6989));   // src/top.v(1198[8] 1265[4])
    defparam i5490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5491_3_lut (.I0(tx_addr_byte[3]), .I1(tx_data_byte[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6990));   // src/top.v(1198[8] 1265[4])
    defparam i5491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5492_3_lut (.I0(tx_addr_byte[2]), .I1(tx_data_byte[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6991));   // src/top.v(1198[8] 1265[4])
    defparam i5492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5493_3_lut (.I0(tx_addr_byte[1]), .I1(tx_data_byte[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n6992));   // src/top.v(1198[8] 1265[4])
    defparam i5493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5494_3_lut (.I0(r_Tx_Data[1]), .I1(fifo_temp_output[1]), .I2(n4435), 
            .I3(GND_net), .O(n6993));   // src/uart_tx.v(38[10] 141[8])
    defparam i5494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5495_3_lut (.I0(r_Tx_Data[2]), .I1(fifo_temp_output[2]), .I2(n4435), 
            .I3(GND_net), .O(n6994));   // src/uart_tx.v(38[10] 141[8])
    defparam i5495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5496_3_lut (.I0(r_Tx_Data[3]), .I1(fifo_temp_output[3]), .I2(n4435), 
            .I3(GND_net), .O(n6995));   // src/uart_tx.v(38[10] 141[8])
    defparam i5496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5497_3_lut (.I0(r_Tx_Data[4]), .I1(fifo_temp_output[4]), .I2(n4435), 
            .I3(GND_net), .O(n6996));   // src/uart_tx.v(38[10] 141[8])
    defparam i5497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5498_3_lut (.I0(r_Tx_Data[5]), .I1(fifo_temp_output[5]), .I2(n4435), 
            .I3(GND_net), .O(n6997));   // src/uart_tx.v(38[10] 141[8])
    defparam i5498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5499_3_lut (.I0(r_Tx_Data[6]), .I1(fifo_temp_output[6]), .I2(n4435), 
            .I3(GND_net), .O(n6998));   // src/uart_tx.v(38[10] 141[8])
    defparam i5499_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF even_byte_flag_89 (.Q(even_byte_flag), .C(SLM_CLK_c), .D(n3414));   // src/top.v(1198[8] 1265[4])
    SB_LUT4 i5500_3_lut (.I0(r_Tx_Data[7]), .I1(fifo_temp_output[7]), .I2(n4435), 
            .I3(GND_net), .O(n6999));   // src/uart_tx.v(38[10] 141[8])
    defparam i5500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5501_3_lut (.I0(rx_shift_reg[1]), .I1(rx_shift_reg[0]), .I2(n5025), 
            .I3(GND_net), .O(n7000));   // src/spi.v(76[8] 221[4])
    defparam i5501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5502_3_lut (.I0(rx_shift_reg[2]), .I1(rx_shift_reg[1]), .I2(n5025), 
            .I3(GND_net), .O(n7001));   // src/spi.v(76[8] 221[4])
    defparam i5502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5503_3_lut (.I0(rx_shift_reg[3]), .I1(rx_shift_reg[2]), .I2(n5025), 
            .I3(GND_net), .O(n7002));   // src/spi.v(76[8] 221[4])
    defparam i5503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5504_3_lut (.I0(rx_shift_reg[4]), .I1(rx_shift_reg[3]), .I2(n5025), 
            .I3(GND_net), .O(n7003));   // src/spi.v(76[8] 221[4])
    defparam i5504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5505_3_lut (.I0(rx_shift_reg[5]), .I1(rx_shift_reg[4]), .I2(n5025), 
            .I3(GND_net), .O(n7004));   // src/spi.v(76[8] 221[4])
    defparam i5505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5506_3_lut (.I0(rx_shift_reg[6]), .I1(rx_shift_reg[5]), .I2(n5025), 
            .I3(GND_net), .O(n7005));   // src/spi.v(76[8] 221[4])
    defparam i5506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5507_3_lut (.I0(rx_shift_reg[7]), .I1(rx_shift_reg[6]), .I2(n5025), 
            .I3(GND_net), .O(n7006));   // src/spi.v(76[8] 221[4])
    defparam i5507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5508_3_lut (.I0(rx_buf_byte[1]), .I1(rx_shift_reg[1]), .I2(n4086), 
            .I3(GND_net), .O(n7007));   // src/spi.v(76[8] 221[4])
    defparam i5508_3_lut.LUT_INIT = 16'hacac;
    SB_DFF led_counter_1466_1542__i0 (.Q(n25_adj_1425), .C(SLM_CLK_c), .D(n130));   // src/top.v(203[20:35])
    SB_LUT4 i5509_3_lut (.I0(rx_buf_byte[2]), .I1(rx_shift_reg[2]), .I2(n4086), 
            .I3(GND_net), .O(n7008));   // src/spi.v(76[8] 221[4])
    defparam i5509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5510_3_lut (.I0(rx_buf_byte[3]), .I1(rx_shift_reg[3]), .I2(n4086), 
            .I3(GND_net), .O(n7009));   // src/spi.v(76[8] 221[4])
    defparam i5510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5511_3_lut (.I0(rx_buf_byte[4]), .I1(rx_shift_reg[4]), .I2(n4086), 
            .I3(GND_net), .O(n7010));   // src/spi.v(76[8] 221[4])
    defparam i5511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4302_3_lut (.I0(\REG.mem_5_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n28), .I3(GND_net), .O(n5801));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4149_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n5648));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4149_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5512_3_lut (.I0(rx_buf_byte[5]), .I1(rx_shift_reg[5]), .I2(n4086), 
            .I3(GND_net), .O(n7011));   // src/spi.v(76[8] 221[4])
    defparam i5512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5513_3_lut (.I0(rx_buf_byte[6]), .I1(rx_shift_reg[6]), .I2(n4086), 
            .I3(GND_net), .O(n7012));   // src/spi.v(76[8] 221[4])
    defparam i5513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut (.I0(state[3]), .I1(n63), .I2(n14692), .I3(GND_net), 
            .O(n5077));   // src/timing_controller.v(153[8] 229[4])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i13896_3_lut_4_lut (.I0(state[3]), .I1(n63), .I2(state[2]), 
            .I3(n9873), .O(n15935));   // src/timing_controller.v(153[8] 229[4])
    defparam i13896_3_lut_4_lut.LUT_INIT = 16'hb000;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[3]), .I1(n63), .I2(state[2]), .I3(state[1]), 
            .O(n14567));   // src/timing_controller.v(153[8] 229[4])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i4303_3_lut (.I0(\REG.mem_5_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n28), .I3(GND_net), .O(n5802));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4304_3_lut (.I0(\REG.mem_5_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n28), .I3(GND_net), .O(n5803));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4304_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_1467__i0 (.Q(reset_clk_counter[0]), .C(SLM_CLK_c), 
           .D(n25));   // src/top.v(259[27:51])
    SB_LUT4 i5514_3_lut (.I0(rx_buf_byte[7]), .I1(rx_shift_reg[7]), .I2(n4086), 
            .I3(GND_net), .O(n7013));   // src/spi.v(76[8] 221[4])
    defparam i5514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5515_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n7014));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5515_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5516_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n7015));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5516_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4305_3_lut (.I0(\REG.mem_5_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n28), .I3(GND_net), .O(n5804));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4306_3_lut (.I0(\REG.mem_5_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n28), .I3(GND_net), .O(n5805));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4307_3_lut (.I0(\REG.mem_5_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n28), .I3(GND_net), .O(n5806));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8271_1_lut (.I0(n2178), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n9752));   // src/timing_controller.v(78[11:16])
    defparam i8271_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4308_3_lut (.I0(\REG.mem_5_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n28), .I3(GND_net), .O(n5807));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5517_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7016));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5517_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4309_3_lut (.I0(\REG.mem_5_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n28), .I3(GND_net), .O(n5808));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4310_3_lut (.I0(\REG.mem_5_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n28), .I3(GND_net), .O(n5809));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4311_3_lut (.I0(\REG.mem_5_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n28), .I3(GND_net), .O(n5810));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4312_3_lut (.I0(\REG.mem_5_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n28), .I3(GND_net), .O(n5811));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5518_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n7017));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5518_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5519_2_lut (.I0(reset_per_frame), .I1(rd_grey_sync_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n7018));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5519_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5520_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n7019));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5520_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5521_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n7020));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5521_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5522_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7021));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5522_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5523_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n7022));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5523_2_lut.LUT_INIT = 16'h4444;
    SB_DFFSR multi_byte_spi_trans_flag_r_86 (.Q(multi_byte_spi_trans_flag_r), 
            .C(SLM_CLK_c), .D(multi_byte_spi_trans_flag_r_N_72), .R(n5418));   // src/top.v(1198[8] 1265[4])
    SB_LUT4 i5524_2_lut (.I0(reset_per_frame), .I1(rp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n7023));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i5524_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5526_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_5__N_573[1]), 
            .I2(GND_net), .I3(GND_net), .O(n7025));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i5526_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4313_3_lut (.I0(\REG.mem_5_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n28), .I3(GND_net), .O(n5812));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5528_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_5__N_573[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7027));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i5528_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5529_2_lut (.I0(reset_per_frame), .I1(rd_addr_nxt_c_5__N_573[4]), 
            .I2(GND_net), .I3(GND_net), .O(n7028));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i5529_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5530_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n7029));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5530_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5531_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n7030));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5531_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5532_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7031));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5532_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5533_2_lut (.I0(reset_per_frame), .I1(wr_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n7032));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5533_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5534_2_lut (.I0(reset_per_frame), .I1(wr_addr_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n7033));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5534_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i12525_4_lut (.I0(rd_addr_p1_w_adj_1507[2]), .I1(rd_addr_p1_w_adj_1507[1]), 
            .I2(wr_addr_r_adj_1502[2]), .I3(wr_addr_r_adj_1502[1]), .O(n14647));
    defparam i12525_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_151 (.I0(rd_addr_r_adj_1505[1]), .I1(rd_addr_r_adj_1505[0]), 
            .I2(wr_addr_r_adj_1502[1]), .I3(wr_addr_r_adj_1502[0]), .O(n32));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_151.LUT_INIT = 16'h8421;
    SB_LUT4 i1_4_lut_adj_152 (.I0(n14647), .I1(reset_all_w), .I2(rd_fifo_en_w_adj_1413), 
            .I3(n4566), .O(n4_adj_1431));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_152.LUT_INIT = 16'hdccc;
    SB_LUT4 i2_4_lut (.I0(is_fifo_empty_flag), .I1(n4_adj_1431), .I2(fifo_write_cmd), 
            .I3(n32), .O(n14096));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i2_4_lut.LUT_INIT = 16'hcecc;
    SB_LUT4 i5535_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n7034));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5535_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5536_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n7035));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5536_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5537_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7036));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5537_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4314_3_lut (.I0(\REG.mem_5_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n28), .I3(GND_net), .O(n5813));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4315_3_lut (.I0(\REG.mem_5_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n28), .I3(GND_net), .O(n5814));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5538_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n7037));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5538_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5539_2_lut (.I0(reset_per_frame), .I1(wp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n7038));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i5539_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4316_3_lut (.I0(\REG.mem_5_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n28), .I3(GND_net), .O(n5815));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4317_3_lut (.I0(\REG.mem_5_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n28), .I3(GND_net), .O(n5816));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5550_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[7]), .I2(\mem_LUT.data_raw_r [7]), 
            .I3(n5207), .O(n7049));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i5550_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i5553_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[6]), .I2(\mem_LUT.data_raw_r [6]), 
            .I3(n5207), .O(n7052));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i5553_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i5556_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[5]), .I2(\mem_LUT.data_raw_r [5]), 
            .I3(n5207), .O(n7055));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i5556_4_lut.LUT_INIT = 16'h5044;
    SB_IO SDAT_pad (.PACKAGE_PIN(SDAT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SDAT_c_15)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SDAT_pad.PIN_TYPE = 6'b011001;
    defparam SDAT_pad.PULLUP = 1'b0;
    defparam SDAT_pad.NEG_TRIGGER = 1'b0;
    defparam SDAT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UPDATE_pad (.PACKAGE_PIN(UPDATE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UPDATE_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UPDATE_pad.PIN_TYPE = 6'b011001;
    defparam UPDATE_pad.PULLUP = 1'b0;
    defparam UPDATE_pad.NEG_TRIGGER = 1'b0;
    defparam UPDATE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO RESET_pad (.PACKAGE_PIN(RESET), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(RESET_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RESET_pad.PIN_TYPE = 6'b011001;
    defparam RESET_pad.PULLUP = 1'b0;
    defparam RESET_pad.NEG_TRIGGER = 1'b0;
    defparam RESET_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SLM_CLK_pad (.PACKAGE_PIN(SLM_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SLM_CLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SLM_CLK_pad.PIN_TYPE = 6'b011001;
    defparam SLM_CLK_pad.PULLUP = 1'b0;
    defparam SLM_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam SLM_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INVERT_pad (.PACKAGE_PIN(INVERT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INVERT_c_4)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INVERT_pad.PIN_TYPE = 6'b011001;
    defparam INVERT_pad.PULLUP = 1'b0;
    defparam INVERT_pad.NEG_TRIGGER = 1'b0;
    defparam INVERT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SYNC_pad (.PACKAGE_PIN(SYNC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SYNC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SYNC_pad.PIN_TYPE = 6'b011001;
    defparam SYNC_pad.PULLUP = 1'b0;
    defparam SYNC_pad.NEG_TRIGGER = 1'b0;
    defparam SYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO VALID_pad (.PACKAGE_PIN(VALID), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam VALID_pad.PIN_TYPE = 6'b011001;
    defparam VALID_pad.PULLUP = 1'b0;
    defparam VALID_pad.NEG_TRIGGER = 1'b0;
    defparam VALID_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA31_pad (.PACKAGE_PIN(DATA31), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA31_c_31));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA31_pad.PIN_TYPE = 6'b011001;
    defparam DATA31_pad.PULLUP = 1'b0;
    defparam DATA31_pad.NEG_TRIGGER = 1'b0;
    defparam DATA31_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA0_pad (.PACKAGE_PIN(DATA0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_8_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA0_pad.PIN_TYPE = 6'b011001;
    defparam DATA0_pad.PULLUP = 1'b0;
    defparam DATA0_pad.NEG_TRIGGER = 1'b0;
    defparam DATA0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA30_pad (.PACKAGE_PIN(DATA30), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA30_c_30));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA30_pad.PIN_TYPE = 6'b011001;
    defparam DATA30_pad.PULLUP = 1'b0;
    defparam DATA30_pad.NEG_TRIGGER = 1'b0;
    defparam DATA30_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA29_pad (.PACKAGE_PIN(DATA29), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA29_c_29));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA29_pad.PIN_TYPE = 6'b011001;
    defparam DATA29_pad.PULLUP = 1'b0;
    defparam DATA29_pad.NEG_TRIGGER = 1'b0;
    defparam DATA29_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA1_pad (.PACKAGE_PIN(DATA1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA1_c_1));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA1_pad.PIN_TYPE = 6'b011001;
    defparam DATA1_pad.PULLUP = 1'b0;
    defparam DATA1_pad.NEG_TRIGGER = 1'b0;
    defparam DATA1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA28_pad (.PACKAGE_PIN(DATA28), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA28_c_28));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA28_pad.PIN_TYPE = 6'b011001;
    defparam DATA28_pad.PULLUP = 1'b0;
    defparam DATA28_pad.NEG_TRIGGER = 1'b0;
    defparam DATA28_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA27_pad (.PACKAGE_PIN(DATA27), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA27_c_27));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA27_pad.PIN_TYPE = 6'b011001;
    defparam DATA27_pad.PULLUP = 1'b0;
    defparam DATA27_pad.NEG_TRIGGER = 1'b0;
    defparam DATA27_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA2_pad (.PACKAGE_PIN(DATA2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA2_c_2));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA2_pad.PIN_TYPE = 6'b011001;
    defparam DATA2_pad.PULLUP = 1'b0;
    defparam DATA2_pad.NEG_TRIGGER = 1'b0;
    defparam DATA2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA26_pad (.PACKAGE_PIN(DATA26), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA26_c_26));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA26_pad.PIN_TYPE = 6'b011001;
    defparam DATA26_pad.PULLUP = 1'b0;
    defparam DATA26_pad.NEG_TRIGGER = 1'b0;
    defparam DATA26_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA25_pad (.PACKAGE_PIN(DATA25), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA25_c_25));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA25_pad.PIN_TYPE = 6'b011001;
    defparam DATA25_pad.PULLUP = 1'b0;
    defparam DATA25_pad.NEG_TRIGGER = 1'b0;
    defparam DATA25_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA3_pad (.PACKAGE_PIN(DATA3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA3_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA3_pad.PIN_TYPE = 6'b011001;
    defparam DATA3_pad.PULLUP = 1'b0;
    defparam DATA3_pad.NEG_TRIGGER = 1'b0;
    defparam DATA3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA24_pad (.PACKAGE_PIN(DATA24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA24_c_24));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA24_pad.PIN_TYPE = 6'b011001;
    defparam DATA24_pad.PULLUP = 1'b0;
    defparam DATA24_pad.NEG_TRIGGER = 1'b0;
    defparam DATA24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA23_pad (.PACKAGE_PIN(DATA23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA23_c_23));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA23_pad.PIN_TYPE = 6'b011001;
    defparam DATA23_pad.PULLUP = 1'b0;
    defparam DATA23_pad.NEG_TRIGGER = 1'b0;
    defparam DATA23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA4_pad (.PACKAGE_PIN(DATA4), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA4_c_4));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA4_pad.PIN_TYPE = 6'b011001;
    defparam DATA4_pad.PULLUP = 1'b0;
    defparam DATA4_pad.NEG_TRIGGER = 1'b0;
    defparam DATA4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA22_pad (.PACKAGE_PIN(DATA22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA22_c_22));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA22_pad.PIN_TYPE = 6'b011001;
    defparam DATA22_pad.PULLUP = 1'b0;
    defparam DATA22_pad.NEG_TRIGGER = 1'b0;
    defparam DATA22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA21_pad (.PACKAGE_PIN(DATA21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA21_c_21));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA21_pad.PIN_TYPE = 6'b011001;
    defparam DATA21_pad.PULLUP = 1'b0;
    defparam DATA21_pad.NEG_TRIGGER = 1'b0;
    defparam DATA21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA5_pad (.PACKAGE_PIN(DATA5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA5_c_5));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA5_pad.PIN_TYPE = 6'b011001;
    defparam DATA5_pad.PULLUP = 1'b0;
    defparam DATA5_pad.NEG_TRIGGER = 1'b0;
    defparam DATA5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA20_pad (.PACKAGE_PIN(DATA20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA20_c_20));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA20_pad.PIN_TYPE = 6'b011001;
    defparam DATA20_pad.PULLUP = 1'b0;
    defparam DATA20_pad.NEG_TRIGGER = 1'b0;
    defparam DATA20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA19_pad (.PACKAGE_PIN(DATA19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA19_c_19));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA19_pad.PIN_TYPE = 6'b011001;
    defparam DATA19_pad.PULLUP = 1'b0;
    defparam DATA19_pad.NEG_TRIGGER = 1'b0;
    defparam DATA19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA6_pad (.PACKAGE_PIN(DATA6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA6_c_6));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA6_pad.PIN_TYPE = 6'b011001;
    defparam DATA6_pad.PULLUP = 1'b0;
    defparam DATA6_pad.NEG_TRIGGER = 1'b0;
    defparam DATA6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA18_pad (.PACKAGE_PIN(DATA18), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA18_c_18));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA18_pad.PIN_TYPE = 6'b011001;
    defparam DATA18_pad.PULLUP = 1'b0;
    defparam DATA18_pad.NEG_TRIGGER = 1'b0;
    defparam DATA18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA17_pad (.PACKAGE_PIN(DATA17), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA17_c_17));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA17_pad.PIN_TYPE = 6'b011001;
    defparam DATA17_pad.PULLUP = 1'b0;
    defparam DATA17_pad.NEG_TRIGGER = 1'b0;
    defparam DATA17_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA7_pad (.PACKAGE_PIN(DATA7), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA7_c_7));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA7_pad.PIN_TYPE = 6'b011001;
    defparam DATA7_pad.PULLUP = 1'b0;
    defparam DATA7_pad.NEG_TRIGGER = 1'b0;
    defparam DATA7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA16_pad (.PACKAGE_PIN(DATA16), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA16_c_16));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA16_pad.PIN_TYPE = 6'b011001;
    defparam DATA16_pad.PULLUP = 1'b0;
    defparam DATA16_pad.NEG_TRIGGER = 1'b0;
    defparam DATA16_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA15_pad (.PACKAGE_PIN(DATA15), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA15_c_15));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA15_pad.PIN_TYPE = 6'b011001;
    defparam DATA15_pad.PULLUP = 1'b0;
    defparam DATA15_pad.NEG_TRIGGER = 1'b0;
    defparam DATA15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA8_pad (.PACKAGE_PIN(DATA8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA8_c_8));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA8_pad.PIN_TYPE = 6'b011001;
    defparam DATA8_pad.PULLUP = 1'b0;
    defparam DATA8_pad.NEG_TRIGGER = 1'b0;
    defparam DATA8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA14_pad (.PACKAGE_PIN(DATA14), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA14_c_14));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA14_pad.PIN_TYPE = 6'b011001;
    defparam DATA14_pad.PULLUP = 1'b0;
    defparam DATA14_pad.NEG_TRIGGER = 1'b0;
    defparam DATA14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA13_pad (.PACKAGE_PIN(DATA13), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA13_c_13));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA13_pad.PIN_TYPE = 6'b011001;
    defparam DATA13_pad.PULLUP = 1'b0;
    defparam DATA13_pad.NEG_TRIGGER = 1'b0;
    defparam DATA13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA12_pad (.PACKAGE_PIN(DATA12), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA12_c_12));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA12_pad.PIN_TYPE = 6'b011001;
    defparam DATA12_pad.PULLUP = 1'b0;
    defparam DATA12_pad.NEG_TRIGGER = 1'b0;
    defparam DATA12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA11_pad (.PACKAGE_PIN(DATA11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA11_c_11));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA11_pad.PIN_TYPE = 6'b011001;
    defparam DATA11_pad.PULLUP = 1'b0;
    defparam DATA11_pad.NEG_TRIGGER = 1'b0;
    defparam DATA11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA9_pad (.PACKAGE_PIN(DATA9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA9_c_9));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA9_pad.PIN_TYPE = 6'b011001;
    defparam DATA9_pad.PULLUP = 1'b0;
    defparam DATA9_pad.NEG_TRIGGER = 1'b0;
    defparam DATA9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA10_pad (.PACKAGE_PIN(DATA10), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA10_c_10));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA10_pad.PIN_TYPE = 6'b011001;
    defparam DATA10_pad.PULLUP = 1'b0;
    defparam DATA10_pad.NEG_TRIGGER = 1'b0;
    defparam DATA10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_OE_pad (.PACKAGE_PIN(FT_OE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_OE_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_OE_pad.PIN_TYPE = 6'b011001;
    defparam FT_OE_pad.PULLUP = 1'b0;
    defparam FT_OE_pad.NEG_TRIGGER = 1'b0;
    defparam FT_OE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_RD_pad (.PACKAGE_PIN(FT_RD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_RD_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_RD_pad.PIN_TYPE = 6'b011001;
    defparam FT_RD_pad.PULLUP = 1'b0;
    defparam FT_RD_pad.NEG_TRIGGER = 1'b0;
    defparam FT_RD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_WR_pad (.PACKAGE_PIN(FT_WR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_WR_pad.PIN_TYPE = 6'b011001;
    defparam FT_WR_pad.PULLUP = 1'b0;
    defparam FT_WR_pad.NEG_TRIGGER = 1'b0;
    defparam FT_WR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_SIWU_pad (.PACKAGE_PIN(FT_SIWU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_SIWU_pad.PIN_TYPE = 6'b011001;
    defparam FT_SIWU_pad.PULLUP = 1'b0;
    defparam FT_SIWU_pad.NEG_TRIGGER = 1'b0;
    defparam FT_SIWU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_0_pad (.PACKAGE_PIN(DEBUG_0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_0_c_24));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_0_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_0_pad.PULLUP = 1'b0;
    defparam DEBUG_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_1_pad (.PACKAGE_PIN(DEBUG_1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_1_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_1_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_1_pad.PULLUP = 1'b0;
    defparam DEBUG_1_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_2_pad (.PACKAGE_PIN(DEBUG_2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_2_c_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_2_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_2_pad.PULLUP = 1'b0;
    defparam DEBUG_2_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_3_pad (.PACKAGE_PIN(DEBUG_3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(\MISC.empty_flag_r )) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_3_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_3_pad.PULLUP = 1'b0;
    defparam DEBUG_3_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_5_pad (.PACKAGE_PIN(DEBUG_5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_5_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_5_pad.PULLUP = 1'b0;
    defparam DEBUG_5_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_6_pad (.PACKAGE_PIN(DEBUG_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_6_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_6_pad.PULLUP = 1'b0;
    defparam DEBUG_6_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_8_pad (.PACKAGE_PIN(DEBUG_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_8_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_8_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_8_pad.PULLUP = 1'b0;
    defparam DEBUG_8_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_9_pad (.PACKAGE_PIN(DEBUG_9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_9_c_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_9_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_9_pad.PULLUP = 1'b0;
    defparam DEBUG_9_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CLK_pad (.PACKAGE_PIN(ICE_CLK), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CLK_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CLK_pad.PULLUP = 1'b0;
    defparam ICE_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CDONE_pad (.PACKAGE_PIN(ICE_CDONE), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CDONE_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CDONE_pad.PULLUP = 1'b0;
    defparam ICE_CDONE_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CDONE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CREST_pad (.PACKAGE_PIN(ICE_CREST), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CREST_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CREST_pad.PULLUP = 1'b0;
    defparam ICE_CREST_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CREST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_SYSCLK_pad (.PACKAGE_PIN(ICE_SYSCLK), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ICE_SYSCLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_SYSCLK_pad.PIN_TYPE = 6'b000001;
    defparam ICE_SYSCLK_pad.PULLUP = 1'b0;
    defparam ICE_SYSCLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_SYSCLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_2_c_pad (.PACKAGE_PIN(UART_RX), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(DEBUG_2_c_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_2_c_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_2_c_pad.PULLUP = 1'b0;
    defparam DEBUG_2_c_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_2_c_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SOUT_pad (.PACKAGE_PIN(SOUT), .OUTPUT_ENABLE(VCC_net), .D_IN_0(SOUT_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SOUT_pad.PIN_TYPE = 6'b000001;
    defparam SOUT_pad.PULLUP = 1'b0;
    defparam SOUT_pad.NEG_TRIGGER = 1'b0;
    defparam SOUT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_9_c_pad (.PACKAGE_PIN(FR_RXF), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(DEBUG_9_c_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_9_c_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_9_c_pad.PULLUP = 1'b0;
    defparam DEBUG_9_c_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_9_c_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D31_pad (.PACKAGE_PIN(FIFO_D31), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D31_c_0));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D31_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D31_pad.PULLUP = 1'b0;
    defparam FIFO_D31_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D31_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D30_pad (.PACKAGE_PIN(FIFO_D30), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D30_c_1));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D30_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D30_pad.PULLUP = 1'b0;
    defparam FIFO_D30_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D30_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D29_pad (.PACKAGE_PIN(FIFO_D29), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D29_c_2));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D29_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D29_pad.PULLUP = 1'b0;
    defparam FIFO_D29_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D29_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D28_pad (.PACKAGE_PIN(FIFO_D28), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D28_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D28_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D28_pad.PULLUP = 1'b0;
    defparam FIFO_D28_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D28_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D27_pad (.PACKAGE_PIN(FIFO_D27), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D27_c_4));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D27_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D27_pad.PULLUP = 1'b0;
    defparam FIFO_D27_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D27_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO FIFO_CLK_pad (.PACKAGE_PIN(FIFO_CLK), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(FIFO_CLK_c));   // src/top.v(84[12:20])
    defparam FIFO_CLK_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_CLK_pad.PULLUP = 1'b0;
    defparam FIFO_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D26_pad (.PACKAGE_PIN(FIFO_D26), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D26_c_5));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D26_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D26_pad.PULLUP = 1'b0;
    defparam FIFO_D26_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D26_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D25_pad (.PACKAGE_PIN(FIFO_D25), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D25_c_6));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D25_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D25_pad.PULLUP = 1'b0;
    defparam FIFO_D25_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D25_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D24_pad (.PACKAGE_PIN(FIFO_D24), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D24_c_7));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D24_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D24_pad.PULLUP = 1'b0;
    defparam FIFO_D24_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D23_pad (.PACKAGE_PIN(FIFO_D23), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D23_c_8));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D23_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D23_pad.PULLUP = 1'b0;
    defparam FIFO_D23_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D22_pad (.PACKAGE_PIN(FIFO_D22), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D22_c_9));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D22_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D22_pad.PULLUP = 1'b0;
    defparam FIFO_D22_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D21_pad (.PACKAGE_PIN(FIFO_D21), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D21_c_10));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D21_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D21_pad.PULLUP = 1'b0;
    defparam FIFO_D21_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D20_pad (.PACKAGE_PIN(FIFO_D20), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D20_c_11));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D20_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D20_pad.PULLUP = 1'b0;
    defparam FIFO_D20_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D19_pad (.PACKAGE_PIN(FIFO_D19), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D19_c_12));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D19_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D19_pad.PULLUP = 1'b0;
    defparam FIFO_D19_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D18_pad (.PACKAGE_PIN(FIFO_D18), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D18_c_13));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D18_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D18_pad.PULLUP = 1'b0;
    defparam FIFO_D18_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D17_pad (.PACKAGE_PIN(FIFO_D17), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D17_c_14));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D17_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D17_pad.PULLUP = 1'b0;
    defparam FIFO_D17_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D17_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D16_pad (.PACKAGE_PIN(FIFO_D16), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D16_c_15));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D16_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D16_pad.PULLUP = 1'b0;
    defparam FIFO_D16_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D16_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D15_pad (.PACKAGE_PIN(FIFO_D15), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D15_c_16));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D15_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D15_pad.PULLUP = 1'b0;
    defparam FIFO_D15_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D14_pad (.PACKAGE_PIN(FIFO_D14), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D14_c_17));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D14_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D14_pad.PULLUP = 1'b0;
    defparam FIFO_D14_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D13_pad (.PACKAGE_PIN(FIFO_D13), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D13_c_18));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D13_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D13_pad.PULLUP = 1'b0;
    defparam FIFO_D13_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D12_pad (.PACKAGE_PIN(FIFO_D12), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D12_c_19));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D12_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D12_pad.PULLUP = 1'b0;
    defparam FIFO_D12_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D11_pad (.PACKAGE_PIN(FIFO_D11), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D11_c_20));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D11_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D11_pad.PULLUP = 1'b0;
    defparam FIFO_D11_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D10_pad (.PACKAGE_PIN(FIFO_D10), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D10_c_21));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D10_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D10_pad.PULLUP = 1'b0;
    defparam FIFO_D10_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D9_pad (.PACKAGE_PIN(FIFO_D9), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D9_c_22));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D9_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D9_pad.PULLUP = 1'b0;
    defparam FIFO_D9_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D8_pad (.PACKAGE_PIN(FIFO_D8), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D8_c_23));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D8_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D8_pad.PULLUP = 1'b0;
    defparam FIFO_D8_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D7_pad (.PACKAGE_PIN(FIFO_D7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D7_c_24));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D7_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D7_pad.PULLUP = 1'b0;
    defparam FIFO_D7_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D6_pad (.PACKAGE_PIN(FIFO_D6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D6_c_25));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D6_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D6_pad.PULLUP = 1'b0;
    defparam FIFO_D6_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D5_pad (.PACKAGE_PIN(FIFO_D5), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D5_c_26));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D5_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D5_pad.PULLUP = 1'b0;
    defparam FIFO_D5_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D4_pad (.PACKAGE_PIN(FIFO_D4), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D4_c_27));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D4_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D4_pad.PULLUP = 1'b0;
    defparam FIFO_D4_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D3_pad (.PACKAGE_PIN(FIFO_D3), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D3_c_28));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D3_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D3_pad.PULLUP = 1'b0;
    defparam FIFO_D3_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D2_pad (.PACKAGE_PIN(FIFO_D2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D2_c_29));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D2_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D2_pad.PULLUP = 1'b0;
    defparam FIFO_D2_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D1_pad (.PACKAGE_PIN(FIFO_D1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D1_c_30));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D1_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D1_pad.PULLUP = 1'b0;
    defparam FIFO_D1_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D0_pad (.PACKAGE_PIN(FIFO_D0), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D0_c_31));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D0_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D0_pad.PULLUP = 1'b0;
    defparam FIFO_D0_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i5559_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[4]), .I2(\mem_LUT.data_raw_r [4]), 
            .I3(n5207), .O(n7058));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i5559_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i5562_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[3]), .I2(\mem_LUT.data_raw_r [3]), 
            .I3(n5207), .O(n7061));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i5562_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i5565_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[2]), .I2(\mem_LUT.data_raw_r [2]), 
            .I3(n5207), .O(n7064));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i5565_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i5568_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[1]), .I2(\mem_LUT.data_raw_r [1]), 
            .I3(n5207), .O(n7067));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i5568_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4318_3_lut (.I0(\REG.mem_5_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n28), .I3(GND_net), .O(n5817));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4319_3_lut (.I0(\REG.mem_5_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n28), .I3(GND_net), .O(n5818));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4320_3_lut (.I0(\REG.mem_5_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n28), .I3(GND_net), .O(n5819));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4321_3_lut (.I0(\REG.mem_5_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n28), .I3(GND_net), .O(n5820));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4322_3_lut (.I0(\REG.mem_5_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n28), .I3(GND_net), .O(n5821));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4323_3_lut (.I0(\REG.mem_5_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n28), .I3(GND_net), .O(n5822));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4324_3_lut (.I0(\REG.mem_5_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n28), .I3(GND_net), .O(n5823));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4325_3_lut (.I0(\REG.mem_5_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n28), .I3(GND_net), .O(n5824));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4326_3_lut (.I0(\REG.mem_5_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n28), .I3(GND_net), .O(n5825));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3794_4_lut (.I0(n63), .I1(n4843), .I2(n10059), .I3(state[3]), 
            .O(n2178));   // src/timing_controller.v(78[11:16])
    defparam i3794_4_lut.LUT_INIT = 16'h0a88;
    SB_LUT4 led_counter_1466_1542_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(DEBUG_0_c_24), .I3(n13776), .O(n106)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1956_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n3414));   // src/top.v(1198[8] 1265[4])
    defparam i1956_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 led_counter_1466_1542_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n2), .I3(n13775), .O(n107)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5002_3_lut (.I0(\REG.mem_27_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n6), .I3(GND_net), .O(n6501));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5003_3_lut (.I0(\REG.mem_27_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n6), .I3(GND_net), .O(n6502));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5004_3_lut (.I0(\REG.mem_27_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n6), .I3(GND_net), .O(n6503));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5005_3_lut (.I0(\REG.mem_27_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n6), .I3(GND_net), .O(n6504));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4327_3_lut (.I0(\REG.mem_5_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n28), .I3(GND_net), .O(n5826));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5006_3_lut (.I0(\REG.mem_27_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n6), .I3(GND_net), .O(n6505));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5007_3_lut (.I0(\REG.mem_27_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n6), .I3(GND_net), .O(n6506));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4328_3_lut (.I0(\REG.mem_5_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n28), .I3(GND_net), .O(n5827));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5008_3_lut (.I0(\REG.mem_27_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n6), .I3(GND_net), .O(n6507));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5009_3_lut (.I0(\REG.mem_27_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n6), .I3(GND_net), .O(n6508));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5010_3_lut (.I0(\REG.mem_27_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n6), .I3(GND_net), .O(n6509));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5011_3_lut (.I0(\REG.mem_27_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n6), .I3(GND_net), .O(n6510));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5012_3_lut (.I0(\REG.mem_27_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n6), .I3(GND_net), .O(n6511));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5012_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1466_1542_add_4_25 (.CI(n13775), .I0(GND_net), 
            .I1(n2), .CO(n13776));
    SB_LUT4 i5013_3_lut (.I0(\REG.mem_27_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n6), .I3(GND_net), .O(n6512));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5014_3_lut (.I0(\REG.mem_27_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n6), .I3(GND_net), .O(n6513));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4329_3_lut (.I0(\REG.mem_5_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n28), .I3(GND_net), .O(n5828));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4330_3_lut (.I0(\REG.mem_6_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n27), .I3(GND_net), .O(n5829));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1466_1542_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3), .I3(n13774), .O(n108)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5015_3_lut (.I0(\REG.mem_27_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n6), .I3(GND_net), .O(n6514));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4331_3_lut (.I0(\REG.mem_6_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n27), .I3(GND_net), .O(n5830));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4332_3_lut (.I0(\REG.mem_6_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n27), .I3(GND_net), .O(n5831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4333_3_lut (.I0(\REG.mem_6_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n27), .I3(GND_net), .O(n5832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5016_3_lut (.I0(\REG.mem_27_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n6), .I3(GND_net), .O(n6515));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5017_3_lut (.I0(\REG.mem_27_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n6), .I3(GND_net), .O(n6516));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5017_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_LUT4 i5018_3_lut (.I0(\REG.mem_27_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n6), .I3(GND_net), .O(n6517));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5019_3_lut (.I0(\REG.mem_27_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n6), .I3(GND_net), .O(n6518));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5020_3_lut (.I0(\REG.mem_27_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n6), .I3(GND_net), .O(n6519));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5021_3_lut (.I0(\REG.mem_27_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n6), .I3(GND_net), .O(n6520));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5022_3_lut (.I0(\REG.mem_27_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n6), .I3(GND_net), .O(n6521));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5023_3_lut (.I0(\REG.mem_27_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n6), .I3(GND_net), .O(n6522));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5024_3_lut (.I0(\REG.mem_27_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n6), .I3(GND_net), .O(n6523));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5025_3_lut (.I0(\REG.mem_27_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n6), .I3(GND_net), .O(n6524));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5026_3_lut (.I0(\REG.mem_27_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n6), .I3(GND_net), .O(n6525));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5027_3_lut (.I0(\REG.mem_27_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n6), .I3(GND_net), .O(n6526));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5028_3_lut (.I0(\REG.mem_27_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n6), .I3(GND_net), .O(n6527));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5029_3_lut (.I0(\REG.mem_27_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n6), .I3(GND_net), .O(n6528));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5030_3_lut (.I0(\REG.mem_27_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n6), .I3(GND_net), .O(n6529));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5030_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1466_1542_add_4_24 (.CI(n13774), .I0(GND_net), 
            .I1(n3), .CO(n13775));
    SB_LUT4 i5031_3_lut (.I0(\REG.mem_27_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n6), .I3(GND_net), .O(n6530));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5032_3_lut (.I0(\REG.mem_27_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n6), .I3(GND_net), .O(n6531));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5033_3_lut (.I0(\REG.mem_27_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n6), .I3(GND_net), .O(n6532));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i5033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4334_3_lut (.I0(\REG.mem_6_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n27), .I3(GND_net), .O(n5833));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11646_2_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_1428));   // src/top.v(259[27:51])
    defparam i11646_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 led_counter_1466_1542_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_1418), .I3(n13773), .O(n109)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_23 (.CI(n13773), .I0(GND_net), 
            .I1(n4_adj_1418), .CO(n13774));
    SB_LUT4 i4335_3_lut (.I0(\REG.mem_6_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n27), .I3(GND_net), .O(n5834));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4336_3_lut (.I0(\REG.mem_6_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n27), .I3(GND_net), .O(n5835));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1466_1542_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5), .I3(n13772), .O(n110)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_22 (.CI(n13772), .I0(GND_net), 
            .I1(n5), .CO(n13773));
    SB_LUT4 led_counter_1466_1542_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_1419), .I3(n13771), .O(n111)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_21 (.CI(n13771), .I0(GND_net), 
            .I1(n6_adj_1419), .CO(n13772));
    SB_LUT4 led_counter_1466_1542_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7), .I3(n13770), .O(n112)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_20 (.CI(n13770), .I0(GND_net), 
            .I1(n7), .CO(n13771));
    SB_LUT4 led_counter_1466_1542_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_1420), .I3(n13769), .O(n113)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_19 (.CI(n13769), .I0(GND_net), 
            .I1(n8_adj_1420), .CO(n13770));
    SB_LUT4 led_counter_1466_1542_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9), .I3(n13768), .O(n114)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_18 (.CI(n13768), .I0(GND_net), 
            .I1(n9), .CO(n13769));
    SB_LUT4 led_counter_1466_1542_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_1421), .I3(n13767), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_17 (.CI(n13767), .I0(GND_net), 
            .I1(n10_adj_1421), .CO(n13768));
    SB_LUT4 led_counter_1466_1542_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_1422), .I3(n13766), .O(n116)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_16 (.CI(n13766), .I0(GND_net), 
            .I1(n11_adj_1422), .CO(n13767));
    SB_LUT4 led_counter_1466_1542_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_1423), .I3(n13765), .O(n117)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_153 (.I0(reset_clk_counter[0]), .I1(reset_clk_counter[2]), 
            .I2(reset_clk_counter[3]), .I3(reset_clk_counter[1]), .O(reset_all_w_N_61));
    defparam i3_4_lut_adj_153.LUT_INIT = 16'hfffe;
    SB_DFF fifo_write_cmd_79 (.Q(fifo_write_cmd), .C(SLM_CLK_c), .D(n5703));   // src/top.v(1013[8] 1022[4])
    SB_LUT4 i4337_3_lut (.I0(\REG.mem_6_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n27), .I3(GND_net), .O(n5836));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4338_3_lut (.I0(\REG.mem_6_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n27), .I3(GND_net), .O(n5837));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4339_3_lut (.I0(\REG.mem_6_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n27), .I3(GND_net), .O(n5838));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4340_3_lut (.I0(\REG.mem_6_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n27), .I3(GND_net), .O(n5839));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4341_3_lut (.I0(\REG.mem_6_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n27), .I3(GND_net), .O(n5840));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4342_3_lut (.I0(\REG.mem_6_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n27), .I3(GND_net), .O(n5841));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4343_3_lut (.I0(\REG.mem_6_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n27), .I3(GND_net), .O(n5842));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4344_3_lut (.I0(\REG.mem_6_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n27), .I3(GND_net), .O(n5843));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4345_3_lut (.I0(\REG.mem_6_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n27), .I3(GND_net), .O(n5844));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4346_3_lut (.I0(\REG.mem_6_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n27), .I3(GND_net), .O(n5845));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4347_3_lut (.I0(\REG.mem_6_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n27), .I3(GND_net), .O(n5846));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4347_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1466_1542_add_4_15 (.CI(n13765), .I0(GND_net), 
            .I1(n12_adj_1423), .CO(n13766));
    SB_LUT4 led_counter_1466_1542_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13), .I3(n13764), .O(n118)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4348_3_lut (.I0(\REG.mem_6_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n27), .I3(GND_net), .O(n5847));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4349_3_lut (.I0(\REG.mem_6_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n27), .I3(GND_net), .O(n5848));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4350_3_lut (.I0(\REG.mem_6_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n27), .I3(GND_net), .O(n5849));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4350_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1466_1542_add_4_14 (.CI(n13764), .I0(GND_net), 
            .I1(n13), .CO(n13765));
    SB_LUT4 led_counter_1466_1542_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14), .I3(n13763), .O(n119)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_13 (.CI(n13763), .I0(GND_net), 
            .I1(n14), .CO(n13764));
    SB_LUT4 i4351_3_lut (.I0(\REG.mem_6_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n27), .I3(GND_net), .O(n5850));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1466_1542_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15), .I3(n13762), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_12 (.CI(n13762), .I0(GND_net), 
            .I1(n15), .CO(n13763));
    SB_LUT4 led_counter_1466_1542_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16), .I3(n13761), .O(n121)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_11 (.CI(n13761), .I0(GND_net), 
            .I1(n16), .CO(n13762));
    SB_LUT4 led_counter_1466_1542_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17), .I3(n13760), .O(n122)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4148_4_lut_4_lut (.I0(wr_fifo_en_w_adj_1412), .I1(reset_all_w), 
            .I2(wr_addr_p1_w_adj_1504[2]), .I3(wr_addr_r_adj_1502[2]), .O(n5647));
    defparam i4148_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4159_4_lut_4_lut_4_lut (.I0(wr_fifo_en_w_adj_1412), .I1(reset_all_w), 
            .I2(wr_addr_r_adj_1502[0]), .I3(wr_addr_r_adj_1502[1]), .O(n5658));
    defparam i4159_4_lut_4_lut_4_lut.LUT_INIT = 16'h1320;
    SB_LUT4 i4352_3_lut (.I0(\REG.mem_6_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n27), .I3(GND_net), .O(n5851));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4353_3_lut (.I0(\REG.mem_6_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n27), .I3(GND_net), .O(n5852));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4353_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1466_1542__i1 (.Q(n24), .C(SLM_CLK_c), .D(n129));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i2 (.Q(n23), .C(SLM_CLK_c), .D(n128));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i3 (.Q(n22_adj_1424), .C(SLM_CLK_c), .D(n127));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i4 (.Q(n21), .C(SLM_CLK_c), .D(n126));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i5 (.Q(n20), .C(SLM_CLK_c), .D(n125));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i6 (.Q(n19), .C(SLM_CLK_c), .D(n124));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i7 (.Q(n18), .C(SLM_CLK_c), .D(n123));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i8 (.Q(n17), .C(SLM_CLK_c), .D(n122));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i9 (.Q(n16), .C(SLM_CLK_c), .D(n121));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i10 (.Q(n15), .C(SLM_CLK_c), .D(n120));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i11 (.Q(n14), .C(SLM_CLK_c), .D(n119));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i12 (.Q(n13), .C(SLM_CLK_c), .D(n118));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i13 (.Q(n12_adj_1423), .C(SLM_CLK_c), 
           .D(n117));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i14 (.Q(n11_adj_1422), .C(SLM_CLK_c), 
           .D(n116));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i15 (.Q(n10_adj_1421), .C(SLM_CLK_c), 
           .D(n115));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i16 (.Q(n9), .C(SLM_CLK_c), .D(n114));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i17 (.Q(n8_adj_1420), .C(SLM_CLK_c), .D(n113));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i18 (.Q(n7), .C(SLM_CLK_c), .D(n112));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i19 (.Q(n6_adj_1419), .C(SLM_CLK_c), .D(n111));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i20 (.Q(n5), .C(SLM_CLK_c), .D(n110));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i21 (.Q(n4_adj_1418), .C(SLM_CLK_c), .D(n109));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i22 (.Q(n3), .C(SLM_CLK_c), .D(n108));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i23 (.Q(n2), .C(SLM_CLK_c), .D(n107));   // src/top.v(203[20:35])
    SB_DFF led_counter_1466_1542__i24 (.Q(DEBUG_0_c_24), .C(SLM_CLK_c), 
           .D(n106));   // src/top.v(203[20:35])
    SB_DFF reset_clk_counter_i3_1467__i1 (.Q(reset_clk_counter[1]), .C(SLM_CLK_c), 
           .D(n13898));   // src/top.v(259[27:51])
    SB_LUT4 i4354_3_lut (.I0(\REG.mem_6_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n27), .I3(GND_net), .O(n5853));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4355_3_lut (.I0(\REG.mem_6_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n27), .I3(GND_net), .O(n5854));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4356_3_lut (.I0(\REG.mem_6_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n27), .I3(GND_net), .O(n5855));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4357_3_lut (.I0(\REG.mem_6_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n27), .I3(GND_net), .O(n5856));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4358_3_lut (.I0(\REG.mem_6_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n27), .I3(GND_net), .O(n5857));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4359_3_lut (.I0(\REG.mem_6_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n27), .I3(GND_net), .O(n5858));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4360_3_lut (.I0(\REG.mem_6_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n27), .I3(GND_net), .O(n5859));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4361_3_lut (.I0(\REG.mem_6_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n27), .I3(GND_net), .O(n5860));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4362_3_lut (.I0(\REG.mem_7_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n26), .I3(GND_net), .O(n5861));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4363_3_lut (.I0(\REG.mem_7_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n26), .I3(GND_net), .O(n5862));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4364_3_lut (.I0(\REG.mem_7_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n26), .I3(GND_net), .O(n5863));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4364_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1466_1542_add_4_10 (.CI(n13760), .I0(GND_net), 
            .I1(n17), .CO(n13761));
    SB_LUT4 i4365_3_lut (.I0(\REG.mem_7_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n26), .I3(GND_net), .O(n5864));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4366_3_lut (.I0(\REG.mem_7_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n26), .I3(GND_net), .O(n5865));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4367_3_lut (.I0(\REG.mem_7_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n26), .I3(GND_net), .O(n5866));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4368_3_lut (.I0(\REG.mem_7_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n26), .I3(GND_net), .O(n5867));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4369_3_lut (.I0(\REG.mem_7_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n26), .I3(GND_net), .O(n5868));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4370_3_lut (.I0(\REG.mem_7_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n26), .I3(GND_net), .O(n5869));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4371_3_lut (.I0(\REG.mem_7_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n26), .I3(GND_net), .O(n5870));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4372_3_lut (.I0(\REG.mem_7_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n26), .I3(GND_net), .O(n5871));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4373_3_lut (.I0(\REG.mem_7_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n26), .I3(GND_net), .O(n5872));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4374_3_lut (.I0(\REG.mem_7_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n26), .I3(GND_net), .O(n5873));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4375_3_lut (.I0(\REG.mem_7_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n26), .I3(GND_net), .O(n5874));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4376_3_lut (.I0(\REG.mem_7_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n26), .I3(GND_net), .O(n5875));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4377_3_lut (.I0(\REG.mem_7_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n26), .I3(GND_net), .O(n5876));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4378_3_lut (.I0(\REG.mem_7_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n26), .I3(GND_net), .O(n5877));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4379_3_lut (.I0(\REG.mem_7_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n26), .I3(GND_net), .O(n5878));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4380_3_lut (.I0(\REG.mem_7_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n26), .I3(GND_net), .O(n5879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4381_3_lut (.I0(\REG.mem_7_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n26), .I3(GND_net), .O(n5880));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4382_3_lut (.I0(\REG.mem_7_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n26), .I3(GND_net), .O(n5881));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4383_3_lut (.I0(\REG.mem_7_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n26), .I3(GND_net), .O(n5882));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4384_3_lut (.I0(\REG.mem_7_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n26), .I3(GND_net), .O(n5883));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut (.I0(reset_clk_counter[1]), .I1(n2_adj_1428), 
            .I2(reset_clk_counter[2]), .I3(reset_clk_counter[3]), .O(n13902));   // src/top.v(259[27:51])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfe01;
    SB_LUT4 i4385_3_lut (.I0(\REG.mem_7_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n26), .I3(GND_net), .O(n5884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4386_3_lut (.I0(\REG.mem_7_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n26), .I3(GND_net), .O(n5885));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4387_3_lut (.I0(\REG.mem_7_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n26), .I3(GND_net), .O(n5886));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4388_3_lut (.I0(\REG.mem_7_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n26), .I3(GND_net), .O(n5887));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4389_3_lut (.I0(\REG.mem_7_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n26), .I3(GND_net), .O(n5888));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4390_3_lut (.I0(\REG.mem_7_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n26), .I3(GND_net), .O(n5889));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4391_3_lut (.I0(\REG.mem_7_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n26), .I3(GND_net), .O(n5890));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4392_3_lut (.I0(\REG.mem_7_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n26), .I3(GND_net), .O(n5891));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4393_3_lut (.I0(\REG.mem_7_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n26), .I3(GND_net), .O(n5892));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1466_1542_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18), .I3(n13759), .O(n123)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_9 (.CI(n13759), .I0(GND_net), .I1(n18), 
            .CO(n13760));
    SB_LUT4 led_counter_1466_1542_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19), .I3(n13758), .O(n124)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_8 (.CI(n13758), .I0(GND_net), .I1(n19), 
            .CO(n13759));
    SB_LUT4 led_counter_1466_1542_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20), .I3(n13757), .O(n125)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF uart_rx_complete_rising_edge_82 (.Q(uart_rx_complete_rising_edge), 
           .C(SLM_CLK_c), .D(n5618));   // src/top.v(1189[8] 1195[4])
    SB_CARRY led_counter_1466_1542_add_4_7 (.CI(n13757), .I0(GND_net), .I1(n20), 
            .CO(n13758));
    SB_LUT4 led_counter_1466_1542_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21), .I3(n13756), .O(n126)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF tx_addr_byte_r_i0_i0 (.Q(tx_addr_byte[0]), .C(SLM_CLK_c), .D(n5614));   // src/top.v(1198[8] 1265[4])
    SB_DFF reset_clk_counter_i3_1467__i2 (.Q(reset_clk_counter[2]), .C(SLM_CLK_c), 
           .D(n13900));   // src/top.v(259[27:51])
    SB_DFF fifo_read_cmd_80 (.Q(fifo_read_cmd), .C(SLM_CLK_c), .D(start_tx_N_64));   // src/top.v(1034[8] 1052[4])
    SB_DFF reset_clk_counter_i3_1467__i3 (.Q(reset_clk_counter[3]), .C(SLM_CLK_c), 
           .D(n13902));   // src/top.v(259[27:51])
    SB_DFF tx_data_byte_r_i0_i0 (.Q(tx_data_byte[0]), .C(SLM_CLK_c), .D(n5597));   // src/top.v(1198[8] 1265[4])
    SB_CARRY led_counter_1466_1542_add_4_6 (.CI(n13756), .I0(GND_net), .I1(n21), 
            .CO(n13757));
    SB_LUT4 i4810_3_lut (.I0(\REG.mem_21_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6309));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4811_3_lut (.I0(\REG.mem_21_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6310));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4812_3_lut (.I0(\REG.mem_21_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6311));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4813_3_lut (.I0(\REG.mem_21_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6312));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4490_3_lut (.I0(\REG.mem_11_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n22), .I3(GND_net), .O(n5989));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1466_1542_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_1424), .I3(n13755), .O(n127)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4491_3_lut (.I0(\REG.mem_11_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n22), .I3(GND_net), .O(n5990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4492_3_lut (.I0(\REG.mem_11_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n22), .I3(GND_net), .O(n5991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4493_3_lut (.I0(\REG.mem_11_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n22), .I3(GND_net), .O(n5992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8388_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n9873));
    defparam i8388_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4494_3_lut (.I0(\REG.mem_11_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n22), .I3(GND_net), .O(n5993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4204_2_lut (.I0(is_tx_fifo_full_flag), .I1(spi_rx_byte_ready), 
            .I2(GND_net), .I3(GND_net), .O(n5703));   // src/top.v(1013[8] 1022[4])
    defparam i4204_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY led_counter_1466_1542_add_4_5 (.CI(n13755), .I0(GND_net), .I1(n22_adj_1424), 
            .CO(n13756));
    SB_LUT4 led_counter_1466_1542_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23), .I3(n13754), .O(n128)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_4 (.CI(n13754), .I0(GND_net), .I1(n23), 
            .CO(n13755));
    SB_LUT4 led_counter_1466_1542_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24), .I3(n13753), .O(n129)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1466_1542_add_4_3 (.CI(n13753), .I0(GND_net), .I1(n24), 
            .CO(n13754));
    SB_LUT4 led_counter_1466_1542_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_1425), .I3(VCC_net), .O(n130)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1466_1542_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4495_3_lut (.I0(\REG.mem_11_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n22), .I3(GND_net), .O(n5994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4496_3_lut (.I0(\REG.mem_11_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n22), .I3(GND_net), .O(n5995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4497_3_lut (.I0(\REG.mem_11_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n22), .I3(GND_net), .O(n5996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4498_3_lut (.I0(\REG.mem_11_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n22), .I3(GND_net), .O(n5997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1214_4_lut (.I0(n2438), .I1(n10059), .I2(state[3]), .I3(n63), 
            .O(n2283));   // src/timing_controller.v(78[11:16])
    defparam i1214_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i4499_3_lut (.I0(\REG.mem_11_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n22), .I3(GND_net), .O(n5998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4500_3_lut (.I0(\REG.mem_11_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n22), .I3(GND_net), .O(n5999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4501_3_lut (.I0(\REG.mem_11_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n22), .I3(GND_net), .O(n6000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4502_3_lut (.I0(\REG.mem_11_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n22), .I3(GND_net), .O(n6001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4503_3_lut (.I0(\REG.mem_11_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n22), .I3(GND_net), .O(n6002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4504_3_lut (.I0(\REG.mem_11_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n22), .I3(GND_net), .O(n6003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4505_3_lut (.I0(\REG.mem_11_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n22), .I3(GND_net), .O(n6004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4506_3_lut (.I0(\REG.mem_11_16 ), .I1(dc32_fifo_data_in[16]), 
            .I2(n22), .I3(GND_net), .O(n6005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4507_3_lut (.I0(\REG.mem_11_17 ), .I1(dc32_fifo_data_in[17]), 
            .I2(n22), .I3(GND_net), .O(n6006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4507_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1466_1542_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(n25_adj_1425), .CO(n13753));
    SB_LUT4 i1_3_lut (.I0(buffer_switch_done_latched), .I1(n989), .I2(n910), 
            .I3(GND_net), .O(n14298));
    defparam i1_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i4508_3_lut (.I0(\REG.mem_11_18 ), .I1(dc32_fifo_data_in[18]), 
            .I2(n22), .I3(GND_net), .O(n6007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4509_3_lut (.I0(\REG.mem_11_19 ), .I1(dc32_fifo_data_in[19]), 
            .I2(n22), .I3(GND_net), .O(n6008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4510_3_lut (.I0(\REG.mem_11_20 ), .I1(dc32_fifo_data_in[20]), 
            .I2(n22), .I3(GND_net), .O(n6009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4511_3_lut (.I0(\REG.mem_11_21 ), .I1(dc32_fifo_data_in[21]), 
            .I2(n22), .I3(GND_net), .O(n6010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4512_3_lut (.I0(\REG.mem_11_22 ), .I1(dc32_fifo_data_in[22]), 
            .I2(n22), .I3(GND_net), .O(n6011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4513_3_lut (.I0(\REG.mem_11_23 ), .I1(dc32_fifo_data_in[23]), 
            .I2(n22), .I3(GND_net), .O(n6012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4514_3_lut (.I0(\REG.mem_11_24 ), .I1(dc32_fifo_data_in[24]), 
            .I2(n22), .I3(GND_net), .O(n6013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4515_3_lut (.I0(\REG.mem_11_25 ), .I1(dc32_fifo_data_in[25]), 
            .I2(n22), .I3(GND_net), .O(n6014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4516_3_lut (.I0(\REG.mem_11_26 ), .I1(dc32_fifo_data_in[26]), 
            .I2(n22), .I3(GND_net), .O(n6015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4517_3_lut (.I0(\REG.mem_11_27 ), .I1(dc32_fifo_data_in[27]), 
            .I2(n22), .I3(GND_net), .O(n6016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4518_3_lut (.I0(\REG.mem_11_28 ), .I1(dc32_fifo_data_in[28]), 
            .I2(n22), .I3(GND_net), .O(n6017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4519_3_lut (.I0(\REG.mem_11_29 ), .I1(dc32_fifo_data_in[29]), 
            .I2(n22), .I3(GND_net), .O(n6018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4520_3_lut (.I0(\REG.mem_11_30 ), .I1(dc32_fifo_data_in[30]), 
            .I2(n22), .I3(GND_net), .O(n6019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4521_3_lut (.I0(\REG.mem_11_31 ), .I1(dc32_fifo_data_in[31]), 
            .I2(n22), .I3(GND_net), .O(n6020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 reset_all_w_I_0_1_lut (.I0(reset_all_w), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(RESET_c));   // src/top.v(295[16:28])
    defparam reset_all_w_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1209_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(n63), 
            .I3(state[2]), .O(n2438));   // src/timing_controller.v(78[11:16])
    defparam i1209_4_lut_4_lut.LUT_INIT = 16'h0806;
    SB_LUT4 i8566_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(n63), 
            .I3(GND_net), .O(n10051));
    defparam i8566_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(reset_clk_counter[1]), .I1(reset_all_w_N_61), 
            .I2(reset_clk_counter[0]), .I3(reset_clk_counter[2]), .O(n13900));   // src/top.v(259[27:51])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfb04;
    SB_LUT4 i1973_2_lut_3_lut_4_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(reset_all_w), .I3(wr_addr_r_adj_1502[0]), .O(n8));
    defparam i1973_2_lut_3_lut_4_lut.LUT_INIT = 16'h0df2;
    fifo_sc_32_lut_gen fifo_sc_32_lut_gen_inst (.n5412(n5412), .GND_net(GND_net), 
            .\sc32_fifo_data_out[0] (sc32_fifo_data_out[0]), .SLM_CLK_c(SLM_CLK_c), 
            .dc32_fifo_data_out({dc32_fifo_data_out}), .\MISC.empty_flag_r (\MISC.empty_flag_r ), 
            .sc32_fifo_almost_empty(sc32_fifo_almost_empty), .reset_all(reset_all), 
            .n5384(n5384), .n5385(n5385), .n5386(n5386), .n5387(n5387), 
            .n5388(n5388), .n5389(n5389), .n5390(n5390), .n5391(n5391), 
            .n5392(n5392), .n5393(n5393), .n5394(n5394), .n5395(n5395), 
            .n5396(n5396), .n5397(n5397), .n5398(n5398), .n5399(n5399), 
            .n5400(n5400), .n5401(n5401), .n5402(n5402), .n5403(n5403), 
            .n5404(n5404), .sc32_fifo_write_enable(sc32_fifo_write_enable), 
            .n5405(n5405), .n5406(n5406), .n5407(n5407), .n5408(n5408), 
            .n5409(n5409), .n5410(n5410), .sc32_fifo_read_enable(sc32_fifo_read_enable), 
            .n5413(n5413), .n5414(n5414), .n5411(n5411)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(653[20] 667[2])
    SB_LUT4 i1_2_lut_3_lut_adj_154 (.I0(reset_clk_counter[1]), .I1(reset_all_w_N_61), 
            .I2(reset_clk_counter[0]), .I3(GND_net), .O(n13898));
    defparam i1_2_lut_3_lut_adj_154.LUT_INIT = 16'ha6a6;
    FIFO_Quad_Word tx_fifo (.\rd_addr_r[1] (rd_addr_r_adj_1505[1]), .\rd_addr_r[0] (rd_addr_r_adj_1505[0]), 
            .SLM_CLK_c(SLM_CLK_c), .reset_all_w(reset_all_w), .wr_addr_r({wr_addr_r_adj_1502}), 
            .rx_buf_byte({rx_buf_byte}), .rd_fifo_en_w(rd_fifo_en_w_adj_1413), 
            .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r [0]), .n8(n8), 
            .n7067(n7067), .VCC_net(VCC_net), .\fifo_temp_output[1] (fifo_temp_output[1]), 
            .n4566(n4566), .GND_net(GND_net), .\wr_addr_p1_w[2] (wr_addr_p1_w_adj_1504[2]), 
            .n13820(n13820), .n7064(n7064), .\fifo_temp_output[2] (fifo_temp_output[2]), 
            .n7061(n7061), .\fifo_temp_output[3] (fifo_temp_output[3]), 
            .n7058(n7058), .\fifo_temp_output[4] (fifo_temp_output[4]), 
            .n7055(n7055), .\fifo_temp_output[5] (fifo_temp_output[5]), 
            .n7052(n7052), .\fifo_temp_output[6] (fifo_temp_output[6]), 
            .n7049(n7049), .\fifo_temp_output[7] (fifo_temp_output[7]), 
            .n5647(n5647), .n5658(n5658), .n6970(n6970), .\fifo_temp_output[0] (fifo_temp_output[0]), 
            .n14076(n14076), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .\rd_addr_p1_w[1] (rd_addr_p1_w_adj_1507[1]), .\rd_addr_p1_w[2] (rd_addr_p1_w_adj_1507[2]), 
            .fifo_write_cmd(fifo_write_cmd), .wr_fifo_en_w(wr_fifo_en_w_adj_1412), 
            .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r [1]), .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r [2]), 
            .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r [3]), .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r [4]), 
            .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r [5]), .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r [6]), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r [7]), .fifo_read_cmd(fifo_read_cmd), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .n5664(n5664), .n14096(n14096), 
            .n5207(n5207)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(1057[16] 1073[2])
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_1451[1]), .I1(r_SM_Main_2__N_1026[1]), 
            .I2(r_SM_Main_adj_1451[0]), .I3(r_SM_Main_adj_1451[2]), .O(n18034));   // src/uart_tx.v(38[10] 141[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i4165_2_lut_3_lut (.I0(reset_all_w), .I1(fifo_read_cmd), .I2(is_fifo_empty_flag), 
            .I3(GND_net), .O(n5664));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    defparam i4165_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i5483_2_lut_3_lut (.I0(sc32_fifo_data_out[0]), .I1(bluejay_data_out_31__N_921), 
            .I2(bluejay_data_out_31__N_922), .I3(GND_net), .O(n6982));   // src/bluejay_data.v(134[8] 156[4])
    defparam i5483_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_4_lut_4_lut (.I0(is_tx_fifo_full_flag), .I1(n14603), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_1429));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5465_3_lut_4_lut (.I0(r_SM_Main_2__N_1029[0]), .I1(fifo_read_cmd), 
            .I2(is_fifo_empty_flag), .I3(tx_uart_active_flag), .O(n6964));   // src/top.v(1034[8] 1052[4])
    defparam i5465_3_lut_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4129_4_lut_4_lut (.I0(tx_uart_active_flag), .I1(r_SM_Main_adj_1451[1]), 
            .I2(r_SM_Main_adj_1451[2]), .I3(n14508), .O(n5628));   // src/uart_tx.v(38[10] 141[8])
    defparam i4129_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i4106_2_lut_4_lut (.I0(reset_per_frame), .I1(wr_addr_r[0]), 
            .I2(wr_addr_p1_w[0]), .I3(wr_fifo_en_w), .O(n5605));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4106_2_lut_4_lut.LUT_INIT = 16'h5044;
    fifo_dc_32_lut_gen2 fifo_dc_32_lut_gen_inst (.dc32_fifo_data_in({dc32_fifo_data_in}), 
            .FIFO_CLK_c(FIFO_CLK_c), .GND_net(GND_net), .\REG.mem_22_29 (\REG.mem_22_29 ), 
            .\REG.mem_23_29 (\REG.mem_23_29 ), .\REG.mem_21_29 (\REG.mem_21_29 ), 
            .\REG.mem_11_15 (\REG.mem_11_15 ), .\REG.mem_11_11 (\REG.mem_11_11 ), 
            .\REG.mem_6_26 (\REG.mem_6_26 ), .\REG.mem_7_26 (\REG.mem_7_26 ), 
            .dc32_fifo_almost_full(dc32_fifo_almost_full), .reset_per_frame(reset_per_frame), 
            .\REG.mem_5_26 (\REG.mem_5_26 ), .rd_fifo_en_w(rd_fifo_en_w), 
            .dc32_fifo_data_out({dc32_fifo_data_out}), .SLM_CLK_c(SLM_CLK_c), 
            .\REG.mem_27_29 (\REG.mem_27_29 ), .\REG.mem_11_8 (\REG.mem_11_8 ), 
            .\REG.mem_22_5 (\REG.mem_22_5 ), .\REG.mem_23_5 (\REG.mem_23_5 ), 
            .rd_grey_sync_r({rd_grey_sync_r}), .\REG.mem_21_5 (\REG.mem_21_5 ), 
            .dc32_fifo_full(dc32_fifo_full), .\REG.mem_6_20 (\REG.mem_6_20 ), 
            .\REG.mem_7_20 (\REG.mem_7_20 ), .empty_nxt_c_N_636(empty_nxt_c_N_636), 
            .dc32_fifo_empty(dc32_fifo_empty), .\REG.mem_5_20 (\REG.mem_5_20 ), 
            .\wr_grey_sync_r[0] (wr_grey_sync_r[0]), .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .\rd_addr_nxt_c_5__N_573[3] (rd_addr_nxt_c_5__N_573[3]), .\rd_addr_nxt_c_5__N_573[1] (rd_addr_nxt_c_5__N_573[1]), 
            .\REG.mem_11_20 (\REG.mem_11_20 ), .\REG.mem_11_21 (\REG.mem_11_21 ), 
            .\REG.mem_27_12 (\REG.mem_27_12 ), .\REG.mem_22_11 (\REG.mem_22_11 ), 
            .\REG.mem_23_11 (\REG.mem_23_11 ), .\REG.mem_21_11 (\REG.mem_21_11 ), 
            .\REG.mem_27_3 (\REG.mem_27_3 ), .\REG.mem_11_10 (\REG.mem_11_10 ), 
            .\REG.mem_22_28 (\REG.mem_22_28 ), .\REG.mem_23_28 (\REG.mem_23_28 ), 
            .\REG.mem_21_28 (\REG.mem_21_28 ), .\REG.mem_27_0 (\REG.mem_27_0 ), 
            .\REG.mem_6_19 (\REG.mem_6_19 ), .\REG.mem_7_19 (\REG.mem_7_19 ), 
            .\REG.mem_5_19 (\REG.mem_5_19 ), .\REG.mem_6_9 (\REG.mem_6_9 ), 
            .\REG.mem_7_9 (\REG.mem_7_9 ), .\REG.mem_11_0 (\REG.mem_11_0 ), 
            .\REG.mem_5_9 (\REG.mem_5_9 ), .\REG.mem_11_13 (\REG.mem_11_13 ), 
            .\REG.mem_6_14 (\REG.mem_6_14 ), .\REG.mem_7_14 (\REG.mem_7_14 ), 
            .\REG.mem_5_14 (\REG.mem_5_14 ), .\REG.mem_22_19 (\REG.mem_22_19 ), 
            .\REG.mem_23_19 (\REG.mem_23_19 ), .\REG.mem_21_19 (\REG.mem_21_19 ), 
            .\REG.mem_27_19 (\REG.mem_27_19 ), .n6(n6), .n22(n22), .\REG.mem_11_14 (\REG.mem_11_14 ), 
            .\REG.mem_22_9 (\REG.mem_22_9 ), .\REG.mem_23_9 (\REG.mem_23_9 ), 
            .\REG.mem_21_9 (\REG.mem_21_9 ), .\REG.mem_6_24 (\REG.mem_6_24 ), 
            .\REG.mem_7_24 (\REG.mem_7_24 ), .\REG.mem_22_1 (\REG.mem_22_1 ), 
            .\REG.mem_23_1 (\REG.mem_23_1 ), .wr_fifo_en_w(wr_fifo_en_w), 
            .\wr_addr_nxt_c[4] (wr_addr_nxt_c[4]), .\wr_addr_nxt_c[2] (wr_addr_nxt_c[2]), 
            .\REG.mem_22_16 (\REG.mem_22_16 ), .\REG.mem_23_16 (\REG.mem_23_16 ), 
            .\REG.mem_21_1 (\REG.mem_21_1 ), .\REG.mem_21_16 (\REG.mem_21_16 ), 
            .\REG.mem_11_12 (\REG.mem_11_12 ), .\REG.mem_5_24 (\REG.mem_5_24 ), 
            .n7038(n7038), .n7037(n7037), .n7036(n7036), .n7035(n7035), 
            .n7034(n7034), .n7033(n7033), .wp_sync1_r({wp_sync1_r}), .n7032(n7032), 
            .n7031(n7031), .n7030(n7030), .n7029(n7029), .n7028(n7028), 
            .n7027(n7027), .n7025(n7025), .n7023(n7023), .n7022(n7022), 
            .n7021(n7021), .n7020(n7020), .n7019(n7019), .n7018(n7018), 
            .rp_sync1_r({rp_sync1_r}), .n7017(n7017), .n7016(n7016), .n7015(n7015), 
            .n7014(n7014), .n6955(n6955), .n6953(n6953), .\wr_addr_r[5] (wr_addr_r[5]), 
            .n6532(n6532), .\REG.mem_27_31 (\REG.mem_27_31 ), .n6531(n6531), 
            .\REG.mem_27_30 (\REG.mem_27_30 ), .n6530(n6530), .n6529(n6529), 
            .\REG.mem_27_28 (\REG.mem_27_28 ), .n6528(n6528), .\REG.mem_27_27 (\REG.mem_27_27 ), 
            .n6527(n6527), .\REG.mem_27_26 (\REG.mem_27_26 ), .n6526(n6526), 
            .\REG.mem_27_25 (\REG.mem_27_25 ), .n6525(n6525), .\REG.mem_27_24 (\REG.mem_27_24 ), 
            .n6524(n6524), .\REG.mem_27_23 (\REG.mem_27_23 ), .n6523(n6523), 
            .\REG.mem_27_22 (\REG.mem_27_22 ), .n6522(n6522), .\REG.mem_27_21 (\REG.mem_27_21 ), 
            .n6521(n6521), .\REG.mem_27_20 (\REG.mem_27_20 ), .n6520(n6520), 
            .n6519(n6519), .\REG.mem_27_18 (\REG.mem_27_18 ), .n6518(n6518), 
            .\REG.mem_27_17 (\REG.mem_27_17 ), .n6517(n6517), .\REG.mem_27_16 (\REG.mem_27_16 ), 
            .n6516(n6516), .\REG.mem_27_15 (\REG.mem_27_15 ), .n6515(n6515), 
            .\REG.mem_27_14 (\REG.mem_27_14 ), .n6514(n6514), .\REG.mem_27_13 (\REG.mem_27_13 ), 
            .n6513(n6513), .n6512(n6512), .\REG.mem_27_11 (\REG.mem_27_11 ), 
            .n6511(n6511), .\REG.mem_27_10 (\REG.mem_27_10 ), .n6510(n6510), 
            .\REG.mem_27_9 (\REG.mem_27_9 ), .n6509(n6509), .\REG.mem_27_8 (\REG.mem_27_8 ), 
            .n6508(n6508), .\REG.mem_27_7 (\REG.mem_27_7 ), .n6507(n6507), 
            .\REG.mem_27_6 (\REG.mem_27_6 ), .n6506(n6506), .\REG.mem_27_5 (\REG.mem_27_5 ), 
            .n6505(n6505), .\REG.mem_27_4 (\REG.mem_27_4 ), .n6504(n6504), 
            .n6503(n6503), .\REG.mem_27_2 (\REG.mem_27_2 ), .n6502(n6502), 
            .\REG.mem_27_1 (\REG.mem_27_1 ), .n6501(n6501), .n6404(n6404), 
            .\REG.mem_23_31 (\REG.mem_23_31 ), .n6403(n6403), .\REG.mem_23_30 (\REG.mem_23_30 ), 
            .n6402(n6402), .n6401(n6401), .n6400(n6400), .\REG.mem_23_27 (\REG.mem_23_27 ), 
            .n6399(n6399), .\REG.mem_23_26 (\REG.mem_23_26 ), .n6398(n6398), 
            .\REG.mem_23_25 (\REG.mem_23_25 ), .n6397(n6397), .\REG.mem_23_24 (\REG.mem_23_24 ), 
            .n6396(n6396), .\REG.mem_23_23 (\REG.mem_23_23 ), .n6395(n6395), 
            .\REG.mem_23_22 (\REG.mem_23_22 ), .n6394(n6394), .\REG.mem_23_21 (\REG.mem_23_21 ), 
            .n6393(n6393), .\REG.mem_23_20 (\REG.mem_23_20 ), .n6392(n6392), 
            .n6391(n6391), .\REG.mem_23_18 (\REG.mem_23_18 ), .n6390(n6390), 
            .\REG.mem_23_17 (\REG.mem_23_17 ), .n6389(n6389), .n6388(n6388), 
            .\REG.mem_23_15 (\REG.mem_23_15 ), .n6387(n6387), .\REG.mem_23_14 (\REG.mem_23_14 ), 
            .n6386(n6386), .\REG.mem_23_13 (\REG.mem_23_13 ), .n6385(n6385), 
            .\REG.mem_23_12 (\REG.mem_23_12 ), .n6384(n6384), .n6383(n6383), 
            .\REG.mem_23_10 (\REG.mem_23_10 ), .n6382(n6382), .n6381(n6381), 
            .\REG.mem_23_8 (\REG.mem_23_8 ), .n6380(n6380), .\REG.mem_23_7 (\REG.mem_23_7 ), 
            .n6379(n6379), .\REG.mem_23_6 (\REG.mem_23_6 ), .n6378(n6378), 
            .n6377(n6377), .\REG.mem_23_4 (\REG.mem_23_4 ), .n6376(n6376), 
            .\REG.mem_23_3 (\REG.mem_23_3 ), .n6375(n6375), .\REG.mem_23_2 (\REG.mem_23_2 ), 
            .n6374(n6374), .n6373(n6373), .\REG.mem_23_0 (\REG.mem_23_0 ), 
            .n6372(n6372), .\REG.mem_22_31 (\REG.mem_22_31 ), .n6371(n6371), 
            .\REG.mem_22_30 (\REG.mem_22_30 ), .n6370(n6370), .n6369(n6369), 
            .n6368(n6368), .\REG.mem_22_27 (\REG.mem_22_27 ), .n6367(n6367), 
            .\REG.mem_22_26 (\REG.mem_22_26 ), .n6366(n6366), .\REG.mem_22_25 (\REG.mem_22_25 ), 
            .n6365(n6365), .\REG.mem_22_24 (\REG.mem_22_24 ), .n6364(n6364), 
            .\REG.mem_22_23 (\REG.mem_22_23 ), .n6363(n6363), .\REG.mem_22_22 (\REG.mem_22_22 ), 
            .n6362(n6362), .\REG.mem_22_21 (\REG.mem_22_21 ), .n6361(n6361), 
            .\REG.mem_22_20 (\REG.mem_22_20 ), .n6360(n6360), .n6359(n6359), 
            .\REG.mem_22_18 (\REG.mem_22_18 ), .n6358(n6358), .\REG.mem_22_17 (\REG.mem_22_17 ), 
            .n6357(n6357), .n6356(n6356), .\REG.mem_22_15 (\REG.mem_22_15 ), 
            .n6355(n6355), .\REG.mem_22_14 (\REG.mem_22_14 ), .n6354(n6354), 
            .\REG.mem_22_13 (\REG.mem_22_13 ), .n6353(n6353), .\REG.mem_22_12 (\REG.mem_22_12 ), 
            .n6352(n6352), .n6351(n6351), .\REG.mem_22_10 (\REG.mem_22_10 ), 
            .n6350(n6350), .n6349(n6349), .\REG.mem_22_8 (\REG.mem_22_8 ), 
            .n6348(n6348), .\REG.mem_22_7 (\REG.mem_22_7 ), .n6347(n6347), 
            .\REG.mem_22_6 (\REG.mem_22_6 ), .n6346(n6346), .n6345(n6345), 
            .\REG.mem_22_4 (\REG.mem_22_4 ), .n6344(n6344), .\REG.mem_22_3 (\REG.mem_22_3 ), 
            .n6343(n6343), .\REG.mem_22_2 (\REG.mem_22_2 ), .n6342(n6342), 
            .n6341(n6341), .\REG.mem_22_0 (\REG.mem_22_0 ), .n6340(n6340), 
            .\REG.mem_21_31 (\REG.mem_21_31 ), .n6339(n6339), .\REG.mem_21_30 (\REG.mem_21_30 ), 
            .n6338(n6338), .n6337(n6337), .n6336(n6336), .\REG.mem_21_27 (\REG.mem_21_27 ), 
            .n6335(n6335), .\REG.mem_21_26 (\REG.mem_21_26 ), .n6334(n6334), 
            .\REG.mem_21_25 (\REG.mem_21_25 ), .n6333(n6333), .\REG.mem_21_24 (\REG.mem_21_24 ), 
            .n6332(n6332), .\REG.mem_21_23 (\REG.mem_21_23 ), .n6331(n6331), 
            .\REG.mem_21_22 (\REG.mem_21_22 ), .n6330(n6330), .\REG.mem_21_21 (\REG.mem_21_21 ), 
            .n6329(n6329), .\REG.mem_21_20 (\REG.mem_21_20 ), .n6328(n6328), 
            .n6327(n6327), .\REG.mem_21_18 (\REG.mem_21_18 ), .n6326(n6326), 
            .\REG.mem_21_17 (\REG.mem_21_17 ), .n6325(n6325), .n6324(n6324), 
            .\REG.mem_21_15 (\REG.mem_21_15 ), .n6323(n6323), .\REG.mem_21_14 (\REG.mem_21_14 ), 
            .n6322(n6322), .\REG.mem_21_13 (\REG.mem_21_13 ), .n6321(n6321), 
            .\REG.mem_21_12 (\REG.mem_21_12 ), .n6320(n6320), .n6319(n6319), 
            .\REG.mem_21_10 (\REG.mem_21_10 ), .n6318(n6318), .n6317(n6317), 
            .\REG.mem_21_8 (\REG.mem_21_8 ), .n6316(n6316), .\REG.mem_21_7 (\REG.mem_21_7 ), 
            .n6315(n6315), .\REG.mem_21_6 (\REG.mem_21_6 ), .n6314(n6314), 
            .n6313(n6313), .\REG.mem_21_4 (\REG.mem_21_4 ), .n6312(n6312), 
            .\REG.mem_21_3 (\REG.mem_21_3 ), .n6311(n6311), .\REG.mem_21_2 (\REG.mem_21_2 ), 
            .n6310(n6310), .n6309(n6309), .\REG.mem_21_0 (\REG.mem_21_0 ), 
            .n12(n12_adj_1415), .n10(n10), .n26(n26), .\rd_addr_nxt_c_5__N_573[4] (rd_addr_nxt_c_5__N_573[4]), 
            .\REG.mem_6_22 (\REG.mem_6_22 ), .\REG.mem_7_22 (\REG.mem_7_22 ), 
            .\REG.mem_6_23 (\REG.mem_6_23 ), .\REG.mem_7_23 (\REG.mem_7_23 ), 
            .\REG.mem_5_23 (\REG.mem_5_23 ), .\REG.mem_5_22 (\REG.mem_5_22 ), 
            .\REG.mem_11_23 (\REG.mem_11_23 ), .\REG.mem_11_18 (\REG.mem_11_18 ), 
            .\REG.mem_6_7 (\REG.mem_6_7 ), .\REG.mem_7_7 (\REG.mem_7_7 ), 
            .\REG.mem_5_7 (\REG.mem_5_7 ), .\REG.mem_11_9 (\REG.mem_11_9 ), 
            .n7(n7_adj_1427), .\REG.mem_6_28 (\REG.mem_6_28 ), .\REG.mem_7_28 (\REG.mem_7_28 ), 
            .\REG.mem_5_28 (\REG.mem_5_28 ), .n8(n8_adj_1426), .\REG.mem_11_28 (\REG.mem_11_28 ), 
            .VCC_net(VCC_net), .n25(n25_adj_1430), .\REG.mem_11_25 (\REG.mem_11_25 ), 
            .\wr_grey_sync_r[1] (wr_grey_sync_r[1]), .\wr_grey_sync_r[2] (wr_grey_sync_r[2]), 
            .\REG.mem_11_5 (\REG.mem_11_5 ), .\wr_grey_sync_r[3] (wr_grey_sync_r[3]), 
            .\wr_grey_sync_r[4] (wr_grey_sync_r[4]), .n6020(n6020), .\REG.mem_11_31 (\REG.mem_11_31 ), 
            .n6019(n6019), .\REG.mem_11_30 (\REG.mem_11_30 ), .n6018(n6018), 
            .\REG.mem_11_29 (\REG.mem_11_29 ), .n6017(n6017), .n6016(n6016), 
            .\REG.mem_11_27 (\REG.mem_11_27 ), .n6015(n6015), .\REG.mem_11_26 (\REG.mem_11_26 ), 
            .n6014(n6014), .n6013(n6013), .\REG.mem_11_24 (\REG.mem_11_24 ), 
            .n6012(n6012), .n6011(n6011), .\REG.mem_11_22 (\REG.mem_11_22 ), 
            .n6010(n6010), .n6009(n6009), .n6008(n6008), .\REG.mem_11_19 (\REG.mem_11_19 ), 
            .n6007(n6007), .\REG.mem_11_6 (\REG.mem_11_6 ), .n6006(n6006), 
            .\REG.mem_11_17 (\REG.mem_11_17 ), .n6005(n6005), .\REG.mem_11_16 (\REG.mem_11_16 ), 
            .n6004(n6004), .n6003(n6003), .n6002(n6002), .n6001(n6001), 
            .n6000(n6000), .n5999(n5999), .n5998(n5998), .\wr_addr_r[0] (wr_addr_r[0]), 
            .DEBUG_5_c(DEBUG_5_c), .\REG.mem_11_2 (\REG.mem_11_2 ), .n5997(n5997), 
            .n5996(n5996), .\REG.mem_11_7 (\REG.mem_11_7 ), .n5995(n5995), 
            .n5994(n5994), .n5993(n5993), .\REG.mem_11_4 (\REG.mem_11_4 ), 
            .\wr_addr_p1_w[0] (wr_addr_p1_w[0]), .n13865(n13865), .n14706(n14706), 
            .n5992(n5992), .\REG.mem_11_3 (\REG.mem_11_3 ), .n5991(n5991), 
            .n5990(n5990), .\REG.mem_11_1 (\REG.mem_11_1 ), .FT_OE_N_496(FT_OE_N_496), 
            .n12_adj_4(n12), .dc32_fifo_read_enable(dc32_fifo_read_enable), 
            .n5989(n5989), .n5892(n5892), .\REG.mem_7_31 (\REG.mem_7_31 ), 
            .n5891(n5891), .\REG.mem_7_30 (\REG.mem_7_30 ), .n5890(n5890), 
            .\REG.mem_7_29 (\REG.mem_7_29 ), .n5889(n5889), .n5888(n5888), 
            .\REG.mem_7_27 (\REG.mem_7_27 ), .n5887(n5887), .n5886(n5886), 
            .\REG.mem_7_25 (\REG.mem_7_25 ), .n5885(n5885), .n5884(n5884), 
            .n5883(n5883), .n5882(n5882), .\REG.mem_7_21 (\REG.mem_7_21 ), 
            .n5881(n5881), .n5880(n5880), .n5879(n5879), .\REG.mem_7_18 (\REG.mem_7_18 ), 
            .n5878(n5878), .\REG.mem_7_17 (\REG.mem_7_17 ), .n5877(n5877), 
            .\REG.mem_7_16 (\REG.mem_7_16 ), .n5876(n5876), .\REG.mem_7_15 (\REG.mem_7_15 ), 
            .n5875(n5875), .n5874(n5874), .\REG.mem_7_13 (\REG.mem_7_13 ), 
            .n5873(n5873), .\REG.mem_7_12 (\REG.mem_7_12 ), .n5872(n5872), 
            .\REG.mem_7_11 (\REG.mem_7_11 ), .n5871(n5871), .\REG.mem_7_10 (\REG.mem_7_10 ), 
            .n5870(n5870), .n5869(n5869), .\REG.mem_7_8 (\REG.mem_7_8 ), 
            .n5868(n5868), .n5867(n5867), .\REG.mem_7_6 (\REG.mem_7_6 ), 
            .n5866(n5866), .\REG.mem_7_5 (\REG.mem_7_5 ), .n5865(n5865), 
            .\REG.mem_7_4 (\REG.mem_7_4 ), .n5864(n5864), .\REG.mem_7_3 (\REG.mem_7_3 ), 
            .n5863(n5863), .\REG.mem_7_2 (\REG.mem_7_2 ), .n5862(n5862), 
            .\REG.mem_7_1 (\REG.mem_7_1 ), .n5861(n5861), .\REG.mem_7_0 (\REG.mem_7_0 ), 
            .n5860(n5860), .\REG.mem_6_31 (\REG.mem_6_31 ), .n5859(n5859), 
            .\REG.mem_6_30 (\REG.mem_6_30 ), .n5858(n5858), .\REG.mem_6_29 (\REG.mem_6_29 ), 
            .n5857(n5857), .n5856(n5856), .\REG.mem_6_27 (\REG.mem_6_27 ), 
            .n5855(n5855), .n5854(n5854), .\REG.mem_6_25 (\REG.mem_6_25 ), 
            .n5853(n5853), .n5852(n5852), .n5851(n5851), .\state[3] (state[3]), 
            .n4843(n4843), .n1224(n1224), .n5850(n5850), .\REG.mem_6_21 (\REG.mem_6_21 ), 
            .n5849(n5849), .n5848(n5848), .n5847(n5847), .\REG.mem_6_18 (\REG.mem_6_18 ), 
            .n5846(n5846), .\REG.mem_6_17 (\REG.mem_6_17 ), .n5845(n5845), 
            .\REG.mem_6_16 (\REG.mem_6_16 ), .n5844(n5844), .\REG.mem_6_15 (\REG.mem_6_15 ), 
            .n5843(n5843), .n5842(n5842), .\REG.mem_6_13 (\REG.mem_6_13 ), 
            .n5841(n5841), .\REG.mem_6_12 (\REG.mem_6_12 ), .n5840(n5840), 
            .\REG.mem_6_11 (\REG.mem_6_11 ), .n5839(n5839), .\REG.mem_6_10 (\REG.mem_6_10 ), 
            .n5838(n5838), .n5837(n5837), .\REG.mem_6_8 (\REG.mem_6_8 ), 
            .n5836(n5836), .n5835(n5835), .\REG.mem_6_6 (\REG.mem_6_6 ), 
            .n5834(n5834), .\REG.mem_6_5 (\REG.mem_6_5 ), .n5833(n5833), 
            .\REG.mem_6_4 (\REG.mem_6_4 ), .\REG.mem_6_2 (\REG.mem_6_2 ), 
            .n5832(n5832), .\REG.mem_6_3 (\REG.mem_6_3 ), .n5831(n5831), 
            .\REG.mem_5_2 (\REG.mem_5_2 ), .n5830(n5830), .\REG.mem_6_1 (\REG.mem_6_1 ), 
            .n5829(n5829), .\REG.mem_6_0 (\REG.mem_6_0 ), .n5828(n5828), 
            .\REG.mem_5_31 (\REG.mem_5_31 ), .n5827(n5827), .\REG.mem_5_30 (\REG.mem_5_30 ), 
            .n5826(n5826), .\REG.mem_5_29 (\REG.mem_5_29 ), .n5825(n5825), 
            .n5824(n5824), .\REG.mem_5_27 (\REG.mem_5_27 ), .n5823(n5823), 
            .n5822(n5822), .\REG.mem_5_25 (\REG.mem_5_25 ), .n5821(n5821), 
            .n5820(n5820), .n5819(n5819), .n5818(n5818), .\REG.mem_5_21 (\REG.mem_5_21 ), 
            .n5817(n5817), .n5816(n5816), .n5815(n5815), .\REG.mem_5_18 (\REG.mem_5_18 ), 
            .n5814(n5814), .\REG.mem_5_17 (\REG.mem_5_17 ), .n5813(n5813), 
            .\REG.mem_5_16 (\REG.mem_5_16 ), .n5812(n5812), .\REG.mem_5_15 (\REG.mem_5_15 ), 
            .n5811(n5811), .n5810(n5810), .\REG.mem_5_13 (\REG.mem_5_13 ), 
            .n5809(n5809), .\REG.mem_5_12 (\REG.mem_5_12 ), .n5808(n5808), 
            .\REG.mem_5_11 (\REG.mem_5_11 ), .n5807(n5807), .\REG.mem_5_10 (\REG.mem_5_10 ), 
            .n5806(n5806), .n5805(n5805), .\REG.mem_5_8 (\REG.mem_5_8 ), 
            .n5804(n5804), .n5803(n5803), .\REG.mem_5_6 (\REG.mem_5_6 ), 
            .n5802(n5802), .\REG.mem_5_5 (\REG.mem_5_5 ), .n5648(n5648), 
            .n5801(n5801), .\REG.mem_5_4 (\REG.mem_5_4 ), .n5800(n5800), 
            .\REG.mem_5_3 (\REG.mem_5_3 ), .n5642(n5642), .n5639(n5639), 
            .n5638(n5638), .n5799(n5799), .n5798(n5798), .\REG.mem_5_1 (\REG.mem_5_1 ), 
            .n5797(n5797), .\REG.mem_5_0 (\REG.mem_5_0 ), .n5605(n5605), 
            .n27(n27), .n11(n11), .n28(n28)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(612[21] 628[2])
    SB_LUT4 i3919_1_lut_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n5418));   // src/top.v(1198[8] 1265[4])
    defparam i3919_1_lut_2_lut.LUT_INIT = 16'h7777;
    clock clock_inst (.GND_net(GND_net), .VCC_net(VCC_net), .ICE_SYSCLK_c(ICE_SYSCLK_c), 
          .pll_clk_unbuf(pll_clk_unbuf)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(222[7] 228[3])
    spi spi0 (.SLM_CLK_c(SLM_CLK_c), .SOUT_c(SOUT_c), .n5025(n5025), .\rx_shift_reg[0] (rx_shift_reg[0]), 
        .n4999(n4999), .SDAT_c_15(SDAT_c_15), .n7013(n7013), .rx_buf_byte({rx_buf_byte}), 
        .n7012(n7012), .n7011(n7011), .n7010(n7010), .n7009(n7009), 
        .n7008(n7008), .n7007(n7007), .n7006(n7006), .\rx_shift_reg[7] (rx_shift_reg[7]), 
        .n7005(n7005), .\rx_shift_reg[6] (rx_shift_reg[6]), .n7004(n7004), 
        .\rx_shift_reg[5] (rx_shift_reg[5]), .n7003(n7003), .\rx_shift_reg[4] (rx_shift_reg[4]), 
        .n7002(n7002), .\rx_shift_reg[3] (rx_shift_reg[3]), .n7001(n7001), 
        .\rx_shift_reg[2] (rx_shift_reg[2]), .n7000(n7000), .\rx_shift_reg[1] (rx_shift_reg[1]), 
        .n14116(n14116), .VCC_net(VCC_net), .\tx_shift_reg[0] (tx_shift_reg[0]), 
        .multi_byte_spi_trans_flag_r(multi_byte_spi_trans_flag_r), .GND_net(GND_net), 
        .n2555(n2555), .spi_start_transfer_r(spi_start_transfer_r), .tx_addr_byte({tx_addr_byte}), 
        .SEN_c_1(SEN_c_1), .spi_rx_byte_ready(spi_rx_byte_ready), .SCK_c_0(SCK_c_0), 
        .n5636(n5636), .\tx_data_byte[7] (tx_data_byte[7]), .\tx_data_byte[6] (tx_data_byte[6]), 
        .\tx_data_byte[5] (tx_data_byte[5]), .\tx_data_byte[4] (tx_data_byte[4]), 
        .\tx_data_byte[3] (tx_data_byte[3]), .\tx_data_byte[2] (tx_data_byte[2]), 
        .\tx_data_byte[1] (tx_data_byte[1]), .n4086(n4086)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(957[5] 981[2])
    \uart_rx(CLKS_PER_BIT=20)  pc_rx (.n14672(n14672), .SLM_CLK_c(SLM_CLK_c), 
            .n14688(n14688), .r_Rx_Data(r_Rx_Data), .DEBUG_2_c_c(DEBUG_2_c_c), 
            .n4935(n4935), .GND_net(GND_net), .n4(n4), .n4_adj_1(n4_adj_1417), 
            .\r_Bit_Index[0] (r_Bit_Index[0]), .n4942(n4942), .n4938(n4938), 
            .n4_adj_2(n4_adj_1416), .n6981(n6981), .pc_data_rx({pc_data_rx}), 
            .VCC_net(VCC_net), .debug_led3(debug_led3), .n6977(n6977), 
            .n5624(n5624), .n5620(n5620), .n5613(n5613), .n5612(n5612), 
            .n5611(n5611), .n5609(n5609), .n5608(n5608)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(823[42] 828[3])
    SB_LUT4 i4814_3_lut (.I0(\REG.mem_21_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n12_adj_1415), .I3(GND_net), .O(n6313));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4814_3_lut.LUT_INIT = 16'hcaca;
    \uart_tx(CLKS_PER_BIT=20)  pc_tx (.n14684(n14684), .SLM_CLK_c(SLM_CLK_c), 
            .n14690(n14690), .DEBUG_1_c(DEBUG_1_c), .r_SM_Main({r_SM_Main_adj_1451}), 
            .\r_SM_Main_2__N_1026[1] (r_SM_Main_2__N_1026[1]), .\r_SM_Main_2__N_1029[0] (r_SM_Main_2__N_1029[0]), 
            .n14508(n14508), .\r_Bit_Index[0] (r_Bit_Index_adj_1453[0]), 
            .r_Tx_Data({r_Tx_Data}), .GND_net(GND_net), .n18034(n18034), 
            .n6999(n6999), .n6998(n6998), .n6997(n6997), .n6996(n6996), 
            .n6995(n6995), .n6994(n6994), .n6993(n6993), .n6974(n6974), 
            .VCC_net(VCC_net), .n4435(n4435), .n5629(n5629), .n5628(n5628), 
            .tx_uart_active_flag(tx_uart_active_flag)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(892[42] 901[3])
    usb3_if usb3_if_inst (.FIFO_CLK_c(FIFO_CLK_c), .reset_per_frame(reset_per_frame), 
            .SLM_CLK_c(SLM_CLK_c), .dc32_fifo_empty(dc32_fifo_empty), .VCC_net(VCC_net), 
            .FT_RD_c(FT_RD_c), .dc32_fifo_data_in({dc32_fifo_data_in}), 
            .DEBUG_5_c(DEBUG_5_c), .buffer_switch_done(buffer_switch_done), 
            .buffer_switch_done_latched(buffer_switch_done_latched), .FT_OE_N_496(FT_OE_N_496), 
            .GND_net(GND_net), .FIFO_D0_c_31(FIFO_D0_c_31), .FIFO_D1_c_30(FIFO_D1_c_30), 
            .FIFO_D2_c_29(FIFO_D2_c_29), .DEBUG_9_c_c(DEBUG_9_c_c), .FIFO_D3_c_28(FIFO_D3_c_28), 
            .FIFO_D4_c_27(FIFO_D4_c_27), .FIFO_D5_c_26(FIFO_D5_c_26), .FIFO_D6_c_25(FIFO_D6_c_25), 
            .FIFO_D7_c_24(FIFO_D7_c_24), .FIFO_D8_c_23(FIFO_D8_c_23), .FIFO_D9_c_22(FIFO_D9_c_22), 
            .FIFO_D10_c_21(FIFO_D10_c_21), .FIFO_D31_c_0(FIFO_D31_c_0), 
            .FIFO_D11_c_20(FIFO_D11_c_20), .FIFO_D12_c_19(FIFO_D12_c_19), 
            .FIFO_D13_c_18(FIFO_D13_c_18), .FIFO_D14_c_17(FIFO_D14_c_17), 
            .FIFO_D15_c_16(FIFO_D15_c_16), .FIFO_D16_c_15(FIFO_D16_c_15), 
            .FIFO_D17_c_14(FIFO_D17_c_14), .FIFO_D18_c_13(FIFO_D18_c_13), 
            .FIFO_D19_c_12(FIFO_D19_c_12), .FIFO_D20_c_11(FIFO_D20_c_11), 
            .FIFO_D21_c_10(FIFO_D21_c_10), .FIFO_D22_c_9(FIFO_D22_c_9), 
            .FT_OE_c(FT_OE_c), .FIFO_D23_c_8(FIFO_D23_c_8), .FIFO_D24_c_7(FIFO_D24_c_7), 
            .FIFO_D25_c_6(FIFO_D25_c_6), .FIFO_D26_c_5(FIFO_D26_c_5), .FIFO_D27_c_4(FIFO_D27_c_4), 
            .n12(n12), .FIFO_D28_c_3(FIFO_D28_c_3), .n14706(n14706), .n13865(n13865), 
            .rd_fifo_en_w(rd_fifo_en_w), .empty_nxt_c_N_636(empty_nxt_c_N_636), 
            .dc32_fifo_almost_full(dc32_fifo_almost_full), .FIFO_D29_c_2(FIFO_D29_c_2), 
            .dc32_fifo_full(dc32_fifo_full), .wr_fifo_en_w(wr_fifo_en_w), 
            .FIFO_D30_c_1(FIFO_D30_c_1)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(577[9] 593[3])
    
endmodule
//
// Verilog Description of module timing_controller
//

module timing_controller (SLM_CLK_c, sc32_fifo_write_enable, sc32_fifo_read_enable, 
            n14567, state, dc32_fifo_read_enable, buffer_switch_done, 
            n5043, GND_net, VCC_net, n2283, n14118, n1224, n63, 
            n5077, line_of_data_available, n2178, INVERT_c_4, n7, 
            n8, \aempty_flag_impl.ae_flag_nxt_w , get_next_word, dc32_fifo_full, 
            reset_all, n9752, n10059, n14542, reset_per_frame, n25, 
            UPDATE_c_3, n14692, n10051, n4843, n910, n989, n1028, 
            buffer_switch_done_latched, n14482, n5529, bluejay_data_out_31__N_920, 
            n5528, bluejay_data_out_31__N_919, n5431) /* synthesis syn_module_defined=1 */ ;
    input SLM_CLK_c;
    output sc32_fifo_write_enable;
    output sc32_fifo_read_enable;
    input n14567;
    output [3:0]state;
    output dc32_fifo_read_enable;
    output buffer_switch_done;
    output n5043;
    input GND_net;
    input VCC_net;
    input n2283;
    input n14118;
    input n1224;
    output n63;
    input n5077;
    output line_of_data_available;
    input n2178;
    output INVERT_c_4;
    input n7;
    input n8;
    output \aempty_flag_impl.ae_flag_nxt_w ;
    input get_next_word;
    input dc32_fifo_full;
    output reset_all;
    input n9752;
    output n10059;
    input n14542;
    output reset_per_frame;
    output n25;
    output UPDATE_c_3;
    output n14692;
    input n10051;
    output n4843;
    input n910;
    input n989;
    output n1028;
    input buffer_switch_done_latched;
    input n14482;
    output n5529;
    input bluejay_data_out_31__N_920;
    output n5528;
    input bluejay_data_out_31__N_919;
    output n5431;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [31:0]n2356;
    
    wire n4989;
    wire [31:0]state_timeout_counter;   // src/timing_controller.v(80[12:33])
    
    wire sc32_fifo_write_enable_N_366, sc32_fifo_read_enable_N_367;
    wire [2:0]fifo_state_2__N_80;
    
    wire n14700;
    wire [2:0]fifo_state;   // src/timing_controller.v(77[11:21])
    wire [3:0]state_3__N_83;
    
    wire dc32_fifo_read_enable_N_359;
    wire [6:0]fifo_state_timeout_counter_5__N_125;
    
    wire n7_c, n14511, n14532, n14533;
    wire [5:0]fifo_state_timeout_counter;   // src/timing_controller.v(79[11:37])
    
    wire n4, n94;
    wire [31:0]n628;
    
    wire n5446, n16071, n13716;
    wire [31:0]n2179;
    wire [31:0]n2284;
    
    wire n15917, n15918, n14494, n14495, n15940, n2355, n9126, 
        n9122, n13147, n15, n5453, n17, n14544, n15916, n15915, 
        n14557, n15914, n13717, n13715, n13687, n13688, n14130, 
        n2, n8104, n13714, n13713, n13686, n15912, n13685, n15913, 
        n13684, n14538, n13683, n13682, n13681;
    wire [4:0]n1114;
    
    wire n13680, n13679, n13678, n13677, n13676, n13675, n13674, 
        n13673, n13697, n13696, n13695, n13672, n13694, n15941, 
        n13671, n13693, n13692, n13670, n13691, n13669, n13690, 
        n13173, n15906, n16, n7_adj_1410, n10029, n18, n14643, 
        n14682, n2437, n6, n14546, n15958, n11, n13689, n13668, 
        n13667, n15900, n5, n38, n52, n56, n54, n55, n53, 
        n50, n58, n62, n49, n15922;
    
    SB_DFFE state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(SLM_CLK_c), 
            .E(n4989), .D(n2356[0]));   // src/timing_controller.v(153[8] 229[4])
    SB_DFF sc32_fifo_write_enable_89 (.Q(sc32_fifo_write_enable), .C(SLM_CLK_c), 
           .D(sc32_fifo_write_enable_N_366));   // src/timing_controller.v(88[8] 150[4])
    SB_DFF sc32_fifo_read_enable_90 (.Q(sc32_fifo_read_enable), .C(SLM_CLK_c), 
           .D(sc32_fifo_read_enable_N_367));   // src/timing_controller.v(88[8] 150[4])
    SB_DFFE fifo_state_i0 (.Q(fifo_state[0]), .C(SLM_CLK_c), .E(n14700), 
            .D(fifo_state_2__N_80[0]));   // src/timing_controller.v(88[8] 150[4])
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n14567), .D(state_3__N_83[0]));   // src/timing_controller.v(153[8] 229[4])
    SB_DFF dc32_fifo_read_enable_88 (.Q(dc32_fifo_read_enable), .C(SLM_CLK_c), 
           .D(dc32_fifo_read_enable_N_359));   // src/timing_controller.v(88[8] 150[4])
    SB_LUT4 i14017_4_lut (.I0(fifo_state[1]), .I1(fifo_state_timeout_counter_5__N_125[3]), 
            .I2(fifo_state[0]), .I3(n7_c), .O(n14511));
    defparam i14017_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 state_3__I_0_103_Mux_2_i15_4_lut (.I0(state[1]), .I1(state[2]), 
            .I2(state[3]), .I3(state[0]), .O(state_3__N_83[2]));   // src/timing_controller.v(159[5] 228[12])
    defparam state_3__I_0_103_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(state[3]), 
            .I3(state[2]), .O(n14532));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_4_lut_adj_136 (.I0(state[0]), .I1(state[1]), .I2(state[3]), 
            .I3(state[2]), .O(n14533));
    defparam i1_2_lut_4_lut_adj_136.LUT_INIT = 16'h0200;
    SB_LUT4 i123_4_lut (.I0(fifo_state[2]), .I1(fifo_state[0]), .I2(fifo_state_timeout_counter[0]), 
            .I3(n4), .O(n94));   // src/timing_controller.v(77[11:21])
    defparam i123_4_lut.LUT_INIT = 16'heece;
    SB_LUT4 i3545_1_lut (.I0(buffer_switch_done), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5043));   // src/timing_controller.v(159[5] 228[12])
    defparam i3545_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR state_timeout_counter_i0_i17 (.Q(state_timeout_counter[17]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[17]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_LUT4 i13947_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n16071));   // src/timing_controller.v(159[5] 228[12])
    defparam i13947_2_lut.LUT_INIT = 16'h9999;
    SB_DFFESR state_timeout_counter_i0_i18 (.Q(state_timeout_counter[18]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[18]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i20 (.Q(state_timeout_counter[20]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[20]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i21 (.Q(state_timeout_counter[21]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[21]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i22 (.Q(state_timeout_counter[22]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[22]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i23 (.Q(state_timeout_counter[23]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[23]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i24 (.Q(state_timeout_counter[24]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[24]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_LUT4 sub_111_add_2_6_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n13716), .O(fifo_state_timeout_counter_5__N_125[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8320_2_lut (.I0(n2179[3]), .I1(n2283), .I2(GND_net), .I3(GND_net), 
            .O(n2284[3]));   // src/timing_controller.v(159[5] 228[12])
    defparam i8320_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mux_1150_i3_3_lut (.I0(n15917), .I1(state[1]), .I2(n2283), 
            .I3(GND_net), .O(n2284[2]));   // src/timing_controller.v(159[5] 228[12])
    defparam mux_1150_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFF invert_98_i2 (.Q(buffer_switch_done), .C(SLM_CLK_c), .D(n14533));   // src/timing_controller.v(159[5] 228[12])
    SB_LUT4 mux_1150_i2_3_lut (.I0(n15918), .I1(state[1]), .I2(n2283), 
            .I3(GND_net), .O(n2284[1]));   // src/timing_controller.v(159[5] 228[12])
    defparam mux_1150_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(VCC_net), .D(n14118));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFE state_timeout_counter_i0_i16 (.Q(state_timeout_counter[16]), .C(SLM_CLK_c), 
            .E(n4989), .D(n2356[16]));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i25 (.Q(state_timeout_counter[25]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[25]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_LUT4 i1_2_lut (.I0(fifo_state[1]), .I1(n14494), .I2(GND_net), .I3(GND_net), 
            .O(n14495));   // src/timing_controller.v(88[8] 150[4])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_DFFESR state_timeout_counter_i0_i26 (.Q(state_timeout_counter[26]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[26]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i27 (.Q(state_timeout_counter[27]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[27]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i28 (.Q(state_timeout_counter[28]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[28]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFE state_timeout_counter_i0_i15 (.Q(state_timeout_counter[15]), .C(SLM_CLK_c), 
            .E(n4989), .D(n2356[15]));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i29 (.Q(state_timeout_counter[29]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[29]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_LUT4 mux_1158_i5_4_lut (.I0(n15940), .I1(state[1]), .I2(n2355), 
            .I3(n2283), .O(n2356[4]));   // src/timing_controller.v(159[5] 228[12])
    defparam mux_1158_i5_4_lut.LUT_INIT = 16'hcfca;
    SB_DFFE state_timeout_counter_i0_i11 (.Q(state_timeout_counter[11]), .C(SLM_CLK_c), 
            .E(n4989), .D(n2356[11]));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFE state_timeout_counter_i0_i8 (.Q(state_timeout_counter[8]), .C(SLM_CLK_c), 
            .E(n4989), .D(n2356[8]));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i30 (.Q(state_timeout_counter[30]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[30]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i31 (.Q(state_timeout_counter[31]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[31]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR fifo_state_timeout_counter_i0_i4 (.Q(fifo_state_timeout_counter[4]), 
            .C(SLM_CLK_c), .E(n9126), .D(fifo_state_timeout_counter_5__N_125[4]), 
            .R(n9122));   // src/timing_controller.v(88[8] 150[4])
    SB_DFFE state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(SLM_CLK_c), 
            .E(n4989), .D(n2356[5]));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFE state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(SLM_CLK_c), 
            .E(n4989), .D(n2356[4]));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESS fifo_state_timeout_counter_i0_i5 (.Q(fifo_state_timeout_counter[5]), 
            .C(SLM_CLK_c), .E(n9126), .D(n14495), .S(n13147));   // src/timing_controller.v(88[8] 150[4])
    SB_LUT4 i1_4_lut (.I0(fifo_state[0]), .I1(n13147), .I2(fifo_state[1]), 
            .I3(n15), .O(n9122));
    defparam i1_4_lut.LUT_INIT = 16'hcdcc;
    SB_DFFESR state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(SLM_CLK_c), 
            .E(n4989), .D(n2284[1]), .R(n5453));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n4989), .D(n2284[2]), .R(n5453));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(SLM_CLK_c), 
            .E(n4989), .D(n2284[3]), .R(n5453));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n4989), .D(n628[6]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(SLM_CLK_c), 
            .E(n4989), .D(n628[7]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_LUT4 i1_2_lut_adj_137 (.I0(fifo_state[2]), .I1(n1224), .I2(GND_net), 
            .I3(GND_net), .O(n17));
    defparam i1_2_lut_adj_137.LUT_INIT = 16'heeee;
    SB_DFFESR state_timeout_counter_i0_i9 (.Q(state_timeout_counter[9]), .C(SLM_CLK_c), 
            .E(n4989), .D(n628[9]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_LUT4 i1_4_lut_adj_138 (.I0(fifo_state[0]), .I1(fifo_state[1]), .I2(n17), 
            .I3(n14544), .O(n9126));
    defparam i1_4_lut_adj_138.LUT_INIT = 16'hba32;
    SB_DFFESR state_timeout_counter_i0_i10 (.Q(state_timeout_counter[10]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[10]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i12 (.Q(state_timeout_counter[12]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[12]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i13 (.Q(state_timeout_counter[13]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[13]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFESR state_timeout_counter_i0_i14 (.Q(state_timeout_counter[14]), 
            .C(SLM_CLK_c), .E(n4989), .D(n628[14]), .R(n5446));   // src/timing_controller.v(153[8] 229[4])
    SB_LUT4 mux_1150_i9_3_lut (.I0(n15916), .I1(state[1]), .I2(n2283), 
            .I3(GND_net), .O(n2284[8]));   // src/timing_controller.v(159[5] 228[12])
    defparam mux_1150_i9_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFESR fifo_state_timeout_counter_i0_i0 (.Q(fifo_state_timeout_counter[0]), 
            .C(SLM_CLK_c), .E(n9126), .D(fifo_state_timeout_counter_5__N_125[0]), 
            .R(n9122));   // src/timing_controller.v(88[8] 150[4])
    SB_DFFESR fifo_state_timeout_counter_i0_i1 (.Q(fifo_state_timeout_counter[1]), 
            .C(SLM_CLK_c), .E(n9126), .D(fifo_state_timeout_counter_5__N_125[1]), 
            .R(n9122));   // src/timing_controller.v(88[8] 150[4])
    SB_DFFESR fifo_state_timeout_counter_i0_i2 (.Q(fifo_state_timeout_counter[2]), 
            .C(SLM_CLK_c), .E(n9126), .D(fifo_state_timeout_counter_5__N_125[2]), 
            .R(n9122));   // src/timing_controller.v(88[8] 150[4])
    SB_LUT4 mux_1150_i12_3_lut (.I0(n15915), .I1(state[1]), .I2(n2283), 
            .I3(GND_net), .O(n2284[11]));   // src/timing_controller.v(159[5] 228[12])
    defparam mux_1150_i12_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFESR fifo_state_timeout_counter_i0_i3 (.Q(fifo_state_timeout_counter[3]), 
            .C(SLM_CLK_c), .E(n9126), .D(n14511), .R(n13147));   // src/timing_controller.v(88[8] 150[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(state[0]), .I1(state[2]), .I2(n63), .I3(GND_net), 
            .O(n14557));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_1150_i16_3_lut (.I0(n15914), .I1(state[1]), .I2(n2283), 
            .I3(GND_net), .O(n2284[15]));   // src/timing_controller.v(159[5] 228[12])
    defparam mux_1150_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n5077), .D(state_3__N_83[2]));   // src/timing_controller.v(153[8] 229[4])
    SB_CARRY sub_111_add_2_6 (.CI(n13716), .I0(fifo_state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n13717));
    SB_LUT4 sub_111_add_2_5_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n13715), .O(fifo_state_timeout_counter_5__N_125[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_23 (.CI(n13687), .I0(state_timeout_counter[21]), 
            .I1(VCC_net), .CO(n13688));
    SB_CARRY sub_111_add_2_5 (.CI(n13715), .I0(fifo_state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n13716));
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n5077), .D(state_3__N_83[1]));   // src/timing_controller.v(153[8] 229[4])
    SB_DFFE fifo_state_i2 (.Q(fifo_state[2]), .C(SLM_CLK_c), .E(n14130), 
            .D(fifo_state_2__N_80[2]));   // src/timing_controller.v(88[8] 150[4])
    SB_DFFSR line_of_data_available_91 (.Q(line_of_data_available), .C(SLM_CLK_c), 
            .D(n2), .R(n8104));   // src/timing_controller.v(88[8] 150[4])
    SB_LUT4 sub_111_add_2_4_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n13714), .O(fifo_state_timeout_counter_5__N_125[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_111_add_2_4 (.CI(n13714), .I0(fifo_state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n13715));
    SB_LUT4 sub_111_add_2_3_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n13713), .O(fifo_state_timeout_counter_5__N_125[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_111_add_2_3 (.CI(n13713), .I0(fifo_state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n13714));
    SB_LUT4 sub_111_add_2_2_lut (.I0(GND_net), .I1(fifo_state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(fifo_state_timeout_counter_5__N_125[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_69_add_2_22_lut (.I0(GND_net), .I1(state_timeout_counter[20]), 
            .I2(VCC_net), .I3(n13686), .O(n628[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_111_add_2_2 (.CI(VCC_net), .I0(fifo_state_timeout_counter[0]), 
            .I1(GND_net), .CO(n13713));
    SB_CARRY sub_69_add_2_22 (.CI(n13686), .I0(state_timeout_counter[20]), 
            .I1(VCC_net), .CO(n13687));
    SB_DFFE fifo_state_i1 (.Q(fifo_state[1]), .C(SLM_CLK_c), .E(n14700), 
            .D(fifo_state_2__N_80[1]));   // src/timing_controller.v(88[8] 150[4])
    SB_DFFE state_timeout_counter_i0_i19 (.Q(state_timeout_counter[19]), .C(SLM_CLK_c), 
            .E(n4989), .D(n2356[19]));   // src/timing_controller.v(153[8] 229[4])
    SB_LUT4 sub_69_add_2_21_lut (.I0(n2178), .I1(state_timeout_counter[19]), 
            .I2(VCC_net), .I3(n13685), .O(n15912)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_21 (.CI(n13685), .I0(state_timeout_counter[19]), 
            .I1(VCC_net), .CO(n13686));
    SB_LUT4 mux_1150_i17_3_lut (.I0(n15913), .I1(state[1]), .I2(n2283), 
            .I3(GND_net), .O(n2284[16]));   // src/timing_controller.v(159[5] 228[12])
    defparam mux_1150_i17_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 sub_69_add_2_20_lut (.I0(GND_net), .I1(state_timeout_counter[18]), 
            .I2(VCC_net), .I3(n13684), .O(n628[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_139 (.I0(n2178), .I1(n2283), .I2(GND_net), .I3(GND_net), 
            .O(n14538));   // src/timing_controller.v(159[5] 228[12])
    defparam i1_2_lut_adj_139.LUT_INIT = 16'h2222;
    SB_CARRY sub_69_add_2_20 (.CI(n13684), .I0(state_timeout_counter[18]), 
            .I1(VCC_net), .CO(n13685));
    SB_LUT4 sub_69_add_2_19_lut (.I0(GND_net), .I1(state_timeout_counter[17]), 
            .I2(VCC_net), .I3(n13683), .O(n628[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_19 (.CI(n13683), .I0(state_timeout_counter[17]), 
            .I1(VCC_net), .CO(n13684));
    SB_LUT4 sub_69_add_2_18_lut (.I0(n2178), .I1(state_timeout_counter[16]), 
            .I2(VCC_net), .I3(n13682), .O(n15913)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_18 (.CI(n13682), .I0(state_timeout_counter[16]), 
            .I1(VCC_net), .CO(n13683));
    SB_LUT4 sub_69_add_2_17_lut (.I0(n2178), .I1(state_timeout_counter[15]), 
            .I2(VCC_net), .I3(n13681), .O(n15914)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_17 (.CI(n13681), .I0(state_timeout_counter[15]), 
            .I1(VCC_net), .CO(n13682));
    SB_DFF invert_98_i4 (.Q(INVERT_c_4), .C(SLM_CLK_c), .D(n1114[4]));   // src/timing_controller.v(159[5] 228[12])
    SB_LUT4 sub_69_add_2_16_lut (.I0(GND_net), .I1(state_timeout_counter[14]), 
            .I2(VCC_net), .I3(n13680), .O(n628[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_16 (.CI(n13680), .I0(state_timeout_counter[14]), 
            .I1(VCC_net), .CO(n13681));
    SB_LUT4 sub_69_add_2_15_lut (.I0(GND_net), .I1(state_timeout_counter[13]), 
            .I2(VCC_net), .I3(n13679), .O(n628[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_15 (.CI(n13679), .I0(state_timeout_counter[13]), 
            .I1(VCC_net), .CO(n13680));
    SB_LUT4 sub_69_add_2_14_lut (.I0(GND_net), .I1(state_timeout_counter[12]), 
            .I2(VCC_net), .I3(n13678), .O(n628[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_14 (.CI(n13678), .I0(state_timeout_counter[12]), 
            .I1(VCC_net), .CO(n13679));
    SB_LUT4 sub_69_add_2_13_lut (.I0(n2178), .I1(state_timeout_counter[11]), 
            .I2(VCC_net), .I3(n13677), .O(n15915)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_13 (.CI(n13677), .I0(state_timeout_counter[11]), 
            .I1(VCC_net), .CO(n13678));
    SB_LUT4 sub_69_add_2_12_lut (.I0(GND_net), .I1(state_timeout_counter[10]), 
            .I2(VCC_net), .I3(n13676), .O(n628[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_12 (.CI(n13676), .I0(state_timeout_counter[10]), 
            .I1(VCC_net), .CO(n13677));
    SB_LUT4 sub_69_add_2_11_lut (.I0(GND_net), .I1(state_timeout_counter[9]), 
            .I2(VCC_net), .I3(n13675), .O(n628[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_11 (.CI(n13675), .I0(state_timeout_counter[9]), 
            .I1(VCC_net), .CO(n13676));
    SB_LUT4 sub_69_add_2_10_lut (.I0(n2178), .I1(state_timeout_counter[8]), 
            .I2(VCC_net), .I3(n13674), .O(n15916)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_10 (.CI(n13674), .I0(state_timeout_counter[8]), 
            .I1(VCC_net), .CO(n13675));
    SB_LUT4 sub_69_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n13673), .O(n628[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_9 (.CI(n13673), .I0(state_timeout_counter[7]), 
            .I1(VCC_net), .CO(n13674));
    SB_LUT4 sub_69_add_2_33_lut (.I0(GND_net), .I1(state_timeout_counter[31]), 
            .I2(VCC_net), .I3(n13697), .O(n628[31])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_69_add_2_32_lut (.I0(GND_net), .I1(state_timeout_counter[30]), 
            .I2(VCC_net), .I3(n13696), .O(n628[30])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_32 (.CI(n13696), .I0(state_timeout_counter[30]), 
            .I1(VCC_net), .CO(n13697));
    SB_LUT4 sub_69_add_2_31_lut (.I0(GND_net), .I1(state_timeout_counter[29]), 
            .I2(VCC_net), .I3(n13695), .O(n628[29])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14026_2_lut (.I0(n7), .I1(n8), .I2(GND_net), .I3(GND_net), 
            .O(\aempty_flag_impl.ae_flag_nxt_w ));
    defparam i14026_2_lut.LUT_INIT = 16'h1111;
    SB_CARRY sub_69_add_2_31 (.CI(n13695), .I0(state_timeout_counter[29]), 
            .I1(VCC_net), .CO(n13696));
    SB_LUT4 sub_69_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n13672), .O(n628[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_69_add_2_30_lut (.I0(GND_net), .I1(state_timeout_counter[28]), 
            .I2(VCC_net), .I3(n13694), .O(n628[28])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_8 (.CI(n13672), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n13673));
    SB_LUT4 sub_69_add_2_7_lut (.I0(n14538), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n13671), .O(n15941)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_30 (.CI(n13694), .I0(state_timeout_counter[28]), 
            .I1(VCC_net), .CO(n13695));
    SB_LUT4 sub_69_add_2_29_lut (.I0(GND_net), .I1(state_timeout_counter[27]), 
            .I2(VCC_net), .I3(n13693), .O(n628[27])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_7 (.CI(n13671), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n13672));
    SB_CARRY sub_69_add_2_29 (.CI(n13693), .I0(state_timeout_counter[27]), 
            .I1(VCC_net), .CO(n13694));
    SB_LUT4 sub_69_add_2_28_lut (.I0(GND_net), .I1(state_timeout_counter[26]), 
            .I2(VCC_net), .I3(n13692), .O(n628[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_28 (.CI(n13692), .I0(state_timeout_counter[26]), 
            .I1(VCC_net), .CO(n13693));
    SB_LUT4 sub_69_add_2_6_lut (.I0(n2178), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n13670), .O(n15940)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_69_add_2_27_lut (.I0(GND_net), .I1(state_timeout_counter[25]), 
            .I2(VCC_net), .I3(n13691), .O(n628[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_6 (.CI(n13670), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n13671));
    SB_LUT4 sub_69_add_2_5_lut (.I0(n2178), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n13669), .O(n2179[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_27 (.CI(n13691), .I0(state_timeout_counter[25]), 
            .I1(VCC_net), .CO(n13692));
    SB_LUT4 sub_69_add_2_26_lut (.I0(GND_net), .I1(state_timeout_counter[24]), 
            .I2(VCC_net), .I3(n13690), .O(n628[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_26 (.CI(n13690), .I0(state_timeout_counter[24]), 
            .I1(VCC_net), .CO(n13691));
    SB_LUT4 i13922_4_lut (.I0(n13173), .I1(fifo_state[2]), .I2(get_next_word), 
            .I3(fifo_state[1]), .O(n15906));
    defparam i13922_4_lut.LUT_INIT = 16'h3011;
    SB_LUT4 i34_4_lut (.I0(n16), .I1(n15906), .I2(fifo_state[0]), .I3(fifo_state[1]), 
            .O(dc32_fifo_read_enable_N_359));
    defparam i34_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 state_3__I_0_103_Mux_0_i7_4_lut (.I0(state[1]), .I1(n63), .I2(state[2]), 
            .I3(state[0]), .O(n7_adj_1410));   // src/timing_controller.v(159[5] 228[12])
    defparam state_3__I_0_103_Mux_0_i7_4_lut.LUT_INIT = 16'hc535;
    SB_LUT4 state_3__I_0_103_Mux_0_i15_4_lut (.I0(n7_adj_1410), .I1(n10029), 
            .I2(state[3]), .I3(state[0]), .O(state_3__N_83[0]));   // src/timing_controller.v(159[5] 228[12])
    defparam state_3__I_0_103_Mux_0_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i37_3_lut (.I0(dc32_fifo_full), .I1(get_next_word), .I2(fifo_state[0]), 
            .I3(GND_net), .O(n18));
    defparam i37_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12577_4_lut (.I0(fifo_state[2]), .I1(n14643), .I2(n18), .I3(fifo_state[1]), 
            .O(n14700));
    defparam i12577_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_4_lut_adj_140 (.I0(fifo_state[2]), .I1(fifo_state[0]), .I2(fifo_state[1]), 
            .I3(n13173), .O(fifo_state_2__N_80[0]));
    defparam i1_4_lut_adj_140.LUT_INIT = 16'h9399;
    SB_LUT4 i1_2_lut_adj_141 (.I0(fifo_state[2]), .I1(get_next_word), .I2(GND_net), 
            .I3(GND_net), .O(n14544));
    defparam i1_2_lut_adj_141.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_142 (.I0(fifo_state[1]), .I1(n13147), .I2(fifo_state[2]), 
            .I3(n14682), .O(sc32_fifo_read_enable_N_367));
    defparam i1_4_lut_adj_142.LUT_INIT = 16'hccdc;
    SB_LUT4 i1208_2_lut_3_lut (.I0(state[0]), .I1(n63), .I2(state[1]), 
            .I3(GND_net), .O(n2437));   // src/timing_controller.v(153[8] 229[4])
    defparam i1208_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2_2_lut (.I0(fifo_state_timeout_counter[1]), .I1(fifo_state_timeout_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // src/timing_controller.v(79[11:37])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mux_1158_i1_3_lut_4_lut (.I0(state[1]), .I1(n14546), .I2(n2355), 
            .I3(n2284[0]), .O(n2356[0]));
    defparam mux_1158_i1_3_lut_4_lut.LUT_INIT = 16'h1f10;
    SB_LUT4 mux_1158_i6_3_lut_4_lut (.I0(state[1]), .I1(n14546), .I2(n2355), 
            .I3(n15941), .O(n2356[5]));
    defparam mux_1158_i6_3_lut_4_lut.LUT_INIT = 16'hefe0;
    SB_LUT4 i1_4_lut_adj_143 (.I0(fifo_state_timeout_counter[5]), .I1(fifo_state_timeout_counter[3]), 
            .I2(n6), .I3(fifo_state_timeout_counter[4]), .O(n4));   // src/timing_controller.v(79[11:37])
    defparam i1_4_lut_adj_143.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_144 (.I0(fifo_state_timeout_counter[0]), .I1(n4), 
            .I2(GND_net), .I3(GND_net), .O(n13173));
    defparam i1_2_lut_adj_144.LUT_INIT = 16'h2222;
    SB_LUT4 i13911_2_lut (.I0(get_next_word), .I1(fifo_state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15958));
    defparam i13911_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i20_4_lut (.I0(n11), .I1(n15958), .I2(fifo_state[0]), .I3(fifo_state[2]), 
            .O(sc32_fifo_write_enable_N_366));
    defparam i20_4_lut.LUT_INIT = 16'h05c0;
    SB_LUT4 sub_69_add_2_25_lut (.I0(GND_net), .I1(state_timeout_counter[23]), 
            .I2(VCC_net), .I3(n13689), .O(n628[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_25 (.CI(n13689), .I0(state_timeout_counter[23]), 
            .I1(VCC_net), .CO(n13690));
    SB_DFF invert_98_i0 (.Q(reset_all), .C(SLM_CLK_c), .D(n14532));   // src/timing_controller.v(159[5] 228[12])
    SB_CARRY sub_69_add_2_5 (.CI(n13669), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n13670));
    SB_LUT4 sub_69_add_2_4_lut (.I0(n9752), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n13668), .O(n15917)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_4_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_69_add_2_4 (.CI(n13668), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n13669));
    SB_LUT4 sub_69_add_2_24_lut (.I0(GND_net), .I1(state_timeout_counter[22]), 
            .I2(VCC_net), .I3(n13688), .O(n628[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_69_add_2_24 (.CI(n13688), .I0(state_timeout_counter[22]), 
            .I1(VCC_net), .CO(n13689));
    SB_LUT4 sub_69_add_2_23_lut (.I0(GND_net), .I1(state_timeout_counter[21]), 
            .I2(VCC_net), .I3(n13687), .O(n628[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_69_add_2_3_lut (.I0(n2178), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n13667), .O(n15918)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_69_add_2_3 (.CI(n13667), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n13668));
    SB_LUT4 i8544_2_lut_3_lut (.I0(state[1]), .I1(state[2]), .I2(n63), 
            .I3(GND_net), .O(n10029));
    defparam i8544_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i8573_2_lut_3_lut (.I0(state[1]), .I1(state[2]), .I2(state[0]), 
            .I3(GND_net), .O(n10059));
    defparam i8573_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF invert_98_i1 (.Q(reset_per_frame), .C(SLM_CLK_c), .D(n14542));   // src/timing_controller.v(159[5] 228[12])
    SB_LUT4 sub_69_add_2_2_lut (.I0(n9752), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n15900)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_69_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i25_1_lut (.I0(dc32_fifo_read_enable), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // src/top.v(483[26:47])
    defparam i25_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR invert_98_i3 (.Q(UPDATE_c_3), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n16071), .R(n5));   // src/timing_controller.v(159[5] 228[12])
    SB_CARRY sub_69_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n13667));
    SB_LUT4 i12570_2_lut_3_lut (.I0(state[0]), .I1(state[2]), .I2(state[1]), 
            .I3(GND_net), .O(n14692));
    defparam i12570_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i14000_2_lut (.I0(state[3]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // src/timing_controller.v(153[8] 229[4])
    defparam i14000_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1219_4_lut (.I0(state[3]), .I1(n2437), .I2(n10051), .I3(state[2]), 
            .O(n2355));   // src/timing_controller.v(153[8] 229[4])
    defparam i1219_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 state_3__I_0_103_Mux_1_i15_4_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[3]), .I3(n14557), .O(state_3__N_83[1]));   // src/timing_controller.v(159[5] 228[12])
    defparam state_3__I_0_103_Mux_1_i15_4_lut_4_lut.LUT_INIT = 16'hc6f6;
    SB_LUT4 i1_3_lut (.I0(state[2]), .I1(state[1]), .I2(state[0]), .I3(GND_net), 
            .O(n4843));   // src/timing_controller.v(159[5] 228[12])
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_2_lut (.I0(state_timeout_counter[9]), .I1(state_timeout_counter[12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // src/timing_controller.v(181[17:45])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut_adj_145 (.I0(state_timeout_counter[17]), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[24]), .I3(state_timeout_counter[4]), 
            .O(n52));   // src/timing_controller.v(181[17:45])
    defparam i20_4_lut_adj_145.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_111_add_2_7_lut (.I0(n94), .I1(fifo_state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n13717), .O(n14494)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_111_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i24_4_lut (.I0(state_timeout_counter[29]), .I1(state_timeout_counter[3]), 
            .I2(state_timeout_counter[13]), .I3(state_timeout_counter[31]), 
            .O(n56));   // src/timing_controller.v(181[17:45])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(state_timeout_counter[19]), .I1(state_timeout_counter[5]), 
            .I2(state_timeout_counter[22]), .I3(state_timeout_counter[6]), 
            .O(n54));   // src/timing_controller.v(181[17:45])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(state_timeout_counter[10]), .I1(state_timeout_counter[15]), 
            .I2(state_timeout_counter[20]), .I3(state_timeout_counter[23]), 
            .O(n55));   // src/timing_controller.v(181[17:45])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(state_timeout_counter[27]), .I1(state_timeout_counter[7]), 
            .I2(state_timeout_counter[30]), .I3(state_timeout_counter[14]), 
            .O(n53));   // src/timing_controller.v(181[17:45])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(state_timeout_counter[8]), .I1(state_timeout_counter[11]), 
            .I2(state_timeout_counter[16]), .I3(state_timeout_counter[21]), 
            .O(n50));   // src/timing_controller.v(181[17:45])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(state_timeout_counter[25]), .I1(n52), .I2(n38), 
            .I3(state_timeout_counter[26]), .O(n58));   // src/timing_controller.v(181[17:45])
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30_4_lut (.I0(n53), .I1(n55), .I2(n54), .I3(n56), .O(n62));   // src/timing_controller.v(181[17:45])
    defparam i30_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(state_timeout_counter[0]), .I1(state_timeout_counter[18]), 
            .I2(state_timeout_counter[28]), .I3(state_timeout_counter[2]), 
            .O(n49));   // src/timing_controller.v(181[17:45])
    defparam i17_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i31_4_lut (.I0(n49), .I1(n62), .I2(n58), .I3(n50), .O(n63));   // src/timing_controller.v(181[17:45])
    defparam i31_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14030_2_lut (.I0(state[3]), .I1(n4843), .I2(GND_net), .I3(GND_net), 
            .O(n4989));
    defparam i14030_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 mux_1150_i1_3_lut (.I0(n15900), .I1(state[1]), .I2(n2283), 
            .I3(GND_net), .O(n2284[0]));   // src/timing_controller.v(159[5] 228[12])
    defparam mux_1150_i1_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1150_i20_3_lut (.I0(n15912), .I1(state[1]), .I2(n2283), 
            .I3(GND_net), .O(n2284[19]));   // src/timing_controller.v(159[5] 228[12])
    defparam mux_1150_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_1158_i9_3_lut_4_lut (.I0(state[1]), .I1(n14546), .I2(n2355), 
            .I3(n2284[8]), .O(n2356[8]));   // src/timing_controller.v(153[8] 229[4])
    defparam mux_1158_i9_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_1158_i17_3_lut_4_lut (.I0(state[1]), .I1(n14546), .I2(n2355), 
            .I3(n2284[16]), .O(n2356[16]));   // src/timing_controller.v(153[8] 229[4])
    defparam mux_1158_i17_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_1158_i16_3_lut_4_lut (.I0(state[1]), .I1(n14546), .I2(n2355), 
            .I3(n2284[15]), .O(n2356[15]));   // src/timing_controller.v(153[8] 229[4])
    defparam mux_1158_i16_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i1_2_lut_3_lut_adj_146 (.I0(line_of_data_available), .I1(n910), 
            .I2(n989), .I3(GND_net), .O(n1028));   // src/timing_controller.v(88[8] 150[4])
    defparam i1_2_lut_3_lut_adj_146.LUT_INIT = 16'h2020;
    SB_LUT4 mux_1158_i12_3_lut_4_lut (.I0(state[1]), .I1(n14546), .I2(n2355), 
            .I3(n2284[11]), .O(n2356[11]));   // src/timing_controller.v(153[8] 229[4])
    defparam mux_1158_i12_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_372_Mux_4_i15_4_lut_4_lut (.I0(state[1]), .I1(state[0]), 
            .I2(state[2]), .I3(state[3]), .O(n1114[4]));   // src/timing_controller.v(159[5] 228[12])
    defparam mux_372_Mux_4_i15_4_lut_4_lut.LUT_INIT = 16'h01a0;
    SB_LUT4 mux_1158_i20_3_lut_4_lut (.I0(state[1]), .I1(n14546), .I2(n2355), 
            .I3(n2284[19]), .O(n2356[19]));   // src/timing_controller.v(153[8] 229[4])
    defparam mux_1158_i20_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i1_2_lut_3_lut_adj_147 (.I0(fifo_state[1]), .I1(fifo_state_timeout_counter[0]), 
            .I2(n4), .I3(GND_net), .O(n11));
    defparam i1_2_lut_3_lut_adj_147.LUT_INIT = 16'haeae;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[0]), .I1(n63), .I2(state[3]), 
            .I3(state[2]), .O(n14546));   // src/timing_controller.v(153[8] 229[4])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i12560_2_lut_3_lut (.I0(fifo_state[0]), .I1(fifo_state_timeout_counter[0]), 
            .I2(n4), .I3(GND_net), .O(n14682));
    defparam i12560_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_3_lut_4_lut (.I0(fifo_state[1]), .I1(fifo_state[0]), .I2(fifo_state[2]), 
            .I3(get_next_word), .O(n13147));   // src/timing_controller.v(88[8] 150[4])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i50_3_lut_4_lut (.I0(n1224), .I1(fifo_state_timeout_counter[0]), 
            .I2(n4), .I3(fifo_state[0]), .O(n14643));
    defparam i50_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i36_3_lut_4_lut (.I0(n1224), .I1(fifo_state_timeout_counter[0]), 
            .I2(n4), .I3(fifo_state[2]), .O(n16));
    defparam i36_3_lut_4_lut.LUT_INIT = 16'hf3aa;
    SB_LUT4 fifo_state_2__I_0_106_Mux_1_i7_3_lut (.I0(fifo_state[0]), .I1(fifo_state[1]), 
            .I2(fifo_state[2]), .I3(GND_net), .O(fifo_state_2__N_80[1]));   // src/timing_controller.v(93[5] 149[12])
    defparam fifo_state_2__I_0_106_Mux_1_i7_3_lut.LUT_INIT = 16'hc6c6;
    SB_LUT4 i13969_3_lut_4_lut (.I0(state[3]), .I1(n4843), .I2(n2355), 
            .I3(n14538), .O(n5446));
    defparam i13969_3_lut_4_lut.LUT_INIT = 16'h7077;
    SB_LUT4 i26_3_lut_4_lut (.I0(n1224), .I1(fifo_state_timeout_counter[0]), 
            .I2(n4), .I3(fifo_state[2]), .O(n15));   // src/timing_controller.v(77[11:21])
    defparam i26_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i3954_2_lut_3_lut (.I0(state[3]), .I1(n4843), .I2(n2355), 
            .I3(GND_net), .O(n5453));   // src/timing_controller.v(153[8] 229[4])
    defparam i3954_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i1_3_lut_3_lut (.I0(buffer_switch_done), .I1(buffer_switch_done_latched), 
            .I2(n14482), .I3(GND_net), .O(n5529));   // src/timing_controller.v(159[5] 228[12])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_2_lut (.I0(buffer_switch_done), .I1(bluejay_data_out_31__N_920), 
            .I2(GND_net), .I3(GND_net), .O(n5528));   // src/timing_controller.v(159[5] 228[12])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_148 (.I0(fifo_state[2]), .I1(fifo_state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n8104));   // src/timing_controller.v(88[8] 150[4])
    defparam i1_2_lut_adj_148.LUT_INIT = 16'hbbbb;
    SB_LUT4 i8334_2_lut (.I0(dc32_fifo_full), .I1(fifo_state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // src/timing_controller.v(93[5] 149[12])
    defparam i8334_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13925_4_lut (.I0(n1224), .I1(n13173), .I2(fifo_state[0]), 
            .I3(fifo_state[2]), .O(n15922));
    defparam i13925_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36_4_lut (.I0(n15922), .I1(n18), .I2(fifo_state[1]), .I3(fifo_state[2]), 
            .O(n14130));
    defparam i36_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_3_lut_3_lut_adj_149 (.I0(buffer_switch_done), .I1(bluejay_data_out_31__N_920), 
            .I2(bluejay_data_out_31__N_919), .I3(GND_net), .O(n5431));   // src/timing_controller.v(159[5] 228[12])
    defparam i1_3_lut_3_lut_adj_149.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_3_lut_adj_150 (.I0(fifo_state[2]), .I1(fifo_state_timeout_counter[0]), 
            .I2(n4), .I3(GND_net), .O(n7_c));
    defparam i1_2_lut_3_lut_adj_150.LUT_INIT = 16'ha2a2;
    SB_LUT4 i12_3_lut (.I0(fifo_state[1]), .I1(fifo_state[2]), .I2(fifo_state[0]), 
            .I3(GND_net), .O(fifo_state_2__N_80[2]));   // src/timing_controller.v(77[11:21])
    defparam i12_3_lut.LUT_INIT = 16'h2c2c;
    
endmodule
//
// Verilog Description of module bluejay_data
//

module bluejay_data (DEBUG_6_c, SLM_CLK_c, buffer_switch_done, buffer_switch_done_latched, 
            GND_net, n910, line_of_data_available, n989, bluejay_data_out_31__N_921, 
            bluejay_data_out_31__N_920, bluejay_data_out_31__N_922, n5043, 
            n14482, n6982, DEBUG_8_c, n5431, VCC_net, DATA10_c_10, 
            n5414, DATA9_c_9, n5413, DATA11_c_11, n5412, DATA12_c_12, 
            n5411, n14298, n1028, bluejay_data_out_31__N_919, SYNC_c, 
            DATA13_c_13, n5410, DATA14_c_14, n5409, DATA8_c_8, n5408, 
            DATA15_c_15, n5407, DATA16_c_16, n5406, DATA7_c_7, n5405, 
            DATA17_c_17, n5404, DATA18_c_18, n5403, DATA6_c_6, n5402, 
            DATA19_c_19, n5401, DATA20_c_20, n5400, DATA5_c_5, n5399, 
            DATA21_c_21, n5398, DATA22_c_22, n5397, DATA4_c_4, n5396, 
            DATA23_c_23, n5395, DATA24_c_24, n5394, n5529, n5528, 
            DATA3_c_3, n5393, get_next_word, DATA25_c_25, n5392, DATA26_c_26, 
            n5391, DATA2_c_2, n5390, DATA27_c_27, n5389, DATA28_c_28, 
            n5388, DATA1_c_1, n5387, DATA29_c_29, n5386, DATA30_c_30, 
            n5385, DATA31_c_31, n5384, sc32_fifo_almost_empty) /* synthesis syn_module_defined=1 */ ;
    output DEBUG_6_c;
    input SLM_CLK_c;
    input buffer_switch_done;
    input buffer_switch_done_latched;
    input GND_net;
    output n910;
    input line_of_data_available;
    output n989;
    output bluejay_data_out_31__N_921;
    output bluejay_data_out_31__N_920;
    output bluejay_data_out_31__N_922;
    input n5043;
    output n14482;
    input n6982;
    output DEBUG_8_c;
    input n5431;
    input VCC_net;
    output DATA10_c_10;
    input n5414;
    output DATA9_c_9;
    input n5413;
    output DATA11_c_11;
    input n5412;
    output DATA12_c_12;
    input n5411;
    input n14298;
    input n1028;
    output bluejay_data_out_31__N_919;
    output SYNC_c;
    output DATA13_c_13;
    input n5410;
    output DATA14_c_14;
    input n5409;
    output DATA8_c_8;
    input n5408;
    output DATA15_c_15;
    input n5407;
    output DATA16_c_16;
    input n5406;
    output DATA7_c_7;
    input n5405;
    output DATA17_c_17;
    input n5404;
    output DATA18_c_18;
    input n5403;
    output DATA6_c_6;
    input n5402;
    output DATA19_c_19;
    input n5401;
    output DATA20_c_20;
    input n5400;
    output DATA5_c_5;
    input n5399;
    output DATA21_c_21;
    input n5398;
    output DATA22_c_22;
    input n5397;
    output DATA4_c_4;
    input n5396;
    output DATA23_c_23;
    input n5395;
    output DATA24_c_24;
    input n5394;
    input n5529;
    input n5528;
    output DATA3_c_3;
    input n5393;
    output get_next_word;
    output DATA25_c_25;
    input n5392;
    output DATA26_c_26;
    input n5391;
    output DATA2_c_2;
    input n5390;
    output DATA27_c_27;
    input n5389;
    output DATA28_c_28;
    input n5388;
    output DATA1_c_1;
    input n5387;
    output DATA29_c_29;
    input n5386;
    output DATA30_c_30;
    input n5385;
    output DATA31_c_31;
    input n5384;
    input sc32_fifo_almost_empty;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire valid_N_925;
    wire [10:0]v_counter_10__N_900;
    
    wire n5132;
    wire [10:0]v_counter;   // src/bluejay_data.v(51[12:21])
    wire [15:0]n974;
    
    wire n45, n6, n14569, n4, n14475;
    wire [7:0]state_timeout_counter;   // src/bluejay_data.v(52[11:32])
    
    wire n6_adj_1401, n14472, n13, n1244, n1528;
    wire [8:0]n74;
    
    wire n5, n14551, n8, n14196, n5625, n5_adj_1402, n8_adj_1403, 
        n14186, n59, n6_adj_1404, n5_adj_1405, n5525, n9, n13811, 
        n5526, n4_adj_1406, n14214, n3, n5527, n14122, n6_adj_1407, 
        n14481, n14050, n3_adj_1408, n5530, n14026, n13652, n13649, 
        n14552, n13651, n13650, n13661, n13648, n13660, n14489, 
        n3546, n3548, n1037, n3550, n1041, n3552, n13647, n13659, 
        n13658, n13645, n13657, n13656, n13646, n13655, n13654, 
        n13653;
    wire [3:0]n99;
    
    wire n102, n13836, n106, n14627, n13985, n2;
    
    SB_DFFN valid_66 (.Q(DEBUG_6_c), .C(SLM_CLK_c), .D(valid_N_925));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFESS v_counter_i10 (.Q(v_counter[10]), .C(SLM_CLK_c), .E(n5132), 
            .D(v_counter_10__N_900[10]), .S(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i9 (.Q(v_counter[9]), .C(SLM_CLK_c), .E(n5132), 
            .D(v_counter_10__N_900[9]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS v_counter_i8 (.Q(v_counter[8]), .C(SLM_CLK_c), .E(n5132), 
            .D(v_counter_10__N_900[8]), .S(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i7 (.Q(v_counter[7]), .C(SLM_CLK_c), .E(n5132), 
            .D(v_counter_10__N_900[7]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i6 (.Q(v_counter[6]), .C(SLM_CLK_c), .E(n5132), 
            .D(v_counter_10__N_900[6]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i5 (.Q(v_counter[5]), .C(SLM_CLK_c), .E(n5132), 
            .D(v_counter_10__N_900[5]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i4 (.Q(v_counter[4]), .C(SLM_CLK_c), .E(n5132), 
            .D(v_counter_10__N_900[4]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i3 (.Q(v_counter[3]), .C(SLM_CLK_c), .E(n5132), 
            .D(v_counter_10__N_900[3]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_LUT4 i1_2_lut (.I0(buffer_switch_done_latched), .I1(n974[2]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_103 (.I0(v_counter[6]), .I1(v_counter[8]), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // src/bluejay_data.v(56[8] 131[4])
    defparam i1_2_lut_adj_103.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(v_counter[3]), .I1(v_counter[7]), .I2(v_counter[5]), 
            .I3(n6), .O(n14569));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(v_counter[4]), .I1(v_counter[0]), .I2(v_counter[2]), 
            .I3(v_counter[1]), .O(n4));
    defparam i1_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i2_3_lut (.I0(v_counter[9]), .I1(n4), .I2(v_counter[10]), 
            .I3(GND_net), .O(n14475));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_104 (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_1401));   // src/bluejay_data.v(107[21:49])
    defparam i1_2_lut_adj_104.LUT_INIT = 16'heeee;
    SB_DFFESR v_counter_i2 (.Q(v_counter[2]), .C(SLM_CLK_c), .E(n5132), 
            .D(v_counter_10__N_900[2]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i1 (.Q(v_counter[1]), .C(SLM_CLK_c), .E(n5132), 
            .D(v_counter_10__N_900[1]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_LUT4 i4_4_lut_adj_105 (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[2]), 
            .I2(state_timeout_counter[4]), .I3(n6_adj_1401), .O(n14472));   // src/bluejay_data.v(107[21:49])
    defparam i4_4_lut_adj_105.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_106 (.I0(state_timeout_counter[6]), .I1(state_timeout_counter[7]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // src/bluejay_data.v(56[8] 131[4])
    defparam i1_2_lut_adj_106.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_107 (.I0(n910), .I1(line_of_data_available), .I2(GND_net), 
            .I3(GND_net), .O(n1244));
    defparam i1_2_lut_adj_107.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_108 (.I0(n974[4]), .I1(n989), .I2(bluejay_data_out_31__N_921), 
            .I3(GND_net), .O(n1528));   // src/bluejay_data.v(43[15:31])
    defparam i2_3_lut_adj_108.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut (.I0(n74[0]), .I1(n5), .I2(n14551), .I3(n8), .O(n14196));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i1_2_lut_adj_109 (.I0(bluejay_data_out_31__N_921), .I1(bluejay_data_out_31__N_920), 
            .I2(GND_net), .I3(GND_net), .O(n5625));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_109.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_110 (.I0(n74[1]), .I1(n5_adj_1402), .I2(n14551), 
            .I3(n8_adj_1403), .O(n14186));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_4_lut_adj_110.LUT_INIT = 16'hffec;
    SB_LUT4 i2_4_lut_adj_111 (.I0(state_timeout_counter[2]), .I1(n59), .I2(n974[2]), 
            .I3(n974[9]), .O(n6_adj_1404));
    defparam i2_4_lut_adj_111.LUT_INIT = 16'heca0;
    SB_LUT4 i1_2_lut_adj_112 (.I0(bluejay_data_out_31__N_922), .I1(buffer_switch_done_latched), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_1405));
    defparam i1_2_lut_adj_112.LUT_INIT = 16'heeee;
    SB_LUT4 i4026_4_lut (.I0(n5043), .I1(bluejay_data_out_31__N_920), .I2(n5_adj_1405), 
            .I3(n6_adj_1404), .O(n5525));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4026_4_lut.LUT_INIT = 16'haaa8;
    SB_LUT4 i3_4_lut (.I0(n1244), .I1(n1528), .I2(n974[5]), .I3(n74[2]), 
            .O(n9));   // src/bluejay_data.v(66[9] 129[16])
    defparam i3_4_lut.LUT_INIT = 16'hfc50;
    SB_LUT4 i4027_4_lut (.I0(n5043), .I1(n74[3]), .I2(n13811), .I3(n1528), 
            .O(n5526));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4027_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_2_lut_adj_113 (.I0(n74[3]), .I1(n4_adj_1406), .I2(GND_net), 
            .I3(GND_net), .O(n14214));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_113.LUT_INIT = 16'h8888;
    SB_LUT4 select_650_Select_4_i3_2_lut (.I0(n74[4]), .I1(n1528), .I2(GND_net), 
            .I3(GND_net), .O(n3));   // src/bluejay_data.v(66[9] 129[16])
    defparam select_650_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4028_4_lut (.I0(n5043), .I1(state_timeout_counter[4]), .I2(n3), 
            .I3(n45), .O(n5527));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4028_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_2_lut_adj_114 (.I0(n74[4]), .I1(n4_adj_1406), .I2(GND_net), 
            .I3(GND_net), .O(n14122));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_114.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_115 (.I0(buffer_switch_done_latched), .I1(n974[2]), 
            .I2(n6_adj_1407), .I3(state_timeout_counter[5]), .O(n14481));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_4_lut_adj_115.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_116 (.I0(n974[2]), .I1(n74[6]), .I2(state_timeout_counter[6]), 
            .I3(n1528), .O(n14482));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_4_lut_adj_116.LUT_INIT = 16'heca0;
    SB_DFFN bluejay_data_out_i1 (.Q(DEBUG_8_c), .C(SLM_CLK_c), .D(n6982));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 i1_2_lut_adj_117 (.I0(n74[6]), .I1(n4_adj_1406), .I2(GND_net), 
            .I3(GND_net), .O(n14050));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_117.LUT_INIT = 16'h8888;
    SB_LUT4 select_650_Select_7_i3_2_lut (.I0(n74[7]), .I1(n1528), .I2(GND_net), 
            .I3(GND_net), .O(n3_adj_1408));   // src/bluejay_data.v(66[9] 129[16])
    defparam select_650_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4031_4_lut (.I0(n5043), .I1(state_timeout_counter[7]), .I2(n3_adj_1408), 
            .I3(n45), .O(n5530));   // src/bluejay_data.v(56[8] 131[4])
    defparam i4031_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_2_lut_adj_118 (.I0(n74[7]), .I1(n4_adj_1406), .I2(GND_net), 
            .I3(GND_net), .O(n14026));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_118.LUT_INIT = 16'h8888;
    SB_DFFESS state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(SLM_CLK_c), 
            .E(n5043), .D(n14196), .S(n5431));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESR v_counter_i0 (.Q(v_counter[0]), .C(SLM_CLK_c), .E(n5132), 
            .D(v_counter_10__N_900[0]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 131[4])
    SB_LUT4 sub_122_add_2_2_lut (.I0(GND_net), .I1(v_counter[0]), .I2(n910), 
            .I3(VCC_net), .O(v_counter_10__N_900[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_2 (.CI(VCC_net), .I0(v_counter[0]), .I1(n910), 
            .CO(n13652));
    SB_DFFNESR bluejay_data_out_i11 (.Q(DATA10_c_10), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5414));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i10 (.Q(DATA9_c_9), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5413));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 sub_120_add_2_7_lut (.I0(n14552), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n13649), .O(n6_adj_1407)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_120_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n13651), .O(n74[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_120_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n13650), .O(n74[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_120_add_2_8 (.CI(n13650), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n13651));
    SB_LUT4 sub_122_add_2_12_lut (.I0(GND_net), .I1(v_counter[10]), .I2(VCC_net), 
            .I3(n13661), .O(v_counter_10__N_900[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_120_add_2_6_lut (.I0(GND_net), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n13648), .O(n74[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_122_add_2_11_lut (.I0(GND_net), .I1(v_counter[9]), .I2(VCC_net), 
            .I3(n13660), .O(v_counter_10__N_900[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFNESR bluejay_data_out_i12 (.Q(DATA11_c_11), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5412));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i13 (.Q(DATA12_c_12), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5411));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFSR state_FSM_i2 (.Q(n989), .C(SLM_CLK_c), .D(n14298), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i3 (.Q(n974[2]), .C(SLM_CLK_c), .D(n14489), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i4 (.Q(bluejay_data_out_31__N_919), .C(SLM_CLK_c), 
            .D(n1028), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i5 (.Q(n974[4]), .C(SLM_CLK_c), .D(n3546), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i6 (.Q(n974[5]), .C(SLM_CLK_c), .D(n3548), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i7 (.Q(bluejay_data_out_31__N_920), .C(SLM_CLK_c), 
            .D(n1037), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i8 (.Q(bluejay_data_out_31__N_921), .C(SLM_CLK_c), 
            .D(n3550), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i9 (.Q(bluejay_data_out_31__N_922), .C(SLM_CLK_c), 
            .D(n1041), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFSR state_FSM_i10 (.Q(n974[9]), .C(SLM_CLK_c), .D(n3552), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 129[16])
    SB_DFFN sync_68 (.Q(SYNC_c), .C(SLM_CLK_c), .D(bluejay_data_out_31__N_919));   // src/bluejay_data.v(134[8] 156[4])
    SB_CARRY sub_122_add_2_11 (.CI(n13660), .I0(v_counter[9]), .I1(VCC_net), 
            .CO(n13661));
    SB_LUT4 sub_120_add_2_5_lut (.I0(GND_net), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n13647), .O(n74[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_122_add_2_10_lut (.I0(GND_net), .I1(v_counter[8]), .I2(VCC_net), 
            .I3(n13659), .O(v_counter_10__N_900[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_10 (.CI(n13659), .I0(v_counter[8]), .I1(VCC_net), 
            .CO(n13660));
    SB_LUT4 sub_122_add_2_9_lut (.I0(GND_net), .I1(v_counter[7]), .I2(VCC_net), 
            .I3(n13658), .O(v_counter_10__N_900[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_120_add_2_7 (.CI(n13649), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n13650));
    SB_LUT4 sub_120_add_2_3_lut (.I0(GND_net), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n13645), .O(n74[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_9 (.CI(n13658), .I0(v_counter[7]), .I1(VCC_net), 
            .CO(n13659));
    SB_LUT4 sub_122_add_2_8_lut (.I0(GND_net), .I1(v_counter[6]), .I2(VCC_net), 
            .I3(n13657), .O(v_counter_10__N_900[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_8 (.CI(n13657), .I0(v_counter[6]), .I1(VCC_net), 
            .CO(n13658));
    SB_LUT4 sub_122_add_2_7_lut (.I0(GND_net), .I1(v_counter[5]), .I2(VCC_net), 
            .I3(n13656), .O(v_counter_10__N_900[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_120_add_2_3 (.CI(n13645), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n13646));
    SB_CARRY sub_120_add_2_5 (.CI(n13647), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n13648));
    SB_CARRY sub_122_add_2_7 (.CI(n13656), .I0(v_counter[5]), .I1(VCC_net), 
            .CO(n13657));
    SB_LUT4 sub_122_add_2_6_lut (.I0(GND_net), .I1(v_counter[4]), .I2(VCC_net), 
            .I3(n13655), .O(v_counter_10__N_900[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_120_add_2_4_lut (.I0(GND_net), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n13646), .O(n74[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_6 (.CI(n13655), .I0(v_counter[4]), .I1(VCC_net), 
            .CO(n13656));
    SB_LUT4 sub_122_add_2_5_lut (.I0(GND_net), .I1(v_counter[3]), .I2(VCC_net), 
            .I3(n13654), .O(v_counter_10__N_900[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_120_add_2_2_lut (.I0(GND_net), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n74[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_120_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_5 (.CI(n13654), .I0(v_counter[3]), .I1(VCC_net), 
            .CO(n13655));
    SB_CARRY sub_120_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n13645));
    SB_CARRY sub_120_add_2_6 (.CI(n13648), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n13649));
    SB_CARRY sub_120_add_2_4 (.CI(n13646), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n13647));
    SB_LUT4 sub_122_add_2_4_lut (.I0(GND_net), .I1(v_counter[2]), .I2(VCC_net), 
            .I3(n13653), .O(v_counter_10__N_900[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_122_add_2_4 (.CI(n13653), .I0(v_counter[2]), .I1(VCC_net), 
            .CO(n13654));
    SB_LUT4 i1_2_lut_adj_119 (.I0(n974[9]), .I1(buffer_switch_done), .I2(GND_net), 
            .I3(GND_net), .O(n5132));
    defparam i1_2_lut_adj_119.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_120 (.I0(bluejay_data_out_31__N_921), .I1(bluejay_data_out_31__N_922), 
            .I2(GND_net), .I3(GND_net), .O(valid_N_925));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_adj_120.LUT_INIT = 16'heeee;
    SB_DFFNESR bluejay_data_out_i14 (.Q(DATA13_c_13), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5410));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i15 (.Q(DATA14_c_14), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5409));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i9 (.Q(DATA8_c_8), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5408));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i16 (.Q(DATA15_c_15), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5407));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i17 (.Q(DATA16_c_16), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5406));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i8 (.Q(DATA7_c_7), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5405));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i18 (.Q(DATA17_c_17), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5404));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i19 (.Q(DATA18_c_18), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5403));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i7 (.Q(DATA6_c_6), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5402));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i20 (.Q(DATA19_c_19), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5401));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i21 (.Q(DATA20_c_20), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5400));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i6 (.Q(DATA5_c_5), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5399));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i22 (.Q(DATA21_c_21), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5398));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 sub_122_add_2_3_lut (.I0(GND_net), .I1(v_counter[1]), .I2(VCC_net), 
            .I3(n13652), .O(v_counter_10__N_900[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_122_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFNESR bluejay_data_out_i23 (.Q(DATA22_c_22), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5397));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i5 (.Q(DATA4_c_4), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5396));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i24 (.Q(DATA23_c_23), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5395));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFESS state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(SLM_CLK_c), 
            .E(n5043), .D(n14026), .S(n5530));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFNESR bluejay_data_out_i25 (.Q(DATA24_c_24), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5394));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFESS state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n5043), .D(n14050), .S(n5529));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(SLM_CLK_c), 
            .E(n5043), .D(n14481), .S(n5528));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(SLM_CLK_c), 
            .E(n5043), .D(n14122), .S(n5527));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(SLM_CLK_c), 
            .E(n5043), .D(n14214), .S(n5526));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFESS state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n5043), .D(n9), .S(n5525));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFNESR bluejay_data_out_i4 (.Q(DATA3_c_3), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5393));   // src/bluejay_data.v(134[8] 156[4])
    SB_CARRY sub_122_add_2_3 (.CI(n13652), .I0(v_counter[1]), .I1(VCC_net), 
            .CO(n13653));
    SB_DFFESS state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(SLM_CLK_c), 
            .E(n5043), .D(n14186), .S(n5431));   // src/bluejay_data.v(56[8] 131[4])
    SB_DFFN get_next_word_67 (.Q(get_next_word), .C(SLM_CLK_c), .D(n5625));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i26 (.Q(DATA25_c_25), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5392));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i27 (.Q(DATA26_c_26), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5391));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i3 (.Q(DATA2_c_2), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5390));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i28 (.Q(DATA27_c_27), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5389));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i29 (.Q(DATA28_c_28), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5388));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i2 (.Q(DATA1_c_1), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5387));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i30 (.Q(DATA29_c_29), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5386));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i31 (.Q(DATA30_c_30), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5385));   // src/bluejay_data.v(134[8] 156[4])
    SB_DFFNESR bluejay_data_out_i32 (.Q(DATA31_c_31), .C(SLM_CLK_c), .E(VCC_net), 
            .D(valid_N_925), .R(n5384));   // src/bluejay_data.v(134[8] 156[4])
    SB_LUT4 i1_2_lut_4_lut (.I0(n99[2]), .I1(n910), .I2(n974[9]), .I3(n14551), 
            .O(n14552));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffd0;
    SB_LUT4 i1_3_lut (.I0(n910), .I1(bluejay_data_out_31__N_921), .I2(sc32_fifo_almost_empty), 
            .I3(GND_net), .O(n1041));   // src/bluejay_data.v(87[17] 89[20])
    defparam i1_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 i1_4_lut_adj_121 (.I0(sc32_fifo_almost_empty), .I1(bluejay_data_out_31__N_920), 
            .I2(n102), .I3(bluejay_data_out_31__N_921), .O(n3550));   // src/bluejay_data.v(62[9] 65[12])
    defparam i1_4_lut_adj_121.LUT_INIT = 16'hdccc;
    SB_LUT4 i1_4_lut_adj_122 (.I0(n910), .I1(n974[5]), .I2(n974[4]), .I3(line_of_data_available), 
            .O(n1037));
    defparam i1_4_lut_adj_122.LUT_INIT = 16'h5450;
    SB_LUT4 i2_4_lut_adj_123 (.I0(buffer_switch_done_latched), .I1(n910), 
            .I2(n974[5]), .I3(line_of_data_available), .O(n13836));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_4_lut_adj_123.LUT_INIT = 16'h4050;
    SB_LUT4 i2068_4_lut (.I0(n13836), .I1(n910), .I2(n99[2]), .I3(n974[9]), 
            .O(n3548));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2068_4_lut.LUT_INIT = 16'hbaaa;
    SB_LUT4 i1_2_lut_adj_124 (.I0(n910), .I1(buffer_switch_done_latched), 
            .I2(GND_net), .I3(GND_net), .O(n102));   // src/bluejay_data.v(62[9] 65[12])
    defparam i1_2_lut_adj_124.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_125 (.I0(n910), .I1(n989), .I2(GND_net), .I3(GND_net), 
            .O(n106));   // src/bluejay_data.v(107[21:49])
    defparam i1_2_lut_adj_125.LUT_INIT = 16'h4444;
    SB_LUT4 i12507_4_lut (.I0(n14472), .I1(n14475), .I2(n14569), .I3(n13), 
            .O(n14627));
    defparam i12507_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_126 (.I0(n14627), .I1(state_timeout_counter[0]), 
            .I2(n974[9]), .I3(GND_net), .O(n13985));
    defparam i2_3_lut_adj_126.LUT_INIT = 16'h4040;
    SB_LUT4 i1_4_lut_adj_127 (.I0(n974[2]), .I1(n13985), .I2(line_of_data_available), 
            .I3(n106), .O(n14489));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_4_lut_adj_127.LUT_INIT = 16'hefee;
    SB_LUT4 i1_3_lut_4_lut (.I0(n99[2]), .I1(n910), .I2(n74[0]), .I3(n974[9]), 
            .O(n8));   // src/bluejay_data.v(107[17] 116[20])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf200;
    SB_LUT4 i1_3_lut_4_lut_adj_128 (.I0(n974[4]), .I1(bluejay_data_out_31__N_919), 
            .I2(n910), .I3(buffer_switch_done_latched), .O(n3546));   // src/bluejay_data.v(62[9] 65[12])
    defparam i1_3_lut_4_lut_adj_128.LUT_INIT = 16'hccec;
    SB_LUT4 i1_3_lut_4_lut_adj_129 (.I0(n974[9]), .I1(bluejay_data_out_31__N_922), 
            .I2(n910), .I3(buffer_switch_done_latched), .O(n3552));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_3_lut_4_lut_adj_129.LUT_INIT = 16'hccec;
    SB_LUT4 i1_2_lut_3_lut (.I0(n99[2]), .I1(n910), .I2(n74[2]), .I3(GND_net), 
            .O(n59));   // src/bluejay_data.v(107[17] 116[20])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_2_lut_3_lut_adj_130 (.I0(n99[2]), .I1(n910), .I2(n974[9]), 
            .I3(GND_net), .O(n2));   // src/bluejay_data.v(107[17] 116[20])
    defparam i1_2_lut_3_lut_adj_130.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_3_lut_4_lut_adj_131 (.I0(n99[2]), .I1(n910), .I2(n74[1]), 
            .I3(n974[9]), .O(n8_adj_1403));   // src/bluejay_data.v(107[17] 116[20])
    defparam i1_3_lut_4_lut_adj_131.LUT_INIT = 16'hf200;
    SB_LUT4 i2_2_lut_3_lut (.I0(state_timeout_counter[3]), .I1(buffer_switch_done_latched), 
            .I2(n974[2]), .I3(GND_net), .O(n13811));   // src/bluejay_data.v(66[9] 129[16])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_3_lut_adj_132 (.I0(state_timeout_counter[1]), .I1(buffer_switch_done_latched), 
            .I2(n974[2]), .I3(GND_net), .O(n5_adj_1402));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_3_lut_adj_132.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_3_lut_adj_133 (.I0(state_timeout_counter[0]), .I1(buffer_switch_done_latched), 
            .I2(n974[2]), .I3(GND_net), .O(n5));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_3_lut_adj_133.LUT_INIT = 16'h2020;
    SB_LUT4 i2_3_lut_4_lut (.I0(state_timeout_counter[6]), .I1(state_timeout_counter[7]), 
            .I2(n14472), .I3(state_timeout_counter[0]), .O(n910));   // src/bluejay_data.v(107[21:49])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_4_lut_adj_134 (.I0(v_counter[9]), .I1(n4), .I2(v_counter[10]), 
            .I3(n14569), .O(n99[2]));   // src/bluejay_data.v(56[8] 131[4])
    defparam i1_2_lut_4_lut_adj_134.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n974[5]), .I1(n910), .I2(line_of_data_available), 
            .I3(n2), .O(n4_adj_1406));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hffa8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_135 (.I0(n974[5]), .I1(n910), .I2(line_of_data_available), 
            .I3(n1528), .O(n14551));   // src/bluejay_data.v(66[9] 129[16])
    defparam i1_2_lut_3_lut_4_lut_adj_135.LUT_INIT = 16'hffa8;
    
endmodule
//
// Verilog Description of module fifo_sc_32_lut_gen
//

module fifo_sc_32_lut_gen (n5412, GND_net, \sc32_fifo_data_out[0] , SLM_CLK_c, 
            dc32_fifo_data_out, \MISC.empty_flag_r , sc32_fifo_almost_empty, 
            reset_all, n5384, n5385, n5386, n5387, n5388, n5389, 
            n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, 
            n5398, n5399, n5400, n5401, n5402, n5403, n5404, sc32_fifo_write_enable, 
            n5405, n5406, n5407, n5408, n5409, n5410, sc32_fifo_read_enable, 
            n5413, n5414, n5411) /* synthesis syn_module_defined=1 */ ;
    output n5412;
    input GND_net;
    output \sc32_fifo_data_out[0] ;
    input SLM_CLK_c;
    input [31:0]dc32_fifo_data_out;
    output \MISC.empty_flag_r ;
    output sc32_fifo_almost_empty;
    input reset_all;
    output n5384;
    output n5385;
    output n5386;
    output n5387;
    output n5388;
    output n5389;
    output n5390;
    output n5391;
    output n5392;
    output n5393;
    output n5394;
    output n5395;
    output n5396;
    output n5397;
    output n5398;
    output n5399;
    output n5400;
    output n5401;
    output n5402;
    output n5403;
    output n5404;
    input sc32_fifo_write_enable;
    output n5405;
    output n5406;
    output n5407;
    output n5408;
    output n5409;
    output n5410;
    input sc32_fifo_read_enable;
    output n5413;
    output n5414;
    output n5411;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    fifo_sc_32_lut_gen_ipgen_lscc_fifo_renamed_due_excessive_length_2 lscc_fifo_inst (.n5412(n5412), 
            .GND_net(GND_net), .\sc32_fifo_data_out[0] (\sc32_fifo_data_out[0] ), 
            .SLM_CLK_c(SLM_CLK_c), .dc32_fifo_data_out({dc32_fifo_data_out}), 
            .\MISC.empty_flag_r (\MISC.empty_flag_r ), .sc32_fifo_almost_empty(sc32_fifo_almost_empty), 
            .reset_all(reset_all), .n5384(n5384), .n5385(n5385), .n5386(n5386), 
            .n5387(n5387), .n5388(n5388), .n5389(n5389), .n5390(n5390), 
            .n5391(n5391), .n5392(n5392), .n5393(n5393), .n5394(n5394), 
            .n5395(n5395), .n5396(n5396), .n5397(n5397), .n5398(n5398), 
            .n5399(n5399), .n5400(n5400), .n5401(n5401), .n5402(n5402), 
            .n5403(n5403), .n5404(n5404), .sc32_fifo_write_enable(sc32_fifo_write_enable), 
            .n5405(n5405), .n5406(n5406), .n5407(n5407), .n5408(n5408), 
            .n5409(n5409), .n5410(n5410), .sc32_fifo_read_enable(sc32_fifo_read_enable), 
            .n5413(n5413), .n5414(n5414), .n5411(n5411)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_sc_32_lut_gen.v(45[37] 59[45])
    
endmodule
//
// Verilog Description of module fifo_sc_32_lut_gen_ipgen_lscc_fifo_renamed_due_excessive_length_2
//

module fifo_sc_32_lut_gen_ipgen_lscc_fifo_renamed_due_excessive_length_2 (n5412, 
            GND_net, \sc32_fifo_data_out[0] , SLM_CLK_c, dc32_fifo_data_out, 
            \MISC.empty_flag_r , sc32_fifo_almost_empty, reset_all, n5384, 
            n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, 
            n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, 
            n5401, n5402, n5403, n5404, sc32_fifo_write_enable, n5405, 
            n5406, n5407, n5408, n5409, n5410, sc32_fifo_read_enable, 
            n5413, n5414, n5411) /* synthesis syn_module_defined=1 */ ;
    output n5412;
    input GND_net;
    output \sc32_fifo_data_out[0] ;
    input SLM_CLK_c;
    input [31:0]dc32_fifo_data_out;
    output \MISC.empty_flag_r ;
    output sc32_fifo_almost_empty;
    input reset_all;
    output n5384;
    output n5385;
    output n5386;
    output n5387;
    output n5388;
    output n5389;
    output n5390;
    output n5391;
    output n5392;
    output n5393;
    output n5394;
    output n5395;
    output n5396;
    output n5397;
    output n5398;
    output n5399;
    output n5400;
    output n5401;
    output n5402;
    output n5403;
    output n5404;
    input sc32_fifo_write_enable;
    output n5405;
    output n5406;
    output n5407;
    output n5408;
    output n5409;
    output n5410;
    input sc32_fifo_read_enable;
    output n5413;
    output n5414;
    output n5411;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [31:0]sc32_fifo_data_out;   // src/top.v(646[12:30])
    wire [31:0]rd_data_o_31__N_759;
    
    wire \MISC.rd_w , n7;
    wire [3:0]wr_addr_r;   // src/fifo_sc_32_lut_gen.v(117[48:57])
    
    wire \mem_REG.mem_0_31 , n6692, \mem_REG.mem_0_30 , n6691, \mem_REG.mem_0_29 , 
        n6690, \mem_REG.mem_0_28 , n6689, \mem_REG.mem_0_27 , n6688, 
        \mem_REG.mem_0_26 , n6687, \mem_REG.mem_0_25 , n6686, \mem_REG.mem_0_24 , 
        n6685, \mem_REG.mem_0_23 , n6684, \mem_REG.mem_0_22 , n6683, 
        \mem_REG.mem_0_21 , n6682, \mem_REG.mem_0_20 , n6681, \mem_REG.mem_0_19 , 
        n6680, \mem_REG.mem_0_18 , n6679, \mem_REG.mem_0_17 , n6678, 
        \mem_REG.mem_0_16 , n6677, \mem_REG.mem_0_15 , n6676, \mem_REG.mem_0_14 , 
        n6675, \mem_REG.mem_0_13 , n6674;
    wire [3:0]wr_addr_r_3__N_690;
    wire [3:0]\MISC.wr_flag_addr_r ;   // src/fifo_sc_32_lut_gen.v(261[56:70])
    wire [3:0]wr_addr_p1_r_3__N_694;
    wire [3:0]\MISC.wr_flag_addr_p1_r ;   // src/fifo_sc_32_lut_gen.v(262[56:73])
    wire [3:0]rd_addr_r_3__N_708;
    wire [3:0]\MISC.rd_flag_addr_r ;   // src/fifo_sc_32_lut_gen.v(263[56:70])
    
    wire \mem_REG.mem_0_12 , n6673, \mem_REG.mem_0_11 , n6672, \mem_REG.mem_0_10 , 
        n6671, \mem_REG.mem_0_9 , n6670;
    wire [3:0]rd_addr_p1_r_3__N_712;
    wire [3:0]\MISC.rd_flag_addr_p1_r ;   // src/fifo_sc_32_lut_gen.v(264[56:73])
    
    wire full_ext_r_N_794, \MISC.full_flag_r , empty_ext_r_N_796, \MISC.AEmpty.almost_empty_nxt_w , 
        \mem_REG.mem_0_8 , n6669, \mem_REG.mem_0_7 , n6668, \mem_REG.mem_0_6 , 
        n6667, \mem_REG.mem_0_5 , n6666, \mem_REG.mem_0_4 , n6665, 
        \mem_REG.mem_0_3 , n6664, \mem_REG.mem_0_2 , n6663, \mem_REG.mem_0_1 , 
        n6662, \mem_REG.mem_0_0 , n6661;
    wire [3:0]rd_addr_r;   // src/fifo_sc_32_lut_gen.v(123[48:57])
    
    wire n15396, n15397, n17031, n15394, n15393, n8, \mem_REG.mem_7_31 , 
        n6916, \mem_REG.mem_7_30 , n6915, \mem_REG.mem_7_29 , n6914, 
        n6913, \mem_REG.mem_7_28 , n6912, \mem_REG.mem_7_27 , n6911, 
        \mem_REG.mem_7_26 , n6910, \mem_REG.mem_7_25 , n6909, \mem_REG.mem_7_24 , 
        n6908, \mem_REG.mem_7_23 , n6907, \mem_REG.mem_7_22 , n6906, 
        \mem_REG.mem_7_21 , n6905, \mem_REG.mem_7_20 , n6904, \mem_REG.mem_7_19 , 
        n6903, \mem_REG.mem_7_18 , n6902, \mem_REG.mem_7_17 , n6901, 
        \mem_REG.mem_7_16 , n6900, \mem_REG.mem_7_15 , n6899, \mem_REG.mem_7_14 , 
        n6898, \mem_REG.mem_7_13 , n6897, \mem_REG.mem_7_12 , n6896, 
        \mem_REG.mem_7_11 , n6895, \mem_REG.mem_7_10 , n6894, \mem_REG.mem_7_9 , 
        n6893, \mem_REG.mem_7_8 , n6892, \mem_REG.mem_7_7 , n6891, 
        \mem_REG.mem_7_6 , n6890, \mem_REG.mem_7_5 , n6889, \mem_REG.mem_7_4 , 
        n6888, \mem_REG.mem_7_3 , n6887, \mem_REG.mem_7_2 , n6886, 
        \mem_REG.mem_7_1 , n6885, \mem_REG.mem_7_0 , n6884, \mem_REG.mem_6_31 , 
        n6883, \mem_REG.mem_6_30 , n6882, \mem_REG.mem_6_29 , n6881, 
        \mem_REG.mem_6_28 , n6880, \mem_REG.mem_6_27 , n6879, \mem_REG.mem_6_26 , 
        n6878, \mem_REG.mem_6_25 , n6877, \mem_REG.mem_6_24 , n6876, 
        \mem_REG.mem_6_23 , n6875, \mem_REG.mem_6_22 , n6874, \mem_REG.mem_6_21 , 
        n6873, \mem_REG.mem_6_20 , n6872, \mem_REG.mem_6_19 , n6871, 
        \mem_REG.mem_6_18 , n6870, \mem_REG.mem_6_17 , n6869, \mem_REG.mem_6_16 , 
        n6868, \mem_REG.mem_6_15 , n6867, \mem_REG.mem_6_14 , n6866, 
        \mem_REG.mem_6_13 , n6865, \mem_REG.mem_6_12 , n6864, \mem_REG.mem_6_11 , 
        n6863, \mem_REG.mem_6_10 , n6862, \mem_REG.mem_6_9 , n6861, 
        \mem_REG.mem_6_8 , n6860, \mem_REG.mem_6_7 , n6859, \mem_REG.mem_6_6 , 
        n6858, \mem_REG.mem_6_5 , n6857, \mem_REG.mem_6_4 , n6856, 
        \mem_REG.mem_6_3 , n6855, \mem_REG.mem_6_2 , n6854, \mem_REG.mem_6_1 , 
        n6853, \mem_REG.mem_6_0 , n6852, \mem_REG.mem_5_31 , n6851, 
        \mem_REG.mem_5_30 , n6850, \mem_REG.mem_5_29 , n6849, \mem_REG.mem_5_28 , 
        n6848, \mem_REG.mem_5_27 , n6847, \mem_REG.mem_5_26 , n6846, 
        \mem_REG.mem_5_25 , n6845, \mem_REG.mem_5_24 , n6844, \mem_REG.mem_5_23 , 
        n6843, \mem_REG.mem_5_22 , n6842, \mem_REG.mem_5_21 , n6841, 
        \mem_REG.mem_5_20 , n6840, \mem_REG.mem_5_19 , n6839, \mem_REG.mem_5_18 , 
        n6838, \mem_REG.mem_5_17 , n6837, \mem_REG.mem_5_16 , n6836, 
        \mem_REG.mem_5_15 , n6835, \mem_REG.mem_5_14 , n6834, \mem_REG.mem_5_13 , 
        n6833, \mem_REG.mem_5_12 , n6832, \mem_REG.mem_5_11 , n6831, 
        \mem_REG.mem_5_10 , n6830, \mem_REG.mem_5_9 , n6829, \mem_REG.mem_5_8 , 
        n6828, \mem_REG.mem_5_7 , n6827, \mem_REG.mem_5_6 , n6826, 
        \mem_REG.mem_5_5 , n6825, \mem_REG.mem_5_4 , n6824, \mem_REG.mem_5_3 , 
        n6823, \mem_REG.mem_5_2 , n6822, \mem_REG.mem_5_1 , n6821, 
        \mem_REG.mem_5_0 , n6820, \mem_REG.mem_4_31 , n6819, \mem_REG.mem_4_30 , 
        n6818, \mem_REG.mem_4_29 , n6817, \mem_REG.mem_4_28 , n6816, 
        \mem_REG.mem_4_27 , n6815, \mem_REG.mem_4_26 , n6814, \mem_REG.mem_4_25 , 
        n6813, \mem_REG.mem_4_24 , n6812, \mem_REG.mem_4_23 , n6811, 
        \mem_REG.mem_4_22 , n6810, \mem_REG.mem_4_21 , n6809, \mem_REG.mem_4_20 , 
        n6808, \mem_REG.mem_4_19 , n6807, \mem_REG.mem_4_18 , n6806, 
        \mem_REG.mem_4_17 , n6805, \mem_REG.mem_4_16 , n6804, \mem_REG.mem_4_15 , 
        n6803, \mem_REG.mem_4_14 , n6802, \mem_REG.mem_4_13 , n6801, 
        \mem_REG.mem_4_12 , n6800, \mem_REG.mem_4_11 , n6799, \mem_REG.mem_4_10 , 
        n6798, \mem_REG.mem_4_9 , n6797, \mem_REG.mem_4_8 , n6796, 
        \mem_REG.mem_4_7 , n6795, \mem_REG.mem_4_6 , n6794, \mem_REG.mem_4_5 , 
        n6793, \mem_REG.mem_4_4 , n6792, \mem_REG.mem_4_3 , n6791, 
        \mem_REG.mem_4_2 , n6790, \mem_REG.mem_4_1 , n6789, \mem_REG.mem_4_0 , 
        n6788, \mem_REG.mem_3_31 , n6787, \mem_REG.mem_3_30 , n6786, 
        \mem_REG.mem_3_29 , n6785, \mem_REG.mem_3_28 , n6784, \mem_REG.mem_3_27 , 
        n6783, \mem_REG.mem_3_26 , n6782, \mem_REG.mem_3_25 , n6781, 
        \mem_REG.mem_3_24 , n6780, \mem_REG.mem_3_23 , n6779, \mem_REG.mem_3_22 , 
        n6778, \mem_REG.mem_3_21 , n6777, \mem_REG.mem_3_20 , n6776, 
        \mem_REG.mem_3_19 , n6775, \mem_REG.mem_3_18 , n6774, \mem_REG.mem_3_17 , 
        n6773, \mem_REG.mem_3_16 , n6772, \mem_REG.mem_3_15 , n6771, 
        \mem_REG.mem_3_14 , n6770, \mem_REG.mem_3_13 , n6769, \mem_REG.mem_3_12 , 
        n6768, \mem_REG.mem_3_11 , n6767, \mem_REG.mem_3_10 , n6766, 
        \mem_REG.mem_3_9 , n6765, \mem_REG.mem_3_8 , n6764, \mem_REG.mem_3_7 , 
        n6763, \mem_REG.mem_3_6 , n6762, \mem_REG.mem_3_5 , n6761, 
        \mem_REG.mem_3_4 , n6760, \mem_REG.mem_3_3 , n6759, \mem_REG.mem_3_2 , 
        n6758, \mem_REG.mem_3_1 , n6757, \mem_REG.mem_3_0 , n6756, 
        \mem_REG.mem_2_31 , n6755, \mem_REG.mem_2_30 , n6754, \mem_REG.mem_2_29 , 
        n6753, \mem_REG.mem_2_28 , n6752, \mem_REG.mem_2_27 , n6751, 
        \mem_REG.mem_2_26 , n6750, \mem_REG.mem_2_25 , n6749, \mem_REG.mem_2_24 , 
        n6748, \mem_REG.mem_2_23 , n6747, \mem_REG.mem_2_22 , n6746, 
        \mem_REG.mem_2_21 , n6745, \mem_REG.mem_2_20 , n6744, \mem_REG.mem_2_19 , 
        n6743, \mem_REG.mem_2_18 , n6742, \mem_REG.mem_2_17 , n6741, 
        \mem_REG.mem_2_16 , n6740, \mem_REG.mem_2_15 , n6739, \mem_REG.mem_2_14 , 
        n6738, \mem_REG.mem_2_13 , n6737, \mem_REG.mem_2_12 , n6736, 
        \mem_REG.mem_2_11 , n6735, \mem_REG.mem_2_10 , n6734, \mem_REG.mem_2_9 , 
        n6733, \mem_REG.mem_2_8 , n6732, \mem_REG.mem_2_7 , n6731, 
        \mem_REG.mem_2_6 , n6730, \mem_REG.mem_2_5 , n6729, \mem_REG.mem_2_4 , 
        n6728, \mem_REG.mem_2_3 , n6727, \mem_REG.mem_2_2 , n6726, 
        \mem_REG.mem_2_1 , n6725, \mem_REG.mem_2_0 , n6724, \mem_REG.mem_1_31 , 
        n6723, \mem_REG.mem_1_30 , n6722, \mem_REG.mem_1_29 , n6721, 
        \mem_REG.mem_1_28 , n6720, \mem_REG.mem_1_27 , n6719, \mem_REG.mem_1_26 , 
        n6718, \mem_REG.mem_1_25 , n6717, \mem_REG.mem_1_24 , n6716, 
        \mem_REG.mem_1_23 , n6715, \mem_REG.mem_1_22 , n6714, \mem_REG.mem_1_21 , 
        n6713, \mem_REG.mem_1_20 , n6712, \mem_REG.mem_1_19 , n6711, 
        \mem_REG.mem_1_18 , n6710, \mem_REG.mem_1_17 , n6709, \mem_REG.mem_1_16 , 
        n6708, \mem_REG.mem_1_15 , n6707, \mem_REG.mem_1_14 , n6706, 
        \mem_REG.mem_1_13 , n6705, \mem_REG.mem_1_12 , n6704, \mem_REG.mem_1_11 , 
        n6703, \mem_REG.mem_1_10 , n6702, \mem_REG.mem_1_9 , n6701, 
        \mem_REG.mem_1_8 , n6700, \mem_REG.mem_1_7 , n6699, \mem_REG.mem_1_6 , 
        n6698, \mem_REG.mem_1_5 , n6697, \mem_REG.mem_1_4 , n6696, 
        \mem_REG.mem_1_3 , n6695, \mem_REG.mem_1_2 , n6694, \mem_REG.mem_1_1 , 
        n6693, \mem_REG.mem_1_0 , n15477, n15478, n16977, n15466, 
        n15465, n17637, n17640, n15555, n15597, n15598, n17577, 
        n15586, n15585, n15556, n15267, n15268, n16881, n15247, 
        n15246, n2495, n3894, n15756, n15757, n16875, n15748, 
        n15747, n17547;
    wire [3:0]wr_addr_p1_r;   // src/fifo_sc_32_lut_gen.v(118[48:60])
    wire [3:0]wr_addr_nxt_w;   // src/fifo_sc_32_lut_gen.v(130[28:41])
    
    wire n17550;
    wire [2:0]wr_cmpaddr_p1_r;   // src/fifo_sc_32_lut_gen.v(122[54:69])
    
    wire n15435, n15436, n16851, n15217, n15216, n15573, n15574, 
        n17535, n14655, n9, n15408, n15409, n15430, n15429, n15186, 
        n15187, n16815, n15157, n15156, n17487, n17490;
    wire [3:0]n2834;
    wire [3:0]rd_addr_p1cmp_r;   // src/fifo_sc_32_lut_gen.v(125[48:63])
    
    wire n3457, n15549, n15550, n17469, n15403, n15402, n3455, 
        n2, n4;
    wire [3:0]wr_addr_p1cmp_r_3__N_698;
    
    wire n3441, n13892, n4_adj_1397, n13894, n6, n17427, n15447, 
        n15448, n16725, n10, full_nxt_w_N_812, empty_nxt_w_N_823, 
        n14653, n17430, n15106, n15105, n4_adj_1398, n6_adj_1399, 
        n14621, full_nxt_w_N_797, n14607, n16713, n16716;
    wire [3:0]rd_addr_nxt_w;   // src/fifo_sc_32_lut_gen.v(133[28:41])
    
    wire n16701, n16704, n6_adj_1400, n15060, n15061, n15067, n15066, 
        n15450, n15451, n16677, n15070, n15069, n15441, n15442, 
        n17391, n17394, n15495, n15496, n17379, n15490, n15489, 
        n17373, n16167, n17376, n16170, n16227, n17349, n17352, 
        n15453, n15454, n17343, n17337, n17331, n17325, n16230, 
        n17328, n17313, n17316, n17301, n17304, n17283, n17286, 
        n17265, n17268, n17241, n17244, n17235, n17238, n17229, 
        n16461, n17232, n16464, n17985, n17988, n17223, n17226, 
        n17199, n17202, n17193, n17196, n17187, n17190, n17175, 
        n17178, n17913, n17916, n16389, n16392, n17889, n17892, 
        n3181, n3152, n16335, n16338, n16329, n16332, n17835, 
        n17838, n17115, n17118, n17106, n17103;
    
    SB_LUT4 i3913_1_lut (.I0(sc32_fifo_data_out[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5412));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3913_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE \mem_REG.data_raw_r_i0_i0  (.Q(\sc32_fifo_data_out[0] ), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[0]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_LUT4 i5193_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[31]), 
            .I3(\mem_REG.mem_0_31 ), .O(n6692));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5193_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5192_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[30]), 
            .I3(\mem_REG.mem_0_30 ), .O(n6691));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5192_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5191_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[29]), 
            .I3(\mem_REG.mem_0_29 ), .O(n6690));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5191_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5190_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[28]), 
            .I3(\mem_REG.mem_0_28 ), .O(n6689));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5190_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5189_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[27]), 
            .I3(\mem_REG.mem_0_27 ), .O(n6688));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5189_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5188_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[26]), 
            .I3(\mem_REG.mem_0_26 ), .O(n6687));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5188_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5187_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[25]), 
            .I3(\mem_REG.mem_0_25 ), .O(n6686));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5187_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5186_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[24]), 
            .I3(\mem_REG.mem_0_24 ), .O(n6685));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5186_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5185_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[23]), 
            .I3(\mem_REG.mem_0_23 ), .O(n6684));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5185_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5184_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[22]), 
            .I3(\mem_REG.mem_0_22 ), .O(n6683));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5184_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5183_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[21]), 
            .I3(\mem_REG.mem_0_21 ), .O(n6682));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5183_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5182_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[20]), 
            .I3(\mem_REG.mem_0_20 ), .O(n6681));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5182_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5181_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[19]), 
            .I3(\mem_REG.mem_0_19 ), .O(n6680));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5181_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5180_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[18]), 
            .I3(\mem_REG.mem_0_18 ), .O(n6679));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5180_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5179_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[17]), 
            .I3(\mem_REG.mem_0_17 ), .O(n6678));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5179_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5178_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[16]), 
            .I3(\mem_REG.mem_0_16 ), .O(n6677));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5178_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5177_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[15]), 
            .I3(\mem_REG.mem_0_15 ), .O(n6676));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5177_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5176_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[14]), 
            .I3(\mem_REG.mem_0_14 ), .O(n6675));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5176_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5175_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[13]), 
            .I3(\mem_REG.mem_0_13 ), .O(n6674));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5175_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF \MISC.wr_flag_addr_r_i0  (.Q(\MISC.wr_flag_addr_r [0]), .C(SLM_CLK_c), 
           .D(wr_addr_r_3__N_690[0]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFF \MISC.wr_flag_addr_p1_r_i0  (.Q(\MISC.wr_flag_addr_p1_r [0]), .C(SLM_CLK_c), 
           .D(wr_addr_p1_r_3__N_694[0]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFF \MISC.rd_flag_addr_r_i0  (.Q(\MISC.rd_flag_addr_r [0]), .C(SLM_CLK_c), 
           .D(rd_addr_r_3__N_708[0]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_LUT4 i5174_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[12]), 
            .I3(\mem_REG.mem_0_12 ), .O(n6673));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5174_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5173_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[11]), 
            .I3(\mem_REG.mem_0_11 ), .O(n6672));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5173_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5172_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[10]), 
            .I3(\mem_REG.mem_0_10 ), .O(n6671));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5172_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5171_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[9]), 
            .I3(\mem_REG.mem_0_9 ), .O(n6670));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5171_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF \MISC.rd_flag_addr_p1_r_i0  (.Q(\MISC.rd_flag_addr_p1_r [0]), .C(SLM_CLK_c), 
           .D(rd_addr_p1_r_3__N_712[0]));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFF \MISC.full_flag_r_143  (.Q(\MISC.full_flag_r ), .C(SLM_CLK_c), 
           .D(full_ext_r_N_794));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFF \MISC.empty_flag_r_144  (.Q(\MISC.empty_flag_r ), .C(SLM_CLK_c), 
           .D(empty_ext_r_N_796));   // src/fifo_sc_32_lut_gen.v(274[25] 296[28])
    SB_DFFSS \MISC.AEmpty.almost_empty_ext_r_147  (.Q(sc32_fifo_almost_empty), 
            .C(SLM_CLK_c), .D(\MISC.AEmpty.almost_empty_nxt_w ), .S(reset_all));   // src/fifo_sc_32_lut_gen.v(403[33] 415[36])
    SB_LUT4 i5170_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[8]), 
            .I3(\mem_REG.mem_0_8 ), .O(n6669));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5170_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5169_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[7]), 
            .I3(\mem_REG.mem_0_7 ), .O(n6668));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5169_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5168_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[6]), 
            .I3(\mem_REG.mem_0_6 ), .O(n6667));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5168_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5167_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[5]), 
            .I3(\mem_REG.mem_0_5 ), .O(n6666));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5167_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5166_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[4]), 
            .I3(\mem_REG.mem_0_4 ), .O(n6665));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5166_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5165_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[3]), 
            .I3(\mem_REG.mem_0_3 ), .O(n6664));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5165_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5164_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[2]), 
            .I3(\mem_REG.mem_0_2 ), .O(n6663));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5164_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5163_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[1]), 
            .I3(\mem_REG.mem_0_1 ), .O(n6662));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5163_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5162_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[0]), 
            .I3(\mem_REG.mem_0_0 ), .O(n6661));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5162_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15007 (.I0(rd_addr_r[1]), .I1(n15396), 
            .I2(n15397), .I3(rd_addr_r[2]), .O(n17031));
    defparam rd_addr_r_1__bdd_4_lut_15007.LUT_INIT = 16'he4aa;
    SB_LUT4 n17031_bdd_4_lut (.I0(n17031), .I1(n15394), .I2(n15393), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[0]));
    defparam n17031_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3885_1_lut (.I0(sc32_fifo_data_out[31]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5384));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3885_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3886_1_lut (.I0(sc32_fifo_data_out[30]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5385));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3886_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3887_1_lut (.I0(sc32_fifo_data_out[29]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5386));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3887_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3888_1_lut (.I0(sc32_fifo_data_out[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5387));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3888_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3889_1_lut (.I0(sc32_fifo_data_out[28]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5388));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3889_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3890_1_lut (.I0(sc32_fifo_data_out[27]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5389));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3890_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3891_1_lut (.I0(sc32_fifo_data_out[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5390));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3891_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3892_1_lut (.I0(sc32_fifo_data_out[26]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5391));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3892_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3893_1_lut (.I0(sc32_fifo_data_out[25]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5392));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3893_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3894_1_lut (.I0(sc32_fifo_data_out[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5393));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3894_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5417_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[31]), 
            .I3(\mem_REG.mem_7_31 ), .O(n6916));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5417_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5416_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[30]), 
            .I3(\mem_REG.mem_7_30 ), .O(n6915));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5416_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5415_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[29]), 
            .I3(\mem_REG.mem_7_29 ), .O(n6914));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5415_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i803_804 (.Q(\mem_REG.mem_7_31 ), .C(SLM_CLK_c), .D(n6916));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i800_801 (.Q(\mem_REG.mem_7_30 ), .C(SLM_CLK_c), .D(n6915));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i797_798 (.Q(\mem_REG.mem_7_29 ), .C(SLM_CLK_c), .D(n6914));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i794_795 (.Q(\mem_REG.mem_7_28 ), .C(SLM_CLK_c), .D(n6913));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i791_792 (.Q(\mem_REG.mem_7_27 ), .C(SLM_CLK_c), .D(n6912));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i788_789 (.Q(\mem_REG.mem_7_26 ), .C(SLM_CLK_c), .D(n6911));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i785_786 (.Q(\mem_REG.mem_7_25 ), .C(SLM_CLK_c), .D(n6910));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i782_783 (.Q(\mem_REG.mem_7_24 ), .C(SLM_CLK_c), .D(n6909));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i779_780 (.Q(\mem_REG.mem_7_23 ), .C(SLM_CLK_c), .D(n6908));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i776_777 (.Q(\mem_REG.mem_7_22 ), .C(SLM_CLK_c), .D(n6907));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i773_774 (.Q(\mem_REG.mem_7_21 ), .C(SLM_CLK_c), .D(n6906));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i770_771 (.Q(\mem_REG.mem_7_20 ), .C(SLM_CLK_c), .D(n6905));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i767_768 (.Q(\mem_REG.mem_7_19 ), .C(SLM_CLK_c), .D(n6904));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i764_765 (.Q(\mem_REG.mem_7_18 ), .C(SLM_CLK_c), .D(n6903));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i761_762 (.Q(\mem_REG.mem_7_17 ), .C(SLM_CLK_c), .D(n6902));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i758_759 (.Q(\mem_REG.mem_7_16 ), .C(SLM_CLK_c), .D(n6901));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i755_756 (.Q(\mem_REG.mem_7_15 ), .C(SLM_CLK_c), .D(n6900));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i752_753 (.Q(\mem_REG.mem_7_14 ), .C(SLM_CLK_c), .D(n6899));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i749_750 (.Q(\mem_REG.mem_7_13 ), .C(SLM_CLK_c), .D(n6898));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i746_747 (.Q(\mem_REG.mem_7_12 ), .C(SLM_CLK_c), .D(n6897));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i743_744 (.Q(\mem_REG.mem_7_11 ), .C(SLM_CLK_c), .D(n6896));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i740_741 (.Q(\mem_REG.mem_7_10 ), .C(SLM_CLK_c), .D(n6895));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i737_738 (.Q(\mem_REG.mem_7_9 ), .C(SLM_CLK_c), .D(n6894));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i734_735 (.Q(\mem_REG.mem_7_8 ), .C(SLM_CLK_c), .D(n6893));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i731_732 (.Q(\mem_REG.mem_7_7 ), .C(SLM_CLK_c), .D(n6892));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i728_729 (.Q(\mem_REG.mem_7_6 ), .C(SLM_CLK_c), .D(n6891));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i725_726 (.Q(\mem_REG.mem_7_5 ), .C(SLM_CLK_c), .D(n6890));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i722_723 (.Q(\mem_REG.mem_7_4 ), .C(SLM_CLK_c), .D(n6889));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i719_720 (.Q(\mem_REG.mem_7_3 ), .C(SLM_CLK_c), .D(n6888));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i716_717 (.Q(\mem_REG.mem_7_2 ), .C(SLM_CLK_c), .D(n6887));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i713_714 (.Q(\mem_REG.mem_7_1 ), .C(SLM_CLK_c), .D(n6886));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i710_711 (.Q(\mem_REG.mem_7_0 ), .C(SLM_CLK_c), .D(n6885));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i707_708 (.Q(\mem_REG.mem_6_31 ), .C(SLM_CLK_c), .D(n6884));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i704_705 (.Q(\mem_REG.mem_6_30 ), .C(SLM_CLK_c), .D(n6883));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i701_702 (.Q(\mem_REG.mem_6_29 ), .C(SLM_CLK_c), .D(n6882));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i698_699 (.Q(\mem_REG.mem_6_28 ), .C(SLM_CLK_c), .D(n6881));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i695_696 (.Q(\mem_REG.mem_6_27 ), .C(SLM_CLK_c), .D(n6880));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i692_693 (.Q(\mem_REG.mem_6_26 ), .C(SLM_CLK_c), .D(n6879));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i689_690 (.Q(\mem_REG.mem_6_25 ), .C(SLM_CLK_c), .D(n6878));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i686_687 (.Q(\mem_REG.mem_6_24 ), .C(SLM_CLK_c), .D(n6877));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i683_684 (.Q(\mem_REG.mem_6_23 ), .C(SLM_CLK_c), .D(n6876));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i680_681 (.Q(\mem_REG.mem_6_22 ), .C(SLM_CLK_c), .D(n6875));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i677_678 (.Q(\mem_REG.mem_6_21 ), .C(SLM_CLK_c), .D(n6874));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i674_675 (.Q(\mem_REG.mem_6_20 ), .C(SLM_CLK_c), .D(n6873));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i671_672 (.Q(\mem_REG.mem_6_19 ), .C(SLM_CLK_c), .D(n6872));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i668_669 (.Q(\mem_REG.mem_6_18 ), .C(SLM_CLK_c), .D(n6871));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i665_666 (.Q(\mem_REG.mem_6_17 ), .C(SLM_CLK_c), .D(n6870));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i662_663 (.Q(\mem_REG.mem_6_16 ), .C(SLM_CLK_c), .D(n6869));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i659_660 (.Q(\mem_REG.mem_6_15 ), .C(SLM_CLK_c), .D(n6868));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i656_657 (.Q(\mem_REG.mem_6_14 ), .C(SLM_CLK_c), .D(n6867));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i653_654 (.Q(\mem_REG.mem_6_13 ), .C(SLM_CLK_c), .D(n6866));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i650_651 (.Q(\mem_REG.mem_6_12 ), .C(SLM_CLK_c), .D(n6865));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i647_648 (.Q(\mem_REG.mem_6_11 ), .C(SLM_CLK_c), .D(n6864));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i644_645 (.Q(\mem_REG.mem_6_10 ), .C(SLM_CLK_c), .D(n6863));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i641_642 (.Q(\mem_REG.mem_6_9 ), .C(SLM_CLK_c), .D(n6862));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i638_639 (.Q(\mem_REG.mem_6_8 ), .C(SLM_CLK_c), .D(n6861));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i635_636 (.Q(\mem_REG.mem_6_7 ), .C(SLM_CLK_c), .D(n6860));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i632_633 (.Q(\mem_REG.mem_6_6 ), .C(SLM_CLK_c), .D(n6859));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i629_630 (.Q(\mem_REG.mem_6_5 ), .C(SLM_CLK_c), .D(n6858));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i626_627 (.Q(\mem_REG.mem_6_4 ), .C(SLM_CLK_c), .D(n6857));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i623_624 (.Q(\mem_REG.mem_6_3 ), .C(SLM_CLK_c), .D(n6856));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i620_621 (.Q(\mem_REG.mem_6_2 ), .C(SLM_CLK_c), .D(n6855));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i617_618 (.Q(\mem_REG.mem_6_1 ), .C(SLM_CLK_c), .D(n6854));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i614_615 (.Q(\mem_REG.mem_6_0 ), .C(SLM_CLK_c), .D(n6853));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i611_612 (.Q(\mem_REG.mem_5_31 ), .C(SLM_CLK_c), .D(n6852));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i608_609 (.Q(\mem_REG.mem_5_30 ), .C(SLM_CLK_c), .D(n6851));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i605_606 (.Q(\mem_REG.mem_5_29 ), .C(SLM_CLK_c), .D(n6850));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i602_603 (.Q(\mem_REG.mem_5_28 ), .C(SLM_CLK_c), .D(n6849));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i599_600 (.Q(\mem_REG.mem_5_27 ), .C(SLM_CLK_c), .D(n6848));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i596_597 (.Q(\mem_REG.mem_5_26 ), .C(SLM_CLK_c), .D(n6847));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i593_594 (.Q(\mem_REG.mem_5_25 ), .C(SLM_CLK_c), .D(n6846));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i590_591 (.Q(\mem_REG.mem_5_24 ), .C(SLM_CLK_c), .D(n6845));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i587_588 (.Q(\mem_REG.mem_5_23 ), .C(SLM_CLK_c), .D(n6844));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i584_585 (.Q(\mem_REG.mem_5_22 ), .C(SLM_CLK_c), .D(n6843));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i581_582 (.Q(\mem_REG.mem_5_21 ), .C(SLM_CLK_c), .D(n6842));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i578_579 (.Q(\mem_REG.mem_5_20 ), .C(SLM_CLK_c), .D(n6841));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i575_576 (.Q(\mem_REG.mem_5_19 ), .C(SLM_CLK_c), .D(n6840));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i572_573 (.Q(\mem_REG.mem_5_18 ), .C(SLM_CLK_c), .D(n6839));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i569_570 (.Q(\mem_REG.mem_5_17 ), .C(SLM_CLK_c), .D(n6838));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i566_567 (.Q(\mem_REG.mem_5_16 ), .C(SLM_CLK_c), .D(n6837));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i563_564 (.Q(\mem_REG.mem_5_15 ), .C(SLM_CLK_c), .D(n6836));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i560_561 (.Q(\mem_REG.mem_5_14 ), .C(SLM_CLK_c), .D(n6835));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i557_558 (.Q(\mem_REG.mem_5_13 ), .C(SLM_CLK_c), .D(n6834));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i554_555 (.Q(\mem_REG.mem_5_12 ), .C(SLM_CLK_c), .D(n6833));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i551_552 (.Q(\mem_REG.mem_5_11 ), .C(SLM_CLK_c), .D(n6832));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i548_549 (.Q(\mem_REG.mem_5_10 ), .C(SLM_CLK_c), .D(n6831));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i545_546 (.Q(\mem_REG.mem_5_9 ), .C(SLM_CLK_c), .D(n6830));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i542_543 (.Q(\mem_REG.mem_5_8 ), .C(SLM_CLK_c), .D(n6829));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i539_540 (.Q(\mem_REG.mem_5_7 ), .C(SLM_CLK_c), .D(n6828));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i536_537 (.Q(\mem_REG.mem_5_6 ), .C(SLM_CLK_c), .D(n6827));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i533_534 (.Q(\mem_REG.mem_5_5 ), .C(SLM_CLK_c), .D(n6826));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i530_531 (.Q(\mem_REG.mem_5_4 ), .C(SLM_CLK_c), .D(n6825));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i527_528 (.Q(\mem_REG.mem_5_3 ), .C(SLM_CLK_c), .D(n6824));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i524_525 (.Q(\mem_REG.mem_5_2 ), .C(SLM_CLK_c), .D(n6823));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i521_522 (.Q(\mem_REG.mem_5_1 ), .C(SLM_CLK_c), .D(n6822));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i518_519 (.Q(\mem_REG.mem_5_0 ), .C(SLM_CLK_c), .D(n6821));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i515_516 (.Q(\mem_REG.mem_4_31 ), .C(SLM_CLK_c), .D(n6820));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i512_513 (.Q(\mem_REG.mem_4_30 ), .C(SLM_CLK_c), .D(n6819));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i509_510 (.Q(\mem_REG.mem_4_29 ), .C(SLM_CLK_c), .D(n6818));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i506_507 (.Q(\mem_REG.mem_4_28 ), .C(SLM_CLK_c), .D(n6817));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i503_504 (.Q(\mem_REG.mem_4_27 ), .C(SLM_CLK_c), .D(n6816));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i500_501 (.Q(\mem_REG.mem_4_26 ), .C(SLM_CLK_c), .D(n6815));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i497_498 (.Q(\mem_REG.mem_4_25 ), .C(SLM_CLK_c), .D(n6814));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i494_495 (.Q(\mem_REG.mem_4_24 ), .C(SLM_CLK_c), .D(n6813));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i491_492 (.Q(\mem_REG.mem_4_23 ), .C(SLM_CLK_c), .D(n6812));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i488_489 (.Q(\mem_REG.mem_4_22 ), .C(SLM_CLK_c), .D(n6811));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i485_486 (.Q(\mem_REG.mem_4_21 ), .C(SLM_CLK_c), .D(n6810));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i482_483 (.Q(\mem_REG.mem_4_20 ), .C(SLM_CLK_c), .D(n6809));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i479_480 (.Q(\mem_REG.mem_4_19 ), .C(SLM_CLK_c), .D(n6808));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i476_477 (.Q(\mem_REG.mem_4_18 ), .C(SLM_CLK_c), .D(n6807));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i473_474 (.Q(\mem_REG.mem_4_17 ), .C(SLM_CLK_c), .D(n6806));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i470_471 (.Q(\mem_REG.mem_4_16 ), .C(SLM_CLK_c), .D(n6805));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i467_468 (.Q(\mem_REG.mem_4_15 ), .C(SLM_CLK_c), .D(n6804));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i464_465 (.Q(\mem_REG.mem_4_14 ), .C(SLM_CLK_c), .D(n6803));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i461_462 (.Q(\mem_REG.mem_4_13 ), .C(SLM_CLK_c), .D(n6802));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i458_459 (.Q(\mem_REG.mem_4_12 ), .C(SLM_CLK_c), .D(n6801));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i455_456 (.Q(\mem_REG.mem_4_11 ), .C(SLM_CLK_c), .D(n6800));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i452_453 (.Q(\mem_REG.mem_4_10 ), .C(SLM_CLK_c), .D(n6799));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i449_450 (.Q(\mem_REG.mem_4_9 ), .C(SLM_CLK_c), .D(n6798));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i446_447 (.Q(\mem_REG.mem_4_8 ), .C(SLM_CLK_c), .D(n6797));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i443_444 (.Q(\mem_REG.mem_4_7 ), .C(SLM_CLK_c), .D(n6796));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i440_441 (.Q(\mem_REG.mem_4_6 ), .C(SLM_CLK_c), .D(n6795));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i437_438 (.Q(\mem_REG.mem_4_5 ), .C(SLM_CLK_c), .D(n6794));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i434_435 (.Q(\mem_REG.mem_4_4 ), .C(SLM_CLK_c), .D(n6793));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i431_432 (.Q(\mem_REG.mem_4_3 ), .C(SLM_CLK_c), .D(n6792));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i428_429 (.Q(\mem_REG.mem_4_2 ), .C(SLM_CLK_c), .D(n6791));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i425_426 (.Q(\mem_REG.mem_4_1 ), .C(SLM_CLK_c), .D(n6790));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i422_423 (.Q(\mem_REG.mem_4_0 ), .C(SLM_CLK_c), .D(n6789));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i419_420 (.Q(\mem_REG.mem_3_31 ), .C(SLM_CLK_c), .D(n6788));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i416_417 (.Q(\mem_REG.mem_3_30 ), .C(SLM_CLK_c), .D(n6787));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i413_414 (.Q(\mem_REG.mem_3_29 ), .C(SLM_CLK_c), .D(n6786));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i410_411 (.Q(\mem_REG.mem_3_28 ), .C(SLM_CLK_c), .D(n6785));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i407_408 (.Q(\mem_REG.mem_3_27 ), .C(SLM_CLK_c), .D(n6784));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i404_405 (.Q(\mem_REG.mem_3_26 ), .C(SLM_CLK_c), .D(n6783));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i401_402 (.Q(\mem_REG.mem_3_25 ), .C(SLM_CLK_c), .D(n6782));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i398_399 (.Q(\mem_REG.mem_3_24 ), .C(SLM_CLK_c), .D(n6781));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i395_396 (.Q(\mem_REG.mem_3_23 ), .C(SLM_CLK_c), .D(n6780));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i392_393 (.Q(\mem_REG.mem_3_22 ), .C(SLM_CLK_c), .D(n6779));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i389_390 (.Q(\mem_REG.mem_3_21 ), .C(SLM_CLK_c), .D(n6778));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i386_387 (.Q(\mem_REG.mem_3_20 ), .C(SLM_CLK_c), .D(n6777));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i383_384 (.Q(\mem_REG.mem_3_19 ), .C(SLM_CLK_c), .D(n6776));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i380_381 (.Q(\mem_REG.mem_3_18 ), .C(SLM_CLK_c), .D(n6775));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i377_378 (.Q(\mem_REG.mem_3_17 ), .C(SLM_CLK_c), .D(n6774));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i374_375 (.Q(\mem_REG.mem_3_16 ), .C(SLM_CLK_c), .D(n6773));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i371_372 (.Q(\mem_REG.mem_3_15 ), .C(SLM_CLK_c), .D(n6772));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i368_369 (.Q(\mem_REG.mem_3_14 ), .C(SLM_CLK_c), .D(n6771));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i365_366 (.Q(\mem_REG.mem_3_13 ), .C(SLM_CLK_c), .D(n6770));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i362_363 (.Q(\mem_REG.mem_3_12 ), .C(SLM_CLK_c), .D(n6769));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i359_360 (.Q(\mem_REG.mem_3_11 ), .C(SLM_CLK_c), .D(n6768));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i356_357 (.Q(\mem_REG.mem_3_10 ), .C(SLM_CLK_c), .D(n6767));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i353_354 (.Q(\mem_REG.mem_3_9 ), .C(SLM_CLK_c), .D(n6766));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i350_351 (.Q(\mem_REG.mem_3_8 ), .C(SLM_CLK_c), .D(n6765));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i347_348 (.Q(\mem_REG.mem_3_7 ), .C(SLM_CLK_c), .D(n6764));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i344_345 (.Q(\mem_REG.mem_3_6 ), .C(SLM_CLK_c), .D(n6763));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i341_342 (.Q(\mem_REG.mem_3_5 ), .C(SLM_CLK_c), .D(n6762));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i338_339 (.Q(\mem_REG.mem_3_4 ), .C(SLM_CLK_c), .D(n6761));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i335_336 (.Q(\mem_REG.mem_3_3 ), .C(SLM_CLK_c), .D(n6760));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i332_333 (.Q(\mem_REG.mem_3_2 ), .C(SLM_CLK_c), .D(n6759));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i329_330 (.Q(\mem_REG.mem_3_1 ), .C(SLM_CLK_c), .D(n6758));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i326_327 (.Q(\mem_REG.mem_3_0 ), .C(SLM_CLK_c), .D(n6757));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i323_324 (.Q(\mem_REG.mem_2_31 ), .C(SLM_CLK_c), .D(n6756));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i320_321 (.Q(\mem_REG.mem_2_30 ), .C(SLM_CLK_c), .D(n6755));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i317_318 (.Q(\mem_REG.mem_2_29 ), .C(SLM_CLK_c), .D(n6754));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i314_315 (.Q(\mem_REG.mem_2_28 ), .C(SLM_CLK_c), .D(n6753));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i311_312 (.Q(\mem_REG.mem_2_27 ), .C(SLM_CLK_c), .D(n6752));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i308_309 (.Q(\mem_REG.mem_2_26 ), .C(SLM_CLK_c), .D(n6751));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i305_306 (.Q(\mem_REG.mem_2_25 ), .C(SLM_CLK_c), .D(n6750));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i302_303 (.Q(\mem_REG.mem_2_24 ), .C(SLM_CLK_c), .D(n6749));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i299_300 (.Q(\mem_REG.mem_2_23 ), .C(SLM_CLK_c), .D(n6748));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i296_297 (.Q(\mem_REG.mem_2_22 ), .C(SLM_CLK_c), .D(n6747));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i293_294 (.Q(\mem_REG.mem_2_21 ), .C(SLM_CLK_c), .D(n6746));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i290_291 (.Q(\mem_REG.mem_2_20 ), .C(SLM_CLK_c), .D(n6745));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i287_288 (.Q(\mem_REG.mem_2_19 ), .C(SLM_CLK_c), .D(n6744));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i284_285 (.Q(\mem_REG.mem_2_18 ), .C(SLM_CLK_c), .D(n6743));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i281_282 (.Q(\mem_REG.mem_2_17 ), .C(SLM_CLK_c), .D(n6742));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i278_279 (.Q(\mem_REG.mem_2_16 ), .C(SLM_CLK_c), .D(n6741));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i275_276 (.Q(\mem_REG.mem_2_15 ), .C(SLM_CLK_c), .D(n6740));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i272_273 (.Q(\mem_REG.mem_2_14 ), .C(SLM_CLK_c), .D(n6739));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i269_270 (.Q(\mem_REG.mem_2_13 ), .C(SLM_CLK_c), .D(n6738));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i266_267 (.Q(\mem_REG.mem_2_12 ), .C(SLM_CLK_c), .D(n6737));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i263_264 (.Q(\mem_REG.mem_2_11 ), .C(SLM_CLK_c), .D(n6736));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i260_261 (.Q(\mem_REG.mem_2_10 ), .C(SLM_CLK_c), .D(n6735));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i257_258 (.Q(\mem_REG.mem_2_9 ), .C(SLM_CLK_c), .D(n6734));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i254_255 (.Q(\mem_REG.mem_2_8 ), .C(SLM_CLK_c), .D(n6733));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i251_252 (.Q(\mem_REG.mem_2_7 ), .C(SLM_CLK_c), .D(n6732));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i248_249 (.Q(\mem_REG.mem_2_6 ), .C(SLM_CLK_c), .D(n6731));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i245_246 (.Q(\mem_REG.mem_2_5 ), .C(SLM_CLK_c), .D(n6730));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i242_243 (.Q(\mem_REG.mem_2_4 ), .C(SLM_CLK_c), .D(n6729));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i239_240 (.Q(\mem_REG.mem_2_3 ), .C(SLM_CLK_c), .D(n6728));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i236_237 (.Q(\mem_REG.mem_2_2 ), .C(SLM_CLK_c), .D(n6727));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i233_234 (.Q(\mem_REG.mem_2_1 ), .C(SLM_CLK_c), .D(n6726));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i230_231 (.Q(\mem_REG.mem_2_0 ), .C(SLM_CLK_c), .D(n6725));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i227_228 (.Q(\mem_REG.mem_1_31 ), .C(SLM_CLK_c), .D(n6724));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i224_225 (.Q(\mem_REG.mem_1_30 ), .C(SLM_CLK_c), .D(n6723));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i221_222 (.Q(\mem_REG.mem_1_29 ), .C(SLM_CLK_c), .D(n6722));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i218_219 (.Q(\mem_REG.mem_1_28 ), .C(SLM_CLK_c), .D(n6721));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i215_216 (.Q(\mem_REG.mem_1_27 ), .C(SLM_CLK_c), .D(n6720));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i212_213 (.Q(\mem_REG.mem_1_26 ), .C(SLM_CLK_c), .D(n6719));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i209_210 (.Q(\mem_REG.mem_1_25 ), .C(SLM_CLK_c), .D(n6718));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i206_207 (.Q(\mem_REG.mem_1_24 ), .C(SLM_CLK_c), .D(n6717));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i203_204 (.Q(\mem_REG.mem_1_23 ), .C(SLM_CLK_c), .D(n6716));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i200_201 (.Q(\mem_REG.mem_1_22 ), .C(SLM_CLK_c), .D(n6715));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i197_198 (.Q(\mem_REG.mem_1_21 ), .C(SLM_CLK_c), .D(n6714));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i194_195 (.Q(\mem_REG.mem_1_20 ), .C(SLM_CLK_c), .D(n6713));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i191_192 (.Q(\mem_REG.mem_1_19 ), .C(SLM_CLK_c), .D(n6712));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i188_189 (.Q(\mem_REG.mem_1_18 ), .C(SLM_CLK_c), .D(n6711));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i185_186 (.Q(\mem_REG.mem_1_17 ), .C(SLM_CLK_c), .D(n6710));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i182_183 (.Q(\mem_REG.mem_1_16 ), .C(SLM_CLK_c), .D(n6709));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i179_180 (.Q(\mem_REG.mem_1_15 ), .C(SLM_CLK_c), .D(n6708));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i176_177 (.Q(\mem_REG.mem_1_14 ), .C(SLM_CLK_c), .D(n6707));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i173_174 (.Q(\mem_REG.mem_1_13 ), .C(SLM_CLK_c), .D(n6706));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i170_171 (.Q(\mem_REG.mem_1_12 ), .C(SLM_CLK_c), .D(n6705));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i167_168 (.Q(\mem_REG.mem_1_11 ), .C(SLM_CLK_c), .D(n6704));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i164_165 (.Q(\mem_REG.mem_1_10 ), .C(SLM_CLK_c), .D(n6703));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i161_162 (.Q(\mem_REG.mem_1_9 ), .C(SLM_CLK_c), .D(n6702));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i158_159 (.Q(\mem_REG.mem_1_8 ), .C(SLM_CLK_c), .D(n6701));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i155_156 (.Q(\mem_REG.mem_1_7 ), .C(SLM_CLK_c), .D(n6700));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i152_153 (.Q(\mem_REG.mem_1_6 ), .C(SLM_CLK_c), .D(n6699));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i149_150 (.Q(\mem_REG.mem_1_5 ), .C(SLM_CLK_c), .D(n6698));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i146_147 (.Q(\mem_REG.mem_1_4 ), .C(SLM_CLK_c), .D(n6697));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i143_144 (.Q(\mem_REG.mem_1_3 ), .C(SLM_CLK_c), .D(n6696));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i140_141 (.Q(\mem_REG.mem_1_2 ), .C(SLM_CLK_c), .D(n6695));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i137_138 (.Q(\mem_REG.mem_1_1 ), .C(SLM_CLK_c), .D(n6694));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i134_135 (.Q(\mem_REG.mem_1_0 ), .C(SLM_CLK_c), .D(n6693));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i131_132 (.Q(\mem_REG.mem_0_31 ), .C(SLM_CLK_c), .D(n6692));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i128_129 (.Q(\mem_REG.mem_0_30 ), .C(SLM_CLK_c), .D(n6691));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i125_126 (.Q(\mem_REG.mem_0_29 ), .C(SLM_CLK_c), .D(n6690));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i122_123 (.Q(\mem_REG.mem_0_28 ), .C(SLM_CLK_c), .D(n6689));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i119_120 (.Q(\mem_REG.mem_0_27 ), .C(SLM_CLK_c), .D(n6688));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i116_117 (.Q(\mem_REG.mem_0_26 ), .C(SLM_CLK_c), .D(n6687));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i113_114 (.Q(\mem_REG.mem_0_25 ), .C(SLM_CLK_c), .D(n6686));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i110_111 (.Q(\mem_REG.mem_0_24 ), .C(SLM_CLK_c), .D(n6685));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i107_108 (.Q(\mem_REG.mem_0_23 ), .C(SLM_CLK_c), .D(n6684));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i104_105 (.Q(\mem_REG.mem_0_22 ), .C(SLM_CLK_c), .D(n6683));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i101_102 (.Q(\mem_REG.mem_0_21 ), .C(SLM_CLK_c), .D(n6682));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i98_99 (.Q(\mem_REG.mem_0_20 ), .C(SLM_CLK_c), .D(n6681));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i95_96 (.Q(\mem_REG.mem_0_19 ), .C(SLM_CLK_c), .D(n6680));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i92_93 (.Q(\mem_REG.mem_0_18 ), .C(SLM_CLK_c), .D(n6679));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i89_90 (.Q(\mem_REG.mem_0_17 ), .C(SLM_CLK_c), .D(n6678));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i86_87 (.Q(\mem_REG.mem_0_16 ), .C(SLM_CLK_c), .D(n6677));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i83_84 (.Q(\mem_REG.mem_0_15 ), .C(SLM_CLK_c), .D(n6676));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i80_81 (.Q(\mem_REG.mem_0_14 ), .C(SLM_CLK_c), .D(n6675));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i77_78 (.Q(\mem_REG.mem_0_13 ), .C(SLM_CLK_c), .D(n6674));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i74_75 (.Q(\mem_REG.mem_0_12 ), .C(SLM_CLK_c), .D(n6673));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i71_72 (.Q(\mem_REG.mem_0_11 ), .C(SLM_CLK_c), .D(n6672));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i68_69 (.Q(\mem_REG.mem_0_10 ), .C(SLM_CLK_c), .D(n6671));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i65_66 (.Q(\mem_REG.mem_0_9 ), .C(SLM_CLK_c), .D(n6670));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i62_63 (.Q(\mem_REG.mem_0_8 ), .C(SLM_CLK_c), .D(n6669));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i59_60 (.Q(\mem_REG.mem_0_7 ), .C(SLM_CLK_c), .D(n6668));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i56_57 (.Q(\mem_REG.mem_0_6 ), .C(SLM_CLK_c), .D(n6667));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i53_54 (.Q(\mem_REG.mem_0_5 ), .C(SLM_CLK_c), .D(n6666));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i50_51 (.Q(\mem_REG.mem_0_4 ), .C(SLM_CLK_c), .D(n6665));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i47_48 (.Q(\mem_REG.mem_0_3 ), .C(SLM_CLK_c), .D(n6664));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i44_45 (.Q(\mem_REG.mem_0_2 ), .C(SLM_CLK_c), .D(n6663));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i41_42 (.Q(\mem_REG.mem_0_1 ), .C(SLM_CLK_c), .D(n6662));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_DFF i38_39 (.Q(\mem_REG.mem_0_0 ), .C(SLM_CLK_c), .D(n6661));   // src/fifo_sc_32_lut_gen.v(604[73:76])
    SB_LUT4 i5414_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[28]), 
            .I3(\mem_REG.mem_7_28 ), .O(n6913));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5414_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14758 (.I0(rd_addr_r[1]), .I1(n15477), 
            .I2(n15478), .I3(rd_addr_r[2]), .O(n16977));
    defparam rd_addr_r_1__bdd_4_lut_14758.LUT_INIT = 16'he4aa;
    SB_LUT4 n16977_bdd_4_lut (.I0(n16977), .I1(n15466), .I2(n15465), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[19]));
    defparam n16977_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3895_1_lut (.I0(sc32_fifo_data_out[24]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5394));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3895_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3896_1_lut (.I0(sc32_fifo_data_out[23]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5395));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3896_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3897_1_lut (.I0(sc32_fifo_data_out[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5396));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3897_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5413_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[27]), 
            .I3(\mem_REG.mem_7_27 ), .O(n6912));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5413_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5412_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[26]), 
            .I3(\mem_REG.mem_7_26 ), .O(n6911));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5412_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5411_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[25]), 
            .I3(\mem_REG.mem_7_25 ), .O(n6910));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5411_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5410_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[24]), 
            .I3(\mem_REG.mem_7_24 ), .O(n6909));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5410_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3898_1_lut (.I0(sc32_fifo_data_out[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5397));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3898_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3899_1_lut (.I0(sc32_fifo_data_out[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5398));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3899_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5409_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[23]), 
            .I3(\mem_REG.mem_7_23 ), .O(n6908));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5409_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3900_1_lut (.I0(sc32_fifo_data_out[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5399));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3900_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3901_1_lut (.I0(sc32_fifo_data_out[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5400));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3901_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3902_1_lut (.I0(sc32_fifo_data_out[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5401));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3902_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_15427  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_2 ), .I2(\mem_REG.mem_3_2 ), .I3(rd_addr_r[1]), 
            .O(n17637));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_15427 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17637_bdd_4_lut (.I0(n17637), .I1(\mem_REG.mem_1_2 ), .I2(\mem_REG.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(n17640));
    defparam n17637_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5408_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[22]), 
            .I3(\mem_REG.mem_7_22 ), .O(n6907));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5408_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5407_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[21]), 
            .I3(\mem_REG.mem_7_21 ), .O(n6906));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5407_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13341_3_lut (.I0(\mem_REG.mem_0_19 ), .I1(\mem_REG.mem_1_19 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15465));
    defparam i13341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13342_3_lut (.I0(\mem_REG.mem_2_19 ), .I1(\mem_REG.mem_3_19 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15466));
    defparam i13342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5406_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[20]), 
            .I3(\mem_REG.mem_7_20 ), .O(n6905));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5406_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13431_3_lut (.I0(\mem_REG.mem_0_23 ), .I1(\mem_REG.mem_1_23 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15555));
    defparam i13431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3903_1_lut (.I0(sc32_fifo_data_out[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5402));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3903_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3904_1_lut (.I0(sc32_fifo_data_out[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5403));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3904_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13354_3_lut (.I0(\mem_REG.mem_6_19 ), .I1(\mem_REG.mem_7_19 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15478));
    defparam i13354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13353_3_lut (.I0(\mem_REG.mem_4_19 ), .I1(\mem_REG.mem_5_19 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15477));
    defparam i13353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut (.I0(rd_addr_r[1]), .I1(n15597), .I2(n15598), 
            .I3(rd_addr_r[2]), .O(n17577));
    defparam rd_addr_r_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n17577_bdd_4_lut (.I0(n17577), .I1(n15586), .I2(n15585), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[24]));
    defparam n17577_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3905_1_lut (.I0(sc32_fifo_data_out[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5404));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3905_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13432_3_lut (.I0(\mem_REG.mem_2_23 ), .I1(\mem_REG.mem_3_23 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15556));
    defparam i13432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14713 (.I0(rd_addr_r[1]), .I1(n15267), 
            .I2(n15268), .I3(rd_addr_r[2]), .O(n16881));
    defparam rd_addr_r_1__bdd_4_lut_14713.LUT_INIT = 16'he4aa;
    SB_LUT4 n16881_bdd_4_lut (.I0(n16881), .I1(n15247), .I2(n15246), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[13]));
    defparam n16881_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2407_3_lut_4_lut (.I0(sc32_fifo_write_enable), .I1(\MISC.full_flag_r ), 
            .I2(\MISC.rd_w ), .I3(n2495), .O(n3894));   // src/fifo_sc_32_lut_gen.v(268[25:51])
    defparam i2407_3_lut_4_lut.LUT_INIT = 16'h00d2;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14633 (.I0(rd_addr_r[1]), .I1(n15756), 
            .I2(n15757), .I3(rd_addr_r[2]), .O(n16875));
    defparam rd_addr_r_1__bdd_4_lut_14633.LUT_INIT = 16'he4aa;
    SB_LUT4 n16875_bdd_4_lut (.I0(n16875), .I1(n15748), .I2(n15747), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[30]));
    defparam n16875_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_15262  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_2 ), .I2(\mem_REG.mem_7_2 ), .I3(rd_addr_r[1]), 
            .O(n17547));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_15262 .LUT_INIT = 16'he4aa;
    SB_LUT4 i3906_1_lut (.I0(sc32_fifo_data_out[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5405));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3906_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 wr_addr_r_3__I_0_i4_3_lut_4_lut (.I0(sc32_fifo_write_enable), 
            .I1(\MISC.full_flag_r ), .I2(wr_addr_p1_r[3]), .I3(wr_addr_r[3]), 
            .O(wr_addr_nxt_w[3]));   // src/fifo_sc_32_lut_gen.v(268[25:51])
    defparam wr_addr_r_3__I_0_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3907_1_lut (.I0(sc32_fifo_data_out[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5406));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3907_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3908_1_lut (.I0(sc32_fifo_data_out[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5407));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3909_1_lut (.I0(sc32_fifo_data_out[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5408));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3909_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n17547_bdd_4_lut (.I0(n17547), .I1(\mem_REG.mem_5_2 ), .I2(\mem_REG.mem_4_2 ), 
            .I3(rd_addr_r[1]), .O(n17550));
    defparam n17547_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_r_3__I_0_i3_3_lut_4_lut (.I0(sc32_fifo_write_enable), 
            .I1(\MISC.full_flag_r ), .I2(wr_cmpaddr_p1_r[2]), .I3(wr_addr_r[2]), 
            .O(wr_addr_nxt_w[2]));   // src/fifo_sc_32_lut_gen.v(268[25:51])
    defparam wr_addr_r_3__I_0_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14628 (.I0(rd_addr_r[1]), .I1(n15435), 
            .I2(n15436), .I3(rd_addr_r[2]), .O(n16851));
    defparam rd_addr_r_1__bdd_4_lut_14628.LUT_INIT = 16'he4aa;
    SB_LUT4 i13269_3_lut (.I0(\mem_REG.mem_0_0 ), .I1(\mem_REG.mem_1_0 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15393));
    defparam i13269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13270_3_lut (.I0(\mem_REG.mem_2_0 ), .I1(\mem_REG.mem_3_0 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15394));
    defparam i13270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13273_3_lut (.I0(\mem_REG.mem_6_0 ), .I1(\mem_REG.mem_7_0 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15397));
    defparam i13273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n16851_bdd_4_lut (.I0(n16851), .I1(n15217), .I2(n15216), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[12]));
    defparam n16851_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13272_3_lut (.I0(\mem_REG.mem_4_0 ), .I1(\mem_REG.mem_5_0 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15396));
    defparam i13272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15212 (.I0(rd_addr_r[1]), .I1(n15573), 
            .I2(n15574), .I3(rd_addr_r[2]), .O(n17535));
    defparam rd_addr_r_1__bdd_4_lut_15212.LUT_INIT = 16'he4aa;
    SB_LUT4 n17535_bdd_4_lut (.I0(n17535), .I1(n15556), .I2(n15555), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[23]));
    defparam n17535_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12533_3_lut_4_lut (.I0(sc32_fifo_write_enable), .I1(\MISC.full_flag_r ), 
            .I2(\MISC.wr_flag_addr_r [0]), .I3(\MISC.rd_flag_addr_p1_r [0]), 
            .O(n14655));   // src/fifo_sc_32_lut_gen.v(268[25:51])
    defparam i12533_3_lut_4_lut.LUT_INIT = 16'h2ff2;
    SB_LUT4 wr_addr_r_3__I_0_i2_3_lut_4_lut (.I0(sc32_fifo_write_enable), 
            .I1(\MISC.full_flag_r ), .I2(wr_cmpaddr_p1_r[1]), .I3(wr_addr_r[1]), 
            .O(wr_addr_nxt_w[1]));   // src/fifo_sc_32_lut_gen.v(268[25:51])
    defparam wr_addr_r_3__I_0_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i9_2_lut_3_lut_4_lut (.I0(sc32_fifo_write_enable), 
            .I1(\MISC.full_flag_r ), .I2(wr_addr_r[1]), .I3(\MISC.wr_flag_addr_r [0]), 
            .O(n9));   // src/fifo_sc_32_lut_gen.v(268[25:51])
    defparam EnabledDecoder_2_i9_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 wr_addr_r_3__I_0_i1_3_lut_4_lut (.I0(sc32_fifo_write_enable), 
            .I1(\MISC.full_flag_r ), .I2(\MISC.wr_flag_addr_p1_r [0]), .I3(\MISC.wr_flag_addr_r [0]), 
            .O(wr_addr_nxt_w[0]));   // src/fifo_sc_32_lut_gen.v(268[25:51])
    defparam wr_addr_r_3__I_0_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5405_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[19]), 
            .I3(\mem_REG.mem_7_19 ), .O(n6904));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5405_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i8_2_lut_3_lut_4_lut (.I0(sc32_fifo_write_enable), 
            .I1(\MISC.full_flag_r ), .I2(wr_addr_r[1]), .I3(\MISC.wr_flag_addr_r [0]), 
            .O(n8));   // src/fifo_sc_32_lut_gen.v(268[25:51])
    defparam EnabledDecoder_2_i8_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i5404_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[18]), 
            .I3(\mem_REG.mem_7_18 ), .O(n6903));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5404_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5403_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[17]), 
            .I3(\mem_REG.mem_7_17 ), .O(n6902));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5403_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3910_1_lut (.I0(sc32_fifo_data_out[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5409));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3910_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE \mem_REG.data_raw_r_i0_i1  (.Q(sc32_fifo_data_out[1]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[1]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_LUT4 i13284_3_lut (.I0(\mem_REG.mem_0_17 ), .I1(\mem_REG.mem_1_17 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15408));
    defparam i13284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13285_3_lut (.I0(\mem_REG.mem_2_17 ), .I1(\mem_REG.mem_3_17 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15409));
    defparam i13285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13306_3_lut (.I0(\mem_REG.mem_6_17 ), .I1(\mem_REG.mem_7_17 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15430));
    defparam i13306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13305_3_lut (.I0(\mem_REG.mem_4_17 ), .I1(\mem_REG.mem_5_17 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15429));
    defparam i13305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3911_1_lut (.I0(sc32_fifo_data_out[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5410));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3911_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5402_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[16]), 
            .I3(\mem_REG.mem_7_16 ), .O(n6901));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5402_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14608 (.I0(rd_addr_r[1]), .I1(n15186), 
            .I2(n15187), .I3(rd_addr_r[2]), .O(n16815));
    defparam rd_addr_r_1__bdd_4_lut_14608.LUT_INIT = 16'he4aa;
    SB_LUT4 i5401_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[15]), 
            .I3(\mem_REG.mem_7_15 ), .O(n6900));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5401_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16815_bdd_4_lut (.I0(n16815), .I1(n15157), .I2(n15156), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[11]));
    defparam n16815_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5400_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[14]), 
            .I3(\mem_REG.mem_7_14 ), .O(n6899));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5400_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_15187  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_3 ), .I2(\mem_REG.mem_3_3 ), .I3(rd_addr_r[1]), 
            .O(n17487));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_15187 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17487_bdd_4_lut (.I0(n17487), .I1(\mem_REG.mem_1_3 ), .I2(\mem_REG.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(n17490));
    defparam n17487_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \mem_REG.data_raw_r_i0_i2  (.Q(sc32_fifo_data_out[2]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[2]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i3  (.Q(sc32_fifo_data_out[3]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[3]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i4  (.Q(sc32_fifo_data_out[4]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[4]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i5  (.Q(sc32_fifo_data_out[5]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[5]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i6  (.Q(sc32_fifo_data_out[6]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[6]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i7  (.Q(sc32_fifo_data_out[7]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[7]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i8  (.Q(sc32_fifo_data_out[8]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[8]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i9  (.Q(sc32_fifo_data_out[9]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[9]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i10  (.Q(sc32_fifo_data_out[10]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[10]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i11  (.Q(sc32_fifo_data_out[11]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[11]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i12  (.Q(sc32_fifo_data_out[12]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[12]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i13  (.Q(sc32_fifo_data_out[13]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[13]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i14  (.Q(sc32_fifo_data_out[14]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[14]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i15  (.Q(sc32_fifo_data_out[15]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[15]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i16  (.Q(sc32_fifo_data_out[16]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[16]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i17  (.Q(sc32_fifo_data_out[17]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[17]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i18  (.Q(sc32_fifo_data_out[18]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[18]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i19  (.Q(sc32_fifo_data_out[19]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[19]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i20  (.Q(sc32_fifo_data_out[20]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[20]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i21  (.Q(sc32_fifo_data_out[21]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[21]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i22  (.Q(sc32_fifo_data_out[22]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[22]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i23  (.Q(sc32_fifo_data_out[23]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[23]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i24  (.Q(sc32_fifo_data_out[24]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[24]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i25  (.Q(sc32_fifo_data_out[25]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[25]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i26  (.Q(sc32_fifo_data_out[26]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[26]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i27  (.Q(sc32_fifo_data_out[27]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[27]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i28  (.Q(sc32_fifo_data_out[28]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[28]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i29  (.Q(sc32_fifo_data_out[29]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[29]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i30  (.Q(sc32_fifo_data_out[30]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[30]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_DFFE \mem_REG.data_raw_r_i0_i31  (.Q(sc32_fifo_data_out[31]), .C(SLM_CLK_c), 
            .E(\MISC.rd_w ), .D(rd_data_o_31__N_759[31]));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    SB_LUT4 i13450_3_lut (.I0(\mem_REG.mem_6_23 ), .I1(\mem_REG.mem_7_23 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15574));
    defparam i13450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13449_3_lut (.I0(\mem_REG.mem_4_23 ), .I1(\mem_REG.mem_5_23 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15573));
    defparam i13449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1458_i3_3_lut (.I0(wr_addr_r[2]), .I1(wr_cmpaddr_p1_r[2]), 
            .I2(n2495), .I3(GND_net), .O(n2834[2]));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam mux_1458_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2410_3_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1cmp_r[2]), .I2(n3894), 
            .I3(GND_net), .O(n3457));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i2410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15177 (.I0(rd_addr_r[1]), .I1(n15549), 
            .I2(n15550), .I3(rd_addr_r[2]), .O(n17469));
    defparam rd_addr_r_1__bdd_4_lut_15177.LUT_INIT = 16'he4aa;
    SB_LUT4 n17469_bdd_4_lut (.I0(n17469), .I1(n15403), .I2(n15402), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[1]));
    defparam n17469_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5399_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[13]), 
            .I3(\mem_REG.mem_7_13 ), .O(n6898));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5399_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1787_3_lut (.I0(n2834[1]), .I1(n3455), .I2(n2), .I3(GND_net), 
            .O(n4));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i1787_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i5398_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[12]), 
            .I3(\mem_REG.mem_7_12 ), .O(n6897));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5398_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF wr_addr_r_i1 (.Q(wr_addr_r[1]), .C(SLM_CLK_c), .D(wr_addr_r_3__N_690[1]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_addr_r_i2 (.Q(wr_addr_r[2]), .C(SLM_CLK_c), .D(wr_addr_r_3__N_690[2]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_addr_r_i3 (.Q(wr_addr_r[3]), .C(SLM_CLK_c), .D(wr_addr_r_3__N_690[3]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_addr_p1_r_i3 (.Q(wr_addr_p1_r[3]), .C(SLM_CLK_c), .D(wr_addr_p1cmp_r_3__N_698[3]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_cmpaddr_p1_r_i1 (.Q(wr_cmpaddr_p1_r[1]), .C(SLM_CLK_c), .D(wr_addr_p1_r_3__N_694[1]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF wr_cmpaddr_p1_r_i2 (.Q(wr_cmpaddr_p1_r[2]), .C(SLM_CLK_c), .D(wr_addr_p1_r_3__N_694[2]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_r_i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(rd_addr_r_3__N_708[1]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_r_i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .D(rd_addr_r_3__N_708[2]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_r_i3 (.Q(rd_addr_r[3]), .C(SLM_CLK_c), .D(rd_addr_r_3__N_708[3]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_p1cmp_r_i1 (.Q(rd_addr_p1cmp_r[1]), .C(SLM_CLK_c), .D(rd_addr_p1_r_3__N_712[1]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_p1cmp_r_i2 (.Q(rd_addr_p1cmp_r[2]), .C(SLM_CLK_c), .D(rd_addr_p1_r_3__N_712[2]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_DFF rd_addr_p1cmp_r_i3 (.Q(rd_addr_p1cmp_r[3]), .C(SLM_CLK_c), .D(rd_addr_p1_r_3__N_712[3]));   // src/fifo_sc_32_lut_gen.v(146[17] 196[20])
    SB_LUT4 mux_1458_i2_3_lut (.I0(wr_addr_r[1]), .I1(wr_cmpaddr_p1_r[1]), 
            .I2(n2495), .I3(GND_net), .O(n2834[1]));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam mux_1458_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2408_3_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1cmp_r[1]), .I2(n3894), 
            .I3(GND_net), .O(n3455));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i2408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2092_3_lut (.I0(\MISC.rd_flag_addr_r [0]), .I1(\MISC.rd_flag_addr_p1_r [0]), 
            .I2(n3894), .I3(GND_net), .O(n3441));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i2092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1779_4_lut (.I0(\MISC.wr_flag_addr_r [0]), .I1(n3441), .I2(\MISC.wr_flag_addr_p1_r [0]), 
            .I3(n2495), .O(n2));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i1779_4_lut.LUT_INIT = 16'hf3bb;
    SB_LUT4 mux_1458_i4_3_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_r[3]), 
            .I2(n2495), .I3(GND_net), .O(n2834[3]));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam mux_1458_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(n2), .I1(n3455), .I2(n2834[1]), .I3(GND_net), 
            .O(n13892));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut (.I0(rd_addr_r[3]), .I1(n2834[3]), .I2(rd_addr_p1cmp_r[3]), 
            .I3(n3894), .O(n4_adj_1397));
    defparam i1_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i2_3_lut_adj_96 (.I0(n4), .I1(n3457), .I2(n2834[2]), .I3(GND_net), 
            .O(n13894));
    defparam i2_3_lut_adj_96.LUT_INIT = 16'h9696;
    SB_LUT4 i5397_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[11]), 
            .I3(\mem_REG.mem_7_11 ), .O(n6896));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5397_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1794_3_lut (.I0(n2834[2]), .I1(n3457), .I2(n4), .I3(GND_net), 
            .O(n6));   // src/fifo_sc_32_lut_gen.v(270[45:108])
    defparam i1794_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i2_4_lut (.I0(n6), .I1(n13894), .I2(n4_adj_1397), .I3(n13892), 
            .O(\MISC.AEmpty.almost_empty_nxt_w ));
    defparam i2_4_lut.LUT_INIT = 16'h4800;
    SB_LUT4 i5396_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[10]), 
            .I3(\mem_REG.mem_7_10 ), .O(n6895));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5396_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_15137  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_25 ), .I2(\mem_REG.mem_3_25 ), .I3(rd_addr_r[1]), 
            .O(n17427));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_15137 .LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14578 (.I0(rd_addr_r[1]), .I1(n15447), 
            .I2(n15448), .I3(rd_addr_r[2]), .O(n16725));
    defparam rd_addr_r_1__bdd_4_lut_14578.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut (.I0(rd_addr_p1cmp_r[1]), .I1(n14655), .I2(\MISC.rd_w ), 
            .I3(wr_addr_r[1]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h2010;
    SB_LUT4 i2_3_lut_adj_97 (.I0(\MISC.empty_flag_r ), .I1(sc32_fifo_write_enable), 
            .I2(full_nxt_w_N_812), .I3(GND_net), .O(empty_nxt_w_N_823));
    defparam i2_3_lut_adj_97.LUT_INIT = 16'h0202;
    SB_LUT4 i12531_4_lut (.I0(rd_addr_p1cmp_r[3]), .I1(rd_addr_p1cmp_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n14653));
    defparam i12531_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_98 (.I0(reset_all), .I1(n14653), .I2(empty_nxt_w_N_823), 
            .I3(n10), .O(empty_ext_r_N_796));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i1_4_lut_adj_98.LUT_INIT = 16'hfbfa;
    SB_LUT4 n17427_bdd_4_lut (.I0(n17427), .I1(\mem_REG.mem_1_25 ), .I2(\mem_REG.mem_0_25 ), 
            .I3(rd_addr_r[1]), .O(n17430));
    defparam n17427_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16725_bdd_4_lut (.I0(n16725), .I1(n15106), .I2(n15105), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[10]));
    defparam n16725_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_99 (.I0(wr_addr_r[2]), .I1(\MISC.wr_flag_addr_r [0]), 
            .I2(rd_addr_r[2]), .I3(\MISC.rd_flag_addr_r [0]), .O(n4_adj_1398));   // src/fifo_sc_32_lut_gen.v(136[186:216])
    defparam i1_4_lut_adj_99.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_3_lut_adj_100 (.I0(wr_addr_r[1]), .I1(n4_adj_1398), .I2(rd_addr_r[1]), 
            .I3(GND_net), .O(full_nxt_w_N_812));   // src/fifo_sc_32_lut_gen.v(136[186:216])
    defparam i2_3_lut_adj_100.LUT_INIT = 16'hdede;
    SB_LUT4 i2_4_lut_adj_101 (.I0(wr_addr_p1_r[3]), .I1(wr_cmpaddr_p1_r[1]), 
            .I2(rd_addr_r[3]), .I3(rd_addr_r[1]), .O(n6_adj_1399));
    defparam i2_4_lut_adj_101.LUT_INIT = 16'h4812;
    SB_LUT4 i12501_4_lut (.I0(\MISC.wr_flag_addr_p1_r [0]), .I1(wr_cmpaddr_p1_r[2]), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(rd_addr_r[2]), .O(n14621));
    defparam i12501_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_3_lut_adj_102 (.I0(n14621), .I1(n2495), .I2(n6_adj_1399), 
            .I3(GND_net), .O(full_nxt_w_N_797));
    defparam i2_3_lut_adj_102.LUT_INIT = 16'h4040;
    SB_LUT4 i8233_4_lut (.I0(full_nxt_w_N_797), .I1(reset_all), .I2(\MISC.full_flag_r ), 
            .I3(n14607), .O(full_ext_r_N_794));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8233_4_lut.LUT_INIT = 16'h2232;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14817  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_27 ), .I2(\mem_REG.mem_7_27 ), .I3(rd_addr_r[1]), 
            .O(n16713));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14817 .LUT_INIT = 16'he4aa;
    SB_LUT4 n16713_bdd_4_lut (.I0(n16713), .I1(\mem_REG.mem_5_27 ), .I2(\mem_REG.mem_4_27 ), 
            .I3(rd_addr_r[1]), .O(n16716));
    defparam n16713_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8238_2_lut (.I0(rd_addr_nxt_w[0]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_addr_p1_r_3__N_712[0]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8238_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i8237_2_lut (.I0(rd_addr_nxt_w[0]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_addr_r_3__N_708[0]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8237_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i8235_2_lut (.I0(wr_addr_nxt_w[0]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_p1_r_3__N_694[0]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8235_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14493  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_14 ), .I2(\mem_REG.mem_3_14 ), .I3(rd_addr_r[1]), 
            .O(n16701));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14493 .LUT_INIT = 16'he4aa;
    SB_LUT4 n16701_bdd_4_lut (.I0(n16701), .I1(\mem_REG.mem_1_14 ), .I2(\mem_REG.mem_0_14 ), 
            .I3(rd_addr_r[1]), .O(n16704));
    defparam n16701_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8232_2_lut (.I0(wr_addr_nxt_w[0]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_r_3__N_690[0]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8232_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5395_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[9]), 
            .I3(\mem_REG.mem_7_9 ), .O(n6894));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5395_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5394_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[8]), 
            .I3(\mem_REG.mem_7_8 ), .O(n6893));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5394_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5385_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[31]), 
            .I3(\mem_REG.mem_6_31 ), .O(n6884));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5385_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5384_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[30]), 
            .I3(\mem_REG.mem_6_30 ), .O(n6883));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5384_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5383_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[29]), 
            .I3(\mem_REG.mem_6_29 ), .O(n6882));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5383_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5382_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[28]), 
            .I3(\mem_REG.mem_6_28 ), .O(n6881));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5382_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5381_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[27]), 
            .I3(\mem_REG.mem_6_27 ), .O(n6880));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5381_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12936_3_lut (.I0(\mem_REG.mem_0_8 ), .I1(\mem_REG.mem_1_8 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15060));
    defparam i12936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12937_3_lut (.I0(\mem_REG.mem_2_8 ), .I1(\mem_REG.mem_3_8 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15061));
    defparam i12937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12943_3_lut (.I0(\mem_REG.mem_6_8 ), .I1(\mem_REG.mem_7_8 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15067));
    defparam i12943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12942_3_lut (.I0(\mem_REG.mem_4_8 ), .I1(\mem_REG.mem_5_8 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15066));
    defparam i12942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14503 (.I0(rd_addr_r[1]), .I1(n15450), 
            .I2(n15451), .I3(rd_addr_r[2]), .O(n16677));
    defparam rd_addr_r_1__bdd_4_lut_14503.LUT_INIT = 16'he4aa;
    SB_LUT4 i5380_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[26]), 
            .I3(\mem_REG.mem_6_26 ), .O(n6879));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5380_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5379_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[25]), 
            .I3(\mem_REG.mem_6_25 ), .O(n6878));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5379_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5378_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[24]), 
            .I3(\mem_REG.mem_6_24 ), .O(n6877));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5378_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5377_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[23]), 
            .I3(\mem_REG.mem_6_23 ), .O(n6876));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5377_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5376_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[22]), 
            .I3(\mem_REG.mem_6_22 ), .O(n6875));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5376_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5375_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[21]), 
            .I3(\mem_REG.mem_6_21 ), .O(n6874));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5375_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5374_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[20]), 
            .I3(\mem_REG.mem_6_20 ), .O(n6873));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5374_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5373_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[19]), 
            .I3(\mem_REG.mem_6_19 ), .O(n6872));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5373_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16677_bdd_4_lut (.I0(n16677), .I1(n15070), .I2(n15069), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[9]));
    defparam n16677_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5372_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[18]), 
            .I3(\mem_REG.mem_6_18 ), .O(n6871));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5372_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5371_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[17]), 
            .I3(\mem_REG.mem_6_17 ), .O(n6870));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5371_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5370_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[16]), 
            .I3(\mem_REG.mem_6_16 ), .O(n6869));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5370_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13317_3_lut (.I0(\mem_REG.mem_0_18 ), .I1(\mem_REG.mem_1_18 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15441));
    defparam i13317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13318_3_lut (.I0(\mem_REG.mem_2_18 ), .I1(\mem_REG.mem_3_18 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15442));
    defparam i13318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5369_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[15]), 
            .I3(\mem_REG.mem_6_15 ), .O(n6868));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5369_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5368_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[14]), 
            .I3(\mem_REG.mem_6_14 ), .O(n6867));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5368_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5367_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[13]), 
            .I3(\mem_REG.mem_6_13 ), .O(n6866));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5367_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5366_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[12]), 
            .I3(\mem_REG.mem_6_12 ), .O(n6865));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5366_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5393_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[7]), 
            .I3(\mem_REG.mem_7_7 ), .O(n6892));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5393_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_15087  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_25 ), .I2(\mem_REG.mem_7_25 ), .I3(rd_addr_r[1]), 
            .O(n17391));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_15087 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17391_bdd_4_lut (.I0(n17391), .I1(\mem_REG.mem_5_25 ), .I2(\mem_REG.mem_4_25 ), 
            .I3(rd_addr_r[1]), .O(n17394));
    defparam n17391_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5365_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[11]), 
            .I3(\mem_REG.mem_6_11 ), .O(n6864));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5365_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5364_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[10]), 
            .I3(\mem_REG.mem_6_10 ), .O(n6863));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5364_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5363_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[9]), 
            .I3(\mem_REG.mem_6_9 ), .O(n6862));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5363_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5362_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[8]), 
            .I3(\mem_REG.mem_6_8 ), .O(n6861));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5362_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5361_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[7]), 
            .I3(\mem_REG.mem_6_7 ), .O(n6860));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5361_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5360_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[6]), 
            .I3(\mem_REG.mem_6_6 ), .O(n6859));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5360_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5359_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[5]), 
            .I3(\mem_REG.mem_6_5 ), .O(n6858));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5359_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5358_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[4]), 
            .I3(\mem_REG.mem_6_4 ), .O(n6857));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5358_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5357_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[3]), 
            .I3(\mem_REG.mem_6_3 ), .O(n6856));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5357_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5356_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[2]), 
            .I3(\mem_REG.mem_6_2 ), .O(n6855));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5356_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5355_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[1]), 
            .I3(\mem_REG.mem_6_1 ), .O(n6854));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5355_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5354_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[0]), 
            .I3(\mem_REG.mem_6_0 ), .O(n6853));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5354_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5353_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[31]), 
            .I3(\mem_REG.mem_5_31 ), .O(n6852));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5353_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5352_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[30]), 
            .I3(\mem_REG.mem_5_30 ), .O(n6851));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5352_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5351_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[29]), 
            .I3(\mem_REG.mem_5_29 ), .O(n6850));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5351_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5350_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[28]), 
            .I3(\mem_REG.mem_5_28 ), .O(n6849));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5350_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5349_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[27]), 
            .I3(\mem_REG.mem_5_27 ), .O(n6848));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5349_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5348_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[26]), 
            .I3(\mem_REG.mem_5_26 ), .O(n6847));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5348_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5347_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[25]), 
            .I3(\mem_REG.mem_5_25 ), .O(n6846));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5347_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5346_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[24]), 
            .I3(\mem_REG.mem_5_24 ), .O(n6845));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5346_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15122 (.I0(rd_addr_r[1]), .I1(n15495), 
            .I2(n15496), .I3(rd_addr_r[2]), .O(n17379));
    defparam rd_addr_r_1__bdd_4_lut_15122.LUT_INIT = 16'he4aa;
    SB_LUT4 i5345_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[23]), 
            .I3(\mem_REG.mem_5_23 ), .O(n6844));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5345_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5344_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[22]), 
            .I3(\mem_REG.mem_5_22 ), .O(n6843));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5344_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17379_bdd_4_lut (.I0(n17379), .I1(n15490), .I2(n15489), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[20]));
    defparam n17379_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5343_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[21]), 
            .I3(\mem_REG.mem_5_21 ), .O(n6842));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5343_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5342_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[20]), 
            .I3(\mem_REG.mem_5_20 ), .O(n6841));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5342_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5341_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[19]), 
            .I3(\mem_REG.mem_5_19 ), .O(n6840));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5341_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_15057  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_4 ), .I2(\mem_REG.mem_3_4 ), .I3(rd_addr_r[1]), 
            .O(n17373));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_15057 .LUT_INIT = 16'he4aa;
    SB_LUT4 i5340_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[18]), 
            .I3(\mem_REG.mem_5_18 ), .O(n6839));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5340_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5392_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[6]), 
            .I3(\mem_REG.mem_7_6 ), .O(n6891));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5392_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5339_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[17]), 
            .I3(\mem_REG.mem_5_17 ), .O(n6838));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5339_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5338_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[16]), 
            .I3(\mem_REG.mem_5_16 ), .O(n6837));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5338_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5337_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[15]), 
            .I3(\mem_REG.mem_5_15 ), .O(n6836));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5337_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5336_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[14]), 
            .I3(\mem_REG.mem_5_14 ), .O(n6835));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5336_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5335_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[13]), 
            .I3(\mem_REG.mem_5_13 ), .O(n6834));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5335_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5334_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[12]), 
            .I3(\mem_REG.mem_5_12 ), .O(n6833));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5334_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5333_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[11]), 
            .I3(\mem_REG.mem_5_11 ), .O(n6832));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5333_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14090  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_16 ), .I2(\mem_REG.mem_7_16 ), .I3(rd_addr_r[1]), 
            .O(n16167));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14090 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17373_bdd_4_lut (.I0(n17373), .I1(\mem_REG.mem_1_4 ), .I2(\mem_REG.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(n17376));
    defparam n17373_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16167_bdd_4_lut (.I0(n16167), .I1(\mem_REG.mem_5_16 ), .I2(\mem_REG.mem_4_16 ), 
            .I3(rd_addr_r[1]), .O(n16170));
    defparam n16167_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5332_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[10]), 
            .I3(\mem_REG.mem_5_10 ), .O(n6831));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5332_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5331_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[9]), 
            .I3(\mem_REG.mem_5_9 ), .O(n6830));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5331_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5330_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[8]), 
            .I3(\mem_REG.mem_5_8 ), .O(n6829));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5330_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5329_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[7]), 
            .I3(\mem_REG.mem_5_7 ), .O(n6828));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5329_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5328_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[6]), 
            .I3(\mem_REG.mem_5_6 ), .O(n6827));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5328_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5327_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[5]), 
            .I3(\mem_REG.mem_5_5 ), .O(n6826));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5327_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5391_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[5]), 
            .I3(\mem_REG.mem_7_5 ), .O(n6890));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5391_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5326_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[4]), 
            .I3(\mem_REG.mem_5_4 ), .O(n6825));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5326_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5325_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[3]), 
            .I3(\mem_REG.mem_5_3 ), .O(n6824));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5325_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5324_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[2]), 
            .I3(\mem_REG.mem_5_2 ), .O(n6823));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5324_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5323_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[1]), 
            .I3(\mem_REG.mem_5_1 ), .O(n6822));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5323_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5390_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[4]), 
            .I3(\mem_REG.mem_7_4 ), .O(n6889));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5390_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_en_i_I_0_181_2_lut (.I0(sc32_fifo_read_enable), .I1(\MISC.empty_flag_r ), 
            .I2(GND_net), .I3(GND_net), .O(\MISC.rd_w ));   // src/fifo_sc_32_lut_gen.v(269[25:52])
    defparam rd_en_i_I_0_181_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5322_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[0]), 
            .I3(\mem_REG.mem_5_0 ), .O(n6821));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5322_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14174  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_16 ), .I2(\mem_REG.mem_3_16 ), .I3(rd_addr_r[1]), 
            .O(n16227));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14174 .LUT_INIT = 16'he4aa;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_15042  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_26 ), .I2(\mem_REG.mem_3_26 ), .I3(rd_addr_r[1]), 
            .O(n17349));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_15042 .LUT_INIT = 16'he4aa;
    SB_LUT4 i5321_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[31]), 
            .I3(\mem_REG.mem_4_31 ), .O(n6820));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5321_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5320_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[30]), 
            .I3(\mem_REG.mem_4_30 ), .O(n6819));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5320_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5319_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[29]), 
            .I3(\mem_REG.mem_4_29 ), .O(n6818));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5319_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5318_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[28]), 
            .I3(\mem_REG.mem_4_28 ), .O(n6817));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5318_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5389_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[3]), 
            .I3(\mem_REG.mem_7_3 ), .O(n6888));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5389_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5317_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[27]), 
            .I3(\mem_REG.mem_4_27 ), .O(n6816));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5317_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5316_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[26]), 
            .I3(\mem_REG.mem_4_26 ), .O(n6815));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5316_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17349_bdd_4_lut (.I0(n17349), .I1(\mem_REG.mem_1_26 ), .I2(\mem_REG.mem_0_26 ), 
            .I3(rd_addr_r[1]), .O(n17352));
    defparam n17349_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5315_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[25]), 
            .I3(\mem_REG.mem_4_25 ), .O(n6814));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5315_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5314_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[24]), 
            .I3(\mem_REG.mem_4_24 ), .O(n6813));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5314_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5313_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[23]), 
            .I3(\mem_REG.mem_4_23 ), .O(n6812));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5313_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5312_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[22]), 
            .I3(\mem_REG.mem_4_22 ), .O(n6811));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5312_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5311_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[21]), 
            .I3(\mem_REG.mem_4_21 ), .O(n6810));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5311_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5310_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[20]), 
            .I3(\mem_REG.mem_4_20 ), .O(n6809));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5310_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5309_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[19]), 
            .I3(\mem_REG.mem_4_19 ), .O(n6808));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5309_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13092_3_lut (.I0(\mem_REG.mem_0_12 ), .I1(\mem_REG.mem_1_12 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15216));
    defparam i13092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5308_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[18]), 
            .I3(\mem_REG.mem_4_18 ), .O(n6807));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5308_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15047 (.I0(rd_addr_r[1]), .I1(n15453), 
            .I2(n15454), .I3(rd_addr_r[2]), .O(n17343));
    defparam rd_addr_r_1__bdd_4_lut_15047.LUT_INIT = 16'he4aa;
    SB_LUT4 i5307_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[17]), 
            .I3(\mem_REG.mem_4_17 ), .O(n6806));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5307_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5306_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[16]), 
            .I3(\mem_REG.mem_4_16 ), .O(n6805));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5306_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5305_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[15]), 
            .I3(\mem_REG.mem_4_15 ), .O(n6804));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5305_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5304_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[14]), 
            .I3(\mem_REG.mem_4_14 ), .O(n6803));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5304_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5303_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[13]), 
            .I3(\mem_REG.mem_4_13 ), .O(n6802));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5303_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5302_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[12]), 
            .I3(\mem_REG.mem_4_12 ), .O(n6801));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5302_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5301_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[11]), 
            .I3(\mem_REG.mem_4_11 ), .O(n6800));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5301_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5300_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[10]), 
            .I3(\mem_REG.mem_4_10 ), .O(n6799));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5300_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5299_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[9]), 
            .I3(\mem_REG.mem_4_9 ), .O(n6798));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5299_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5298_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[8]), 
            .I3(\mem_REG.mem_4_8 ), .O(n6797));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5298_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17343_bdd_4_lut (.I0(n17343), .I1(n15442), .I2(n15441), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[18]));
    defparam n17343_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5297_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[7]), 
            .I3(\mem_REG.mem_4_7 ), .O(n6796));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5297_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5296_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[6]), 
            .I3(\mem_REG.mem_4_6 ), .O(n6795));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5296_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15017 (.I0(rd_addr_r[1]), .I1(n15066), 
            .I2(n15067), .I3(rd_addr_r[2]), .O(n17337));
    defparam rd_addr_r_1__bdd_4_lut_15017.LUT_INIT = 16'he4aa;
    SB_LUT4 n17337_bdd_4_lut (.I0(n17337), .I1(n15061), .I2(n15060), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[8]));
    defparam n17337_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5295_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[5]), 
            .I3(\mem_REG.mem_4_5 ), .O(n6794));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5295_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5294_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[4]), 
            .I3(\mem_REG.mem_4_4 ), .O(n6793));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5294_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13093_3_lut (.I0(\mem_REG.mem_2_12 ), .I1(\mem_REG.mem_3_12 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15217));
    defparam i13093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5293_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[3]), 
            .I3(\mem_REG.mem_4_3 ), .O(n6792));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5293_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5292_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[2]), 
            .I3(\mem_REG.mem_4_2 ), .O(n6791));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5292_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5291_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[1]), 
            .I3(\mem_REG.mem_4_1 ), .O(n6790));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5291_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5290_3_lut_4_lut (.I0(n7), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[0]), 
            .I3(\mem_REG.mem_4_0 ), .O(n6789));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5290_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15012 (.I0(rd_addr_r[1]), .I1(n15429), 
            .I2(n15430), .I3(rd_addr_r[2]), .O(n17331));
    defparam rd_addr_r_1__bdd_4_lut_15012.LUT_INIT = 16'he4aa;
    SB_LUT4 n17331_bdd_4_lut (.I0(n17331), .I1(n15409), .I2(n15408), .I3(rd_addr_r[2]), 
            .O(rd_data_o_31__N_759[17]));
    defparam n17331_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_15022  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_26 ), .I2(\mem_REG.mem_7_26 ), .I3(rd_addr_r[1]), 
            .O(n17325));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_15022 .LUT_INIT = 16'he4aa;
    SB_LUT4 n16227_bdd_4_lut (.I0(n16227), .I1(\mem_REG.mem_1_16 ), .I2(\mem_REG.mem_0_16 ), 
            .I3(rd_addr_r[1]), .O(n16230));
    defparam n16227_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17325_bdd_4_lut (.I0(n17325), .I1(\mem_REG.mem_5_26 ), .I2(\mem_REG.mem_4_26 ), 
            .I3(rd_addr_r[1]), .O(n17328));
    defparam n17325_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5388_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[2]), 
            .I3(\mem_REG.mem_7_2 ), .O(n6887));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5388_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5289_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[31]), 
            .I3(\mem_REG.mem_3_31 ), .O(n6788));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5289_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5288_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[30]), 
            .I3(\mem_REG.mem_3_30 ), .O(n6787));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5288_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5287_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[29]), 
            .I3(\mem_REG.mem_3_29 ), .O(n6786));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5287_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5286_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[28]), 
            .I3(\mem_REG.mem_3_28 ), .O(n6785));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5286_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5285_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[27]), 
            .I3(\mem_REG.mem_3_27 ), .O(n6784));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5285_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5284_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[26]), 
            .I3(\mem_REG.mem_3_26 ), .O(n6783));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5284_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5283_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[25]), 
            .I3(\mem_REG.mem_3_25 ), .O(n6782));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5283_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5282_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[24]), 
            .I3(\mem_REG.mem_3_24 ), .O(n6781));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5282_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5281_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[23]), 
            .I3(\mem_REG.mem_3_23 ), .O(n6780));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5281_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5280_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[22]), 
            .I3(\mem_REG.mem_3_22 ), .O(n6779));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5280_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5279_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[21]), 
            .I3(\mem_REG.mem_3_21 ), .O(n6778));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5279_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5278_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[20]), 
            .I3(\mem_REG.mem_3_20 ), .O(n6777));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5278_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_15002  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_4 ), .I2(\mem_REG.mem_7_4 ), .I3(rd_addr_r[1]), 
            .O(n17313));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_15002 .LUT_INIT = 16'he4aa;
    SB_LUT4 i5277_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[19]), 
            .I3(\mem_REG.mem_3_19 ), .O(n6776));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5277_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5387_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[1]), 
            .I3(\mem_REG.mem_7_1 ), .O(n6886));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5387_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17313_bdd_4_lut (.I0(n17313), .I1(\mem_REG.mem_5_4 ), .I2(\mem_REG.mem_4_4 ), 
            .I3(rd_addr_r[1]), .O(n17316));
    defparam n17313_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5276_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[18]), 
            .I3(\mem_REG.mem_3_18 ), .O(n6775));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5276_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5275_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[17]), 
            .I3(\mem_REG.mem_3_17 ), .O(n6774));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5275_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5274_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[16]), 
            .I3(\mem_REG.mem_3_16 ), .O(n6773));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5274_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5273_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[15]), 
            .I3(\mem_REG.mem_3_15 ), .O(n6772));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5273_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5272_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[14]), 
            .I3(\mem_REG.mem_3_14 ), .O(n6771));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5272_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5271_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[13]), 
            .I3(\mem_REG.mem_3_13 ), .O(n6770));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5271_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5270_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[12]), 
            .I3(\mem_REG.mem_3_12 ), .O(n6769));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5270_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5269_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[11]), 
            .I3(\mem_REG.mem_3_11 ), .O(n6768));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5269_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5268_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[10]), 
            .I3(\mem_REG.mem_3_10 ), .O(n6767));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5268_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5267_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[9]), 
            .I3(\mem_REG.mem_3_9 ), .O(n6766));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5267_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14992  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_27 ), .I2(\mem_REG.mem_3_27 ), .I3(rd_addr_r[1]), 
            .O(n17301));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14992 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17301_bdd_4_lut (.I0(n17301), .I1(\mem_REG.mem_1_27 ), .I2(\mem_REG.mem_0_27 ), 
            .I3(rd_addr_r[1]), .O(n17304));
    defparam n17301_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5266_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[8]), 
            .I3(\mem_REG.mem_3_8 ), .O(n6765));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5266_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5265_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[7]), 
            .I3(\mem_REG.mem_3_7 ), .O(n6764));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5265_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5264_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[6]), 
            .I3(\mem_REG.mem_3_6 ), .O(n6763));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5264_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5263_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[5]), 
            .I3(\mem_REG.mem_3_5 ), .O(n6762));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5263_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5262_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[4]), 
            .I3(\mem_REG.mem_3_4 ), .O(n6761));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5262_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5261_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[3]), 
            .I3(\mem_REG.mem_3_3 ), .O(n6760));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5261_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5260_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[2]), 
            .I3(\mem_REG.mem_3_2 ), .O(n6759));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5260_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5259_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[1]), 
            .I3(\mem_REG.mem_3_1 ), .O(n6758));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5259_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5258_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[0]), 
            .I3(\mem_REG.mem_3_0 ), .O(n6757));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5258_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5257_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[31]), 
            .I3(\mem_REG.mem_2_31 ), .O(n6756));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5257_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5256_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[30]), 
            .I3(\mem_REG.mem_2_30 ), .O(n6755));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5256_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5255_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[29]), 
            .I3(\mem_REG.mem_2_29 ), .O(n6754));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5255_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5254_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[28]), 
            .I3(\mem_REG.mem_2_28 ), .O(n6753));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5254_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5253_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[27]), 
            .I3(\mem_REG.mem_2_27 ), .O(n6752));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5253_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5252_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[26]), 
            .I3(\mem_REG.mem_2_26 ), .O(n6751));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5252_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5251_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[25]), 
            .I3(\mem_REG.mem_2_25 ), .O(n6750));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5251_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5250_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[24]), 
            .I3(\mem_REG.mem_2_24 ), .O(n6749));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5250_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5249_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[23]), 
            .I3(\mem_REG.mem_2_23 ), .O(n6748));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5249_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5248_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[22]), 
            .I3(\mem_REG.mem_2_22 ), .O(n6747));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5248_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5247_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[21]), 
            .I3(\mem_REG.mem_2_21 ), .O(n6746));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5247_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5246_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[20]), 
            .I3(\mem_REG.mem_2_20 ), .O(n6745));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5246_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5245_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[19]), 
            .I3(\mem_REG.mem_2_19 ), .O(n6744));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5245_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5244_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[18]), 
            .I3(\mem_REG.mem_2_18 ), .O(n6743));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5244_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5243_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[17]), 
            .I3(\mem_REG.mem_2_17 ), .O(n6742));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5243_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5242_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[16]), 
            .I3(\mem_REG.mem_2_16 ), .O(n6741));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5242_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5241_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[15]), 
            .I3(\mem_REG.mem_2_15 ), .O(n6740));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5241_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5240_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[14]), 
            .I3(\mem_REG.mem_2_14 ), .O(n6739));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5240_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5239_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[13]), 
            .I3(\mem_REG.mem_2_13 ), .O(n6738));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5239_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5386_3_lut_4_lut (.I0(n8), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[0]), 
            .I3(\mem_REG.mem_7_0 ), .O(n6885));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5386_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5238_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[12]), 
            .I3(\mem_REG.mem_2_12 ), .O(n6737));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5238_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5237_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[11]), 
            .I3(\mem_REG.mem_2_11 ), .O(n6736));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5237_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5236_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[10]), 
            .I3(\mem_REG.mem_2_10 ), .O(n6735));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5236_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5235_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[9]), 
            .I3(\mem_REG.mem_2_9 ), .O(n6734));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5235_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13312_3_lut (.I0(\mem_REG.mem_6_12 ), .I1(\mem_REG.mem_7_12 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15436));
    defparam i13312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5234_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[8]), 
            .I3(\mem_REG.mem_2_8 ), .O(n6733));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5234_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14982  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_5 ), .I2(\mem_REG.mem_3_5 ), .I3(rd_addr_r[1]), 
            .O(n17283));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14982 .LUT_INIT = 16'he4aa;
    SB_LUT4 i13311_3_lut (.I0(\mem_REG.mem_4_12 ), .I1(\mem_REG.mem_5_12 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15435));
    defparam i13311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17283_bdd_4_lut (.I0(n17283), .I1(\mem_REG.mem_1_5 ), .I2(\mem_REG.mem_0_5 ), 
            .I3(rd_addr_r[1]), .O(n17286));
    defparam n17283_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5233_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[7]), 
            .I3(\mem_REG.mem_2_7 ), .O(n6732));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5233_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5232_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[6]), 
            .I3(\mem_REG.mem_2_6 ), .O(n6731));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5232_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5231_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[5]), 
            .I3(\mem_REG.mem_2_5 ), .O(n6730));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5231_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5230_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[4]), 
            .I3(\mem_REG.mem_2_4 ), .O(n6729));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5230_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5229_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[3]), 
            .I3(\mem_REG.mem_2_3 ), .O(n6728));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5229_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5228_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[2]), 
            .I3(\mem_REG.mem_2_2 ), .O(n6727));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5228_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5227_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[1]), 
            .I3(\mem_REG.mem_2_1 ), .O(n6726));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5227_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5226_3_lut_4_lut (.I0(n6_adj_1400), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[0]), 
            .I3(\mem_REG.mem_2_0 ), .O(n6725));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5226_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14967  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_28 ), .I2(\mem_REG.mem_3_28 ), .I3(rd_addr_r[1]), 
            .O(n17265));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14967 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17265_bdd_4_lut (.I0(n17265), .I1(\mem_REG.mem_1_28 ), .I2(\mem_REG.mem_0_28 ), 
            .I3(rd_addr_r[1]), .O(n17268));
    defparam n17265_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14952  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_28 ), .I2(\mem_REG.mem_7_28 ), .I3(rd_addr_r[1]), 
            .O(n17241));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14952 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17241_bdd_4_lut (.I0(n17241), .I1(\mem_REG.mem_5_28 ), .I2(\mem_REG.mem_4_28 ), 
            .I3(rd_addr_r[1]), .O(n17244));
    defparam n17241_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14932  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_5 ), .I2(\mem_REG.mem_7_5 ), .I3(rd_addr_r[1]), 
            .O(n17235));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14932 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17235_bdd_4_lut (.I0(n17235), .I1(\mem_REG.mem_5_5 ), .I2(\mem_REG.mem_4_5 ), 
            .I3(rd_addr_r[1]), .O(n17238));
    defparam n17235_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13330_3_lut (.I0(\mem_REG.mem_6_18 ), .I1(\mem_REG.mem_7_18 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15454));
    defparam i13330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13329_3_lut (.I0(\mem_REG.mem_4_18 ), .I1(\mem_REG.mem_5_18 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15453));
    defparam i13329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14927  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_29 ), .I2(\mem_REG.mem_3_29 ), .I3(rd_addr_r[1]), 
            .O(n17229));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14927 .LUT_INIT = 16'he4aa;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14483  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_15 ), .I2(\mem_REG.mem_3_15 ), .I3(rd_addr_r[1]), 
            .O(n16461));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14483 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17229_bdd_4_lut (.I0(n17229), .I1(\mem_REG.mem_1_29 ), .I2(\mem_REG.mem_0_29 ), 
            .I3(rd_addr_r[1]), .O(n17232));
    defparam n17229_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16461_bdd_4_lut (.I0(n16461), .I1(\mem_REG.mem_1_15 ), .I2(\mem_REG.mem_0_15 ), 
            .I3(rd_addr_r[1]), .O(n16464));
    defparam n16461_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_14 ), .I2(\mem_REG.mem_7_14 ), .I3(rd_addr_r[1]), 
            .O(n17985));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut .LUT_INIT = 16'he4aa;
    SB_LUT4 n17985_bdd_4_lut (.I0(n17985), .I1(\mem_REG.mem_5_14 ), .I2(\mem_REG.mem_4_14 ), 
            .I3(rd_addr_r[1]), .O(n17988));
    defparam n17985_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14922  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_29 ), .I2(\mem_REG.mem_7_29 ), .I3(rd_addr_r[1]), 
            .O(n17223));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14922 .LUT_INIT = 16'he4aa;
    SB_LUT4 i13365_3_lut (.I0(\mem_REG.mem_0_20 ), .I1(\mem_REG.mem_1_20 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15489));
    defparam i13365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13366_3_lut (.I0(\mem_REG.mem_2_20 ), .I1(\mem_REG.mem_3_20 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15490));
    defparam i13366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13372_3_lut (.I0(\mem_REG.mem_6_20 ), .I1(\mem_REG.mem_7_20 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15496));
    defparam i13372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13371_3_lut (.I0(\mem_REG.mem_4_20 ), .I1(\mem_REG.mem_5_20 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15495));
    defparam i13371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17223_bdd_4_lut (.I0(n17223), .I1(\mem_REG.mem_5_29 ), .I2(\mem_REG.mem_4_29 ), 
            .I3(rd_addr_r[1]), .O(n17226));
    defparam n17223_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12945_3_lut (.I0(\mem_REG.mem_0_9 ), .I1(\mem_REG.mem_1_9 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15069));
    defparam i12945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12946_3_lut (.I0(\mem_REG.mem_2_9 ), .I1(\mem_REG.mem_3_9 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15070));
    defparam i12946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13623_3_lut (.I0(\mem_REG.mem_0_30 ), .I1(\mem_REG.mem_1_30 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15747));
    defparam i13623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13624_3_lut (.I0(\mem_REG.mem_2_30 ), .I1(\mem_REG.mem_3_30 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15748));
    defparam i13624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13633_3_lut (.I0(\mem_REG.mem_6_30 ), .I1(\mem_REG.mem_7_30 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15757));
    defparam i13633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13632_3_lut (.I0(\mem_REG.mem_4_30 ), .I1(\mem_REG.mem_5_30 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15756));
    defparam i13632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13122_3_lut (.I0(\mem_REG.mem_0_13 ), .I1(\mem_REG.mem_1_13 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15246));
    defparam i13122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13123_3_lut (.I0(\mem_REG.mem_2_13 ), .I1(\mem_REG.mem_3_13 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15247));
    defparam i13123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13144_3_lut (.I0(\mem_REG.mem_6_13 ), .I1(\mem_REG.mem_7_13 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15268));
    defparam i13144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13143_3_lut (.I0(\mem_REG.mem_4_13 ), .I1(\mem_REG.mem_5_13 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15267));
    defparam i13143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14917  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_6 ), .I2(\mem_REG.mem_3_6 ), .I3(rd_addr_r[1]), 
            .O(n17199));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14917 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17199_bdd_4_lut (.I0(n17199), .I1(\mem_REG.mem_1_6 ), .I2(\mem_REG.mem_0_6 ), 
            .I3(rd_addr_r[1]), .O(n17202));
    defparam n17199_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13327_3_lut (.I0(\mem_REG.mem_6_9 ), .I1(\mem_REG.mem_7_9 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15451));
    defparam i13327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13326_3_lut (.I0(\mem_REG.mem_4_9 ), .I1(\mem_REG.mem_5_9 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15450));
    defparam i13326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14897  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_6 ), .I2(\mem_REG.mem_7_6 ), .I3(rd_addr_r[1]), 
            .O(n17193));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14897 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17193_bdd_4_lut (.I0(n17193), .I1(\mem_REG.mem_5_6 ), .I2(\mem_REG.mem_4_6 ), 
            .I3(rd_addr_r[1]), .O(n17196));
    defparam n17193_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14892  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_31 ), .I2(\mem_REG.mem_3_31 ), .I3(rd_addr_r[1]), 
            .O(n17187));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14892 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17187_bdd_4_lut (.I0(n17187), .I1(\mem_REG.mem_1_31 ), .I2(\mem_REG.mem_0_31 ), 
            .I3(rd_addr_r[1]), .O(n17190));
    defparam n17187_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14887  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_31 ), .I2(\mem_REG.mem_7_31 ), .I3(rd_addr_r[1]), 
            .O(n17175));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14887 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17175_bdd_4_lut (.I0(n17175), .I1(\mem_REG.mem_5_31 ), .I2(\mem_REG.mem_4_31 ), 
            .I3(rd_addr_r[1]), .O(n17178));
    defparam n17175_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5225_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[31]), 
            .I3(\mem_REG.mem_1_31 ), .O(n6724));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5225_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5224_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[30]), 
            .I3(\mem_REG.mem_1_30 ), .O(n6723));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5224_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5223_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[29]), 
            .I3(\mem_REG.mem_1_29 ), .O(n6722));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5223_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5222_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[28]), 
            .I3(\mem_REG.mem_1_28 ), .O(n6721));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5222_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5221_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[27]), 
            .I3(\mem_REG.mem_1_27 ), .O(n6720));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5221_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5220_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[26]), 
            .I3(\mem_REG.mem_1_26 ), .O(n6719));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5220_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5219_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[25]), 
            .I3(\mem_REG.mem_1_25 ), .O(n6718));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5219_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5218_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[24]), 
            .I3(\mem_REG.mem_1_24 ), .O(n6717));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5218_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5217_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[23]), 
            .I3(\mem_REG.mem_1_23 ), .O(n6716));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5217_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5216_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[22]), 
            .I3(\mem_REG.mem_1_22 ), .O(n6715));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5216_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5215_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[21]), 
            .I3(\mem_REG.mem_1_21 ), .O(n6714));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5215_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_15552  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_3 ), .I2(\mem_REG.mem_7_3 ), .I3(rd_addr_r[1]), 
            .O(n17913));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_15552 .LUT_INIT = 16'he4aa;
    SB_LUT4 n17913_bdd_4_lut (.I0(n17913), .I1(\mem_REG.mem_5_3 ), .I2(\mem_REG.mem_4_3 ), 
            .I3(rd_addr_r[1]), .O(n17916));
    defparam n17913_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5214_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[20]), 
            .I3(\mem_REG.mem_1_20 ), .O(n6713));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5214_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5213_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[19]), 
            .I3(\mem_REG.mem_1_19 ), .O(n6712));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5213_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5212_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[18]), 
            .I3(\mem_REG.mem_1_18 ), .O(n6711));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5212_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5211_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[17]), 
            .I3(\mem_REG.mem_1_17 ), .O(n6710));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5211_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5210_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[16]), 
            .I3(\mem_REG.mem_1_16 ), .O(n6709));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5210_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5209_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[15]), 
            .I3(\mem_REG.mem_1_15 ), .O(n6708));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5209_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14284  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_15 ), .I2(\mem_REG.mem_7_15 ), .I3(rd_addr_r[1]), 
            .O(n16389));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14284 .LUT_INIT = 16'he4aa;
    SB_LUT4 n16389_bdd_4_lut (.I0(n16389), .I1(\mem_REG.mem_5_15 ), .I2(\mem_REG.mem_4_15 ), 
            .I3(rd_addr_r[1]), .O(n16392));
    defparam n16389_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5208_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[14]), 
            .I3(\mem_REG.mem_1_14 ), .O(n6707));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5208_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5207_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[13]), 
            .I3(\mem_REG.mem_1_13 ), .O(n6706));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5207_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5206_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[12]), 
            .I3(\mem_REG.mem_1_12 ), .O(n6705));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5206_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5205_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[11]), 
            .I3(\mem_REG.mem_1_11 ), .O(n6704));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5205_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5204_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[10]), 
            .I3(\mem_REG.mem_1_10 ), .O(n6703));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5204_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5203_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[9]), 
            .I3(\mem_REG.mem_1_9 ), .O(n6702));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5203_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5202_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[8]), 
            .I3(\mem_REG.mem_1_8 ), .O(n6701));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5202_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5201_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[7]), 
            .I3(\mem_REG.mem_1_7 ), .O(n6700));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5201_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5200_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[6]), 
            .I3(\mem_REG.mem_1_6 ), .O(n6699));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5200_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5199_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[5]), 
            .I3(\mem_REG.mem_1_5 ), .O(n6698));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5199_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_15492  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_21 ), .I2(\mem_REG.mem_3_21 ), .I3(rd_addr_r[1]), 
            .O(n17889));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_15492 .LUT_INIT = 16'he4aa;
    SB_LUT4 i5198_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[4]), 
            .I3(\mem_REG.mem_1_4 ), .O(n6697));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5198_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17889_bdd_4_lut (.I0(n17889), .I1(\mem_REG.mem_1_21 ), .I2(\mem_REG.mem_0_21 ), 
            .I3(rd_addr_r[1]), .O(n17892));
    defparam n17889_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5197_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[3]), 
            .I3(\mem_REG.mem_1_3 ), .O(n6696));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5197_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12981_3_lut (.I0(\mem_REG.mem_0_10 ), .I1(\mem_REG.mem_1_10 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15105));
    defparam i12981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12982_3_lut (.I0(\mem_REG.mem_2_10 ), .I1(\mem_REG.mem_3_10 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15106));
    defparam i12982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13324_3_lut (.I0(\mem_REG.mem_6_10 ), .I1(\mem_REG.mem_7_10 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15448));
    defparam i13324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13323_3_lut (.I0(\mem_REG.mem_4_10 ), .I1(\mem_REG.mem_5_10 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15447));
    defparam i13323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5196_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[2]), 
            .I3(\mem_REG.mem_1_2 ), .O(n6695));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5196_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5195_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[1]), 
            .I3(\mem_REG.mem_1_1 ), .O(n6694));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5195_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5194_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(dc32_fifo_data_out[0]), 
            .I3(\mem_REG.mem_1_0 ), .O(n6693));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam i5194_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i6_2_lut_4_lut (.I0(sc32_fifo_write_enable), 
            .I1(\MISC.full_flag_r ), .I2(\MISC.wr_flag_addr_r [0]), .I3(wr_addr_r[1]), 
            .O(n6_adj_1400));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam EnabledDecoder_2_i6_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i8375_3_lut_4_lut (.I0(wr_addr_nxt_w[2]), .I1(reset_all), .I2(wr_addr_nxt_w[1]), 
            .I3(wr_addr_nxt_w[0]), .O(wr_addr_p1_r_3__N_694[2]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8375_3_lut_4_lut.LUT_INIT = 16'h1222;
    SB_LUT4 rd_addr_r_3__I_0_i2_3_lut_4_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1cmp_r[1]), 
            .I2(sc32_fifo_read_enable), .I3(\MISC.empty_flag_r ), .O(rd_addr_nxt_w[1]));   // src/fifo_sc_32_lut_gen.v(133[44:95])
    defparam rd_addr_r_3__I_0_i2_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 rd_addr_r_3__I_0_i3_3_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1cmp_r[2]), 
            .I2(sc32_fifo_read_enable), .I3(\MISC.empty_flag_r ), .O(rd_addr_nxt_w[2]));   // src/fifo_sc_32_lut_gen.v(133[44:95])
    defparam rd_addr_r_3__I_0_i3_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 rd_addr_r_3__I_0_i4_3_lut_4_lut (.I0(rd_addr_r[3]), .I1(rd_addr_p1cmp_r[3]), 
            .I2(sc32_fifo_read_enable), .I3(\MISC.empty_flag_r ), .O(rd_addr_nxt_w[3]));   // src/fifo_sc_32_lut_gen.v(133[44:95])
    defparam rd_addr_r_3__I_0_i4_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i8380_3_lut_4_lut (.I0(rd_addr_nxt_w[2]), .I1(reset_all), .I2(rd_addr_nxt_w[1]), 
            .I3(rd_addr_nxt_w[0]), .O(rd_addr_p1_r_3__N_712[2]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8380_3_lut_4_lut.LUT_INIT = 16'h1222;
    SB_LUT4 i8381_4_lut (.I0(rd_addr_nxt_w[3]), .I1(reset_all), .I2(rd_addr_nxt_w[2]), 
            .I3(n3181), .O(rd_addr_p1_r_3__N_712[3]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8381_4_lut.LUT_INIT = 16'h1222;
    SB_LUT4 i1711_2_lut (.I0(rd_addr_nxt_w[1]), .I1(rd_addr_nxt_w[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3181));   // src/fifo_sc_32_lut_gen.v(134[47:69])
    defparam i1711_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8379_3_lut (.I0(rd_addr_nxt_w[1]), .I1(reset_all), .I2(rd_addr_nxt_w[0]), 
            .I3(GND_net), .O(rd_addr_p1_r_3__N_712[1]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8379_3_lut.LUT_INIT = 16'h1212;
    SB_LUT4 i8378_2_lut (.I0(rd_addr_nxt_w[3]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_addr_r_3__N_708[3]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8378_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i8377_2_lut (.I0(rd_addr_nxt_w[2]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_addr_r_3__N_708[2]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8377_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i8376_2_lut (.I0(rd_addr_nxt_w[1]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(rd_addr_r_3__N_708[1]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8376_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i8374_3_lut (.I0(wr_addr_nxt_w[1]), .I1(reset_all), .I2(wr_addr_nxt_w[0]), 
            .I3(GND_net), .O(wr_addr_p1_r_3__N_694[1]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8374_3_lut.LUT_INIT = 16'h1212;
    SB_LUT4 i1682_2_lut (.I0(wr_addr_nxt_w[1]), .I1(wr_addr_nxt_w[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3152));   // src/fifo_sc_32_lut_gen.v(131[47:69])
    defparam i1682_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8236_4_lut (.I0(wr_addr_nxt_w[3]), .I1(reset_all), .I2(wr_addr_nxt_w[2]), 
            .I3(n3152), .O(wr_addr_p1cmp_r_3__N_698[3]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8236_4_lut.LUT_INIT = 16'h1222;
    SB_LUT4 i3914_1_lut (.I0(sc32_fifo_data_out[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5413));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3914_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 EnabledDecoder_2_i7_2_lut_4_lut (.I0(sc32_fifo_write_enable), 
            .I1(\MISC.full_flag_r ), .I2(\MISC.wr_flag_addr_r [0]), .I3(wr_addr_r[1]), 
            .O(n7));   // src/fifo_sc_32_lut_gen.v(613[33:45])
    defparam EnabledDecoder_2_i7_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14224  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_22 ), .I2(\mem_REG.mem_3_22 ), .I3(rd_addr_r[1]), 
            .O(n16335));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14224 .LUT_INIT = 16'he4aa;
    SB_LUT4 n16335_bdd_4_lut (.I0(n16335), .I1(\mem_REG.mem_1_22 ), .I2(\mem_REG.mem_0_22 ), 
            .I3(rd_addr_r[1]), .O(n16338));
    defparam n16335_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14179  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_21 ), .I2(\mem_REG.mem_7_21 ), .I3(rd_addr_r[1]), 
            .O(n16329));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14179 .LUT_INIT = 16'he4aa;
    SB_LUT4 n16329_bdd_4_lut (.I0(n16329), .I1(\mem_REG.mem_5_21 ), .I2(\mem_REG.mem_4_21 ), 
            .I3(rd_addr_r[1]), .O(n16332));
    defparam n16329_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8373_2_lut (.I0(wr_addr_nxt_w[3]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_r_3__N_690[3]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8373_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i8372_2_lut (.I0(wr_addr_nxt_w[2]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_r_3__N_690[2]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8372_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i8371_2_lut (.I0(wr_addr_nxt_w[1]), .I1(reset_all), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_r_3__N_690[1]));   // src/fifo_sc_32_lut_gen.v(176[25] 195[28])
    defparam i8371_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13278_3_lut (.I0(\mem_REG.mem_0_1 ), .I1(\mem_REG.mem_1_1 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15402));
    defparam i13278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13279_3_lut (.I0(\mem_REG.mem_2_1 ), .I1(\mem_REG.mem_3_1 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15403));
    defparam i13279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13426_3_lut (.I0(\mem_REG.mem_6_1 ), .I1(\mem_REG.mem_7_1 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15550));
    defparam i13426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13425_3_lut (.I0(\mem_REG.mem_4_1 ), .I1(\mem_REG.mem_5_1 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15549));
    defparam i13425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_3__I_0_i1_3_lut_4_lut (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\MISC.rd_flag_addr_p1_r [0]), .I2(sc32_fifo_read_enable), 
            .I3(\MISC.empty_flag_r ), .O(rd_addr_nxt_w[0]));   // src/fifo_sc_32_lut_gen.v(133[44:95])
    defparam rd_addr_r_3__I_0_i1_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i12487_2_lut_4_lut (.I0(sc32_fifo_read_enable), .I1(wr_addr_r[1]), 
            .I2(n4_adj_1398), .I3(rd_addr_r[1]), .O(n14607));
    defparam i12487_2_lut_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 i3915_1_lut (.I0(sc32_fifo_data_out[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5414));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3915_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13461_3_lut (.I0(\mem_REG.mem_0_24 ), .I1(\mem_REG.mem_1_24 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15585));
    defparam i13461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_15472  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_22 ), .I2(\mem_REG.mem_7_22 ), .I3(rd_addr_r[1]), 
            .O(n17835));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_15472 .LUT_INIT = 16'he4aa;
    SB_LUT4 i13462_3_lut (.I0(\mem_REG.mem_2_24 ), .I1(\mem_REG.mem_3_24 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15586));
    defparam i13462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17835_bdd_4_lut (.I0(n17835), .I1(\mem_REG.mem_5_22 ), .I2(\mem_REG.mem_4_22 ), 
            .I3(rd_addr_r[1]), .O(n17838));
    defparam n17835_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1254_2_lut_3_lut_4_lut (.I0(sc32_fifo_write_enable), .I1(\MISC.full_flag_r ), 
            .I2(sc32_fifo_read_enable), .I3(\MISC.empty_flag_r ), .O(n2495));   // src/fifo_sc_32_lut_gen.v(268[25:51])
    defparam i1254_2_lut_3_lut_4_lut.LUT_INIT = 16'h2202;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14877  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_2_7 ), .I2(\mem_REG.mem_3_7 ), .I3(rd_addr_r[1]), 
            .O(n17115));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14877 .LUT_INIT = 16'he4aa;
    SB_LUT4 i9046253_i1_3_lut (.I0(n17190), .I1(n17178), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[31]));
    defparam i9046253_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9034247_i1_3_lut (.I0(n17232), .I1(n17226), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[29]));
    defparam i9034247_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9028244_i1_3_lut (.I0(n17268), .I1(n17244), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[28]));
    defparam i9028244_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9022241_i1_3_lut (.I0(n17304), .I1(n16716), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[27]));
    defparam i9022241_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9016238_i1_3_lut (.I0(n17352), .I1(n17328), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[26]));
    defparam i9016238_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9010235_i1_3_lut (.I0(n17430), .I1(n17394), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[25]));
    defparam i9010235_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8968214_i1_3_lut (.I0(n16338), .I1(n17838), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[22]));
    defparam i8968214_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8962211_i1_3_lut (.I0(n17892), .I1(n16332), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[21]));
    defparam i8962211_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8932196_i1_3_lut (.I0(n16230), .I1(n16170), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[16]));
    defparam i8932196_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17115_bdd_4_lut (.I0(n17115), .I1(\mem_REG.mem_1_7 ), .I2(\mem_REG.mem_0_7 ), 
            .I3(rd_addr_r[1]), .O(n17118));
    defparam n17115_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8926193_i1_3_lut (.I0(n16464), .I1(n16392), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[15]));
    defparam i8926193_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8920190_i1_3_lut (.I0(n16704), .I1(n17988), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[14]));
    defparam i8920190_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8854157_i1_3_lut (.I0(n17118), .I1(n17106), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[7]));
    defparam i8854157_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8848154_i1_3_lut (.I0(n17202), .I1(n17196), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[6]));
    defparam i8848154_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8842151_i1_3_lut (.I0(n17286), .I1(n17238), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[5]));
    defparam i8842151_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8836148_i1_3_lut (.I0(n17376), .I1(n17316), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[4]));
    defparam i8836148_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13474_3_lut (.I0(\mem_REG.mem_6_24 ), .I1(\mem_REG.mem_7_24 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15598));
    defparam i13474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13473_3_lut (.I0(\mem_REG.mem_4_24 ), .I1(\mem_REG.mem_5_24 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15597));
    defparam i13473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8830145_i1_3_lut (.I0(n17490), .I1(n17916), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[3]));
    defparam i8830145_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8824142_i1_3_lut (.I0(n17640), .I1(n17550), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(rd_data_o_31__N_759[2]));
    defparam i8824142_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \MISC.rd_flag_addr_r_0__bdd_4_lut_14827  (.I0(\MISC.rd_flag_addr_r [0]), 
            .I1(\mem_REG.mem_6_7 ), .I2(\mem_REG.mem_7_7 ), .I3(rd_addr_r[1]), 
            .O(n17103));
    defparam \MISC.rd_flag_addr_r_0__bdd_4_lut_14827 .LUT_INIT = 16'he4aa;
    SB_LUT4 i3912_1_lut (.I0(sc32_fifo_data_out[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n5411));   // src/fifo_sc_32_lut_gen.v(617[21] 623[24])
    defparam i3912_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13032_3_lut (.I0(\mem_REG.mem_0_11 ), .I1(\mem_REG.mem_1_11 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15156));
    defparam i13032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13033_3_lut (.I0(\mem_REG.mem_2_11 ), .I1(\mem_REG.mem_3_11 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15157));
    defparam i13033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13063_3_lut (.I0(\mem_REG.mem_6_11 ), .I1(\mem_REG.mem_7_11 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15187));
    defparam i13063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13062_3_lut (.I0(\mem_REG.mem_4_11 ), .I1(\mem_REG.mem_5_11 ), 
            .I2(\MISC.rd_flag_addr_r [0]), .I3(GND_net), .O(n15186));
    defparam i13062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17103_bdd_4_lut (.I0(n17103), .I1(\mem_REG.mem_5_7 ), .I2(\mem_REG.mem_4_7 ), 
            .I3(rd_addr_r[1]), .O(n17106));
    defparam n17103_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word
//

module FIFO_Quad_Word (\rd_addr_r[1] , \rd_addr_r[0] , SLM_CLK_c, reset_all_w, 
            wr_addr_r, rx_buf_byte, rd_fifo_en_w, \mem_LUT.data_raw_r[0] , 
            n8, n7067, VCC_net, \fifo_temp_output[1] , n4566, GND_net, 
            \wr_addr_p1_w[2] , n13820, n7064, \fifo_temp_output[2] , 
            n7061, \fifo_temp_output[3] , n7058, \fifo_temp_output[4] , 
            n7055, \fifo_temp_output[5] , n7052, \fifo_temp_output[6] , 
            n7049, \fifo_temp_output[7] , n5647, n5658, n6970, \fifo_temp_output[0] , 
            n14076, is_tx_fifo_full_flag, \rd_addr_p1_w[1] , \rd_addr_p1_w[2] , 
            fifo_write_cmd, wr_fifo_en_w, \mem_LUT.data_raw_r[1] , \mem_LUT.data_raw_r[2] , 
            \mem_LUT.data_raw_r[3] , \mem_LUT.data_raw_r[4] , \mem_LUT.data_raw_r[5] , 
            \mem_LUT.data_raw_r[6] , \mem_LUT.data_raw_r[7] , fifo_read_cmd, 
            is_fifo_empty_flag, n5664, n14096, n5207) /* synthesis syn_module_defined=1 */ ;
    output \rd_addr_r[1] ;
    output \rd_addr_r[0] ;
    input SLM_CLK_c;
    input reset_all_w;
    output [2:0]wr_addr_r;
    input [7:0]rx_buf_byte;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[0] ;
    input n8;
    input n7067;
    input VCC_net;
    output \fifo_temp_output[1] ;
    output n4566;
    input GND_net;
    output \wr_addr_p1_w[2] ;
    output n13820;
    input n7064;
    output \fifo_temp_output[2] ;
    input n7061;
    output \fifo_temp_output[3] ;
    input n7058;
    output \fifo_temp_output[4] ;
    input n7055;
    output \fifo_temp_output[5] ;
    input n7052;
    output \fifo_temp_output[6] ;
    input n7049;
    output \fifo_temp_output[7] ;
    input n5647;
    input n5658;
    input n6970;
    output \fifo_temp_output[0] ;
    input n14076;
    output is_tx_fifo_full_flag;
    output \rd_addr_p1_w[1] ;
    output \rd_addr_p1_w[2] ;
    input fifo_write_cmd;
    output wr_fifo_en_w;
    output \mem_LUT.data_raw_r[1] ;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[3] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[7] ;
    input fifo_read_cmd;
    output is_fifo_empty_flag;
    input n5664;
    input n14096;
    output n5207;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_3 lscc_fifo_inst (.rd_addr_r({Open_0, 
            \rd_addr_r[1] , \rd_addr_r[0] }), .SLM_CLK_c(SLM_CLK_c), .reset_all_w(reset_all_w), 
            .wr_addr_r({wr_addr_r}), .rx_buf_byte({rx_buf_byte}), .rd_fifo_en_w(rd_fifo_en_w), 
            .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r[0] ), .n8(n8), 
            .n7067(n7067), .VCC_net(VCC_net), .\fifo_temp_output[1] (\fifo_temp_output[1] ), 
            .n4566(n4566), .GND_net(GND_net), .\wr_addr_p1_w[2] (\wr_addr_p1_w[2] ), 
            .n13820(n13820), .n7064(n7064), .\fifo_temp_output[2] (\fifo_temp_output[2] ), 
            .n7061(n7061), .\fifo_temp_output[3] (\fifo_temp_output[3] ), 
            .n7058(n7058), .\fifo_temp_output[4] (\fifo_temp_output[4] ), 
            .n7055(n7055), .\fifo_temp_output[5] (\fifo_temp_output[5] ), 
            .n7052(n7052), .\fifo_temp_output[6] (\fifo_temp_output[6] ), 
            .n7049(n7049), .\fifo_temp_output[7] (\fifo_temp_output[7] ), 
            .n5647(n5647), .n5658(n5658), .n6970(n6970), .\fifo_temp_output[0] (\fifo_temp_output[0] ), 
            .n14076(n14076), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .\rd_addr_p1_w[1] (\rd_addr_p1_w[1] ), .\rd_addr_p1_w[2] (\rd_addr_p1_w[2] ), 
            .fifo_write_cmd(fifo_write_cmd), .wr_fifo_en_w(wr_fifo_en_w), 
            .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r[1] ), .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r[2] ), 
            .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r[3] ), .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r[4] ), 
            .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r[5] ), .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r[6] ), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r[7] ), .fifo_read_cmd(fifo_read_cmd), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .n5664(n5664), .n14096(n14096), 
            .n5207(n5207)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_quad_word_mod.v(20[37:380])
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_3
//

module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_3 (rd_addr_r, 
            SLM_CLK_c, reset_all_w, wr_addr_r, rx_buf_byte, rd_fifo_en_w, 
            \mem_LUT.data_raw_r[0] , n8, n7067, VCC_net, \fifo_temp_output[1] , 
            n4566, GND_net, \wr_addr_p1_w[2] , n13820, n7064, \fifo_temp_output[2] , 
            n7061, \fifo_temp_output[3] , n7058, \fifo_temp_output[4] , 
            n7055, \fifo_temp_output[5] , n7052, \fifo_temp_output[6] , 
            n7049, \fifo_temp_output[7] , n5647, n5658, n6970, \fifo_temp_output[0] , 
            n14076, is_tx_fifo_full_flag, \rd_addr_p1_w[1] , \rd_addr_p1_w[2] , 
            fifo_write_cmd, wr_fifo_en_w, \mem_LUT.data_raw_r[1] , \mem_LUT.data_raw_r[2] , 
            \mem_LUT.data_raw_r[3] , \mem_LUT.data_raw_r[4] , \mem_LUT.data_raw_r[5] , 
            \mem_LUT.data_raw_r[6] , \mem_LUT.data_raw_r[7] , fifo_read_cmd, 
            is_fifo_empty_flag, n5664, n14096, n5207) /* synthesis syn_module_defined=1 */ ;
    output [2:0]rd_addr_r;
    input SLM_CLK_c;
    input reset_all_w;
    output [2:0]wr_addr_r;
    input [7:0]rx_buf_byte;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[0] ;
    input n8;
    input n7067;
    input VCC_net;
    output \fifo_temp_output[1] ;
    output n4566;
    input GND_net;
    output \wr_addr_p1_w[2] ;
    output n13820;
    input n7064;
    output \fifo_temp_output[2] ;
    input n7061;
    output \fifo_temp_output[3] ;
    input n7058;
    output \fifo_temp_output[4] ;
    input n7055;
    output \fifo_temp_output[5] ;
    input n7052;
    output \fifo_temp_output[6] ;
    input n7049;
    output \fifo_temp_output[7] ;
    input n5647;
    input n5658;
    input n6970;
    output \fifo_temp_output[0] ;
    input n14076;
    output is_tx_fifo_full_flag;
    output \rd_addr_p1_w[1] ;
    output \rd_addr_p1_w[2] ;
    input fifo_write_cmd;
    output wr_fifo_en_w;
    output \mem_LUT.data_raw_r[1] ;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[3] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[7] ;
    input fifo_read_cmd;
    output is_fifo_empty_flag;
    input n5664;
    input n14096;
    output n5207;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n16311, \mem_LUT.mem_1_2 , \mem_LUT.mem_0_2 ;
    wire [31:0]\mem_LUT.data_raw_r_31__N_1269 ;
    wire [2:0]n12;
    
    wire n4, \mem_LUT.mem_0_7 , n6924, \mem_LUT.mem_2_1 , \mem_LUT.mem_3_1 , 
        n16305, \mem_LUT.mem_0_6 , n6923, \mem_LUT.mem_1_1 , \mem_LUT.mem_0_1 , 
        \mem_LUT.mem_0_5 , n6922, \mem_LUT.mem_0_4 , n6921, \mem_LUT.mem_0_3 , 
        n6920, n6919, n6918, n2;
    wire [2:0]rd_addr_r_c;   // src/fifo_quad_word_mod.v(69[31:40])
    
    wire \mem_LUT.mem_0_0 , n6917, n5692, n5698, n6951, \mem_LUT.mem_3_7 , 
        n6950, \mem_LUT.mem_3_6 , n6949, \mem_LUT.mem_3_5 , n6948, 
        \mem_LUT.mem_3_4 , n6947, \mem_LUT.mem_3_3 , n6946, \mem_LUT.mem_3_2 , 
        n6945, n6944, \mem_LUT.mem_3_0 , n6940, \mem_LUT.mem_2_7 , 
        n6939, \mem_LUT.mem_2_6 , n6938, \mem_LUT.mem_2_5 , n6937, 
        \mem_LUT.mem_2_4 , n6936, \mem_LUT.mem_2_3 , n6935, \mem_LUT.mem_2_2 , 
        n6934, n6933, \mem_LUT.mem_2_0 , n6932, \mem_LUT.mem_1_7 , 
        n6931, \mem_LUT.mem_1_6 , n6930, \mem_LUT.mem_1_5 , n6929, 
        \mem_LUT.mem_1_4 , n6928, \mem_LUT.mem_1_3 , n6927, n6926, 
        n6925, \mem_LUT.mem_1_0 , n16257, n3, rd_fifo_en_prev_r, n16509, 
        n16491, n16485, n16467, n16443;
    
    SB_LUT4 n16311_bdd_4_lut (.I0(n16311), .I1(\mem_LUT.mem_1_2 ), .I2(\mem_LUT.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [2]));
    defparam n16311_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n12[0]), 
            .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i5425_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_0_7 ), .O(n6924));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5425_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14159 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_1 ), 
            .I2(\mem_LUT.mem_3_1 ), .I3(rd_addr_r[1]), .O(n16305));
    defparam rd_addr_r_0__bdd_4_lut_14159.LUT_INIT = 16'he4aa;
    SB_LUT4 i5424_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_0_6 ), .O(n6923));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5424_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \mem_LUT.data_raw_r__i1  (.Q(\mem_LUT.data_raw_r[0] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [0]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 n16305_bdd_4_lut (.I0(n16305), .I1(\mem_LUT.mem_1_1 ), .I2(\mem_LUT.mem_0_1 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [1]));
    defparam n16305_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(SLM_CLK_c), .D(n8), .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i5423_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_0_5 ), .O(n6922));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5423_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5422_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_0_4 ), .O(n6921));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5422_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5421_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_0_3 ), .O(n6920));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5421_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5420_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_0_2 ), .O(n6919));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5420_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5419_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_0_1 ), .O(n6918));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5419_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \mem_LUT.data_buff_r__i1  (.Q(\fifo_temp_output[1] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n7067));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 i1_2_lut (.I0(wr_addr_r[0]), .I1(rd_addr_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4566));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(n4566), .I1(\wr_addr_p1_w[2] ), .I2(n2), .I3(rd_addr_r_c[2]), 
            .O(n13820));
    defparam i1_4_lut.LUT_INIT = 16'h0208;
    SB_LUT4 i5418_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_0_0 ), .O(n6917));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5418_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \mem_LUT.data_buff_r__i2  (.Q(\fifo_temp_output[2] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n7064));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_buff_r__i3  (.Q(\fifo_temp_output[3] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n7061));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_buff_r__i4  (.Q(\fifo_temp_output[4] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n7058));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_buff_r__i5  (.Q(\fifo_temp_output[5] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n7055));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_buff_r__i6  (.Q(\fifo_temp_output[6] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n7052));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_buff_r__i7  (.Q(\fifo_temp_output[7] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n7049));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(SLM_CLK_c), .D(n5647));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(SLM_CLK_c), .D(n5658));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r_c[2]), .C(SLM_CLK_c), .D(n5692));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(n5698));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFE \mem_LUT.data_buff_r__i0  (.Q(\fifo_temp_output[0] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n6970));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE full_r_84 (.Q(is_tx_fifo_full_flag), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n14076));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF i347_348 (.Q(\mem_LUT.mem_3_7 ), .C(SLM_CLK_c), .D(n6951));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i344_345 (.Q(\mem_LUT.mem_3_6 ), .C(SLM_CLK_c), .D(n6950));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i341_342 (.Q(\mem_LUT.mem_3_5 ), .C(SLM_CLK_c), .D(n6949));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i338_339 (.Q(\mem_LUT.mem_3_4 ), .C(SLM_CLK_c), .D(n6948));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i335_336 (.Q(\mem_LUT.mem_3_3 ), .C(SLM_CLK_c), .D(n6947));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i332_333 (.Q(\mem_LUT.mem_3_2 ), .C(SLM_CLK_c), .D(n6946));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i329_330 (.Q(\mem_LUT.mem_3_1 ), .C(SLM_CLK_c), .D(n6945));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i326_327 (.Q(\mem_LUT.mem_3_0 ), .C(SLM_CLK_c), .D(n6944));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i251_252 (.Q(\mem_LUT.mem_2_7 ), .C(SLM_CLK_c), .D(n6940));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i248_249 (.Q(\mem_LUT.mem_2_6 ), .C(SLM_CLK_c), .D(n6939));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i245_246 (.Q(\mem_LUT.mem_2_5 ), .C(SLM_CLK_c), .D(n6938));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i242_243 (.Q(\mem_LUT.mem_2_4 ), .C(SLM_CLK_c), .D(n6937));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i239_240 (.Q(\mem_LUT.mem_2_3 ), .C(SLM_CLK_c), .D(n6936));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i236_237 (.Q(\mem_LUT.mem_2_2 ), .C(SLM_CLK_c), .D(n6935));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i233_234 (.Q(\mem_LUT.mem_2_1 ), .C(SLM_CLK_c), .D(n6934));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i230_231 (.Q(\mem_LUT.mem_2_0 ), .C(SLM_CLK_c), .D(n6933));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i155_156 (.Q(\mem_LUT.mem_1_7 ), .C(SLM_CLK_c), .D(n6932));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i152_153 (.Q(\mem_LUT.mem_1_6 ), .C(SLM_CLK_c), .D(n6931));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i149_150 (.Q(\mem_LUT.mem_1_5 ), .C(SLM_CLK_c), .D(n6930));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i146_147 (.Q(\mem_LUT.mem_1_4 ), .C(SLM_CLK_c), .D(n6929));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i143_144 (.Q(\mem_LUT.mem_1_3 ), .C(SLM_CLK_c), .D(n6928));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i140_141 (.Q(\mem_LUT.mem_1_2 ), .C(SLM_CLK_c), .D(n6927));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i137_138 (.Q(\mem_LUT.mem_1_1 ), .C(SLM_CLK_c), .D(n6926));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i134_135 (.Q(\mem_LUT.mem_1_0 ), .C(SLM_CLK_c), .D(n6925));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i59_60 (.Q(\mem_LUT.mem_0_7 ), .C(SLM_CLK_c), .D(n6924));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i56_57 (.Q(\mem_LUT.mem_0_6 ), .C(SLM_CLK_c), .D(n6923));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i53_54 (.Q(\mem_LUT.mem_0_5 ), .C(SLM_CLK_c), .D(n6922));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i50_51 (.Q(\mem_LUT.mem_0_4 ), .C(SLM_CLK_c), .D(n6921));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i47_48 (.Q(\mem_LUT.mem_0_3 ), .C(SLM_CLK_c), .D(n6920));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i44_45 (.Q(\mem_LUT.mem_0_2 ), .C(SLM_CLK_c), .D(n6919));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i41_42 (.Q(\mem_LUT.mem_0_1 ), .C(SLM_CLK_c), .D(n6918));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i38_39 (.Q(\mem_LUT.mem_0_0 ), .C(SLM_CLK_c), .D(n6917));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 i4199_4_lut_4_lut (.I0(rd_fifo_en_w), .I1(reset_all_w), .I2(\rd_addr_p1_w[1] ), 
            .I3(rd_addr_r[1]), .O(n5698));   // src/fifo_quad_word_mod.v(155[29] 160[32])
    defparam i4199_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4193_4_lut_4_lut (.I0(rd_fifo_en_w), .I1(reset_all_w), .I2(\rd_addr_p1_w[2] ), 
            .I3(rd_addr_r_c[2]), .O(n5692));   // src/fifo_quad_word_mod.v(155[29] 160[32])
    defparam i4193_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14154 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_0 ), 
            .I2(\mem_LUT.mem_3_0 ), .I3(rd_addr_r[1]), .O(n16257));
    defparam rd_addr_r_0__bdd_4_lut_14154.LUT_INIT = 16'he4aa;
    SB_LUT4 n16257_bdd_4_lut (.I0(n16257), .I1(\mem_LUT.mem_1_0 ), .I2(\mem_LUT.mem_0_0 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [0]));
    defparam n16257_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1760_2_lut (.I0(rd_addr_r[1]), .I1(rd_addr_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(\rd_addr_p1_w[1] ));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1760_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1767_3_lut (.I0(rd_addr_r_c[2]), .I1(rd_addr_r[1]), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(\rd_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1767_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1745_3_lut (.I0(wr_addr_r[2]), .I1(wr_addr_r[1]), .I2(wr_addr_r[0]), 
            .I3(GND_net), .O(\wr_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam i1745_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 wr_en_i_I_0_2_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(GND_net), .I3(GND_net), .O(wr_fifo_en_w));   // src/fifo_quad_word_mod.v(103[21:60])
    defparam wr_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5452_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_3_7 ), .O(n6951));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5452_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5451_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_3_6 ), .O(n6950));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5451_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE \mem_LUT.data_raw_r__i2  (.Q(\mem_LUT.data_raw_r[1] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [1]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i3  (.Q(\mem_LUT.data_raw_r[2] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [2]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i4  (.Q(\mem_LUT.data_raw_r[3] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [3]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i5  (.Q(\mem_LUT.data_raw_r[4] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [4]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i6  (.Q(\mem_LUT.data_raw_r[5] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [5]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i7  (.Q(\mem_LUT.data_raw_r[6] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [6]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i8  (.Q(\mem_LUT.data_raw_r[7] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1269 [7]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 i5450_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_3_5 ), .O(n6949));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5450_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5449_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_3_4 ), .O(n6948));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5449_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5448_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_3_3 ), .O(n6947));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5448_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5447_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_3_2 ), .O(n6946));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5447_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5446_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_3_1 ), .O(n6945));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5446_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5445_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_3_0 ), .O(n6944));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5445_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_en_i_I_0_2_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(GND_net), .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_quad_word_mod.v(62[29:51])
    defparam rd_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_DFF rd_fifo_en_prev_r_86 (.Q(rd_fifo_en_prev_r), .C(SLM_CLK_c), .D(n5664));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    SB_DFF empty_r_85 (.Q(is_fifo_empty_flag), .C(SLM_CLK_c), .D(n14096));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_7 ), 
            .I2(\mem_LUT.mem_3_7 ), .I3(rd_addr_r[1]), .O(n16509));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n16509_bdd_4_lut (.I0(n16509), .I1(\mem_LUT.mem_1_7 ), .I2(\mem_LUT.mem_0_7 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [7]));
    defparam n16509_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14324 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_6 ), 
            .I2(\mem_LUT.mem_3_6 ), .I3(rd_addr_r[1]), .O(n16491));
    defparam rd_addr_r_0__bdd_4_lut_14324.LUT_INIT = 16'he4aa;
    SB_LUT4 n16491_bdd_4_lut (.I0(n16491), .I1(\mem_LUT.mem_1_6 ), .I2(\mem_LUT.mem_0_6 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [6]));
    defparam n16491_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14309 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_5 ), 
            .I2(\mem_LUT.mem_3_5 ), .I3(rd_addr_r[1]), .O(n16485));
    defparam rd_addr_r_0__bdd_4_lut_14309.LUT_INIT = 16'he4aa;
    SB_LUT4 n16485_bdd_4_lut (.I0(n16485), .I1(\mem_LUT.mem_1_5 ), .I2(\mem_LUT.mem_0_5 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [5]));
    defparam n16485_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14304 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_4 ), 
            .I2(\mem_LUT.mem_3_4 ), .I3(rd_addr_r[1]), .O(n16467));
    defparam rd_addr_r_0__bdd_4_lut_14304.LUT_INIT = 16'he4aa;
    SB_LUT4 n16467_bdd_4_lut (.I0(n16467), .I1(\mem_LUT.mem_1_4 ), .I2(\mem_LUT.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [4]));
    defparam n16467_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14289 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_3 ), 
            .I2(\mem_LUT.mem_3_3 ), .I3(rd_addr_r[1]), .O(n16443));
    defparam rd_addr_r_0__bdd_4_lut_14289.LUT_INIT = 16'he4aa;
    SB_LUT4 n16443_bdd_4_lut (.I0(n16443), .I1(\mem_LUT.mem_1_3 ), .I2(\mem_LUT.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1269 [3]));
    defparam n16443_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5441_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_2_7 ), .O(n6940));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5441_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5440_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_2_6 ), .O(n6939));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5440_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5439_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_2_5 ), .O(n6938));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5439_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5438_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_2_4 ), .O(n6937));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5438_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5437_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_2_3 ), .O(n6936));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5437_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5436_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_2_2 ), .O(n6935));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5436_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5435_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_2_1 ), .O(n6934));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5435_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5434_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_2_0 ), .O(n6933));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5434_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5433_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_1_7 ), .O(n6932));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5433_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_p1_w_1__I_0_i2_2_lut_3_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[0]), 
            .I2(rd_addr_r[1]), .I3(GND_net), .O(n2));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam wr_addr_p1_w_1__I_0_i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5432_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_1_6 ), .O(n6931));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5432_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5431_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_1_5 ), .O(n6930));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5431_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5430_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_1_4 ), .O(n6929));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5430_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5429_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_1_3 ), .O(n6928));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5429_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5428_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_1_2 ), .O(n6927));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5428_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5427_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_1_1 ), .O(n6926));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5427_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14269 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_2 ), 
            .I2(\mem_LUT.mem_3_2 ), .I3(rd_addr_r[1]), .O(n16311));
    defparam rd_addr_r_0__bdd_4_lut_14269.LUT_INIT = 16'he4aa;
    SB_LUT4 i5426_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_1_0 ), .O(n6925));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i5426_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1970_2_lut_3_lut_4_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(reset_all_w), .I3(rd_addr_r[0]), .O(n12[0]));   // src/fifo_quad_word_mod.v(155[29] 160[32])
    defparam i1970_2_lut_3_lut_4_lut.LUT_INIT = 16'h0df2;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(reset_all_w), .I3(rd_fifo_en_prev_r), .O(n5207));   // src/fifo_quad_word_mod.v(155[29] 160[32])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff2;
    SB_LUT4 EnabledDecoder_2_i3_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n3));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i3_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i4_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n4));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i4_2_lut_3_lut.LUT_INIT = 16'h0202;
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen2
//

module fifo_dc_32_lut_gen2 (dc32_fifo_data_in, FIFO_CLK_c, GND_net, \REG.mem_22_29 , 
            \REG.mem_23_29 , \REG.mem_21_29 , \REG.mem_11_15 , \REG.mem_11_11 , 
            \REG.mem_6_26 , \REG.mem_7_26 , dc32_fifo_almost_full, reset_per_frame, 
            \REG.mem_5_26 , rd_fifo_en_w, dc32_fifo_data_out, SLM_CLK_c, 
            \REG.mem_27_29 , \REG.mem_11_8 , \REG.mem_22_5 , \REG.mem_23_5 , 
            rd_grey_sync_r, \REG.mem_21_5 , dc32_fifo_full, \REG.mem_6_20 , 
            \REG.mem_7_20 , empty_nxt_c_N_636, dc32_fifo_empty, \REG.mem_5_20 , 
            \wr_grey_sync_r[0] , \aempty_flag_impl.ae_flag_nxt_w , \rd_addr_nxt_c_5__N_573[3] , 
            \rd_addr_nxt_c_5__N_573[1] , \REG.mem_11_20 , \REG.mem_11_21 , 
            \REG.mem_27_12 , \REG.mem_22_11 , \REG.mem_23_11 , \REG.mem_21_11 , 
            \REG.mem_27_3 , \REG.mem_11_10 , \REG.mem_22_28 , \REG.mem_23_28 , 
            \REG.mem_21_28 , \REG.mem_27_0 , \REG.mem_6_19 , \REG.mem_7_19 , 
            \REG.mem_5_19 , \REG.mem_6_9 , \REG.mem_7_9 , \REG.mem_11_0 , 
            \REG.mem_5_9 , \REG.mem_11_13 , \REG.mem_6_14 , \REG.mem_7_14 , 
            \REG.mem_5_14 , \REG.mem_22_19 , \REG.mem_23_19 , \REG.mem_21_19 , 
            \REG.mem_27_19 , n6, n22, \REG.mem_11_14 , \REG.mem_22_9 , 
            \REG.mem_23_9 , \REG.mem_21_9 , \REG.mem_6_24 , \REG.mem_7_24 , 
            \REG.mem_22_1 , \REG.mem_23_1 , wr_fifo_en_w, \wr_addr_nxt_c[4] , 
            \wr_addr_nxt_c[2] , \REG.mem_22_16 , \REG.mem_23_16 , \REG.mem_21_1 , 
            \REG.mem_21_16 , \REG.mem_11_12 , \REG.mem_5_24 , n7038, 
            n7037, n7036, n7035, n7034, n7033, wp_sync1_r, n7032, 
            n7031, n7030, n7029, n7028, n7027, n7025, n7023, n7022, 
            n7021, n7020, n7019, n7018, rp_sync1_r, n7017, n7016, 
            n7015, n7014, n6955, n6953, \wr_addr_r[5] , n6532, \REG.mem_27_31 , 
            n6531, \REG.mem_27_30 , n6530, n6529, \REG.mem_27_28 , 
            n6528, \REG.mem_27_27 , n6527, \REG.mem_27_26 , n6526, 
            \REG.mem_27_25 , n6525, \REG.mem_27_24 , n6524, \REG.mem_27_23 , 
            n6523, \REG.mem_27_22 , n6522, \REG.mem_27_21 , n6521, 
            \REG.mem_27_20 , n6520, n6519, \REG.mem_27_18 , n6518, 
            \REG.mem_27_17 , n6517, \REG.mem_27_16 , n6516, \REG.mem_27_15 , 
            n6515, \REG.mem_27_14 , n6514, \REG.mem_27_13 , n6513, 
            n6512, \REG.mem_27_11 , n6511, \REG.mem_27_10 , n6510, 
            \REG.mem_27_9 , n6509, \REG.mem_27_8 , n6508, \REG.mem_27_7 , 
            n6507, \REG.mem_27_6 , n6506, \REG.mem_27_5 , n6505, \REG.mem_27_4 , 
            n6504, n6503, \REG.mem_27_2 , n6502, \REG.mem_27_1 , n6501, 
            n6404, \REG.mem_23_31 , n6403, \REG.mem_23_30 , n6402, 
            n6401, n6400, \REG.mem_23_27 , n6399, \REG.mem_23_26 , 
            n6398, \REG.mem_23_25 , n6397, \REG.mem_23_24 , n6396, 
            \REG.mem_23_23 , n6395, \REG.mem_23_22 , n6394, \REG.mem_23_21 , 
            n6393, \REG.mem_23_20 , n6392, n6391, \REG.mem_23_18 , 
            n6390, \REG.mem_23_17 , n6389, n6388, \REG.mem_23_15 , 
            n6387, \REG.mem_23_14 , n6386, \REG.mem_23_13 , n6385, 
            \REG.mem_23_12 , n6384, n6383, \REG.mem_23_10 , n6382, 
            n6381, \REG.mem_23_8 , n6380, \REG.mem_23_7 , n6379, \REG.mem_23_6 , 
            n6378, n6377, \REG.mem_23_4 , n6376, \REG.mem_23_3 , n6375, 
            \REG.mem_23_2 , n6374, n6373, \REG.mem_23_0 , n6372, \REG.mem_22_31 , 
            n6371, \REG.mem_22_30 , n6370, n6369, n6368, \REG.mem_22_27 , 
            n6367, \REG.mem_22_26 , n6366, \REG.mem_22_25 , n6365, 
            \REG.mem_22_24 , n6364, \REG.mem_22_23 , n6363, \REG.mem_22_22 , 
            n6362, \REG.mem_22_21 , n6361, \REG.mem_22_20 , n6360, 
            n6359, \REG.mem_22_18 , n6358, \REG.mem_22_17 , n6357, 
            n6356, \REG.mem_22_15 , n6355, \REG.mem_22_14 , n6354, 
            \REG.mem_22_13 , n6353, \REG.mem_22_12 , n6352, n6351, 
            \REG.mem_22_10 , n6350, n6349, \REG.mem_22_8 , n6348, 
            \REG.mem_22_7 , n6347, \REG.mem_22_6 , n6346, n6345, \REG.mem_22_4 , 
            n6344, \REG.mem_22_3 , n6343, \REG.mem_22_2 , n6342, n6341, 
            \REG.mem_22_0 , n6340, \REG.mem_21_31 , n6339, \REG.mem_21_30 , 
            n6338, n6337, n6336, \REG.mem_21_27 , n6335, \REG.mem_21_26 , 
            n6334, \REG.mem_21_25 , n6333, \REG.mem_21_24 , n6332, 
            \REG.mem_21_23 , n6331, \REG.mem_21_22 , n6330, \REG.mem_21_21 , 
            n6329, \REG.mem_21_20 , n6328, n6327, \REG.mem_21_18 , 
            n6326, \REG.mem_21_17 , n6325, n6324, \REG.mem_21_15 , 
            n6323, \REG.mem_21_14 , n6322, \REG.mem_21_13 , n6321, 
            \REG.mem_21_12 , n6320, n6319, \REG.mem_21_10 , n6318, 
            n6317, \REG.mem_21_8 , n6316, \REG.mem_21_7 , n6315, \REG.mem_21_6 , 
            n6314, n6313, \REG.mem_21_4 , n6312, \REG.mem_21_3 , n6311, 
            \REG.mem_21_2 , n6310, n6309, \REG.mem_21_0 , n12, n10, 
            n26, \rd_addr_nxt_c_5__N_573[4] , \REG.mem_6_22 , \REG.mem_7_22 , 
            \REG.mem_6_23 , \REG.mem_7_23 , \REG.mem_5_23 , \REG.mem_5_22 , 
            \REG.mem_11_23 , \REG.mem_11_18 , \REG.mem_6_7 , \REG.mem_7_7 , 
            \REG.mem_5_7 , \REG.mem_11_9 , n7, \REG.mem_6_28 , \REG.mem_7_28 , 
            \REG.mem_5_28 , n8, \REG.mem_11_28 , VCC_net, n25, \REG.mem_11_25 , 
            \wr_grey_sync_r[1] , \wr_grey_sync_r[2] , \REG.mem_11_5 , 
            \wr_grey_sync_r[3] , \wr_grey_sync_r[4] , n6020, \REG.mem_11_31 , 
            n6019, \REG.mem_11_30 , n6018, \REG.mem_11_29 , n6017, 
            n6016, \REG.mem_11_27 , n6015, \REG.mem_11_26 , n6014, 
            n6013, \REG.mem_11_24 , n6012, n6011, \REG.mem_11_22 , 
            n6010, n6009, n6008, \REG.mem_11_19 , n6007, \REG.mem_11_6 , 
            n6006, \REG.mem_11_17 , n6005, \REG.mem_11_16 , n6004, 
            n6003, n6002, n6001, n6000, n5999, n5998, \wr_addr_r[0] , 
            DEBUG_5_c, \REG.mem_11_2 , n5997, n5996, \REG.mem_11_7 , 
            n5995, n5994, n5993, \REG.mem_11_4 , \wr_addr_p1_w[0] , 
            n13865, n14706, n5992, \REG.mem_11_3 , n5991, n5990, 
            \REG.mem_11_1 , FT_OE_N_496, n12_adj_4, dc32_fifo_read_enable, 
            n5989, n5892, \REG.mem_7_31 , n5891, \REG.mem_7_30 , n5890, 
            \REG.mem_7_29 , n5889, n5888, \REG.mem_7_27 , n5887, n5886, 
            \REG.mem_7_25 , n5885, n5884, n5883, n5882, \REG.mem_7_21 , 
            n5881, n5880, n5879, \REG.mem_7_18 , n5878, \REG.mem_7_17 , 
            n5877, \REG.mem_7_16 , n5876, \REG.mem_7_15 , n5875, n5874, 
            \REG.mem_7_13 , n5873, \REG.mem_7_12 , n5872, \REG.mem_7_11 , 
            n5871, \REG.mem_7_10 , n5870, n5869, \REG.mem_7_8 , n5868, 
            n5867, \REG.mem_7_6 , n5866, \REG.mem_7_5 , n5865, \REG.mem_7_4 , 
            n5864, \REG.mem_7_3 , n5863, \REG.mem_7_2 , n5862, \REG.mem_7_1 , 
            n5861, \REG.mem_7_0 , n5860, \REG.mem_6_31 , n5859, \REG.mem_6_30 , 
            n5858, \REG.mem_6_29 , n5857, n5856, \REG.mem_6_27 , n5855, 
            n5854, \REG.mem_6_25 , n5853, n5852, n5851, \state[3] , 
            n4843, n1224, n5850, \REG.mem_6_21 , n5849, n5848, n5847, 
            \REG.mem_6_18 , n5846, \REG.mem_6_17 , n5845, \REG.mem_6_16 , 
            n5844, \REG.mem_6_15 , n5843, n5842, \REG.mem_6_13 , n5841, 
            \REG.mem_6_12 , n5840, \REG.mem_6_11 , n5839, \REG.mem_6_10 , 
            n5838, n5837, \REG.mem_6_8 , n5836, n5835, \REG.mem_6_6 , 
            n5834, \REG.mem_6_5 , n5833, \REG.mem_6_4 , \REG.mem_6_2 , 
            n5832, \REG.mem_6_3 , n5831, \REG.mem_5_2 , n5830, \REG.mem_6_1 , 
            n5829, \REG.mem_6_0 , n5828, \REG.mem_5_31 , n5827, \REG.mem_5_30 , 
            n5826, \REG.mem_5_29 , n5825, n5824, \REG.mem_5_27 , n5823, 
            n5822, \REG.mem_5_25 , n5821, n5820, n5819, n5818, \REG.mem_5_21 , 
            n5817, n5816, n5815, \REG.mem_5_18 , n5814, \REG.mem_5_17 , 
            n5813, \REG.mem_5_16 , n5812, \REG.mem_5_15 , n5811, n5810, 
            \REG.mem_5_13 , n5809, \REG.mem_5_12 , n5808, \REG.mem_5_11 , 
            n5807, \REG.mem_5_10 , n5806, n5805, \REG.mem_5_8 , n5804, 
            n5803, \REG.mem_5_6 , n5802, \REG.mem_5_5 , n5648, n5801, 
            \REG.mem_5_4 , n5800, \REG.mem_5_3 , n5642, n5639, n5638, 
            n5799, n5798, \REG.mem_5_1 , n5797, \REG.mem_5_0 , n5605, 
            n27, n11, n28) /* synthesis syn_module_defined=1 */ ;
    input [31:0]dc32_fifo_data_in;
    input FIFO_CLK_c;
    input GND_net;
    output \REG.mem_22_29 ;
    output \REG.mem_23_29 ;
    output \REG.mem_21_29 ;
    output \REG.mem_11_15 ;
    output \REG.mem_11_11 ;
    output \REG.mem_6_26 ;
    output \REG.mem_7_26 ;
    output dc32_fifo_almost_full;
    input reset_per_frame;
    output \REG.mem_5_26 ;
    output rd_fifo_en_w;
    output [31:0]dc32_fifo_data_out;
    input SLM_CLK_c;
    output \REG.mem_27_29 ;
    output \REG.mem_11_8 ;
    output \REG.mem_22_5 ;
    output \REG.mem_23_5 ;
    output [5:0]rd_grey_sync_r;
    output \REG.mem_21_5 ;
    output dc32_fifo_full;
    output \REG.mem_6_20 ;
    output \REG.mem_7_20 ;
    input empty_nxt_c_N_636;
    output dc32_fifo_empty;
    output \REG.mem_5_20 ;
    output \wr_grey_sync_r[0] ;
    input \aempty_flag_impl.ae_flag_nxt_w ;
    output \rd_addr_nxt_c_5__N_573[3] ;
    output \rd_addr_nxt_c_5__N_573[1] ;
    output \REG.mem_11_20 ;
    output \REG.mem_11_21 ;
    output \REG.mem_27_12 ;
    output \REG.mem_22_11 ;
    output \REG.mem_23_11 ;
    output \REG.mem_21_11 ;
    output \REG.mem_27_3 ;
    output \REG.mem_11_10 ;
    output \REG.mem_22_28 ;
    output \REG.mem_23_28 ;
    output \REG.mem_21_28 ;
    output \REG.mem_27_0 ;
    output \REG.mem_6_19 ;
    output \REG.mem_7_19 ;
    output \REG.mem_5_19 ;
    output \REG.mem_6_9 ;
    output \REG.mem_7_9 ;
    output \REG.mem_11_0 ;
    output \REG.mem_5_9 ;
    output \REG.mem_11_13 ;
    output \REG.mem_6_14 ;
    output \REG.mem_7_14 ;
    output \REG.mem_5_14 ;
    output \REG.mem_22_19 ;
    output \REG.mem_23_19 ;
    output \REG.mem_21_19 ;
    output \REG.mem_27_19 ;
    output n6;
    output n22;
    output \REG.mem_11_14 ;
    output \REG.mem_22_9 ;
    output \REG.mem_23_9 ;
    output \REG.mem_21_9 ;
    output \REG.mem_6_24 ;
    output \REG.mem_7_24 ;
    output \REG.mem_22_1 ;
    output \REG.mem_23_1 ;
    input wr_fifo_en_w;
    output \wr_addr_nxt_c[4] ;
    output \wr_addr_nxt_c[2] ;
    output \REG.mem_22_16 ;
    output \REG.mem_23_16 ;
    output \REG.mem_21_1 ;
    output \REG.mem_21_16 ;
    output \REG.mem_11_12 ;
    output \REG.mem_5_24 ;
    input n7038;
    input n7037;
    input n7036;
    input n7035;
    input n7034;
    input n7033;
    output [5:0]wp_sync1_r;
    input n7032;
    input n7031;
    input n7030;
    input n7029;
    input n7028;
    input n7027;
    input n7025;
    input n7023;
    input n7022;
    input n7021;
    input n7020;
    input n7019;
    input n7018;
    output [5:0]rp_sync1_r;
    input n7017;
    input n7016;
    input n7015;
    input n7014;
    input n6955;
    input n6953;
    output \wr_addr_r[5] ;
    input n6532;
    output \REG.mem_27_31 ;
    input n6531;
    output \REG.mem_27_30 ;
    input n6530;
    input n6529;
    output \REG.mem_27_28 ;
    input n6528;
    output \REG.mem_27_27 ;
    input n6527;
    output \REG.mem_27_26 ;
    input n6526;
    output \REG.mem_27_25 ;
    input n6525;
    output \REG.mem_27_24 ;
    input n6524;
    output \REG.mem_27_23 ;
    input n6523;
    output \REG.mem_27_22 ;
    input n6522;
    output \REG.mem_27_21 ;
    input n6521;
    output \REG.mem_27_20 ;
    input n6520;
    input n6519;
    output \REG.mem_27_18 ;
    input n6518;
    output \REG.mem_27_17 ;
    input n6517;
    output \REG.mem_27_16 ;
    input n6516;
    output \REG.mem_27_15 ;
    input n6515;
    output \REG.mem_27_14 ;
    input n6514;
    output \REG.mem_27_13 ;
    input n6513;
    input n6512;
    output \REG.mem_27_11 ;
    input n6511;
    output \REG.mem_27_10 ;
    input n6510;
    output \REG.mem_27_9 ;
    input n6509;
    output \REG.mem_27_8 ;
    input n6508;
    output \REG.mem_27_7 ;
    input n6507;
    output \REG.mem_27_6 ;
    input n6506;
    output \REG.mem_27_5 ;
    input n6505;
    output \REG.mem_27_4 ;
    input n6504;
    input n6503;
    output \REG.mem_27_2 ;
    input n6502;
    output \REG.mem_27_1 ;
    input n6501;
    input n6404;
    output \REG.mem_23_31 ;
    input n6403;
    output \REG.mem_23_30 ;
    input n6402;
    input n6401;
    input n6400;
    output \REG.mem_23_27 ;
    input n6399;
    output \REG.mem_23_26 ;
    input n6398;
    output \REG.mem_23_25 ;
    input n6397;
    output \REG.mem_23_24 ;
    input n6396;
    output \REG.mem_23_23 ;
    input n6395;
    output \REG.mem_23_22 ;
    input n6394;
    output \REG.mem_23_21 ;
    input n6393;
    output \REG.mem_23_20 ;
    input n6392;
    input n6391;
    output \REG.mem_23_18 ;
    input n6390;
    output \REG.mem_23_17 ;
    input n6389;
    input n6388;
    output \REG.mem_23_15 ;
    input n6387;
    output \REG.mem_23_14 ;
    input n6386;
    output \REG.mem_23_13 ;
    input n6385;
    output \REG.mem_23_12 ;
    input n6384;
    input n6383;
    output \REG.mem_23_10 ;
    input n6382;
    input n6381;
    output \REG.mem_23_8 ;
    input n6380;
    output \REG.mem_23_7 ;
    input n6379;
    output \REG.mem_23_6 ;
    input n6378;
    input n6377;
    output \REG.mem_23_4 ;
    input n6376;
    output \REG.mem_23_3 ;
    input n6375;
    output \REG.mem_23_2 ;
    input n6374;
    input n6373;
    output \REG.mem_23_0 ;
    input n6372;
    output \REG.mem_22_31 ;
    input n6371;
    output \REG.mem_22_30 ;
    input n6370;
    input n6369;
    input n6368;
    output \REG.mem_22_27 ;
    input n6367;
    output \REG.mem_22_26 ;
    input n6366;
    output \REG.mem_22_25 ;
    input n6365;
    output \REG.mem_22_24 ;
    input n6364;
    output \REG.mem_22_23 ;
    input n6363;
    output \REG.mem_22_22 ;
    input n6362;
    output \REG.mem_22_21 ;
    input n6361;
    output \REG.mem_22_20 ;
    input n6360;
    input n6359;
    output \REG.mem_22_18 ;
    input n6358;
    output \REG.mem_22_17 ;
    input n6357;
    input n6356;
    output \REG.mem_22_15 ;
    input n6355;
    output \REG.mem_22_14 ;
    input n6354;
    output \REG.mem_22_13 ;
    input n6353;
    output \REG.mem_22_12 ;
    input n6352;
    input n6351;
    output \REG.mem_22_10 ;
    input n6350;
    input n6349;
    output \REG.mem_22_8 ;
    input n6348;
    output \REG.mem_22_7 ;
    input n6347;
    output \REG.mem_22_6 ;
    input n6346;
    input n6345;
    output \REG.mem_22_4 ;
    input n6344;
    output \REG.mem_22_3 ;
    input n6343;
    output \REG.mem_22_2 ;
    input n6342;
    input n6341;
    output \REG.mem_22_0 ;
    input n6340;
    output \REG.mem_21_31 ;
    input n6339;
    output \REG.mem_21_30 ;
    input n6338;
    input n6337;
    input n6336;
    output \REG.mem_21_27 ;
    input n6335;
    output \REG.mem_21_26 ;
    input n6334;
    output \REG.mem_21_25 ;
    input n6333;
    output \REG.mem_21_24 ;
    input n6332;
    output \REG.mem_21_23 ;
    input n6331;
    output \REG.mem_21_22 ;
    input n6330;
    output \REG.mem_21_21 ;
    input n6329;
    output \REG.mem_21_20 ;
    input n6328;
    input n6327;
    output \REG.mem_21_18 ;
    input n6326;
    output \REG.mem_21_17 ;
    input n6325;
    input n6324;
    output \REG.mem_21_15 ;
    input n6323;
    output \REG.mem_21_14 ;
    input n6322;
    output \REG.mem_21_13 ;
    input n6321;
    output \REG.mem_21_12 ;
    input n6320;
    input n6319;
    output \REG.mem_21_10 ;
    input n6318;
    input n6317;
    output \REG.mem_21_8 ;
    input n6316;
    output \REG.mem_21_7 ;
    input n6315;
    output \REG.mem_21_6 ;
    input n6314;
    input n6313;
    output \REG.mem_21_4 ;
    input n6312;
    output \REG.mem_21_3 ;
    input n6311;
    output \REG.mem_21_2 ;
    input n6310;
    input n6309;
    output \REG.mem_21_0 ;
    output n12;
    output n10;
    output n26;
    output \rd_addr_nxt_c_5__N_573[4] ;
    output \REG.mem_6_22 ;
    output \REG.mem_7_22 ;
    output \REG.mem_6_23 ;
    output \REG.mem_7_23 ;
    output \REG.mem_5_23 ;
    output \REG.mem_5_22 ;
    output \REG.mem_11_23 ;
    output \REG.mem_11_18 ;
    output \REG.mem_6_7 ;
    output \REG.mem_7_7 ;
    output \REG.mem_5_7 ;
    output \REG.mem_11_9 ;
    output n7;
    output \REG.mem_6_28 ;
    output \REG.mem_7_28 ;
    output \REG.mem_5_28 ;
    output n8;
    output \REG.mem_11_28 ;
    input VCC_net;
    input n25;
    output \REG.mem_11_25 ;
    output \wr_grey_sync_r[1] ;
    output \wr_grey_sync_r[2] ;
    output \REG.mem_11_5 ;
    output \wr_grey_sync_r[3] ;
    output \wr_grey_sync_r[4] ;
    input n6020;
    output \REG.mem_11_31 ;
    input n6019;
    output \REG.mem_11_30 ;
    input n6018;
    output \REG.mem_11_29 ;
    input n6017;
    input n6016;
    output \REG.mem_11_27 ;
    input n6015;
    output \REG.mem_11_26 ;
    input n6014;
    input n6013;
    output \REG.mem_11_24 ;
    input n6012;
    input n6011;
    output \REG.mem_11_22 ;
    input n6010;
    input n6009;
    input n6008;
    output \REG.mem_11_19 ;
    input n6007;
    output \REG.mem_11_6 ;
    input n6006;
    output \REG.mem_11_17 ;
    input n6005;
    output \REG.mem_11_16 ;
    input n6004;
    input n6003;
    input n6002;
    input n6001;
    input n6000;
    input n5999;
    input n5998;
    output \wr_addr_r[0] ;
    input DEBUG_5_c;
    output \REG.mem_11_2 ;
    input n5997;
    input n5996;
    output \REG.mem_11_7 ;
    input n5995;
    input n5994;
    input n5993;
    output \REG.mem_11_4 ;
    output \wr_addr_p1_w[0] ;
    output n13865;
    output n14706;
    input n5992;
    output \REG.mem_11_3 ;
    input n5991;
    input n5990;
    output \REG.mem_11_1 ;
    input FT_OE_N_496;
    output n12_adj_4;
    input dc32_fifo_read_enable;
    input n5989;
    input n5892;
    output \REG.mem_7_31 ;
    input n5891;
    output \REG.mem_7_30 ;
    input n5890;
    output \REG.mem_7_29 ;
    input n5889;
    input n5888;
    output \REG.mem_7_27 ;
    input n5887;
    input n5886;
    output \REG.mem_7_25 ;
    input n5885;
    input n5884;
    input n5883;
    input n5882;
    output \REG.mem_7_21 ;
    input n5881;
    input n5880;
    input n5879;
    output \REG.mem_7_18 ;
    input n5878;
    output \REG.mem_7_17 ;
    input n5877;
    output \REG.mem_7_16 ;
    input n5876;
    output \REG.mem_7_15 ;
    input n5875;
    input n5874;
    output \REG.mem_7_13 ;
    input n5873;
    output \REG.mem_7_12 ;
    input n5872;
    output \REG.mem_7_11 ;
    input n5871;
    output \REG.mem_7_10 ;
    input n5870;
    input n5869;
    output \REG.mem_7_8 ;
    input n5868;
    input n5867;
    output \REG.mem_7_6 ;
    input n5866;
    output \REG.mem_7_5 ;
    input n5865;
    output \REG.mem_7_4 ;
    input n5864;
    output \REG.mem_7_3 ;
    input n5863;
    output \REG.mem_7_2 ;
    input n5862;
    output \REG.mem_7_1 ;
    input n5861;
    output \REG.mem_7_0 ;
    input n5860;
    output \REG.mem_6_31 ;
    input n5859;
    output \REG.mem_6_30 ;
    input n5858;
    output \REG.mem_6_29 ;
    input n5857;
    input n5856;
    output \REG.mem_6_27 ;
    input n5855;
    input n5854;
    output \REG.mem_6_25 ;
    input n5853;
    input n5852;
    input n5851;
    input \state[3] ;
    input n4843;
    output n1224;
    input n5850;
    output \REG.mem_6_21 ;
    input n5849;
    input n5848;
    input n5847;
    output \REG.mem_6_18 ;
    input n5846;
    output \REG.mem_6_17 ;
    input n5845;
    output \REG.mem_6_16 ;
    input n5844;
    output \REG.mem_6_15 ;
    input n5843;
    input n5842;
    output \REG.mem_6_13 ;
    input n5841;
    output \REG.mem_6_12 ;
    input n5840;
    output \REG.mem_6_11 ;
    input n5839;
    output \REG.mem_6_10 ;
    input n5838;
    input n5837;
    output \REG.mem_6_8 ;
    input n5836;
    input n5835;
    output \REG.mem_6_6 ;
    input n5834;
    output \REG.mem_6_5 ;
    input n5833;
    output \REG.mem_6_4 ;
    output \REG.mem_6_2 ;
    input n5832;
    output \REG.mem_6_3 ;
    input n5831;
    output \REG.mem_5_2 ;
    input n5830;
    output \REG.mem_6_1 ;
    input n5829;
    output \REG.mem_6_0 ;
    input n5828;
    output \REG.mem_5_31 ;
    input n5827;
    output \REG.mem_5_30 ;
    input n5826;
    output \REG.mem_5_29 ;
    input n5825;
    input n5824;
    output \REG.mem_5_27 ;
    input n5823;
    input n5822;
    output \REG.mem_5_25 ;
    input n5821;
    input n5820;
    input n5819;
    input n5818;
    output \REG.mem_5_21 ;
    input n5817;
    input n5816;
    input n5815;
    output \REG.mem_5_18 ;
    input n5814;
    output \REG.mem_5_17 ;
    input n5813;
    output \REG.mem_5_16 ;
    input n5812;
    output \REG.mem_5_15 ;
    input n5811;
    input n5810;
    output \REG.mem_5_13 ;
    input n5809;
    output \REG.mem_5_12 ;
    input n5808;
    output \REG.mem_5_11 ;
    input n5807;
    output \REG.mem_5_10 ;
    input n5806;
    input n5805;
    output \REG.mem_5_8 ;
    input n5804;
    input n5803;
    output \REG.mem_5_6 ;
    input n5802;
    output \REG.mem_5_5 ;
    input n5648;
    input n5801;
    output \REG.mem_5_4 ;
    input n5800;
    output \REG.mem_5_3 ;
    input n5642;
    input n5639;
    input n5638;
    input n5799;
    input n5798;
    output \REG.mem_5_1 ;
    input n5797;
    output \REG.mem_5_0 ;
    input n5605;
    output n27;
    output n11;
    output n28;
    
    wire FIFO_CLK_c /* synthesis SET_AS_NETWORK=FIFO_CLK_c, is_clock=1 */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 lscc_fifo_dc_inst (.dc32_fifo_data_in({dc32_fifo_data_in}), 
            .FIFO_CLK_c(FIFO_CLK_c), .GND_net(GND_net), .\REG.mem_22_29 (\REG.mem_22_29 ), 
            .\REG.mem_23_29 (\REG.mem_23_29 ), .\REG.mem_21_29 (\REG.mem_21_29 ), 
            .\REG.mem_11_15 (\REG.mem_11_15 ), .\REG.mem_11_11 (\REG.mem_11_11 ), 
            .\REG.mem_6_26 (\REG.mem_6_26 ), .\REG.mem_7_26 (\REG.mem_7_26 ), 
            .dc32_fifo_almost_full(dc32_fifo_almost_full), .reset_per_frame(reset_per_frame), 
            .\REG.mem_5_26 (\REG.mem_5_26 ), .rd_fifo_en_w(rd_fifo_en_w), 
            .dc32_fifo_data_out({dc32_fifo_data_out}), .SLM_CLK_c(SLM_CLK_c), 
            .\REG.mem_27_29 (\REG.mem_27_29 ), .\REG.mem_11_8 (\REG.mem_11_8 ), 
            .\REG.mem_22_5 (\REG.mem_22_5 ), .\REG.mem_23_5 (\REG.mem_23_5 ), 
            .rd_grey_sync_r({rd_grey_sync_r}), .\REG.mem_21_5 (\REG.mem_21_5 ), 
            .dc32_fifo_full(dc32_fifo_full), .\REG.mem_6_20 (\REG.mem_6_20 ), 
            .\REG.mem_7_20 (\REG.mem_7_20 ), .empty_nxt_c_N_636(empty_nxt_c_N_636), 
            .dc32_fifo_empty(dc32_fifo_empty), .\REG.mem_5_20 (\REG.mem_5_20 ), 
            .\wr_grey_sync_r[0] (\wr_grey_sync_r[0] ), .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .\rd_addr_nxt_c_5__N_573[3] (\rd_addr_nxt_c_5__N_573[3] ), .\rd_addr_nxt_c_5__N_573[1] (\rd_addr_nxt_c_5__N_573[1] ), 
            .\REG.mem_11_20 (\REG.mem_11_20 ), .\REG.mem_11_21 (\REG.mem_11_21 ), 
            .\REG.mem_27_12 (\REG.mem_27_12 ), .\REG.mem_22_11 (\REG.mem_22_11 ), 
            .\REG.mem_23_11 (\REG.mem_23_11 ), .\REG.mem_21_11 (\REG.mem_21_11 ), 
            .\REG.mem_27_3 (\REG.mem_27_3 ), .\REG.mem_11_10 (\REG.mem_11_10 ), 
            .\REG.mem_22_28 (\REG.mem_22_28 ), .\REG.mem_23_28 (\REG.mem_23_28 ), 
            .\REG.mem_21_28 (\REG.mem_21_28 ), .\REG.mem_27_0 (\REG.mem_27_0 ), 
            .\REG.mem_6_19 (\REG.mem_6_19 ), .\REG.mem_7_19 (\REG.mem_7_19 ), 
            .\REG.mem_5_19 (\REG.mem_5_19 ), .\REG.mem_6_9 (\REG.mem_6_9 ), 
            .\REG.mem_7_9 (\REG.mem_7_9 ), .\REG.mem_11_0 (\REG.mem_11_0 ), 
            .\REG.mem_5_9 (\REG.mem_5_9 ), .\REG.mem_11_13 (\REG.mem_11_13 ), 
            .\REG.mem_6_14 (\REG.mem_6_14 ), .\REG.mem_7_14 (\REG.mem_7_14 ), 
            .\REG.mem_5_14 (\REG.mem_5_14 ), .\REG.mem_22_19 (\REG.mem_22_19 ), 
            .\REG.mem_23_19 (\REG.mem_23_19 ), .\REG.mem_21_19 (\REG.mem_21_19 ), 
            .\REG.mem_27_19 (\REG.mem_27_19 ), .n6(n6), .n22(n22), .\REG.mem_11_14 (\REG.mem_11_14 ), 
            .\REG.mem_22_9 (\REG.mem_22_9 ), .\REG.mem_23_9 (\REG.mem_23_9 ), 
            .\REG.mem_21_9 (\REG.mem_21_9 ), .\REG.mem_6_24 (\REG.mem_6_24 ), 
            .\REG.mem_7_24 (\REG.mem_7_24 ), .\REG.mem_22_1 (\REG.mem_22_1 ), 
            .\REG.mem_23_1 (\REG.mem_23_1 ), .wr_fifo_en_w(wr_fifo_en_w), 
            .\wr_addr_nxt_c[4] (\wr_addr_nxt_c[4] ), .\wr_addr_nxt_c[2] (\wr_addr_nxt_c[2] ), 
            .\REG.mem_22_16 (\REG.mem_22_16 ), .\REG.mem_23_16 (\REG.mem_23_16 ), 
            .\REG.mem_21_1 (\REG.mem_21_1 ), .\REG.mem_21_16 (\REG.mem_21_16 ), 
            .\REG.mem_11_12 (\REG.mem_11_12 ), .\REG.mem_5_24 (\REG.mem_5_24 ), 
            .n7038(n7038), .n7037(n7037), .n7036(n7036), .n7035(n7035), 
            .n7034(n7034), .n7033(n7033), .wp_sync1_r({wp_sync1_r}), .n7032(n7032), 
            .n7031(n7031), .n7030(n7030), .n7029(n7029), .n7028(n7028), 
            .n7027(n7027), .n7025(n7025), .n7023(n7023), .n7022(n7022), 
            .n7021(n7021), .n7020(n7020), .n7019(n7019), .n7018(n7018), 
            .rp_sync1_r({rp_sync1_r}), .n7017(n7017), .n7016(n7016), .n7015(n7015), 
            .n7014(n7014), .n6955(n6955), .n6953(n6953), .\wr_addr_r[5] (\wr_addr_r[5] ), 
            .n6532(n6532), .\REG.mem_27_31 (\REG.mem_27_31 ), .n6531(n6531), 
            .\REG.mem_27_30 (\REG.mem_27_30 ), .n6530(n6530), .n6529(n6529), 
            .\REG.mem_27_28 (\REG.mem_27_28 ), .n6528(n6528), .\REG.mem_27_27 (\REG.mem_27_27 ), 
            .n6527(n6527), .\REG.mem_27_26 (\REG.mem_27_26 ), .n6526(n6526), 
            .\REG.mem_27_25 (\REG.mem_27_25 ), .n6525(n6525), .\REG.mem_27_24 (\REG.mem_27_24 ), 
            .n6524(n6524), .\REG.mem_27_23 (\REG.mem_27_23 ), .n6523(n6523), 
            .\REG.mem_27_22 (\REG.mem_27_22 ), .n6522(n6522), .\REG.mem_27_21 (\REG.mem_27_21 ), 
            .n6521(n6521), .\REG.mem_27_20 (\REG.mem_27_20 ), .n6520(n6520), 
            .n6519(n6519), .\REG.mem_27_18 (\REG.mem_27_18 ), .n6518(n6518), 
            .\REG.mem_27_17 (\REG.mem_27_17 ), .n6517(n6517), .\REG.mem_27_16 (\REG.mem_27_16 ), 
            .n6516(n6516), .\REG.mem_27_15 (\REG.mem_27_15 ), .n6515(n6515), 
            .\REG.mem_27_14 (\REG.mem_27_14 ), .n6514(n6514), .\REG.mem_27_13 (\REG.mem_27_13 ), 
            .n6513(n6513), .n6512(n6512), .\REG.mem_27_11 (\REG.mem_27_11 ), 
            .n6511(n6511), .\REG.mem_27_10 (\REG.mem_27_10 ), .n6510(n6510), 
            .\REG.mem_27_9 (\REG.mem_27_9 ), .n6509(n6509), .\REG.mem_27_8 (\REG.mem_27_8 ), 
            .n6508(n6508), .\REG.mem_27_7 (\REG.mem_27_7 ), .n6507(n6507), 
            .\REG.mem_27_6 (\REG.mem_27_6 ), .n6506(n6506), .\REG.mem_27_5 (\REG.mem_27_5 ), 
            .n6505(n6505), .\REG.mem_27_4 (\REG.mem_27_4 ), .n6504(n6504), 
            .n6503(n6503), .\REG.mem_27_2 (\REG.mem_27_2 ), .n6502(n6502), 
            .\REG.mem_27_1 (\REG.mem_27_1 ), .n6501(n6501), .n6404(n6404), 
            .\REG.mem_23_31 (\REG.mem_23_31 ), .n6403(n6403), .\REG.mem_23_30 (\REG.mem_23_30 ), 
            .n6402(n6402), .n6401(n6401), .n6400(n6400), .\REG.mem_23_27 (\REG.mem_23_27 ), 
            .n6399(n6399), .\REG.mem_23_26 (\REG.mem_23_26 ), .n6398(n6398), 
            .\REG.mem_23_25 (\REG.mem_23_25 ), .n6397(n6397), .\REG.mem_23_24 (\REG.mem_23_24 ), 
            .n6396(n6396), .\REG.mem_23_23 (\REG.mem_23_23 ), .n6395(n6395), 
            .\REG.mem_23_22 (\REG.mem_23_22 ), .n6394(n6394), .\REG.mem_23_21 (\REG.mem_23_21 ), 
            .n6393(n6393), .\REG.mem_23_20 (\REG.mem_23_20 ), .n6392(n6392), 
            .n6391(n6391), .\REG.mem_23_18 (\REG.mem_23_18 ), .n6390(n6390), 
            .\REG.mem_23_17 (\REG.mem_23_17 ), .n6389(n6389), .n6388(n6388), 
            .\REG.mem_23_15 (\REG.mem_23_15 ), .n6387(n6387), .\REG.mem_23_14 (\REG.mem_23_14 ), 
            .n6386(n6386), .\REG.mem_23_13 (\REG.mem_23_13 ), .n6385(n6385), 
            .\REG.mem_23_12 (\REG.mem_23_12 ), .n6384(n6384), .n6383(n6383), 
            .\REG.mem_23_10 (\REG.mem_23_10 ), .n6382(n6382), .n6381(n6381), 
            .\REG.mem_23_8 (\REG.mem_23_8 ), .n6380(n6380), .\REG.mem_23_7 (\REG.mem_23_7 ), 
            .n6379(n6379), .\REG.mem_23_6 (\REG.mem_23_6 ), .n6378(n6378), 
            .n6377(n6377), .\REG.mem_23_4 (\REG.mem_23_4 ), .n6376(n6376), 
            .\REG.mem_23_3 (\REG.mem_23_3 ), .n6375(n6375), .\REG.mem_23_2 (\REG.mem_23_2 ), 
            .n6374(n6374), .n6373(n6373), .\REG.mem_23_0 (\REG.mem_23_0 ), 
            .n6372(n6372), .\REG.mem_22_31 (\REG.mem_22_31 ), .n6371(n6371), 
            .\REG.mem_22_30 (\REG.mem_22_30 ), .n6370(n6370), .n6369(n6369), 
            .n6368(n6368), .\REG.mem_22_27 (\REG.mem_22_27 ), .n6367(n6367), 
            .\REG.mem_22_26 (\REG.mem_22_26 ), .n6366(n6366), .\REG.mem_22_25 (\REG.mem_22_25 ), 
            .n6365(n6365), .\REG.mem_22_24 (\REG.mem_22_24 ), .n6364(n6364), 
            .\REG.mem_22_23 (\REG.mem_22_23 ), .n6363(n6363), .\REG.mem_22_22 (\REG.mem_22_22 ), 
            .n6362(n6362), .\REG.mem_22_21 (\REG.mem_22_21 ), .n6361(n6361), 
            .\REG.mem_22_20 (\REG.mem_22_20 ), .n6360(n6360), .n6359(n6359), 
            .\REG.mem_22_18 (\REG.mem_22_18 ), .n6358(n6358), .\REG.mem_22_17 (\REG.mem_22_17 ), 
            .n6357(n6357), .n6356(n6356), .\REG.mem_22_15 (\REG.mem_22_15 ), 
            .n6355(n6355), .\REG.mem_22_14 (\REG.mem_22_14 ), .n6354(n6354), 
            .\REG.mem_22_13 (\REG.mem_22_13 ), .n6353(n6353), .\REG.mem_22_12 (\REG.mem_22_12 ), 
            .n6352(n6352), .n6351(n6351), .\REG.mem_22_10 (\REG.mem_22_10 ), 
            .n6350(n6350), .n6349(n6349), .\REG.mem_22_8 (\REG.mem_22_8 ), 
            .n6348(n6348), .\REG.mem_22_7 (\REG.mem_22_7 ), .n6347(n6347), 
            .\REG.mem_22_6 (\REG.mem_22_6 ), .n6346(n6346), .n6345(n6345), 
            .\REG.mem_22_4 (\REG.mem_22_4 ), .n6344(n6344), .\REG.mem_22_3 (\REG.mem_22_3 ), 
            .n6343(n6343), .\REG.mem_22_2 (\REG.mem_22_2 ), .n6342(n6342), 
            .n6341(n6341), .\REG.mem_22_0 (\REG.mem_22_0 ), .n6340(n6340), 
            .\REG.mem_21_31 (\REG.mem_21_31 ), .n6339(n6339), .\REG.mem_21_30 (\REG.mem_21_30 ), 
            .n6338(n6338), .n6337(n6337), .n6336(n6336), .\REG.mem_21_27 (\REG.mem_21_27 ), 
            .n6335(n6335), .\REG.mem_21_26 (\REG.mem_21_26 ), .n6334(n6334), 
            .\REG.mem_21_25 (\REG.mem_21_25 ), .n6333(n6333), .\REG.mem_21_24 (\REG.mem_21_24 ), 
            .n6332(n6332), .\REG.mem_21_23 (\REG.mem_21_23 ), .n6331(n6331), 
            .\REG.mem_21_22 (\REG.mem_21_22 ), .n6330(n6330), .\REG.mem_21_21 (\REG.mem_21_21 ), 
            .n6329(n6329), .\REG.mem_21_20 (\REG.mem_21_20 ), .n6328(n6328), 
            .n6327(n6327), .\REG.mem_21_18 (\REG.mem_21_18 ), .n6326(n6326), 
            .\REG.mem_21_17 (\REG.mem_21_17 ), .n6325(n6325), .n6324(n6324), 
            .\REG.mem_21_15 (\REG.mem_21_15 ), .n6323(n6323), .\REG.mem_21_14 (\REG.mem_21_14 ), 
            .n6322(n6322), .\REG.mem_21_13 (\REG.mem_21_13 ), .n6321(n6321), 
            .\REG.mem_21_12 (\REG.mem_21_12 ), .n6320(n6320), .n6319(n6319), 
            .\REG.mem_21_10 (\REG.mem_21_10 ), .n6318(n6318), .n6317(n6317), 
            .\REG.mem_21_8 (\REG.mem_21_8 ), .n6316(n6316), .\REG.mem_21_7 (\REG.mem_21_7 ), 
            .n6315(n6315), .\REG.mem_21_6 (\REG.mem_21_6 ), .n6314(n6314), 
            .n6313(n6313), .\REG.mem_21_4 (\REG.mem_21_4 ), .n6312(n6312), 
            .\REG.mem_21_3 (\REG.mem_21_3 ), .n6311(n6311), .\REG.mem_21_2 (\REG.mem_21_2 ), 
            .n6310(n6310), .n6309(n6309), .\REG.mem_21_0 (\REG.mem_21_0 ), 
            .n12(n12), .n10(n10), .n26(n26), .\rd_addr_nxt_c_5__N_573[4] (\rd_addr_nxt_c_5__N_573[4] ), 
            .\REG.mem_6_22 (\REG.mem_6_22 ), .\REG.mem_7_22 (\REG.mem_7_22 ), 
            .\REG.mem_6_23 (\REG.mem_6_23 ), .\REG.mem_7_23 (\REG.mem_7_23 ), 
            .\REG.mem_5_23 (\REG.mem_5_23 ), .\REG.mem_5_22 (\REG.mem_5_22 ), 
            .\REG.mem_11_23 (\REG.mem_11_23 ), .\REG.mem_11_18 (\REG.mem_11_18 ), 
            .\REG.mem_6_7 (\REG.mem_6_7 ), .\REG.mem_7_7 (\REG.mem_7_7 ), 
            .\REG.mem_5_7 (\REG.mem_5_7 ), .\REG.mem_11_9 (\REG.mem_11_9 ), 
            .n7(n7), .\REG.mem_6_28 (\REG.mem_6_28 ), .\REG.mem_7_28 (\REG.mem_7_28 ), 
            .\REG.mem_5_28 (\REG.mem_5_28 ), .n8(n8), .\REG.mem_11_28 (\REG.mem_11_28 ), 
            .VCC_net(VCC_net), .n25(n25), .\REG.mem_11_25 (\REG.mem_11_25 ), 
            .\wr_grey_sync_r[1] (\wr_grey_sync_r[1] ), .\wr_grey_sync_r[2] (\wr_grey_sync_r[2] ), 
            .\REG.mem_11_5 (\REG.mem_11_5 ), .\wr_grey_sync_r[3] (\wr_grey_sync_r[3] ), 
            .\wr_grey_sync_r[4] (\wr_grey_sync_r[4] ), .n6020(n6020), .\REG.mem_11_31 (\REG.mem_11_31 ), 
            .n6019(n6019), .\REG.mem_11_30 (\REG.mem_11_30 ), .n6018(n6018), 
            .\REG.mem_11_29 (\REG.mem_11_29 ), .n6017(n6017), .n6016(n6016), 
            .\REG.mem_11_27 (\REG.mem_11_27 ), .n6015(n6015), .\REG.mem_11_26 (\REG.mem_11_26 ), 
            .n6014(n6014), .n6013(n6013), .\REG.mem_11_24 (\REG.mem_11_24 ), 
            .n6012(n6012), .n6011(n6011), .\REG.mem_11_22 (\REG.mem_11_22 ), 
            .n6010(n6010), .n6009(n6009), .n6008(n6008), .\REG.mem_11_19 (\REG.mem_11_19 ), 
            .n6007(n6007), .\REG.mem_11_6 (\REG.mem_11_6 ), .n6006(n6006), 
            .\REG.mem_11_17 (\REG.mem_11_17 ), .n6005(n6005), .\REG.mem_11_16 (\REG.mem_11_16 ), 
            .n6004(n6004), .n6003(n6003), .n6002(n6002), .n6001(n6001), 
            .n6000(n6000), .n5999(n5999), .n5998(n5998), .\wr_addr_r[0] (\wr_addr_r[0] ), 
            .DEBUG_5_c(DEBUG_5_c), .\REG.mem_11_2 (\REG.mem_11_2 ), .n5997(n5997), 
            .n5996(n5996), .\REG.mem_11_7 (\REG.mem_11_7 ), .n5995(n5995), 
            .n5994(n5994), .n5993(n5993), .\REG.mem_11_4 (\REG.mem_11_4 ), 
            .\wr_addr_p1_w[0] (\wr_addr_p1_w[0] ), .n13865(n13865), .n14706(n14706), 
            .n5992(n5992), .\REG.mem_11_3 (\REG.mem_11_3 ), .n5991(n5991), 
            .n5990(n5990), .\REG.mem_11_1 (\REG.mem_11_1 ), .FT_OE_N_496(FT_OE_N_496), 
            .n12_adj_3(n12_adj_4), .dc32_fifo_read_enable(dc32_fifo_read_enable), 
            .n5989(n5989), .n5892(n5892), .\REG.mem_7_31 (\REG.mem_7_31 ), 
            .n5891(n5891), .\REG.mem_7_30 (\REG.mem_7_30 ), .n5890(n5890), 
            .\REG.mem_7_29 (\REG.mem_7_29 ), .n5889(n5889), .n5888(n5888), 
            .\REG.mem_7_27 (\REG.mem_7_27 ), .n5887(n5887), .n5886(n5886), 
            .\REG.mem_7_25 (\REG.mem_7_25 ), .n5885(n5885), .n5884(n5884), 
            .n5883(n5883), .n5882(n5882), .\REG.mem_7_21 (\REG.mem_7_21 ), 
            .n5881(n5881), .n5880(n5880), .n5879(n5879), .\REG.mem_7_18 (\REG.mem_7_18 ), 
            .n5878(n5878), .\REG.mem_7_17 (\REG.mem_7_17 ), .n5877(n5877), 
            .\REG.mem_7_16 (\REG.mem_7_16 ), .n5876(n5876), .\REG.mem_7_15 (\REG.mem_7_15 ), 
            .n5875(n5875), .n5874(n5874), .\REG.mem_7_13 (\REG.mem_7_13 ), 
            .n5873(n5873), .\REG.mem_7_12 (\REG.mem_7_12 ), .n5872(n5872), 
            .\REG.mem_7_11 (\REG.mem_7_11 ), .n5871(n5871), .\REG.mem_7_10 (\REG.mem_7_10 ), 
            .n5870(n5870), .n5869(n5869), .\REG.mem_7_8 (\REG.mem_7_8 ), 
            .n5868(n5868), .n5867(n5867), .\REG.mem_7_6 (\REG.mem_7_6 ), 
            .n5866(n5866), .\REG.mem_7_5 (\REG.mem_7_5 ), .n5865(n5865), 
            .\REG.mem_7_4 (\REG.mem_7_4 ), .n5864(n5864), .\REG.mem_7_3 (\REG.mem_7_3 ), 
            .n5863(n5863), .\REG.mem_7_2 (\REG.mem_7_2 ), .n5862(n5862), 
            .\REG.mem_7_1 (\REG.mem_7_1 ), .n5861(n5861), .\REG.mem_7_0 (\REG.mem_7_0 ), 
            .n5860(n5860), .\REG.mem_6_31 (\REG.mem_6_31 ), .n5859(n5859), 
            .\REG.mem_6_30 (\REG.mem_6_30 ), .n5858(n5858), .\REG.mem_6_29 (\REG.mem_6_29 ), 
            .n5857(n5857), .n5856(n5856), .\REG.mem_6_27 (\REG.mem_6_27 ), 
            .n5855(n5855), .n5854(n5854), .\REG.mem_6_25 (\REG.mem_6_25 ), 
            .n5853(n5853), .n5852(n5852), .n5851(n5851), .\state[3] (\state[3] ), 
            .n4843(n4843), .n1224(n1224), .n5850(n5850), .\REG.mem_6_21 (\REG.mem_6_21 ), 
            .n5849(n5849), .n5848(n5848), .n5847(n5847), .\REG.mem_6_18 (\REG.mem_6_18 ), 
            .n5846(n5846), .\REG.mem_6_17 (\REG.mem_6_17 ), .n5845(n5845), 
            .\REG.mem_6_16 (\REG.mem_6_16 ), .n5844(n5844), .\REG.mem_6_15 (\REG.mem_6_15 ), 
            .n5843(n5843), .n5842(n5842), .\REG.mem_6_13 (\REG.mem_6_13 ), 
            .n5841(n5841), .\REG.mem_6_12 (\REG.mem_6_12 ), .n5840(n5840), 
            .\REG.mem_6_11 (\REG.mem_6_11 ), .n5839(n5839), .\REG.mem_6_10 (\REG.mem_6_10 ), 
            .n5838(n5838), .n5837(n5837), .\REG.mem_6_8 (\REG.mem_6_8 ), 
            .n5836(n5836), .n5835(n5835), .\REG.mem_6_6 (\REG.mem_6_6 ), 
            .n5834(n5834), .\REG.mem_6_5 (\REG.mem_6_5 ), .n5833(n5833), 
            .\REG.mem_6_4 (\REG.mem_6_4 ), .\REG.mem_6_2 (\REG.mem_6_2 ), 
            .n5832(n5832), .\REG.mem_6_3 (\REG.mem_6_3 ), .n5831(n5831), 
            .\REG.mem_5_2 (\REG.mem_5_2 ), .n5830(n5830), .\REG.mem_6_1 (\REG.mem_6_1 ), 
            .n5829(n5829), .\REG.mem_6_0 (\REG.mem_6_0 ), .n5828(n5828), 
            .\REG.mem_5_31 (\REG.mem_5_31 ), .n5827(n5827), .\REG.mem_5_30 (\REG.mem_5_30 ), 
            .n5826(n5826), .\REG.mem_5_29 (\REG.mem_5_29 ), .n5825(n5825), 
            .n5824(n5824), .\REG.mem_5_27 (\REG.mem_5_27 ), .n5823(n5823), 
            .n5822(n5822), .\REG.mem_5_25 (\REG.mem_5_25 ), .n5821(n5821), 
            .n5820(n5820), .n5819(n5819), .n5818(n5818), .\REG.mem_5_21 (\REG.mem_5_21 ), 
            .n5817(n5817), .n5816(n5816), .n5815(n5815), .\REG.mem_5_18 (\REG.mem_5_18 ), 
            .n5814(n5814), .\REG.mem_5_17 (\REG.mem_5_17 ), .n5813(n5813), 
            .\REG.mem_5_16 (\REG.mem_5_16 ), .n5812(n5812), .\REG.mem_5_15 (\REG.mem_5_15 ), 
            .n5811(n5811), .n5810(n5810), .\REG.mem_5_13 (\REG.mem_5_13 ), 
            .n5809(n5809), .\REG.mem_5_12 (\REG.mem_5_12 ), .n5808(n5808), 
            .\REG.mem_5_11 (\REG.mem_5_11 ), .n5807(n5807), .\REG.mem_5_10 (\REG.mem_5_10 ), 
            .n5806(n5806), .n5805(n5805), .\REG.mem_5_8 (\REG.mem_5_8 ), 
            .n5804(n5804), .n5803(n5803), .\REG.mem_5_6 (\REG.mem_5_6 ), 
            .n5802(n5802), .\REG.mem_5_5 (\REG.mem_5_5 ), .n5648(n5648), 
            .n5801(n5801), .\REG.mem_5_4 (\REG.mem_5_4 ), .n5800(n5800), 
            .\REG.mem_5_3 (\REG.mem_5_3 ), .n5642(n5642), .n5639(n5639), 
            .n5638(n5638), .n5799(n5799), .n5798(n5798), .\REG.mem_5_1 (\REG.mem_5_1 ), 
            .n5797(n5797), .\REG.mem_5_0 (\REG.mem_5_0 ), .n5605(n5605), 
            .n27(n27), .n11(n11), .n28(n28)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_dc_32_lut_gen.v(53[33] 72[34])
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1
//

module fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 (dc32_fifo_data_in, 
            FIFO_CLK_c, GND_net, \REG.mem_22_29 , \REG.mem_23_29 , \REG.mem_21_29 , 
            \REG.mem_11_15 , \REG.mem_11_11 , \REG.mem_6_26 , \REG.mem_7_26 , 
            dc32_fifo_almost_full, reset_per_frame, \REG.mem_5_26 , rd_fifo_en_w, 
            dc32_fifo_data_out, SLM_CLK_c, \REG.mem_27_29 , \REG.mem_11_8 , 
            \REG.mem_22_5 , \REG.mem_23_5 , rd_grey_sync_r, \REG.mem_21_5 , 
            dc32_fifo_full, \REG.mem_6_20 , \REG.mem_7_20 , empty_nxt_c_N_636, 
            dc32_fifo_empty, \REG.mem_5_20 , \wr_grey_sync_r[0] , \aempty_flag_impl.ae_flag_nxt_w , 
            \rd_addr_nxt_c_5__N_573[3] , \rd_addr_nxt_c_5__N_573[1] , \REG.mem_11_20 , 
            \REG.mem_11_21 , \REG.mem_27_12 , \REG.mem_22_11 , \REG.mem_23_11 , 
            \REG.mem_21_11 , \REG.mem_27_3 , \REG.mem_11_10 , \REG.mem_22_28 , 
            \REG.mem_23_28 , \REG.mem_21_28 , \REG.mem_27_0 , \REG.mem_6_19 , 
            \REG.mem_7_19 , \REG.mem_5_19 , \REG.mem_6_9 , \REG.mem_7_9 , 
            \REG.mem_11_0 , \REG.mem_5_9 , \REG.mem_11_13 , \REG.mem_6_14 , 
            \REG.mem_7_14 , \REG.mem_5_14 , \REG.mem_22_19 , \REG.mem_23_19 , 
            \REG.mem_21_19 , \REG.mem_27_19 , n6, n22, \REG.mem_11_14 , 
            \REG.mem_22_9 , \REG.mem_23_9 , \REG.mem_21_9 , \REG.mem_6_24 , 
            \REG.mem_7_24 , \REG.mem_22_1 , \REG.mem_23_1 , wr_fifo_en_w, 
            \wr_addr_nxt_c[4] , \wr_addr_nxt_c[2] , \REG.mem_22_16 , \REG.mem_23_16 , 
            \REG.mem_21_1 , \REG.mem_21_16 , \REG.mem_11_12 , \REG.mem_5_24 , 
            n7038, n7037, n7036, n7035, n7034, n7033, wp_sync1_r, 
            n7032, n7031, n7030, n7029, n7028, n7027, n7025, n7023, 
            n7022, n7021, n7020, n7019, n7018, rp_sync1_r, n7017, 
            n7016, n7015, n7014, n6955, n6953, \wr_addr_r[5] , n6532, 
            \REG.mem_27_31 , n6531, \REG.mem_27_30 , n6530, n6529, 
            \REG.mem_27_28 , n6528, \REG.mem_27_27 , n6527, \REG.mem_27_26 , 
            n6526, \REG.mem_27_25 , n6525, \REG.mem_27_24 , n6524, 
            \REG.mem_27_23 , n6523, \REG.mem_27_22 , n6522, \REG.mem_27_21 , 
            n6521, \REG.mem_27_20 , n6520, n6519, \REG.mem_27_18 , 
            n6518, \REG.mem_27_17 , n6517, \REG.mem_27_16 , n6516, 
            \REG.mem_27_15 , n6515, \REG.mem_27_14 , n6514, \REG.mem_27_13 , 
            n6513, n6512, \REG.mem_27_11 , n6511, \REG.mem_27_10 , 
            n6510, \REG.mem_27_9 , n6509, \REG.mem_27_8 , n6508, \REG.mem_27_7 , 
            n6507, \REG.mem_27_6 , n6506, \REG.mem_27_5 , n6505, \REG.mem_27_4 , 
            n6504, n6503, \REG.mem_27_2 , n6502, \REG.mem_27_1 , n6501, 
            n6404, \REG.mem_23_31 , n6403, \REG.mem_23_30 , n6402, 
            n6401, n6400, \REG.mem_23_27 , n6399, \REG.mem_23_26 , 
            n6398, \REG.mem_23_25 , n6397, \REG.mem_23_24 , n6396, 
            \REG.mem_23_23 , n6395, \REG.mem_23_22 , n6394, \REG.mem_23_21 , 
            n6393, \REG.mem_23_20 , n6392, n6391, \REG.mem_23_18 , 
            n6390, \REG.mem_23_17 , n6389, n6388, \REG.mem_23_15 , 
            n6387, \REG.mem_23_14 , n6386, \REG.mem_23_13 , n6385, 
            \REG.mem_23_12 , n6384, n6383, \REG.mem_23_10 , n6382, 
            n6381, \REG.mem_23_8 , n6380, \REG.mem_23_7 , n6379, \REG.mem_23_6 , 
            n6378, n6377, \REG.mem_23_4 , n6376, \REG.mem_23_3 , n6375, 
            \REG.mem_23_2 , n6374, n6373, \REG.mem_23_0 , n6372, \REG.mem_22_31 , 
            n6371, \REG.mem_22_30 , n6370, n6369, n6368, \REG.mem_22_27 , 
            n6367, \REG.mem_22_26 , n6366, \REG.mem_22_25 , n6365, 
            \REG.mem_22_24 , n6364, \REG.mem_22_23 , n6363, \REG.mem_22_22 , 
            n6362, \REG.mem_22_21 , n6361, \REG.mem_22_20 , n6360, 
            n6359, \REG.mem_22_18 , n6358, \REG.mem_22_17 , n6357, 
            n6356, \REG.mem_22_15 , n6355, \REG.mem_22_14 , n6354, 
            \REG.mem_22_13 , n6353, \REG.mem_22_12 , n6352, n6351, 
            \REG.mem_22_10 , n6350, n6349, \REG.mem_22_8 , n6348, 
            \REG.mem_22_7 , n6347, \REG.mem_22_6 , n6346, n6345, \REG.mem_22_4 , 
            n6344, \REG.mem_22_3 , n6343, \REG.mem_22_2 , n6342, n6341, 
            \REG.mem_22_0 , n6340, \REG.mem_21_31 , n6339, \REG.mem_21_30 , 
            n6338, n6337, n6336, \REG.mem_21_27 , n6335, \REG.mem_21_26 , 
            n6334, \REG.mem_21_25 , n6333, \REG.mem_21_24 , n6332, 
            \REG.mem_21_23 , n6331, \REG.mem_21_22 , n6330, \REG.mem_21_21 , 
            n6329, \REG.mem_21_20 , n6328, n6327, \REG.mem_21_18 , 
            n6326, \REG.mem_21_17 , n6325, n6324, \REG.mem_21_15 , 
            n6323, \REG.mem_21_14 , n6322, \REG.mem_21_13 , n6321, 
            \REG.mem_21_12 , n6320, n6319, \REG.mem_21_10 , n6318, 
            n6317, \REG.mem_21_8 , n6316, \REG.mem_21_7 , n6315, \REG.mem_21_6 , 
            n6314, n6313, \REG.mem_21_4 , n6312, \REG.mem_21_3 , n6311, 
            \REG.mem_21_2 , n6310, n6309, \REG.mem_21_0 , n12, n10, 
            n26, \rd_addr_nxt_c_5__N_573[4] , \REG.mem_6_22 , \REG.mem_7_22 , 
            \REG.mem_6_23 , \REG.mem_7_23 , \REG.mem_5_23 , \REG.mem_5_22 , 
            \REG.mem_11_23 , \REG.mem_11_18 , \REG.mem_6_7 , \REG.mem_7_7 , 
            \REG.mem_5_7 , \REG.mem_11_9 , n7, \REG.mem_6_28 , \REG.mem_7_28 , 
            \REG.mem_5_28 , n8, \REG.mem_11_28 , VCC_net, n25, \REG.mem_11_25 , 
            \wr_grey_sync_r[1] , \wr_grey_sync_r[2] , \REG.mem_11_5 , 
            \wr_grey_sync_r[3] , \wr_grey_sync_r[4] , n6020, \REG.mem_11_31 , 
            n6019, \REG.mem_11_30 , n6018, \REG.mem_11_29 , n6017, 
            n6016, \REG.mem_11_27 , n6015, \REG.mem_11_26 , n6014, 
            n6013, \REG.mem_11_24 , n6012, n6011, \REG.mem_11_22 , 
            n6010, n6009, n6008, \REG.mem_11_19 , n6007, \REG.mem_11_6 , 
            n6006, \REG.mem_11_17 , n6005, \REG.mem_11_16 , n6004, 
            n6003, n6002, n6001, n6000, n5999, n5998, \wr_addr_r[0] , 
            DEBUG_5_c, \REG.mem_11_2 , n5997, n5996, \REG.mem_11_7 , 
            n5995, n5994, n5993, \REG.mem_11_4 , \wr_addr_p1_w[0] , 
            n13865, n14706, n5992, \REG.mem_11_3 , n5991, n5990, 
            \REG.mem_11_1 , FT_OE_N_496, n12_adj_3, dc32_fifo_read_enable, 
            n5989, n5892, \REG.mem_7_31 , n5891, \REG.mem_7_30 , n5890, 
            \REG.mem_7_29 , n5889, n5888, \REG.mem_7_27 , n5887, n5886, 
            \REG.mem_7_25 , n5885, n5884, n5883, n5882, \REG.mem_7_21 , 
            n5881, n5880, n5879, \REG.mem_7_18 , n5878, \REG.mem_7_17 , 
            n5877, \REG.mem_7_16 , n5876, \REG.mem_7_15 , n5875, n5874, 
            \REG.mem_7_13 , n5873, \REG.mem_7_12 , n5872, \REG.mem_7_11 , 
            n5871, \REG.mem_7_10 , n5870, n5869, \REG.mem_7_8 , n5868, 
            n5867, \REG.mem_7_6 , n5866, \REG.mem_7_5 , n5865, \REG.mem_7_4 , 
            n5864, \REG.mem_7_3 , n5863, \REG.mem_7_2 , n5862, \REG.mem_7_1 , 
            n5861, \REG.mem_7_0 , n5860, \REG.mem_6_31 , n5859, \REG.mem_6_30 , 
            n5858, \REG.mem_6_29 , n5857, n5856, \REG.mem_6_27 , n5855, 
            n5854, \REG.mem_6_25 , n5853, n5852, n5851, \state[3] , 
            n4843, n1224, n5850, \REG.mem_6_21 , n5849, n5848, n5847, 
            \REG.mem_6_18 , n5846, \REG.mem_6_17 , n5845, \REG.mem_6_16 , 
            n5844, \REG.mem_6_15 , n5843, n5842, \REG.mem_6_13 , n5841, 
            \REG.mem_6_12 , n5840, \REG.mem_6_11 , n5839, \REG.mem_6_10 , 
            n5838, n5837, \REG.mem_6_8 , n5836, n5835, \REG.mem_6_6 , 
            n5834, \REG.mem_6_5 , n5833, \REG.mem_6_4 , \REG.mem_6_2 , 
            n5832, \REG.mem_6_3 , n5831, \REG.mem_5_2 , n5830, \REG.mem_6_1 , 
            n5829, \REG.mem_6_0 , n5828, \REG.mem_5_31 , n5827, \REG.mem_5_30 , 
            n5826, \REG.mem_5_29 , n5825, n5824, \REG.mem_5_27 , n5823, 
            n5822, \REG.mem_5_25 , n5821, n5820, n5819, n5818, \REG.mem_5_21 , 
            n5817, n5816, n5815, \REG.mem_5_18 , n5814, \REG.mem_5_17 , 
            n5813, \REG.mem_5_16 , n5812, \REG.mem_5_15 , n5811, n5810, 
            \REG.mem_5_13 , n5809, \REG.mem_5_12 , n5808, \REG.mem_5_11 , 
            n5807, \REG.mem_5_10 , n5806, n5805, \REG.mem_5_8 , n5804, 
            n5803, \REG.mem_5_6 , n5802, \REG.mem_5_5 , n5648, n5801, 
            \REG.mem_5_4 , n5800, \REG.mem_5_3 , n5642, n5639, n5638, 
            n5799, n5798, \REG.mem_5_1 , n5797, \REG.mem_5_0 , n5605, 
            n27, n11, n28) /* synthesis syn_module_defined=1 */ ;
    input [31:0]dc32_fifo_data_in;
    input FIFO_CLK_c;
    input GND_net;
    output \REG.mem_22_29 ;
    output \REG.mem_23_29 ;
    output \REG.mem_21_29 ;
    output \REG.mem_11_15 ;
    output \REG.mem_11_11 ;
    output \REG.mem_6_26 ;
    output \REG.mem_7_26 ;
    output dc32_fifo_almost_full;
    input reset_per_frame;
    output \REG.mem_5_26 ;
    output rd_fifo_en_w;
    output [31:0]dc32_fifo_data_out;
    input SLM_CLK_c;
    output \REG.mem_27_29 ;
    output \REG.mem_11_8 ;
    output \REG.mem_22_5 ;
    output \REG.mem_23_5 ;
    output [5:0]rd_grey_sync_r;
    output \REG.mem_21_5 ;
    output dc32_fifo_full;
    output \REG.mem_6_20 ;
    output \REG.mem_7_20 ;
    input empty_nxt_c_N_636;
    output dc32_fifo_empty;
    output \REG.mem_5_20 ;
    output \wr_grey_sync_r[0] ;
    input \aempty_flag_impl.ae_flag_nxt_w ;
    output \rd_addr_nxt_c_5__N_573[3] ;
    output \rd_addr_nxt_c_5__N_573[1] ;
    output \REG.mem_11_20 ;
    output \REG.mem_11_21 ;
    output \REG.mem_27_12 ;
    output \REG.mem_22_11 ;
    output \REG.mem_23_11 ;
    output \REG.mem_21_11 ;
    output \REG.mem_27_3 ;
    output \REG.mem_11_10 ;
    output \REG.mem_22_28 ;
    output \REG.mem_23_28 ;
    output \REG.mem_21_28 ;
    output \REG.mem_27_0 ;
    output \REG.mem_6_19 ;
    output \REG.mem_7_19 ;
    output \REG.mem_5_19 ;
    output \REG.mem_6_9 ;
    output \REG.mem_7_9 ;
    output \REG.mem_11_0 ;
    output \REG.mem_5_9 ;
    output \REG.mem_11_13 ;
    output \REG.mem_6_14 ;
    output \REG.mem_7_14 ;
    output \REG.mem_5_14 ;
    output \REG.mem_22_19 ;
    output \REG.mem_23_19 ;
    output \REG.mem_21_19 ;
    output \REG.mem_27_19 ;
    output n6;
    output n22;
    output \REG.mem_11_14 ;
    output \REG.mem_22_9 ;
    output \REG.mem_23_9 ;
    output \REG.mem_21_9 ;
    output \REG.mem_6_24 ;
    output \REG.mem_7_24 ;
    output \REG.mem_22_1 ;
    output \REG.mem_23_1 ;
    input wr_fifo_en_w;
    output \wr_addr_nxt_c[4] ;
    output \wr_addr_nxt_c[2] ;
    output \REG.mem_22_16 ;
    output \REG.mem_23_16 ;
    output \REG.mem_21_1 ;
    output \REG.mem_21_16 ;
    output \REG.mem_11_12 ;
    output \REG.mem_5_24 ;
    input n7038;
    input n7037;
    input n7036;
    input n7035;
    input n7034;
    input n7033;
    output [5:0]wp_sync1_r;
    input n7032;
    input n7031;
    input n7030;
    input n7029;
    input n7028;
    input n7027;
    input n7025;
    input n7023;
    input n7022;
    input n7021;
    input n7020;
    input n7019;
    input n7018;
    output [5:0]rp_sync1_r;
    input n7017;
    input n7016;
    input n7015;
    input n7014;
    input n6955;
    input n6953;
    output \wr_addr_r[5] ;
    input n6532;
    output \REG.mem_27_31 ;
    input n6531;
    output \REG.mem_27_30 ;
    input n6530;
    input n6529;
    output \REG.mem_27_28 ;
    input n6528;
    output \REG.mem_27_27 ;
    input n6527;
    output \REG.mem_27_26 ;
    input n6526;
    output \REG.mem_27_25 ;
    input n6525;
    output \REG.mem_27_24 ;
    input n6524;
    output \REG.mem_27_23 ;
    input n6523;
    output \REG.mem_27_22 ;
    input n6522;
    output \REG.mem_27_21 ;
    input n6521;
    output \REG.mem_27_20 ;
    input n6520;
    input n6519;
    output \REG.mem_27_18 ;
    input n6518;
    output \REG.mem_27_17 ;
    input n6517;
    output \REG.mem_27_16 ;
    input n6516;
    output \REG.mem_27_15 ;
    input n6515;
    output \REG.mem_27_14 ;
    input n6514;
    output \REG.mem_27_13 ;
    input n6513;
    input n6512;
    output \REG.mem_27_11 ;
    input n6511;
    output \REG.mem_27_10 ;
    input n6510;
    output \REG.mem_27_9 ;
    input n6509;
    output \REG.mem_27_8 ;
    input n6508;
    output \REG.mem_27_7 ;
    input n6507;
    output \REG.mem_27_6 ;
    input n6506;
    output \REG.mem_27_5 ;
    input n6505;
    output \REG.mem_27_4 ;
    input n6504;
    input n6503;
    output \REG.mem_27_2 ;
    input n6502;
    output \REG.mem_27_1 ;
    input n6501;
    input n6404;
    output \REG.mem_23_31 ;
    input n6403;
    output \REG.mem_23_30 ;
    input n6402;
    input n6401;
    input n6400;
    output \REG.mem_23_27 ;
    input n6399;
    output \REG.mem_23_26 ;
    input n6398;
    output \REG.mem_23_25 ;
    input n6397;
    output \REG.mem_23_24 ;
    input n6396;
    output \REG.mem_23_23 ;
    input n6395;
    output \REG.mem_23_22 ;
    input n6394;
    output \REG.mem_23_21 ;
    input n6393;
    output \REG.mem_23_20 ;
    input n6392;
    input n6391;
    output \REG.mem_23_18 ;
    input n6390;
    output \REG.mem_23_17 ;
    input n6389;
    input n6388;
    output \REG.mem_23_15 ;
    input n6387;
    output \REG.mem_23_14 ;
    input n6386;
    output \REG.mem_23_13 ;
    input n6385;
    output \REG.mem_23_12 ;
    input n6384;
    input n6383;
    output \REG.mem_23_10 ;
    input n6382;
    input n6381;
    output \REG.mem_23_8 ;
    input n6380;
    output \REG.mem_23_7 ;
    input n6379;
    output \REG.mem_23_6 ;
    input n6378;
    input n6377;
    output \REG.mem_23_4 ;
    input n6376;
    output \REG.mem_23_3 ;
    input n6375;
    output \REG.mem_23_2 ;
    input n6374;
    input n6373;
    output \REG.mem_23_0 ;
    input n6372;
    output \REG.mem_22_31 ;
    input n6371;
    output \REG.mem_22_30 ;
    input n6370;
    input n6369;
    input n6368;
    output \REG.mem_22_27 ;
    input n6367;
    output \REG.mem_22_26 ;
    input n6366;
    output \REG.mem_22_25 ;
    input n6365;
    output \REG.mem_22_24 ;
    input n6364;
    output \REG.mem_22_23 ;
    input n6363;
    output \REG.mem_22_22 ;
    input n6362;
    output \REG.mem_22_21 ;
    input n6361;
    output \REG.mem_22_20 ;
    input n6360;
    input n6359;
    output \REG.mem_22_18 ;
    input n6358;
    output \REG.mem_22_17 ;
    input n6357;
    input n6356;
    output \REG.mem_22_15 ;
    input n6355;
    output \REG.mem_22_14 ;
    input n6354;
    output \REG.mem_22_13 ;
    input n6353;
    output \REG.mem_22_12 ;
    input n6352;
    input n6351;
    output \REG.mem_22_10 ;
    input n6350;
    input n6349;
    output \REG.mem_22_8 ;
    input n6348;
    output \REG.mem_22_7 ;
    input n6347;
    output \REG.mem_22_6 ;
    input n6346;
    input n6345;
    output \REG.mem_22_4 ;
    input n6344;
    output \REG.mem_22_3 ;
    input n6343;
    output \REG.mem_22_2 ;
    input n6342;
    input n6341;
    output \REG.mem_22_0 ;
    input n6340;
    output \REG.mem_21_31 ;
    input n6339;
    output \REG.mem_21_30 ;
    input n6338;
    input n6337;
    input n6336;
    output \REG.mem_21_27 ;
    input n6335;
    output \REG.mem_21_26 ;
    input n6334;
    output \REG.mem_21_25 ;
    input n6333;
    output \REG.mem_21_24 ;
    input n6332;
    output \REG.mem_21_23 ;
    input n6331;
    output \REG.mem_21_22 ;
    input n6330;
    output \REG.mem_21_21 ;
    input n6329;
    output \REG.mem_21_20 ;
    input n6328;
    input n6327;
    output \REG.mem_21_18 ;
    input n6326;
    output \REG.mem_21_17 ;
    input n6325;
    input n6324;
    output \REG.mem_21_15 ;
    input n6323;
    output \REG.mem_21_14 ;
    input n6322;
    output \REG.mem_21_13 ;
    input n6321;
    output \REG.mem_21_12 ;
    input n6320;
    input n6319;
    output \REG.mem_21_10 ;
    input n6318;
    input n6317;
    output \REG.mem_21_8 ;
    input n6316;
    output \REG.mem_21_7 ;
    input n6315;
    output \REG.mem_21_6 ;
    input n6314;
    input n6313;
    output \REG.mem_21_4 ;
    input n6312;
    output \REG.mem_21_3 ;
    input n6311;
    output \REG.mem_21_2 ;
    input n6310;
    input n6309;
    output \REG.mem_21_0 ;
    output n12;
    output n10;
    output n26;
    output \rd_addr_nxt_c_5__N_573[4] ;
    output \REG.mem_6_22 ;
    output \REG.mem_7_22 ;
    output \REG.mem_6_23 ;
    output \REG.mem_7_23 ;
    output \REG.mem_5_23 ;
    output \REG.mem_5_22 ;
    output \REG.mem_11_23 ;
    output \REG.mem_11_18 ;
    output \REG.mem_6_7 ;
    output \REG.mem_7_7 ;
    output \REG.mem_5_7 ;
    output \REG.mem_11_9 ;
    output n7;
    output \REG.mem_6_28 ;
    output \REG.mem_7_28 ;
    output \REG.mem_5_28 ;
    output n8;
    output \REG.mem_11_28 ;
    input VCC_net;
    input n25;
    output \REG.mem_11_25 ;
    output \wr_grey_sync_r[1] ;
    output \wr_grey_sync_r[2] ;
    output \REG.mem_11_5 ;
    output \wr_grey_sync_r[3] ;
    output \wr_grey_sync_r[4] ;
    input n6020;
    output \REG.mem_11_31 ;
    input n6019;
    output \REG.mem_11_30 ;
    input n6018;
    output \REG.mem_11_29 ;
    input n6017;
    input n6016;
    output \REG.mem_11_27 ;
    input n6015;
    output \REG.mem_11_26 ;
    input n6014;
    input n6013;
    output \REG.mem_11_24 ;
    input n6012;
    input n6011;
    output \REG.mem_11_22 ;
    input n6010;
    input n6009;
    input n6008;
    output \REG.mem_11_19 ;
    input n6007;
    output \REG.mem_11_6 ;
    input n6006;
    output \REG.mem_11_17 ;
    input n6005;
    output \REG.mem_11_16 ;
    input n6004;
    input n6003;
    input n6002;
    input n6001;
    input n6000;
    input n5999;
    input n5998;
    output \wr_addr_r[0] ;
    input DEBUG_5_c;
    output \REG.mem_11_2 ;
    input n5997;
    input n5996;
    output \REG.mem_11_7 ;
    input n5995;
    input n5994;
    input n5993;
    output \REG.mem_11_4 ;
    output \wr_addr_p1_w[0] ;
    output n13865;
    output n14706;
    input n5992;
    output \REG.mem_11_3 ;
    input n5991;
    input n5990;
    output \REG.mem_11_1 ;
    input FT_OE_N_496;
    output n12_adj_3;
    input dc32_fifo_read_enable;
    input n5989;
    input n5892;
    output \REG.mem_7_31 ;
    input n5891;
    output \REG.mem_7_30 ;
    input n5890;
    output \REG.mem_7_29 ;
    input n5889;
    input n5888;
    output \REG.mem_7_27 ;
    input n5887;
    input n5886;
    output \REG.mem_7_25 ;
    input n5885;
    input n5884;
    input n5883;
    input n5882;
    output \REG.mem_7_21 ;
    input n5881;
    input n5880;
    input n5879;
    output \REG.mem_7_18 ;
    input n5878;
    output \REG.mem_7_17 ;
    input n5877;
    output \REG.mem_7_16 ;
    input n5876;
    output \REG.mem_7_15 ;
    input n5875;
    input n5874;
    output \REG.mem_7_13 ;
    input n5873;
    output \REG.mem_7_12 ;
    input n5872;
    output \REG.mem_7_11 ;
    input n5871;
    output \REG.mem_7_10 ;
    input n5870;
    input n5869;
    output \REG.mem_7_8 ;
    input n5868;
    input n5867;
    output \REG.mem_7_6 ;
    input n5866;
    output \REG.mem_7_5 ;
    input n5865;
    output \REG.mem_7_4 ;
    input n5864;
    output \REG.mem_7_3 ;
    input n5863;
    output \REG.mem_7_2 ;
    input n5862;
    output \REG.mem_7_1 ;
    input n5861;
    output \REG.mem_7_0 ;
    input n5860;
    output \REG.mem_6_31 ;
    input n5859;
    output \REG.mem_6_30 ;
    input n5858;
    output \REG.mem_6_29 ;
    input n5857;
    input n5856;
    output \REG.mem_6_27 ;
    input n5855;
    input n5854;
    output \REG.mem_6_25 ;
    input n5853;
    input n5852;
    input n5851;
    input \state[3] ;
    input n4843;
    output n1224;
    input n5850;
    output \REG.mem_6_21 ;
    input n5849;
    input n5848;
    input n5847;
    output \REG.mem_6_18 ;
    input n5846;
    output \REG.mem_6_17 ;
    input n5845;
    output \REG.mem_6_16 ;
    input n5844;
    output \REG.mem_6_15 ;
    input n5843;
    input n5842;
    output \REG.mem_6_13 ;
    input n5841;
    output \REG.mem_6_12 ;
    input n5840;
    output \REG.mem_6_11 ;
    input n5839;
    output \REG.mem_6_10 ;
    input n5838;
    input n5837;
    output \REG.mem_6_8 ;
    input n5836;
    input n5835;
    output \REG.mem_6_6 ;
    input n5834;
    output \REG.mem_6_5 ;
    input n5833;
    output \REG.mem_6_4 ;
    output \REG.mem_6_2 ;
    input n5832;
    output \REG.mem_6_3 ;
    input n5831;
    output \REG.mem_5_2 ;
    input n5830;
    output \REG.mem_6_1 ;
    input n5829;
    output \REG.mem_6_0 ;
    input n5828;
    output \REG.mem_5_31 ;
    input n5827;
    output \REG.mem_5_30 ;
    input n5826;
    output \REG.mem_5_29 ;
    input n5825;
    input n5824;
    output \REG.mem_5_27 ;
    input n5823;
    input n5822;
    output \REG.mem_5_25 ;
    input n5821;
    input n5820;
    input n5819;
    input n5818;
    output \REG.mem_5_21 ;
    input n5817;
    input n5816;
    input n5815;
    output \REG.mem_5_18 ;
    input n5814;
    output \REG.mem_5_17 ;
    input n5813;
    output \REG.mem_5_16 ;
    input n5812;
    output \REG.mem_5_15 ;
    input n5811;
    input n5810;
    output \REG.mem_5_13 ;
    input n5809;
    output \REG.mem_5_12 ;
    input n5808;
    output \REG.mem_5_11 ;
    input n5807;
    output \REG.mem_5_10 ;
    input n5806;
    input n5805;
    output \REG.mem_5_8 ;
    input n5804;
    input n5803;
    output \REG.mem_5_6 ;
    input n5802;
    output \REG.mem_5_5 ;
    input n5648;
    input n5801;
    output \REG.mem_5_4 ;
    input n5800;
    output \REG.mem_5_3 ;
    input n5642;
    input n5639;
    input n5638;
    input n5799;
    input n5798;
    output \REG.mem_5_1 ;
    input n5797;
    output \REG.mem_5_0 ;
    input n5605;
    output n27;
    output n11;
    output n28;
    
    wire FIFO_CLK_c /* synthesis SET_AS_NETWORK=FIFO_CLK_c, is_clock=1 */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n20;
    wire [5:0]wr_addr_r;   // src/fifo_dc_32_lut_gen.v(196[29:38])
    
    wire \REG.mem_8_31 , n5924, \REG.mem_8_30 , n5923, n22_c, \REG.mem_25_11 , 
        n6448, \REG.mem_8_29 , n5922, \REG.mem_8_28 , n5921, \REG.mem_8_27 , 
        n5920, \REG.mem_8_26 , n5919, \REG.mem_8_25 , n5918, \REG.mem_8_24 , 
        n5917;
    wire [5:0]rd_addr_r;   // src/fifo_dc_32_lut_gen.v(217[29:38])
    
    wire \REG.mem_14_1 , \REG.mem_15_1 , n17091, \REG.mem_25_10 , n6447, 
        \REG.mem_25_9 , n6446, n17811, \REG.mem_1_20 , \REG.mem_0_20 , 
        n15080, n5753, \REG.mem_3_20 , n5752, \REG.mem_3_19 ;
    wire [5:0]n1;
    wire [5:0]wp_sync2_r;   // src/fifo_dc_32_lut_gen.v(223[37:47])
    wire [5:0]wp_sync_w;   // src/fifo_dc_32_lut_gen.v(226[30:39])
    
    wire \REG.mem_16_29 , \REG.mem_17_29 , n14739, \REG.mem_18_29 , 
        \REG.mem_19_29 , n14740, n14719, \REG.mem_8_23 , n5916, \REG.mem_20_29 , 
        n14718, \REG.mem_8_22 , n5915, \REG.mem_25_8 , n6445, \REG.mem_8_21 , 
        n5914, \REG.mem_18_3 , \REG.mem_19_3 , n17805, \REG.mem_13_1 , 
        \REG.mem_12_1 , n15797, \REG.mem_17_3 , \REG.mem_16_3 , n15566, 
        \REG.mem_25_7 , n6444, \REG.mem_10_15 , n17085, \REG.mem_8_20 , 
        n5913, \REG.mem_8_19 , n5912, \REG.mem_8_18 , n5911, \REG.mem_8_17 , 
        n5910, \REG.mem_0_26 , \REG.mem_1_26 , n15498, \REG.mem_8_16 , 
        n5909, \REG.mem_8_15 , n5908, n5751, \REG.mem_3_18 , \REG.mem_9_15 , 
        n15800, \REG.mem_8_11 , \REG.mem_9_11 , n15114, \REG.mem_2_26 , 
        \REG.mem_3_26 , n15499, \REG.mem_25_6 , n6443, \REG.mem_30_26 , 
        \REG.mem_31_26 , n17079, \REG.mem_29_26 , \REG.mem_28_26 , n17082, 
        \REG.mem_8_14 , n5907, \REG.mem_10_11 , n15115, n15571, \REG.mem_25_5 , 
        n6442, \afull_flag_impl.af_flag_nxt_w , \REG.mem_4_26 , n15570, 
        \REG.mem_8_13 , n5906, \REG.mem_2_18 , n17799, \REG.mem_1_18 , 
        \REG.mem_0_18 , n15569, \REG.mem_18_1 , \REG.mem_19_1 , n17073, 
        \REG.mem_25_4 , n6441;
    wire [31:0]rd_data_o_31__N_598;
    
    wire \REG.mem_16_5 , \REG.mem_17_5 , n15063, \REG.mem_8_12 , n5905, 
        \REG.mem_18_5 , \REG.mem_19_5 , n15064, \REG.mem_17_1 , \REG.mem_16_1 , 
        n15806, n5904, \REG.mem_8_10 , n5903, \REG.mem_14_16 , \REG.mem_15_16 , 
        n17793, \REG.mem_13_16 , \REG.mem_12_16 , n15083, \REG.mem_8_9 , 
        n5902, \REG.mem_26_29 , n17067, \REG.mem_8_8 , n5901, \REG.mem_25_3 , 
        n6440, \REG.mem_25_29 , \REG.mem_24_29 , n17070, \REG.mem_14_15 , 
        \REG.mem_15_15 , n17061, \REG.mem_10_8 , n17787, \REG.mem_8_7 , 
        n5900, \REG.mem_25_2 , n6439, \REG.mem_8_6 , n5899, \REG.mem_9_8 , 
        n17790, \REG.mem_13_15 , \REG.mem_12_15 , n15809, n15471, 
        n15472, n17781, n15433, n15432, n15580, \REG.mem_8_5 , n5898, 
        \REG.mem_8_4 , n5897, \REG.mem_8_3 , n5896, n15457, \REG.mem_8_2 , 
        n5895, \REG.mem_8_1 , n5894, \REG.mem_25_1 , n6438, \REG.mem_8_0 , 
        n5893, \REG.mem_25_0 , n6437;
    wire [5:0]rd_grey_w;   // src/fifo_dc_32_lut_gen.v(224[38:47])
    
    wire \REG.mem_2_15 , \REG.mem_3_15 , n17055, \REG.mem_1_15 , \REG.mem_0_15 , 
        n15254, \REG.mem_20_5 , n15456, full_nxt_c_N_633, n5750, \REG.mem_3_17 , 
        n17775, \REG.mem_4_20 , n15095;
    wire [5:0]wr_grey_w;   // src/fifo_dc_32_lut_gen.v(203[38:47])
    
    wire dc32_fifo_almost_empty, n5749, \REG.mem_3_16 , n16398, n17142, 
        n5748, n16236, n17280, n17418, n16458, \REG.mem_30_24 , 
        \REG.mem_31_24 , n17769, \REG.mem_29_24 , \REG.mem_28_24 , n17772, 
        n17496, n17442, n16380, n16212, n15177, n15178, n17049, 
        \REG.mem_18_16 , \REG.mem_19_16 , n17763;
    wire [5:0]rd_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(221[30:42])
    
    wire \REG.mem_17_16 , \REG.mem_16_16 , n15098, n5747, \REG.mem_3_14 , 
        n5746, \REG.mem_3_13 , n16812, n16770, n16950, n17160, n16284, 
        n17904, n15151, n15150, n17052, n27_c, n16248, n16932, 
        n16974, n16944, n15226, \REG.mem_24_12 , \REG.mem_25_12 , 
        n15039, \REG.mem_10_20 , n17757, \REG.mem_9_20 , n15101, \REG.mem_10_21 , 
        n17751, \REG.mem_9_21 , n15104, n16842, n15227, n16908, 
        \REG.mem_26_12 , n15040, \REG.mem_30_12 , \REG.mem_31_12 , n15046, 
        \REG.mem_28_12 , \REG.mem_29_12 , n15045, n16758, n16740, 
        n14953, n16548, n14954, n17742, n15553, n16872, n17826, 
        n15415, n16176, \REG.mem_16_11 , \REG.mem_17_11 , n15135, 
        \REG.mem_18_11 , \REG.mem_19_11 , n15136, n15142, \REG.mem_20_11 , 
        n15141, \REG.mem_26_3 , n17745, \REG.mem_9_10 , n15207, \REG.mem_10_10 , 
        n15208, \REG.mem_14_10 , \REG.mem_15_10 , n15214, \REG.mem_12_10 , 
        \REG.mem_13_10 , n15213, \REG.mem_16_28 , \REG.mem_17_28 , n14757, 
        \REG.mem_3_12 , n5745, \REG.mem_18_28 , \REG.mem_19_28 , n14758, 
        n14761, \REG.mem_20_28 , n14760, \REG.mem_3_11 , n5744, \REG.mem_24_0 , 
        n15000, \REG.mem_26_0 , n15001, \REG.mem_3_10 , n5743, \REG.mem_30_0 , 
        \REG.mem_31_0 , n15010, \REG.mem_3_9 , n5742, \REG.mem_3_8 , 
        n5741, \REG.mem_24_3 , n15590, \REG.mem_28_0 , \REG.mem_29_0 , 
        n15009, \REG.mem_14_8 , \REG.mem_15_8 , n17739, \REG.mem_13_8 , 
        \REG.mem_12_8 , \REG.mem_0_19 , \REG.mem_1_19 , n14772, \REG.mem_2_22 , 
        \REG.mem_3_22 , n17037, \REG.mem_2_19 , n14773, n14779, \REG.mem_3_7 , 
        n5740, \REG.mem_3_6 , n5739, \REG.mem_1_22 , \REG.mem_0_22 , 
        n17040, \REG.mem_3_5 , n5738, \REG.mem_4_19 , n14778, n17733, 
        \REG.mem_9_0 , n14970, \REG.mem_10_0 , n14971, \REG.mem_3_4 , 
        n5737, \REG.mem_14_0 , \REG.mem_15_0 , n14974, \REG.mem_12_0 , 
        \REG.mem_13_0 , n14973, \REG.mem_3_3 , n5736, \REG.mem_4_9 , 
        n14777, n17448, n17406, n15481, n7026, \REG.mem_9_13 , n14985, 
        \REG.mem_10_13 , n14986, \REG.mem_3_2 , n5735, \REG.mem_3_1 , 
        n5734, \REG.mem_3_0 , n5733, n32, \REG.mem_14_31 , n6116, 
        \REG.mem_14_13 , \REG.mem_15_13 , n14989, \REG.mem_12_13 , \REG.mem_13_13 , 
        n14988, n15483, n15484, n17727, n17016, n16938, n15595, 
        n17604, n17028, n15594, n16962, n15897, \REG.mem_3_31 , 
        n5764, n16848, n16824, n14755, \REG.mem_0_14 , \REG.mem_1_14 , 
        n15849, n6_c, n13666;
    wire [5:0]rd_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(233[30:44])
    
    wire \REG.mem_3_30 , n5763, \REG.mem_2_14 , n15850, n15460, n15459, 
        n15592, n15862, \REG.mem_3_29 , n5762, n17358, n15482, n16986, 
        \REG.mem_14_30 , n6115, n16272, n17946, \REG.mem_4_14 , n15861, 
        \REG.mem_3_28 , n5761, n16200, n16578, n14731, \REG.mem_3_27 , 
        n5760, n17592, n17526, n17025, n5759, n14751, n14752, 
        n17721, \REG.mem_3_25 , n5758, \REG.mem_18_7 , \REG.mem_19_7 , 
        n16299, n16914, n17208, n14746, n14745, n14782, \REG.mem_14_29 , 
        n6114, \REG.mem_20_19 , \REG.mem_14_28 , n6113, \REG.mem_3_24 , 
        n5757, \REG.mem_14_27 , n6112, \REG.mem_3_23 , n5756, n5755, 
        n14769, n14770, n17019, \REG.mem_3_21 , n5754, n14767, n14766, 
        n14809, \REG.mem_2_17 , n17715, \REG.mem_14_11 , \REG.mem_15_11 , 
        n15127, \REG.mem_26_19 , n17013, \REG.mem_12_11 , \REG.mem_13_11 , 
        n15126, \REG.mem_14_26 , n6111, n10_c, \REG.mem_19_31 , n6276, 
        \REG.mem_17_7 , \REG.mem_16_7 , n16302, \REG.mem_19_30 , n6275, 
        \REG.mem_14_25 , n6110, \REG.mem_14_24 , n6109, n14742, n14743, 
        n16293, n6274, n6273, \REG.mem_25_19 , \REG.mem_24_19 , \REG.mem_9_14 , 
        n15867, \REG.mem_19_27 , n6272, \REG.mem_14_23 , n6108, \REG.mem_19_26 , 
        n6271, \REG.mem_10_14 , n15868, \REG.mem_1_17 , \REG.mem_0_17 , 
        n15119, n16890, n16836, \REG.mem_19_25 , n6270, \REG.mem_14_14 , 
        \REG.mem_15_14 , n15880, \REG.mem_12_14 , \REG.mem_13_14 , n15879, 
        \REG.mem_16_9 , \REG.mem_17_9 , n14814, \REG.mem_18_9 , \REG.mem_19_9 , 
        n14815, n15601, \REG.mem_20_9 , n15600, \REG.mem_19_24 , n6269, 
        \REG.mem_19_23 , n6268, \REG.mem_19_22 , n6267, n16992, n15661, 
        \REG.mem_19_21 , n6266, \REG.mem_0_29 , \REG.mem_1_29 , n14928, 
        \REG.mem_2_29 , n14929, \REG.mem_19_20 , n6265, \REG.mem_16_10 , 
        \REG.mem_17_10 , n15219, \REG.mem_18_10 , \REG.mem_19_10 , n15220, 
        \REG.mem_19_19 , n6264, \REG.mem_19_18 , n6263, \REG.mem_0_24 , 
        \REG.mem_1_24 , n14829, \REG.mem_2_24 , n14830, n14839, n17007, 
        \REG.mem_19_17 , n6262;
    wire [5:0]wr_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(200[30:42])
    
    wire n6261, \REG.mem_19_15 , n6260, \REG.mem_19_14 , n6259, \REG.mem_19_13 , 
        n6258, \REG.mem_14_22 , n6107, n16185, \REG.mem_13_24 , \REG.mem_12_24 , 
        n16188, \REG.mem_19_12 , n6257, n6256, n6255, n17709, \REG.mem_14_21 , 
        n6106, n14734, n14733, n16296, \REG.mem_20_1 , n15818, \REG.mem_20_16 , 
        n15122, \REG.mem_14_20 , n6105, n6254, \REG.mem_19_8 , n6253, 
        n6252, \REG.mem_14_19 , n6104, \REG.mem_10_12 , n17703, \REG.mem_19_6 , 
        n6251, \REG.mem_2_4 , n17001, \REG.mem_9_12 , n17706, \REG.mem_4_24 , 
        n14838, n6250, \REG.mem_19_4 , n6249, n6248, \REG.mem_1_4 , 
        \REG.mem_0_4 , n15260, \REG.mem_19_2 , n6247, \REG.mem_14_18 , 
        n6103, \REG.mem_14_17 , n6102, n6246, \REG.mem_2_1 , n16995, 
        \REG.mem_19_0 , n6245, n34, \REG.mem_31_31 , n6660, n6101, 
        \REG.mem_31_30 , n6659, \REG.mem_1_1 , \REG.mem_0_1 , n15263, 
        \REG.mem_31_29 , n6658, \REG.mem_2_3 , n16287, \REG.mem_31_28 , 
        n6657, \REG.mem_30_29 , n16989, \REG.mem_29_29 , \REG.mem_28_29 , 
        \REG.mem_15_20 , n17697, n6100, \REG.mem_1_3 , \REG.mem_0_3 , 
        n16290, \REG.mem_31_27 , n6656, n6655, \REG.mem_31_25 , n6654, 
        n6099, \REG.mem_13_20 , \REG.mem_12_20 , n15131, n15746, n15488, 
        n16983, n7024;
    wire [5:0]rp_sync2_r;   // src/fifo_dc_32_lut_gen.v(202[37:47])
    
    wire n6653, \REG.mem_30_3 , \REG.mem_31_3 , n17691, n6098, \REG.mem_29_3 , 
        \REG.mem_28_3 , n15605, n6956, n6954, n6952, n6652, \REG.mem_31_23 , 
        n6651, \REG.mem_31_22 , n6650, \REG.mem_31_21 , n6649, \REG.mem_31_20 , 
        n6648, \REG.mem_31_19 , n6647, \REG.mem_31_18 , n6646, \REG.mem_31_17 , 
        n6645, \REG.mem_31_16 , n6644, \REG.mem_31_15 , n6643, \REG.mem_31_14 , 
        n6642, \REG.mem_31_13 , n6641, n6640, \REG.mem_31_11 , n6639, 
        \REG.mem_31_10 , n6638, \REG.mem_31_9 , n6637, \REG.mem_31_8 , 
        n6636, \REG.mem_31_7 , n6635, \REG.mem_31_6 , n6634, \REG.mem_31_5 , 
        n6633, \REG.mem_31_4 , n6632, n6631, \REG.mem_31_2 , n6630, 
        \REG.mem_31_1 , n6629, n6628, \REG.mem_30_31 , n6627, \REG.mem_30_30 , 
        n6626, n6625, \REG.mem_30_28 , n6624, \REG.mem_30_27 , n6623, 
        n6622, \REG.mem_30_25 , n6621, n6620, \REG.mem_30_23 , n6619, 
        \REG.mem_30_22 , n6618, \REG.mem_30_21 , n6617, \REG.mem_30_20 , 
        n6616, \REG.mem_30_19 , n6615, \REG.mem_30_18 , n6614, \REG.mem_30_17 , 
        n6613, \REG.mem_30_16 , n6612, \REG.mem_30_15 , n6611, \REG.mem_30_14 , 
        n6610, \REG.mem_30_13 , n6609, n6608, \REG.mem_30_11 , n6607, 
        \REG.mem_30_10 , n6606, \REG.mem_30_9 , n6605, \REG.mem_30_8 , 
        n6604, \REG.mem_30_7 , n6603, \REG.mem_30_6 , n6602, \REG.mem_30_5 , 
        n6601, \REG.mem_30_4 , n6600, n6599, \REG.mem_30_2 , n6598, 
        \REG.mem_30_1 , n6597, n6596, \REG.mem_29_31 , n6595, \REG.mem_29_30 , 
        n6594, n6593, \REG.mem_29_28 , n6592, \REG.mem_29_27 , n6591, 
        n6590, \REG.mem_29_25 , n6589, n6588, \REG.mem_29_23 , n6587, 
        \REG.mem_29_22 , n6586, \REG.mem_29_21 , n6585, \REG.mem_29_20 , 
        n6584, \REG.mem_29_19 , n6583, \REG.mem_29_18 , n6582, \REG.mem_29_17 , 
        n6581, \REG.mem_29_16 , n6580, \REG.mem_29_15 , n6579, \REG.mem_29_14 , 
        n6578, \REG.mem_29_13 , n6577, n6576, \REG.mem_29_11 , n6575, 
        \REG.mem_29_10 , n6574, \REG.mem_29_9 , n6573, \REG.mem_29_8 , 
        n6572, \REG.mem_29_7 , n6571, \REG.mem_29_6 , n6570, \REG.mem_29_5 , 
        n6569, \REG.mem_29_4 , n6568, n6567, \REG.mem_29_2 , n6566, 
        \REG.mem_29_1 , n6565, n6564, \REG.mem_28_31 , n6563, \REG.mem_28_30 , 
        n6562, n6561, \REG.mem_28_28 , n6560, \REG.mem_28_27 , n6559, 
        n6558, \REG.mem_28_25 , n6557, n6556, \REG.mem_28_23 , n6555, 
        \REG.mem_28_22 , n6554, \REG.mem_28_21 , n6553, \REG.mem_28_20 , 
        n6552, \REG.mem_28_19 , n6551, \REG.mem_28_18 , n6550, \REG.mem_28_17 , 
        n6549, \REG.mem_28_16 , n6548, \REG.mem_28_15 , n6547, \REG.mem_28_14 , 
        n6546, \REG.mem_28_13 , n6545, n6544, \REG.mem_28_11 , n6543, 
        \REG.mem_28_10 , n6542, \REG.mem_28_9 , n6541, \REG.mem_28_8 , 
        n6540, \REG.mem_28_7 , n6539, \REG.mem_28_6 , n6538, \REG.mem_28_5 , 
        n6537, \REG.mem_28_4 , n6536, n6535, \REG.mem_28_2 , n6534, 
        \REG.mem_28_1 , n6533, n6500, \REG.mem_26_31 , n6499, \REG.mem_26_30 , 
        n6498, n6497, \REG.mem_26_28 , n6496, \REG.mem_26_27 , n6495, 
        \REG.mem_26_26 , n6494, \REG.mem_26_25 , n6493, \REG.mem_26_24 , 
        n6492, \REG.mem_26_23 , n6491, \REG.mem_26_22 , n6490, \REG.mem_26_21 , 
        n6489, \REG.mem_26_20 , n6488, n6487, \REG.mem_26_18 , n6486, 
        \REG.mem_26_17 , n6485, \REG.mem_26_16 , n6484, \REG.mem_26_15 , 
        n6483, \REG.mem_26_14 , n6482, \REG.mem_26_13 , n6481, n6480, 
        \REG.mem_26_11 , n6479, \REG.mem_26_10 , n6478, \REG.mem_26_9 , 
        n6477, \REG.mem_26_8 , n6476, \REG.mem_26_7 , n6475, \REG.mem_26_6 , 
        n6474, \REG.mem_26_5 , n6473, \REG.mem_26_4 , n6472, n6471, 
        \REG.mem_26_2 , n6470, \REG.mem_26_1 , n6469, n6468, \REG.mem_25_31 , 
        n6467, \REG.mem_25_30 , n6466, n6465, \REG.mem_25_28 , n6464, 
        \REG.mem_25_27 , n6463, \REG.mem_25_26 , n6462, \REG.mem_25_25 , 
        n6461, \REG.mem_25_24 , n6460, \REG.mem_25_23 , n6459, \REG.mem_25_22 , 
        n6458, \REG.mem_25_21 , n6457, \REG.mem_25_20 , n6456, n6455, 
        \REG.mem_25_18 , n6454, \REG.mem_25_17 , n6453, \REG.mem_25_16 , 
        n6452, \REG.mem_25_15 , n6451, \REG.mem_25_14 , n6450, \REG.mem_25_13 , 
        n6449, n6436, \REG.mem_24_31 , n6435, \REG.mem_24_30 , n6434, 
        n6433, \REG.mem_24_28 , n6432, \REG.mem_24_27 , n6431, \REG.mem_24_26 , 
        n6430, \REG.mem_24_25 , n6429, \REG.mem_24_24 , n6428, \REG.mem_24_23 , 
        n6427, \REG.mem_24_22 , n6426, \REG.mem_24_21 , n6425, \REG.mem_24_20 , 
        n6424, n6423, \REG.mem_24_18 , n6422, \REG.mem_24_17 , n6421, 
        \REG.mem_24_16 , n6420, \REG.mem_24_15 , n6419, \REG.mem_24_14 , 
        n6418, \REG.mem_24_13 , n6417, n6416, \REG.mem_24_11 , n6415, 
        \REG.mem_24_10 , n6414, \REG.mem_24_9 , n6413, \REG.mem_24_8 , 
        n6412, \REG.mem_24_7 , n6411, \REG.mem_24_6 , n6410, \REG.mem_24_5 , 
        n6409, \REG.mem_24_4 , n6408, n6407, \REG.mem_24_2 , n6406, 
        \REG.mem_24_1 , n6405, n6308, \REG.mem_20_31 , n6307, \REG.mem_20_30 , 
        n6306, n6305, n6304, \REG.mem_20_27 , n6303, \REG.mem_20_26 , 
        n6302, \REG.mem_20_25 , n6301, \REG.mem_20_24 , n6300, \REG.mem_20_23 , 
        n6299, \REG.mem_20_22 , n6298, \REG.mem_20_21 , n6297, \REG.mem_20_20 , 
        n6296, n6295, \REG.mem_20_18 , n6294, \REG.mem_20_17 , n6293, 
        n6292, \REG.mem_20_15 , n6291, \REG.mem_20_14 , n6290, \REG.mem_20_13 , 
        n6289, \REG.mem_20_12 , n6288, n6287, \REG.mem_20_10 , n6286, 
        n6285, \REG.mem_20_8 , n6284, \REG.mem_20_7 , n6283, \REG.mem_20_6 , 
        n6282, n6281, \REG.mem_20_4 , n6280, \REG.mem_20_3 , n6279, 
        \REG.mem_20_2 , n6278, n6277, \REG.mem_20_0 , n6244, \REG.mem_18_31 , 
        n6243, \REG.mem_18_30 , n6242, n6241, n6240, \REG.mem_18_27 , 
        n6239, \REG.mem_18_26 , n6238, \REG.mem_18_25 , n6237, \REG.mem_18_24 , 
        n6236, \REG.mem_18_23 , n6235, \REG.mem_18_22 , n6234, \REG.mem_18_21 , 
        n6233, \REG.mem_18_20 , n6232, \REG.mem_18_19 , n6231, \REG.mem_18_18 , 
        n6230, \REG.mem_18_17 , n6229, n6228, \REG.mem_18_15 , n6227, 
        \REG.mem_18_14 , n6226, \REG.mem_18_13 , n6225, \REG.mem_18_12 , 
        n6224, n6223, n6222, n6221, \REG.mem_18_8 , n6220, n6219, 
        \REG.mem_18_6 , n6218, n6217, \REG.mem_18_4 , n6216, n6215, 
        \REG.mem_18_2 , n6214, n6213, \REG.mem_18_0 , n6212, \REG.mem_17_31 , 
        n6211, \REG.mem_17_30 , n6210, n6209, n6208, \REG.mem_17_27 , 
        n6207, \REG.mem_17_26 , n6206, \REG.mem_17_25 , n6205, \REG.mem_17_24 , 
        n6204, \REG.mem_17_23 , n6203, \REG.mem_17_22 , n6202, \REG.mem_17_21 , 
        n6201, \REG.mem_17_20 , n6200, \REG.mem_17_19 , n6199, \REG.mem_17_18 , 
        n6198, \REG.mem_17_17 , n6197, n6196, \REG.mem_17_15 , n6195, 
        \REG.mem_17_14 , n6194, \REG.mem_17_13 , n6193, \REG.mem_17_12 , 
        n6192, n6191, n6190, n6189, \REG.mem_17_8 , n6188, n6187, 
        \REG.mem_17_6 , n6186, n6185, \REG.mem_17_4 , n6184, n6183, 
        \REG.mem_17_2 , n6182, n6181, \REG.mem_17_0 , n6180, \REG.mem_16_31 , 
        n6179, \REG.mem_16_30 , n6178, n6177, n6176, \REG.mem_16_27 , 
        n6175, \REG.mem_16_26 , n6174, \REG.mem_16_25 , n6173, \REG.mem_16_24 , 
        n6172, \REG.mem_16_23 , n6171, \REG.mem_16_22 , n6170, \REG.mem_16_21 , 
        n6169, \REG.mem_16_20 , n6168, \REG.mem_16_19 , n6167, \REG.mem_16_18 , 
        n6166, \REG.mem_16_17 , n6165, n6164, \REG.mem_16_15 , n6163, 
        \REG.mem_16_14 , n6162, \REG.mem_16_13 , n6161, \REG.mem_16_12 , 
        n6160, n6159, n6158, n6157, \REG.mem_16_8 , n6156, n6155, 
        \REG.mem_16_6 , n6154, n6153, \REG.mem_16_4 , n6152, n6151, 
        \REG.mem_16_2 , n6150, n6149, \REG.mem_16_0 , n6148, \REG.mem_15_31 , 
        n6147, \REG.mem_15_30 , n6146, \REG.mem_15_29 , n6145, \REG.mem_15_28 , 
        n6144, \REG.mem_15_27 , n6143, \REG.mem_15_26 , n6142, \REG.mem_15_25 , 
        n15728, n15503, n15239, n15296, n16281, \REG.mem_14_12 , 
        n6097, n6141, \REG.mem_15_24 , n6140, \REG.mem_15_23 , n6139, 
        \REG.mem_15_22 , n6138, \REG.mem_15_21 , n6137, n6136, \REG.mem_15_19 , 
        n6135, \REG.mem_15_18 , n6134, \REG.mem_15_17 , n6133, n6132, 
        n6131, n6130, n6129, \REG.mem_15_12 , n6128, n6127, n6126, 
        \REG.mem_15_9 , n6125, n16197, \REG.mem_9_29 , n17685, \REG.mem_13_21 , 
        \REG.mem_12_21 , n15134, n15813, n6124, \REG.mem_15_7 , n6123, 
        \REG.mem_15_6 , n6122, \REG.mem_15_5 , n14, n15006, n15007, 
        n17679, n6096, n6121, \REG.mem_15_4 , n6120, \REG.mem_15_3 , 
        n6119, \REG.mem_15_2 , n6118, n6117, n15440, n6095, \REG.mem_14_9 , 
        n6094, n6093, \REG.mem_14_7 , n6092, n15004, n15003, n15139, 
        n16971, \REG.mem_2_23 , n17673, \REG.mem_1_23 , \REG.mem_0_23 , 
        n15608, \REG.mem_14_6 , n6091, \REG.mem_14_5 , n6090, n16965, 
        n16275, n17667, n16278, n15314, n15326, n16269, \REG.mem_14_4 , 
        n6089, \REG.mem_14_3 , n6088, \REG.mem_14_2 , n6087, n6086, 
        n15146, n6085, n15266, n25_c, n16959, n15428, n15814, 
        n17661, \REG.mem_4_23 , n15614, n16263, n14943, n6084, \REG.mem_13_31 , 
        n6083, \REG.mem_13_30 , n6082, \REG.mem_13_29 , n6081, \REG.mem_13_28 , 
        \REG.mem_4_22 , n14944, n14950, \REG.mem_10_23 , n17655, n6080, 
        \REG.mem_13_27 , n6079, \REG.mem_13_26 , n14949, n6078, \REG.mem_13_25 , 
        n6077, \REG.mem_9_23 , n15617, n6076, \REG.mem_13_23 , n6075, 
        \REG.mem_13_22 , n17649, n6074, n15149, n16266, n6073, n6072, 
        \REG.mem_13_19 , n6071, \REG.mem_13_18 , n17643, n16953, n15885, 
        n15833, n6070, \REG.mem_13_17 , n15823, \REG.mem_10_18 , n17631, 
        n15822, \REG.mem_9_18 , n15623, n6069, n6068, n17625, n6067, 
        n15650, n16947, n6066, \REG.mem_4_7 , n17628, n15852, n6065, 
        \REG.mem_13_12 , n6064, n15853, n6063, n17619, \REG.mem_12_23 , 
        n15626, n16428, n6062, \REG.mem_13_9 , n6061, n6060, \REG.mem_13_7 , 
        n16941, n6059, \REG.mem_13_6 , \REG.mem_10_9 , n17613, \REG.mem_9_9 , 
        n14789, n17607, n15660, n16935, n17601, n15176, n15200, 
        n16929, n7_c, n24, n13665, n46, n17595, n5641, n16923, 
        n15842, \REG.mem_12_9 , n14798, n14790, n14791, n16917, 
        n6058, \REG.mem_13_5 ;
    wire [5:0]wr_addr_nxt_c;   // src/fifo_dc_32_lut_gen.v(198[29:42])
    
    wire n15536, n16368, n17589, n30, n15527, n14785, n14784, 
        n14821, n15680, n15692, n16911, n16596, n15665, n13664, 
        n17400, n15520, n17583, n17556, n16905, n15794, n16899, 
        n15278, n17571, n15164, n6057, \REG.mem_13_4 , n17565, n15635, 
        n16893, n15281, n6056, \REG.mem_13_3 , n6055, \REG.mem_13_2 , 
        n6054, n6053, n17559, n15170, n5732, \REG.mem_2_31 , n15788, 
        n16887, n15782, n15444, n15445, n17553, n15412, n15411, 
        \REG.mem_0_28 , \REG.mem_1_28 , \REG.mem_2_28 , n6_adj_1378, 
        n23, \REG.mem_4_28 , n5731, \REG.mem_2_30 , n5730, n5729, 
        n5728, \REG.mem_2_27 , n5727, n16869, n15864, n15865, n16251, 
        n16776, n17964, n15172, n16164, n14722, n16863, n15241, 
        n16860, n15195, n15196, n16857, n15193, n15192, n13663, 
        \REG.mem_9_28 , \REG.mem_10_28 , n13662, n49, \REG.mem_12_28 , 
        \REG.mem_9_25 , n17541, \REG.mem_10_25 , n5726, \REG.mem_2_25 , 
        n5725, n5724, n5723, n5722, \REG.mem_2_21 , n5721, \REG.mem_2_20 , 
        n5720, n5719, n5718, n16845, n6052, \REG.mem_12_31 , n16254, 
        \REG.mem_12_25 , n17529, n15050, n16245, n16839, n15641, 
        n5717, \REG.mem_2_16 , n5716, n17523, n16404, n17517, n15044, 
        n15035, n16833, n5715, n16827, n6051, \REG.mem_12_30 , n6050, 
        \REG.mem_12_29 , n16239, n16830, n16242, n15181, n17511, 
        n6049, n6048, \REG.mem_12_27 , n6047, \REG.mem_12_26 , n6046, 
        n6045, n6044, n6043, \REG.mem_12_22 , n16821, n6042, n15647, 
        n17505, n5714, \REG.mem_2_13 , n6041, \REG.mem_12_18 , n16809, 
        n17499, n16386, n14800, n16803, n16800, n6040, \REG.mem_12_19 , 
        n6039, n6038, \REG.mem_12_17 , n6037, n15185, n17493, n15108, 
        n15109, n16797, n15091, n15090, n6036, n6035, n6034, n6033, 
        \REG.mem_12_12 , n6032, n6031, n6030, n6029, n6028, \REG.mem_12_7 , 
        n6027, \REG.mem_12_6 , n6026, \REG.mem_12_5 , n6025, \REG.mem_12_4 , 
        n15651, n15652, n16791, n14763, n14764, n17481, n15610, 
        n15609, n15886, n16785, n14749, n14748, n15190, n5713, 
        \REG.mem_2_12 , n5712, \REG.mem_2_11 , n16788, n15576, n15577, 
        n17475, n15876, n15877, n16779, n15859, n15858, n16782, 
        n14965, n14964, n15552, \REG.mem_10_5 , n16773, \REG.mem_2_2 , 
        n17463, n28_c, \REG.mem_1_2 , \REG.mem_0_2 , \REG.mem_9_5 , 
        n17457, n16767, n15668, n6024, \REG.mem_12_3 , n6023, \REG.mem_12_2 , 
        n15846, n15847, n16761, n15475, n15474, n15898, n16755, 
        n6022, n6021, n15165, n15166, n17451, n15160, n15159, 
        n16749, n15293, \REG.mem_10_6 , n17445, \REG.mem_9_6 , n16743, 
        n16536, n17439, n16737, n14909, n14912, n16233, n17433, 
        n14997, n14998, n16731, n14995, n14994, n15138;
    wire [5:0]n1_adj_1394;
    
    wire n13702, n13844, n8_adj_1383;
    wire [5:0]rp_sync_w;   // src/fifo_dc_32_lut_gen.v(205[30:39])
    
    wire n13701, n6_adj_1384, n13700;
    wire [5:0]wr_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(212[30:44])
    
    wire n7_adj_1385, n13699, n14_adj_1386, n13698, n16179, n16719, 
        n16722, n15579, n17421, n15547, n15546, n13727, n13726, 
        n13725, n16707, n14960, n15077, n17415, \REG.mem_1_27 , 
        \REG.mem_0_27 , n16710, n14948, n13724, n13723, \REG.mem_10_2 , 
        n17409, n16695, n5711, \REG.mem_2_10 , n29, \REG.mem_4_31 , 
        n5796, n5710, \REG.mem_2_9 , n5709, \REG.mem_2_8 , n5708, 
        \REG.mem_2_7 , n5707, \REG.mem_2_6 , n5706, \REG.mem_0_11 , 
        n5705, \REG.mem_0_12 , n5704, \REG.mem_0_13 , n5702, \REG.mem_4_30 , 
        n5795, \REG.mem_9_2 , \REG.mem_4_29 , n5794, n16698, n17403, 
        n5701, n5700, \REG.mem_0_16 , n15528, n15529, n17397, n16689, 
        n4962, \REG.mem_1_7 , \REG.mem_0_7 , n16692, n16683, n13722, 
        n16686, n15514, n15513, n8_adj_1387, n7_adj_1388, n9, n16182, 
        n16173, n14625, n15251, n14670, n5793, n16656, n15058, 
        n16671, \REG.mem_4_27 , n5792, n5791, n17370, n15189, n21, 
        n13721, n16566, n14968, n16665, n13720, n13719, n15087, 
        n15088, n17385, n13718, n14962, n16560, n15073, n15072, 
        n15205, n14649, n16650, n15055, n16659, n14663, n8_adj_1389, 
        n15052, n16644, n14593, n15492, n15493, n16653, n14906, 
        n14903, n15697, n15696, n14613, n14704, n15036, n15037, 
        n16647, n15904, n15031, n15030, n16, \REG.mem_4_25 , n5790, 
        n15024, n15025, n16641, n15019, n15018, n16632, n15022, 
        n16635, n5789, n5788, n15016, n16620, n14931, n14932, 
        n16191, n14991, n14992, n16629, \REG.mem_10_29 , n14983, 
        n14982, n17367, n16623, n5787, \REG.mem_4_21 , n5786, n5785, 
        n5784, \REG.mem_4_18 , n5783, n17361, \REG.mem_4_17 , n5782, 
        \REG.mem_4_16 , n5781, n15013, n16614, n5685, \REG.mem_2_0 , 
        n5687, \REG.mem_4_15 , n5780, n14802, n14803, n16617, n15895, 
        n15894, n15507, n15508, n17355, n15628, n15627, \REG.mem_2_5 , 
        n5681, n5599, n5623, n14979, n14980, n16611, n5603, n5779, 
        n14977, n14976, \REG.mem_4_13 , n5778, \REG.mem_4_12 , n5777, 
        \REG.mem_4_11 , n5776, n15222, n15223, n16161, n5988, \REG.mem_10_31 , 
        n5987, \REG.mem_10_30 , n5986, n5985, n5984, \REG.mem_10_27 , 
        n5983, \REG.mem_10_26 , n5982, n5981, \REG.mem_10_24 , n5980, 
        n5979, \REG.mem_10_22 , n5978, n5977, n5976, \REG.mem_10_19 , 
        n5975, n5974, \REG.mem_10_17 , n5973, \REG.mem_10_16 , n5972, 
        n5971, n5970, n5969, n5968, n5967, n5966, n5965, n5964, 
        \REG.mem_10_7 , n5963, n5962, n5961, \REG.mem_10_4 , n5960, 
        \REG.mem_10_3 , n5959, n5958, \REG.mem_10_1 , n5957, n5956, 
        \REG.mem_9_31 , n5955, \REG.mem_9_30 , n5954, n5953, n5952, 
        \REG.mem_9_27 , n5951, \REG.mem_9_26 , n5950, n5949, \REG.mem_9_24 , 
        n5948, n5947, \REG.mem_9_22 , n5946, n5945, n5944, \REG.mem_9_19 , 
        n5943, n5942, \REG.mem_9_17 , n5941, \REG.mem_9_16 , n5940, 
        n5939, n5938, n5937, n5936, n5935, n5934, n5933, n5932, 
        \REG.mem_9_7 , n5931, n5930, n5929, \REG.mem_9_4 , n5928, 
        \REG.mem_9_3 , n5927, n5926, \REG.mem_9_1 , n5925, \REG.mem_4_10 , 
        n5775, n16605, n5699, n5695, n5694, n5693, n16542, n16482, 
        n5689, \REG.mem_0_21 , n5688, n5686, n5684, n5683, \REG.mem_0_25 , 
        n5682, n5774, \REG.mem_4_8 , n5773, n5772, \REG.mem_4_6 , 
        n5771, \REG.mem_0_0 , n5676, n5679, n16599, n5680, \REG.mem_4_5 , 
        n5770, \REG.mem_4_4 , n5769, n16593, \REG.mem_4_2 , \REG.mem_4_3 , 
        n5768, n17319, n5767, \REG.mem_4_1 , n5766, n16587, \REG.mem_0_10 , 
        n5621, \REG.mem_0_9 , n5622, \REG.mem_0_8 , n5626, n16590, 
        n5627, \REG.mem_0_6 , n5632, n5678, \REG.mem_0_5 , n5633, 
        n5663, n5669, \REG.mem_4_0 , n5765, \REG.mem_0_31 , n5671, 
        n5672, n5675, n16581, n5677, \REG.mem_0_30 , n16584, n5670, 
        \REG.mem_1_0 , n5668, n5667, n5666, n5665, n5662, n5660, 
        n5659, \REG.mem_1_31 , n16575, n5655, n17307, n5654, \REG.mem_1_5 , 
        n16569, n14879, n5653, \REG.mem_1_6 , n16563, n5652, n16221, 
        n5651, \REG.mem_1_8 , n5650, \REG.mem_1_9 , n15707, n5649, 
        \REG.mem_1_10 , n16224, n16557, n5644, \REG.mem_1_30 , n5643, 
        \REG.mem_1_25 , n17295, n5640, \REG.mem_1_21 , n16194, n5637, 
        \REG.mem_1_11 , n5635, \REG.mem_1_12 , n5634, \REG.mem_1_13 , 
        n16215, n15713, n5630, n16551, n5619, n5616, n17289, n5615, 
        \REG.mem_1_16 , n15230, n14882, n16545, n16539, n5610, n5607, 
        n5606, n5602, n5601, n5600, n5598, n16533, n17277, n16326, 
        n16344, n16527, n14885, n12_adj_1391, n17271, n16521, n15722, 
        n16524, n18027, n15392, n16515, n16518, n16503, n18021, 
        n16506, n17259, n18015, n16497, n17256, n17214, n15401, 
        n17253, n18009, n15407, n17247, n15731, n18003, n16479, 
        n18006, n16473, n17997, n15419, n17991, n16455, n16449, 
        n17979, n17217, n15425, n17211, n16422, n17973, n17928, 
        n17148, n17967, n16437, n16440, n17205, n17961, n16410, 
        n16431, n16425, n17955, n17949, n16419, n16206, n17943, 
        n17937, n16413, n16416, n17931, n17181, n17925, n16407, 
        n16401, n17919, n16209, n16395, n17169, n17907, n16383, 
        n17901, n16320, n17163, n17895, n15518, n16377, n15542, 
        n16371, n17154, n17157, n17883, n17880, n17151, n17877, 
        n16365, n17145, n16359, n17871, n17865, n17139, n16353, 
        n17859, n17862, n16347, n17853, n16341, n17847, n17127, 
        n16323, n17841, n17121, n16317, n17829, n17109, n17832, 
        n16203, n17823, n17817, n17097;
    
    SB_LUT4 i4425_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_8_31 ), .O(n5924));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4425_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4424_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_8_30 ), .O(n5923));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4424_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4949_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_25_11 ), .O(n6448));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4949_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4423_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_8_29 ), .O(n5922));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4423_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4422_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_8_28 ), .O(n5921));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4422_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4421_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_8_27 ), .O(n5920));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4421_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4420_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_8_26 ), .O(n5919));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4420_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4419_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_8_25 ), .O(n5918));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4419_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4418_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_8_24 ), .O(n5917));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4418_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14812 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_1 ), 
            .I2(\REG.mem_15_1 ), .I3(rd_addr_r[1]), .O(n17091));
    defparam rd_addr_r_0__bdd_4_lut_14812.LUT_INIT = 16'he4aa;
    SB_LUT4 i4948_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_25_10 ), .O(n6447));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4948_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4947_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_25_9 ), .O(n6446));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4947_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17811_bdd_4_lut (.I0(n17811), .I1(\REG.mem_1_20 ), .I2(\REG.mem_0_20 ), 
            .I3(rd_addr_r[1]), .O(n15080));
    defparam n17811_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i386_387 (.Q(\REG.mem_3_20 ), .C(FIFO_CLK_c), .D(n5753));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i383_384 (.Q(\REG.mem_3_19 ), .C(FIFO_CLK_c), .D(n5752));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i5_1_lut (.I0(rd_addr_r[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 wp_sync2_r_5__I_0_130_i1_2_lut (.I0(wp_sync2_r[4]), .I1(wp_sync2_r[5]), 
            .I2(GND_net), .I3(GND_net), .O(wp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam wp_sync2_r_5__I_0_130_i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12615_3_lut (.I0(\REG.mem_16_29 ), .I1(\REG.mem_17_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14739));
    defparam i12615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12616_3_lut (.I0(\REG.mem_18_29 ), .I1(\REG.mem_19_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14740));
    defparam i12616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12595_3_lut (.I0(\REG.mem_22_29 ), .I1(\REG.mem_23_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14719));
    defparam i12595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4417_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_8_23 ), .O(n5916));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4417_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12594_3_lut (.I0(\REG.mem_20_29 ), .I1(\REG.mem_21_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14718));
    defparam i12594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4416_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_8_22 ), .O(n5915));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4416_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4946_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_25_8 ), .O(n6445));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4946_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4415_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_8_21 ), .O(n5914));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4415_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15407 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_3 ), 
            .I2(\REG.mem_19_3 ), .I3(rd_addr_r[1]), .O(n17805));
    defparam rd_addr_r_0__bdd_4_lut_15407.LUT_INIT = 16'he4aa;
    SB_LUT4 n17091_bdd_4_lut (.I0(n17091), .I1(\REG.mem_13_1 ), .I2(\REG.mem_12_1 ), 
            .I3(rd_addr_r[1]), .O(n15797));
    defparam n17091_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17805_bdd_4_lut (.I0(n17805), .I1(\REG.mem_17_3 ), .I2(\REG.mem_16_3 ), 
            .I3(rd_addr_r[1]), .O(n15566));
    defparam n17805_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4945_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_25_7 ), .O(n6444));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4945_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14807 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_15 ), 
            .I2(\REG.mem_11_15 ), .I3(rd_addr_r[1]), .O(n17085));
    defparam rd_addr_r_0__bdd_4_lut_14807.LUT_INIT = 16'he4aa;
    SB_LUT4 i4414_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_8_20 ), .O(n5913));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4414_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4413_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_8_19 ), .O(n5912));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4413_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4412_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_8_18 ), .O(n5911));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4412_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4411_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_8_17 ), .O(n5910));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4411_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13374_3_lut (.I0(\REG.mem_0_26 ), .I1(\REG.mem_1_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15498));
    defparam i13374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4410_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_8_16 ), .O(n5909));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4410_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4409_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_8_15 ), .O(n5908));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4409_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i380_381 (.Q(\REG.mem_3_18 ), .C(FIFO_CLK_c), .D(n5751));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n17085_bdd_4_lut (.I0(n17085), .I1(\REG.mem_9_15 ), .I2(\REG.mem_8_15 ), 
            .I3(rd_addr_r[1]), .O(n15800));
    defparam n17085_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12990_3_lut (.I0(\REG.mem_8_11 ), .I1(\REG.mem_9_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15114));
    defparam i12990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13375_3_lut (.I0(\REG.mem_2_26 ), .I1(\REG.mem_3_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15499));
    defparam i13375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4944_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_25_6 ), .O(n6443));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4944_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14802 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_26 ), 
            .I2(\REG.mem_31_26 ), .I3(rd_addr_r[1]), .O(n17079));
    defparam rd_addr_r_0__bdd_4_lut_14802.LUT_INIT = 16'he4aa;
    SB_LUT4 n17079_bdd_4_lut (.I0(n17079), .I1(\REG.mem_29_26 ), .I2(\REG.mem_28_26 ), 
            .I3(rd_addr_r[1]), .O(n17082));
    defparam n17079_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4408_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_8_14 ), .O(n5907));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4408_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12991_3_lut (.I0(\REG.mem_10_11 ), .I1(\REG.mem_11_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15115));
    defparam i12991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13447_3_lut (.I0(\REG.mem_6_26 ), .I1(\REG.mem_7_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15571));
    defparam i13447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4943_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_25_5 ), .O(n6442));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4943_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFSR \afull_flag_impl.af_flag_ext_r_111  (.Q(dc32_fifo_almost_full), 
            .C(FIFO_CLK_c), .D(\afull_flag_impl.af_flag_nxt_w ), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    SB_LUT4 i13446_3_lut (.I0(\REG.mem_4_26 ), .I1(\REG.mem_5_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15570));
    defparam i13446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4407_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_8_13 ), .O(n5906));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4407_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15402 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_18 ), 
            .I2(\REG.mem_3_18 ), .I3(rd_addr_r[1]), .O(n17799));
    defparam rd_addr_r_0__bdd_4_lut_15402.LUT_INIT = 16'he4aa;
    SB_LUT4 n17799_bdd_4_lut (.I0(n17799), .I1(\REG.mem_1_18 ), .I2(\REG.mem_0_18 ), 
            .I3(rd_addr_r[1]), .O(n15569));
    defparam n17799_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14797 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_1 ), 
            .I2(\REG.mem_19_1 ), .I3(rd_addr_r[1]), .O(n17073));
    defparam rd_addr_r_0__bdd_4_lut_14797.LUT_INIT = 16'he4aa;
    SB_LUT4 i4942_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_25_4 ), .O(n6441));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4942_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE \REG.out_raw_i0_i0  (.Q(dc32_fifo_data_out[0]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[0]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 i12939_3_lut (.I0(\REG.mem_16_5 ), .I1(\REG.mem_17_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15063));
    defparam i12939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4406_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_8_12 ), .O(n5905));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4406_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12940_3_lut (.I0(\REG.mem_18_5 ), .I1(\REG.mem_19_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15064));
    defparam i12940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17073_bdd_4_lut (.I0(n17073), .I1(\REG.mem_17_1 ), .I2(\REG.mem_16_1 ), 
            .I3(rd_addr_r[1]), .O(n15806));
    defparam n17073_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4405_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_8_11 ), .O(n5904));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4405_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4404_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_8_10 ), .O(n5903));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4404_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15397 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_16 ), 
            .I2(\REG.mem_15_16 ), .I3(rd_addr_r[1]), .O(n17793));
    defparam rd_addr_r_0__bdd_4_lut_15397.LUT_INIT = 16'he4aa;
    SB_LUT4 n17793_bdd_4_lut (.I0(n17793), .I1(\REG.mem_13_16 ), .I2(\REG.mem_12_16 ), 
            .I3(rd_addr_r[1]), .O(n15083));
    defparam n17793_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4403_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_8_9 ), .O(n5902));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4403_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14792 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_29 ), 
            .I2(\REG.mem_27_29 ), .I3(rd_addr_r[1]), .O(n17067));
    defparam rd_addr_r_0__bdd_4_lut_14792.LUT_INIT = 16'he4aa;
    SB_LUT4 i4402_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_8_8 ), .O(n5901));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4402_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4941_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_25_3 ), .O(n6440));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4941_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17067_bdd_4_lut (.I0(n17067), .I1(\REG.mem_25_29 ), .I2(\REG.mem_24_29 ), 
            .I3(rd_addr_r[1]), .O(n17070));
    defparam n17067_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14787 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_15 ), 
            .I2(\REG.mem_15_15 ), .I3(rd_addr_r[1]), .O(n17061));
    defparam rd_addr_r_0__bdd_4_lut_14787.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15392 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_8 ), 
            .I2(\REG.mem_11_8 ), .I3(rd_addr_r[1]), .O(n17787));
    defparam rd_addr_r_0__bdd_4_lut_15392.LUT_INIT = 16'he4aa;
    SB_LUT4 i4401_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_8_7 ), .O(n5900));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4401_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4940_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_25_2 ), .O(n6439));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4940_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4400_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_8_6 ), .O(n5899));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4400_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17787_bdd_4_lut (.I0(n17787), .I1(\REG.mem_9_8 ), .I2(\REG.mem_8_8 ), 
            .I3(rd_addr_r[1]), .O(n17790));
    defparam n17787_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17061_bdd_4_lut (.I0(n17061), .I1(\REG.mem_13_15 ), .I2(\REG.mem_12_15 ), 
            .I3(rd_addr_r[1]), .O(n15809));
    defparam n17061_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15437 (.I0(rd_addr_r[1]), .I1(n15471), 
            .I2(n15472), .I3(rd_addr_r[2]), .O(n17781));
    defparam rd_addr_r_1__bdd_4_lut_15437.LUT_INIT = 16'he4aa;
    SB_LUT4 n17781_bdd_4_lut (.I0(n17781), .I1(n15433), .I2(n15432), .I3(rd_addr_r[2]), 
            .O(n15580));
    defparam n17781_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4399_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_8_5 ), .O(n5898));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4399_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4398_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_8_4 ), .O(n5897));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4398_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4397_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_8_3 ), .O(n5896));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4397_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13333_3_lut (.I0(\REG.mem_22_5 ), .I1(\REG.mem_23_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15457));
    defparam i13333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4396_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_8_2 ), .O(n5895));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4396_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4395_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_8_1 ), .O(n5894));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4395_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4939_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_25_1 ), .O(n6438));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4939_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4394_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_8_0 ), .O(n5893));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4394_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4938_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_25_0 ), .O(n6437));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4938_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFSR rd_grey_sync_r__i0 (.Q(rd_grey_sync_r[0]), .C(SLM_CLK_c), .D(rd_grey_w[0]), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14782 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_15 ), 
            .I2(\REG.mem_3_15 ), .I3(rd_addr_r[1]), .O(n17055));
    defparam rd_addr_r_0__bdd_4_lut_14782.LUT_INIT = 16'he4aa;
    SB_LUT4 n17055_bdd_4_lut (.I0(n17055), .I1(\REG.mem_1_15 ), .I2(\REG.mem_0_15 ), 
            .I3(rd_addr_r[1]), .O(n15254));
    defparam n17055_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13332_3_lut (.I0(\REG.mem_20_5 ), .I1(\REG.mem_21_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15456));
    defparam i13332_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR full_ext_r_107 (.Q(dc32_fifo_full), .C(FIFO_CLK_c), .D(full_nxt_c_N_633), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i377_378 (.Q(\REG.mem_3_17 ), .C(FIFO_CLK_c), .D(n5750));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15387 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_20 ), 
            .I2(\REG.mem_7_20 ), .I3(rd_addr_r[1]), .O(n17775));
    defparam rd_addr_r_0__bdd_4_lut_15387.LUT_INIT = 16'he4aa;
    SB_DFFSS empty_ext_r_114 (.Q(dc32_fifo_empty), .C(SLM_CLK_c), .D(empty_nxt_c_N_636), 
            .S(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_LUT4 n17775_bdd_4_lut (.I0(n17775), .I1(\REG.mem_5_20 ), .I2(\REG.mem_4_20 ), 
            .I3(rd_addr_r[1]), .O(n15095));
    defparam n17775_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR wr_grey_sync_r__i0 (.Q(\wr_grey_sync_r[0] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[0]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFS \aempty_flag_impl.ae_flag_ext_r_120  (.Q(dc32_fifo_almost_empty), 
            .C(SLM_CLK_c), .D(\aempty_flag_impl.ae_flag_nxt_w ), .S(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(669[37] 672[40])
    SB_DFF i374_375 (.Q(\REG.mem_3_16 ), .C(FIFO_CLK_c), .D(n5749));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9484472_i1_3_lut (.I0(n16398), .I1(n17142), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[31]));
    defparam i9484472_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i371_372 (.Q(\REG.mem_3_15 ), .C(FIFO_CLK_c), .D(n5748));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9508484_i1_3_lut (.I0(n16236), .I1(n17280), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[30]));
    defparam i9508484_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9580520_i1_3_lut (.I0(n17418), .I1(n16458), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[27]));
    defparam i9580520_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15377 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_24 ), 
            .I2(\REG.mem_31_24 ), .I3(rd_addr_r[1]), .O(n17769));
    defparam rd_addr_r_0__bdd_4_lut_15377.LUT_INIT = 16'he4aa;
    SB_LUT4 n17769_bdd_4_lut (.I0(n17769), .I1(\REG.mem_29_24 ), .I2(\REG.mem_28_24 ), 
            .I3(rd_addr_r[1]), .O(n17772));
    defparam n17769_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9004232_i1_3_lut (.I0(n17496), .I1(n17442), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[23]));
    defparam i9004232_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8794127_i1_3_lut (.I0(n16380), .I1(n16212), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[21]));
    defparam i8794127_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14872 (.I0(rd_addr_r[1]), .I1(n15177), 
            .I2(n15178), .I3(rd_addr_r[2]), .O(n17049));
    defparam rd_addr_r_1__bdd_4_lut_14872.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15372 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_16 ), 
            .I2(\REG.mem_19_16 ), .I3(rd_addr_r[1]), .O(n17763));
    defparam rd_addr_r_0__bdd_4_lut_15372.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i3_2_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_5__N_573[3] ), .O(rd_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i3_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n17763_bdd_4_lut (.I0(n17763), .I1(\REG.mem_17_16 ), .I2(\REG.mem_16_16 ), 
            .I3(rd_addr_r[1]), .O(n15098));
    defparam n17763_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i368_369 (.Q(\REG.mem_3_14 ), .C(FIFO_CLK_c), .D(n5747));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i2_2_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_5__N_573[1] ), .O(rd_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_DFF i365_366 (.Q(\REG.mem_3_13 ), .C(FIFO_CLK_c), .D(n5746));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i8758109_i1_3_lut (.I0(n16812), .I1(n16770), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[20]));
    defparam i8758109_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9652556_i1_3_lut (.I0(n16950), .I1(n17160), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[18]));
    defparam i9652556_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9628544_i1_3_lut (.I0(n16284), .I1(n17904), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[17]));
    defparam i9628544_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17049_bdd_4_lut (.I0(n17049), .I1(n15151), .I2(n15150), .I3(rd_addr_r[2]), 
            .O(n17052));
    defparam n17049_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4254_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_3_20 ), .O(n5753));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4254_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9460460_i1_3_lut (.I0(n16248), .I1(n16932), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[16]));
    defparam i9460460_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4253_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_3_19 ), .O(n5752));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4253_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13102_3_lut (.I0(n16974), .I1(n16944), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15226));
    defparam i13102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4252_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_3_18 ), .O(n5751));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4252_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4251_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_3_17 ), .O(n5750));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4251_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12915_3_lut (.I0(\REG.mem_24_12 ), .I1(\REG.mem_25_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15039));
    defparam i12915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4250_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_3_16 ), .O(n5749));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4250_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15367 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_20 ), 
            .I2(\REG.mem_11_20 ), .I3(rd_addr_r[1]), .O(n17757));
    defparam rd_addr_r_0__bdd_4_lut_15367.LUT_INIT = 16'he4aa;
    SB_LUT4 n17757_bdd_4_lut (.I0(n17757), .I1(\REG.mem_9_20 ), .I2(\REG.mem_8_20 ), 
            .I3(rd_addr_r[1]), .O(n15101));
    defparam n17757_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15362 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_21 ), 
            .I2(\REG.mem_11_21 ), .I3(rd_addr_r[1]), .O(n17751));
    defparam rd_addr_r_0__bdd_4_lut_15362.LUT_INIT = 16'he4aa;
    SB_LUT4 n17751_bdd_4_lut (.I0(n17751), .I1(\REG.mem_9_21 ), .I2(\REG.mem_8_21 ), 
            .I3(rd_addr_r[1]), .O(n15104));
    defparam n17751_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13103_3_lut (.I0(n16842), .I1(n15226), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n15227));
    defparam i13103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9076268_i1_3_lut (.I0(n16908), .I1(n15227), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[15]));
    defparam i9076268_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12916_3_lut (.I0(\REG.mem_26_12 ), .I1(\REG.mem_27_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15040));
    defparam i12916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12922_3_lut (.I0(\REG.mem_30_12 ), .I1(\REG.mem_31_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15046));
    defparam i12922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12921_3_lut (.I0(\REG.mem_28_12 ), .I1(\REG.mem_29_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15045));
    defparam i12921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4249_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_3_15 ), .O(n5748));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4249_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12829_3_lut (.I0(n16758), .I1(n16740), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n14953));
    defparam i12829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12830_3_lut (.I0(n16548), .I1(n14953), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n14954));
    defparam i12830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13429_3_lut (.I0(n17790), .I1(n17742), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15553));
    defparam i13429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13291_3_lut (.I0(n16872), .I1(n17826), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15415));
    defparam i13291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9220340_i1_3_lut (.I0(n16176), .I1(n14954), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[9]));
    defparam i9220340_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13011_3_lut (.I0(\REG.mem_16_11 ), .I1(\REG.mem_17_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15135));
    defparam i13011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13012_3_lut (.I0(\REG.mem_18_11 ), .I1(\REG.mem_19_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15136));
    defparam i13012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4248_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_3_14 ), .O(n5747));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4248_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13018_3_lut (.I0(\REG.mem_22_11 ), .I1(\REG.mem_23_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15142));
    defparam i13018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13017_3_lut (.I0(\REG.mem_20_11 ), .I1(\REG.mem_21_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15141));
    defparam i13017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4247_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_3_13 ), .O(n5746));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4247_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15357 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_3 ), 
            .I2(\REG.mem_27_3 ), .I3(rd_addr_r[1]), .O(n17745));
    defparam rd_addr_r_0__bdd_4_lut_15357.LUT_INIT = 16'he4aa;
    SB_LUT4 i13083_3_lut (.I0(\REG.mem_8_10 ), .I1(\REG.mem_9_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15207));
    defparam i13083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13084_3_lut (.I0(\REG.mem_10_10 ), .I1(\REG.mem_11_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15208));
    defparam i13084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13090_3_lut (.I0(\REG.mem_14_10 ), .I1(\REG.mem_15_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15214));
    defparam i13090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13089_3_lut (.I0(\REG.mem_12_10 ), .I1(\REG.mem_13_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15213));
    defparam i13089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12633_3_lut (.I0(\REG.mem_16_28 ), .I1(\REG.mem_17_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14757));
    defparam i12633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4246_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_3_12 ), .O(n5745));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4246_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12634_3_lut (.I0(\REG.mem_18_28 ), .I1(\REG.mem_19_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14758));
    defparam i12634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12637_3_lut (.I0(\REG.mem_22_28 ), .I1(\REG.mem_23_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14761));
    defparam i12637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12636_3_lut (.I0(\REG.mem_20_28 ), .I1(\REG.mem_21_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14760));
    defparam i12636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4245_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_3_11 ), .O(n5744));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4245_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12876_3_lut (.I0(\REG.mem_24_0 ), .I1(\REG.mem_25_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15000));
    defparam i12876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12877_3_lut (.I0(\REG.mem_26_0 ), .I1(\REG.mem_27_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15001));
    defparam i12877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4244_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_3_10 ), .O(n5743));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4244_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12886_3_lut (.I0(\REG.mem_30_0 ), .I1(\REG.mem_31_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15010));
    defparam i12886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4243_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_3_9 ), .O(n5742));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4243_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4242_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_3_8 ), .O(n5741));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4242_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17745_bdd_4_lut (.I0(n17745), .I1(\REG.mem_25_3 ), .I2(\REG.mem_24_3 ), 
            .I3(rd_addr_r[1]), .O(n15590));
    defparam n17745_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12885_3_lut (.I0(\REG.mem_28_0 ), .I1(\REG.mem_29_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15009));
    defparam i12885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15352 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_8 ), 
            .I2(\REG.mem_15_8 ), .I3(rd_addr_r[1]), .O(n17739));
    defparam rd_addr_r_0__bdd_4_lut_15352.LUT_INIT = 16'he4aa;
    SB_LUT4 n17739_bdd_4_lut (.I0(n17739), .I1(\REG.mem_13_8 ), .I2(\REG.mem_12_8 ), 
            .I3(rd_addr_r[1]), .O(n17742));
    defparam n17739_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12648_3_lut (.I0(\REG.mem_0_19 ), .I1(\REG.mem_1_19 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14772));
    defparam i12648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14777 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_22 ), 
            .I2(\REG.mem_3_22 ), .I3(rd_addr_r[1]), .O(n17037));
    defparam rd_addr_r_0__bdd_4_lut_14777.LUT_INIT = 16'he4aa;
    SB_LUT4 i12649_3_lut (.I0(\REG.mem_2_19 ), .I1(\REG.mem_3_19 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14773));
    defparam i12649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12655_3_lut (.I0(\REG.mem_6_19 ), .I1(\REG.mem_7_19 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14779));
    defparam i12655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4241_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_3_7 ), .O(n5740));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4241_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4240_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_3_6 ), .O(n5739));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4240_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17037_bdd_4_lut (.I0(n17037), .I1(\REG.mem_1_22 ), .I2(\REG.mem_0_22 ), 
            .I3(rd_addr_r[1]), .O(n17040));
    defparam n17037_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4239_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_3_5 ), .O(n5738));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4239_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12654_3_lut (.I0(\REG.mem_4_19 ), .I1(\REG.mem_5_19 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14778));
    defparam i12654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15347 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_9 ), 
            .I2(\REG.mem_7_9 ), .I3(rd_addr_r[1]), .O(n17733));
    defparam rd_addr_r_0__bdd_4_lut_15347.LUT_INIT = 16'he4aa;
    SB_LUT4 i12846_3_lut (.I0(\REG.mem_8_0 ), .I1(\REG.mem_9_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14970));
    defparam i12846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12847_3_lut (.I0(\REG.mem_10_0 ), .I1(\REG.mem_11_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14971));
    defparam i12847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4238_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_3_4 ), .O(n5737));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4238_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12850_3_lut (.I0(\REG.mem_14_0 ), .I1(\REG.mem_15_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14974));
    defparam i12850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12849_3_lut (.I0(\REG.mem_12_0 ), .I1(\REG.mem_13_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14973));
    defparam i12849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4237_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_3_3 ), .O(n5736));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4237_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17733_bdd_4_lut (.I0(n17733), .I1(\REG.mem_5_9 ), .I2(\REG.mem_4_9 ), 
            .I3(rd_addr_r[1]), .O(n14777));
    defparam n17733_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13357_3_lut (.I0(n17448), .I1(n17406), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15481));
    defparam i13357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5527_2_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n7026));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i5527_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i12861_3_lut (.I0(\REG.mem_8_13 ), .I1(\REG.mem_9_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14985));
    defparam i12861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12862_3_lut (.I0(\REG.mem_10_13 ), .I1(\REG.mem_11_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14986));
    defparam i12862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4236_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_3_2 ), .O(n5735));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4236_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4235_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_3_1 ), .O(n5734));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4235_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4234_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_3_0 ), .O(n5733));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4234_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4617_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_14_31 ), .O(n6116));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4617_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12865_3_lut (.I0(\REG.mem_14_13 ), .I1(\REG.mem_15_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14989));
    defparam i12865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12864_3_lut (.I0(\REG.mem_12_13 ), .I1(\REG.mem_13_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14988));
    defparam i12864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15382 (.I0(rd_addr_r[1]), .I1(n15483), 
            .I2(n15484), .I3(rd_addr_r[2]), .O(n17727));
    defparam rd_addr_r_1__bdd_4_lut_15382.LUT_INIT = 16'he4aa;
    SB_LUT4 i13471_3_lut (.I0(n17016), .I1(n16938), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15595));
    defparam i13471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13470_3_lut (.I0(n17604), .I1(n17028), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15594));
    defparam i13470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13773_3_lut (.I0(n17040), .I1(n16962), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15897));
    defparam i13773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4265_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_3_31 ), .O(n5764));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4265_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i362_363 (.Q(\REG.mem_3_12 ), .C(FIFO_CLK_c), .D(n5745));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i12631_3_lut (.I0(n16848), .I1(n16824), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n14755));
    defparam i12631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13725_3_lut (.I0(\REG.mem_0_14 ), .I1(\REG.mem_1_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15849));
    defparam i13725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_7_lut (.I0(rd_sig_diff0_w[3]), .I1(wp_sync2_r[5]), 
            .I2(n1[5]), .I3(n13666), .O(n6_c)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i4264_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_3_30 ), .O(n5763));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4264_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i359_360 (.Q(\REG.mem_3_11 ), .C(FIFO_CLK_c), .D(n5744));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i13726_3_lut (.I0(\REG.mem_2_14 ), .I1(\REG.mem_3_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15850));
    defparam i13726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17727_bdd_4_lut (.I0(n17727), .I1(n15460), .I2(n15459), .I3(rd_addr_r[2]), 
            .O(n15592));
    defparam n17727_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13738_3_lut (.I0(\REG.mem_6_14 ), .I1(\REG.mem_7_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15862));
    defparam i13738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4263_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_3_29 ), .O(n5762));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4263_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13358_3_lut (.I0(n17358), .I1(n15481), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n15482));
    defparam i13358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9292376_i1_3_lut (.I0(n15482), .I1(n16986), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[6]));
    defparam i9292376_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4616_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_14_30 ), .O(n6115));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4616_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9340400_i1_3_lut (.I0(n16272), .I1(n17946), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[4]));
    defparam i9340400_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13737_3_lut (.I0(\REG.mem_4_14 ), .I1(\REG.mem_5_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15861));
    defparam i13737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4262_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_3_28 ), .O(n5761));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4262_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12607_3_lut (.I0(n16200), .I1(n16578), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n14731));
    defparam i12607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4261_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_3_27 ), .O(n5760));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4261_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9364412_i1_3_lut (.I0(n17592), .I1(n17526), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[3]));
    defparam i9364412_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14763 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_19 ), 
            .I2(\REG.mem_23_19 ), .I3(rd_addr_r[1]), .O(n17025));
    defparam rd_addr_r_0__bdd_4_lut_14763.LUT_INIT = 16'he4aa;
    SB_LUT4 i4260_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_3_26 ), .O(n5759));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4260_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15337 (.I0(rd_addr_r[1]), .I1(n14751), 
            .I2(n14752), .I3(rd_addr_r[2]), .O(n17721));
    defparam rd_addr_r_1__bdd_4_lut_15337.LUT_INIT = 16'he4aa;
    SB_LUT4 i4259_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_3_25 ), .O(n5758));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4259_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14164 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_7 ), 
            .I2(\REG.mem_19_7 ), .I3(rd_addr_r[1]), .O(n16299));
    defparam rd_addr_r_0__bdd_4_lut_14164.LUT_INIT = 16'he4aa;
    SB_LUT4 i9388424_i1_3_lut (.I0(n16914), .I1(n17208), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[2]));
    defparam i9388424_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17721_bdd_4_lut (.I0(n17721), .I1(n14746), .I2(n14745), .I3(rd_addr_r[2]), 
            .O(n14782));
    defparam n17721_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4615_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_14_29 ), .O(n6114));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4615_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17025_bdd_4_lut (.I0(n17025), .I1(\REG.mem_21_19 ), .I2(\REG.mem_20_19 ), 
            .I3(rd_addr_r[1]), .O(n17028));
    defparam n17025_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4614_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_14_28 ), .O(n6113));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4614_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4258_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_3_24 ), .O(n5757));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4258_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4613_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_14_27 ), .O(n6112));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4613_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4257_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_3_23 ), .O(n5756));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4257_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4256_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_3_22 ), .O(n5755));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4256_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14772 (.I0(rd_addr_r[1]), .I1(n14769), 
            .I2(n14770), .I3(rd_addr_r[2]), .O(n17019));
    defparam rd_addr_r_1__bdd_4_lut_14772.LUT_INIT = 16'he4aa;
    SB_LUT4 i4255_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_3_21 ), .O(n5754));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4255_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17019_bdd_4_lut (.I0(n17019), .I1(n14767), .I2(n14766), .I3(rd_addr_r[2]), 
            .O(n14809));
    defparam n17019_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15342 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_17 ), 
            .I2(\REG.mem_3_17 ), .I3(rd_addr_r[1]), .O(n17715));
    defparam rd_addr_r_0__bdd_4_lut_15342.LUT_INIT = 16'he4aa;
    SB_LUT4 i13003_3_lut (.I0(\REG.mem_14_11 ), .I1(\REG.mem_15_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15127));
    defparam i13003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14753 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_19 ), 
            .I2(\REG.mem_27_19 ), .I3(rd_addr_r[1]), .O(n17013));
    defparam rd_addr_r_0__bdd_4_lut_14753.LUT_INIT = 16'he4aa;
    SB_LUT4 i13002_3_lut (.I0(\REG.mem_12_11 ), .I1(\REG.mem_13_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15126));
    defparam i13002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4612_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_14_26 ), .O(n6111));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4612_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i58_2_lut_3_lut_4_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n6));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i58_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i59_2_lut_3_lut_4_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n22));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i59_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i4777_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_19_31 ), .O(n6276));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4777_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16299_bdd_4_lut (.I0(n16299), .I1(\REG.mem_17_7 ), .I2(\REG.mem_16_7 ), 
            .I3(rd_addr_r[1]), .O(n16302));
    defparam n16299_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4776_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_19_30 ), .O(n6275));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4776_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4611_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_14_25 ), .O(n6110));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4611_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4610_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_14_24 ), .O(n6109));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4610_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14219 (.I0(rd_addr_r[1]), .I1(n14742), 
            .I2(n14743), .I3(rd_addr_r[2]), .O(n16293));
    defparam rd_addr_r_1__bdd_4_lut_14219.LUT_INIT = 16'he4aa;
    SB_LUT4 i4775_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_19_29 ), .O(n6274));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4775_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4774_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_19_28 ), .O(n6273));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4774_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17013_bdd_4_lut (.I0(n17013), .I1(\REG.mem_25_19 ), .I2(\REG.mem_24_19 ), 
            .I3(rd_addr_r[1]), .O(n17016));
    defparam n17013_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13743_3_lut (.I0(\REG.mem_8_14 ), .I1(\REG.mem_9_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15867));
    defparam i13743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4773_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_19_27 ), .O(n6272));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4773_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4609_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_14_23 ), .O(n6108));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4609_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4772_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_19_26 ), .O(n6271));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4772_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13744_3_lut (.I0(\REG.mem_10_14 ), .I1(\REG.mem_11_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15868));
    defparam i13744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17715_bdd_4_lut (.I0(n17715), .I1(\REG.mem_1_17 ), .I2(\REG.mem_0_17 ), 
            .I3(rd_addr_r[1]), .O(n15119));
    defparam n17715_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9412436_i1_3_lut (.I0(n16890), .I1(n16836), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(rd_data_o_31__N_598[1]));
    defparam i9412436_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4771_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_19_25 ), .O(n6270));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4771_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13756_3_lut (.I0(\REG.mem_14_14 ), .I1(\REG.mem_15_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15880));
    defparam i13756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13755_3_lut (.I0(\REG.mem_12_14 ), .I1(\REG.mem_13_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15879));
    defparam i13755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12690_3_lut (.I0(\REG.mem_16_9 ), .I1(\REG.mem_17_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14814));
    defparam i12690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12691_3_lut (.I0(\REG.mem_18_9 ), .I1(\REG.mem_19_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14815));
    defparam i12691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13477_3_lut (.I0(\REG.mem_22_9 ), .I1(\REG.mem_23_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15601));
    defparam i13477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13476_3_lut (.I0(\REG.mem_20_9 ), .I1(\REG.mem_21_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15600));
    defparam i13476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4770_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_19_24 ), .O(n6269));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4770_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4769_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_19_23 ), .O(n6268));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4769_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4768_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_19_22 ), .O(n6267));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4768_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13537_3_lut (.I0(n17070), .I1(n16992), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15661));
    defparam i13537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4767_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_19_21 ), .O(n6266));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4767_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12804_3_lut (.I0(\REG.mem_0_29 ), .I1(\REG.mem_1_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14928));
    defparam i12804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12805_3_lut (.I0(\REG.mem_2_29 ), .I1(\REG.mem_3_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14929));
    defparam i12805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4766_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_19_20 ), .O(n6265));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4766_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13095_3_lut (.I0(\REG.mem_16_10 ), .I1(\REG.mem_17_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15219));
    defparam i13095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13096_3_lut (.I0(\REG.mem_18_10 ), .I1(\REG.mem_19_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15220));
    defparam i13096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4765_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_19_19 ), .O(n6264));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4765_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4764_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_19_18 ), .O(n6263));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4764_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12705_3_lut (.I0(\REG.mem_0_24 ), .I1(\REG.mem_1_24 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14829));
    defparam i12705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12706_3_lut (.I0(\REG.mem_2_24 ), .I1(\REG.mem_3_24 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14830));
    defparam i12706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12715_3_lut (.I0(\REG.mem_6_24 ), .I1(\REG.mem_7_24 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14839));
    defparam i12715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14743 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_1 ), 
            .I2(\REG.mem_23_1 ), .I3(rd_addr_r[1]), .O(n17007));
    defparam rd_addr_r_0__bdd_4_lut_14743.LUT_INIT = 16'he4aa;
    SB_LUT4 i4763_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_19_17 ), .O(n6262));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4763_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_r_5__I_0_123_i5_3_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(wr_fifo_en_w), .I3(GND_net), .O(\wr_addr_nxt_c[4] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_5__I_0_123_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4762_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_19_16 ), .O(n6261));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4762_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4761_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_19_15 ), .O(n6260));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4761_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_r_5__I_0_123_i3_3_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(wr_fifo_en_w), .I3(GND_net), .O(\wr_addr_nxt_c[2] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_5__I_0_123_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4760_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_19_14 ), .O(n6259));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4760_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4759_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_19_13 ), .O(n6258));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4759_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4608_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_14_22 ), .O(n6107));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4608_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16185_bdd_4_lut (.I0(n16185), .I1(\REG.mem_13_24 ), .I2(\REG.mem_12_24 ), 
            .I3(rd_addr_r[1]), .O(n16188));
    defparam n16185_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4758_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_19_12 ), .O(n6257));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4758_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4757_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_19_11 ), .O(n6256));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4757_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4756_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_19_10 ), .O(n6255));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4756_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15327 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_16 ), 
            .I2(\REG.mem_23_16 ), .I3(rd_addr_r[1]), .O(n17709));
    defparam rd_addr_r_0__bdd_4_lut_15327.LUT_INIT = 16'he4aa;
    SB_LUT4 i4607_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_14_21 ), .O(n6106));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4607_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16293_bdd_4_lut (.I0(n16293), .I1(n14734), .I2(n14733), .I3(rd_addr_r[2]), 
            .O(n16296));
    defparam n16293_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17007_bdd_4_lut (.I0(n17007), .I1(\REG.mem_21_1 ), .I2(\REG.mem_20_1 ), 
            .I3(rd_addr_r[1]), .O(n15818));
    defparam n17007_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17709_bdd_4_lut (.I0(n17709), .I1(\REG.mem_21_16 ), .I2(\REG.mem_20_16 ), 
            .I3(rd_addr_r[1]), .O(n15122));
    defparam n17709_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4606_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_14_20 ), .O(n6105));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4606_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4755_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_19_9 ), .O(n6254));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4755_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4754_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_19_8 ), .O(n6253));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4754_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4753_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_19_7 ), .O(n6252));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4753_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4605_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_14_19 ), .O(n6104));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4605_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15322 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_12 ), 
            .I2(\REG.mem_11_12 ), .I3(rd_addr_r[1]), .O(n17703));
    defparam rd_addr_r_0__bdd_4_lut_15322.LUT_INIT = 16'he4aa;
    SB_LUT4 i4752_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_19_6 ), .O(n6251));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4752_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14738 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_4 ), 
            .I2(\REG.mem_3_4 ), .I3(rd_addr_r[1]), .O(n17001));
    defparam rd_addr_r_0__bdd_4_lut_14738.LUT_INIT = 16'he4aa;
    SB_LUT4 n17703_bdd_4_lut (.I0(n17703), .I1(\REG.mem_9_12 ), .I2(\REG.mem_8_12 ), 
            .I3(rd_addr_r[1]), .O(n17706));
    defparam n17703_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12714_3_lut (.I0(\REG.mem_4_24 ), .I1(\REG.mem_5_24 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14838));
    defparam i12714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4751_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_19_5 ), .O(n6250));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4751_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4750_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_19_4 ), .O(n6249));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4750_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4749_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_19_3 ), .O(n6248));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4749_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17001_bdd_4_lut (.I0(n17001), .I1(\REG.mem_1_4 ), .I2(\REG.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(n15260));
    defparam n17001_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4748_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_19_2 ), .O(n6247));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4748_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4604_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_14_18 ), .O(n6103));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4604_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4603_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_14_17 ), .O(n6102));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4603_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4747_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_19_1 ), .O(n6246));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4747_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14733 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_1 ), 
            .I2(\REG.mem_3_1 ), .I3(rd_addr_r[1]), .O(n16995));
    defparam rd_addr_r_0__bdd_4_lut_14733.LUT_INIT = 16'he4aa;
    SB_LUT4 i4746_3_lut_4_lut (.I0(n27_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_19_0 ), .O(n6245));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4746_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5161_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_31_31 ), .O(n6660));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5161_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4602_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_14_16 ), .O(n6101));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4602_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5160_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_31_30 ), .O(n6659));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5160_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16995_bdd_4_lut (.I0(n16995), .I1(\REG.mem_1_1 ), .I2(\REG.mem_0_1 ), 
            .I3(rd_addr_r[1]), .O(n15263));
    defparam n16995_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5159_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_31_29 ), .O(n6658));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5159_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14149 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_3 ), 
            .I2(\REG.mem_3_3 ), .I3(rd_addr_r[1]), .O(n16287));
    defparam rd_addr_r_0__bdd_4_lut_14149.LUT_INIT = 16'he4aa;
    SB_LUT4 i5158_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_31_28 ), .O(n6657));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5158_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14728 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_29 ), 
            .I2(\REG.mem_31_29 ), .I3(rd_addr_r[1]), .O(n16989));
    defparam rd_addr_r_0__bdd_4_lut_14728.LUT_INIT = 16'he4aa;
    SB_LUT4 n16989_bdd_4_lut (.I0(n16989), .I1(\REG.mem_29_29 ), .I2(\REG.mem_28_29 ), 
            .I3(rd_addr_r[1]), .O(n16992));
    defparam n16989_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15317 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_20 ), 
            .I2(\REG.mem_15_20 ), .I3(rd_addr_r[1]), .O(n17697));
    defparam rd_addr_r_0__bdd_4_lut_15317.LUT_INIT = 16'he4aa;
    SB_LUT4 i4601_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_14_15 ), .O(n6100));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4601_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16287_bdd_4_lut (.I0(n16287), .I1(\REG.mem_1_3 ), .I2(\REG.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(n16290));
    defparam n16287_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5157_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_31_27 ), .O(n6656));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5157_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5156_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_31_26 ), .O(n6655));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5156_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5155_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_31_25 ), .O(n6654));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5155_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4600_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_14_14 ), .O(n6099));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4600_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17697_bdd_4_lut (.I0(n17697), .I1(\REG.mem_13_20 ), .I2(\REG.mem_12_20 ), 
            .I3(rd_addr_r[1]), .O(n15131));
    defparam n17697_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14847 (.I0(rd_addr_r[2]), .I1(n15746), 
            .I2(n15488), .I3(rd_addr_r[3]), .O(n16983));
    defparam rd_addr_r_2__bdd_4_lut_14847.LUT_INIT = 16'he4aa;
    SB_DFF wp_sync2_r__i5 (.Q(wp_sync2_r[5]), .C(SLM_CLK_c), .D(n7038));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i4 (.Q(wp_sync2_r[4]), .C(SLM_CLK_c), .D(n7037));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i3 (.Q(wp_sync2_r[3]), .C(SLM_CLK_c), .D(n7036));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i2 (.Q(wp_sync2_r[2]), .C(SLM_CLK_c), .D(n7035));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i1 (.Q(wp_sync2_r[1]), .C(SLM_CLK_c), .D(n7034));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i5 (.Q(wp_sync1_r[5]), .C(SLM_CLK_c), .D(n7033));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i4 (.Q(wp_sync1_r[4]), .C(SLM_CLK_c), .D(n7032));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i3 (.Q(wp_sync1_r[3]), .C(SLM_CLK_c), .D(n7031));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i2 (.Q(wp_sync1_r[2]), .C(SLM_CLK_c), .D(n7030));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i1 (.Q(wp_sync1_r[1]), .C(SLM_CLK_c), .D(n7029));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF rd_addr_r__i4 (.Q(rd_addr_r[4]), .C(SLM_CLK_c), .D(n7028));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i3 (.Q(rd_addr_r[3]), .C(SLM_CLK_c), .D(n7027));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .D(n7026));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(n7025));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_grey_sync_r__i5 (.Q(rd_grey_sync_r[5]), .C(SLM_CLK_c), .D(n7024));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFF rp_sync2_r__i5 (.Q(rp_sync2_r[5]), .C(FIFO_CLK_c), .D(n7023));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i4 (.Q(rp_sync2_r[4]), .C(FIFO_CLK_c), .D(n7022));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i3 (.Q(rp_sync2_r[3]), .C(FIFO_CLK_c), .D(n7021));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i2 (.Q(rp_sync2_r[2]), .C(FIFO_CLK_c), .D(n7020));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i1 (.Q(rp_sync2_r[1]), .C(FIFO_CLK_c), .D(n7019));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i5 (.Q(rp_sync1_r[5]), .C(FIFO_CLK_c), .D(n7018));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i4 (.Q(rp_sync1_r[4]), .C(FIFO_CLK_c), .D(n7017));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i3 (.Q(rp_sync1_r[3]), .C(FIFO_CLK_c), .D(n7016));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i2 (.Q(rp_sync1_r[2]), .C(FIFO_CLK_c), .D(n7015));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i1 (.Q(rp_sync1_r[1]), .C(FIFO_CLK_c), .D(n7014));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_LUT4 i5154_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_31_24 ), .O(n6653));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5154_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15312 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_3 ), 
            .I2(\REG.mem_31_3 ), .I3(rd_addr_r[1]), .O(n17691));
    defparam rd_addr_r_0__bdd_4_lut_15312.LUT_INIT = 16'he4aa;
    SB_LUT4 i4599_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_14_13 ), .O(n6098));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4599_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17691_bdd_4_lut (.I0(n17691), .I1(\REG.mem_29_3 ), .I2(\REG.mem_28_3 ), 
            .I3(rd_addr_r[1]), .O(n15605));
    defparam n17691_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(FIFO_CLK_c), .D(n6956));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(FIFO_CLK_c), .D(n6955));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i3 (.Q(wr_addr_r[3]), .C(FIFO_CLK_c), .D(n6954));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i4 (.Q(wr_addr_r[4]), .C(FIFO_CLK_c), .D(n6953));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i5 (.Q(\wr_addr_r[5] ), .C(FIFO_CLK_c), .D(n6952));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i3107_3108 (.Q(\REG.mem_31_31 ), .C(FIFO_CLK_c), .D(n6660));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3104_3105 (.Q(\REG.mem_31_30 ), .C(FIFO_CLK_c), .D(n6659));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3101_3102 (.Q(\REG.mem_31_29 ), .C(FIFO_CLK_c), .D(n6658));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3098_3099 (.Q(\REG.mem_31_28 ), .C(FIFO_CLK_c), .D(n6657));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3095_3096 (.Q(\REG.mem_31_27 ), .C(FIFO_CLK_c), .D(n6656));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3092_3093 (.Q(\REG.mem_31_26 ), .C(FIFO_CLK_c), .D(n6655));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3089_3090 (.Q(\REG.mem_31_25 ), .C(FIFO_CLK_c), .D(n6654));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3086_3087 (.Q(\REG.mem_31_24 ), .C(FIFO_CLK_c), .D(n6653));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3083_3084 (.Q(\REG.mem_31_23 ), .C(FIFO_CLK_c), .D(n6652));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3080_3081 (.Q(\REG.mem_31_22 ), .C(FIFO_CLK_c), .D(n6651));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3077_3078 (.Q(\REG.mem_31_21 ), .C(FIFO_CLK_c), .D(n6650));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3074_3075 (.Q(\REG.mem_31_20 ), .C(FIFO_CLK_c), .D(n6649));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3071_3072 (.Q(\REG.mem_31_19 ), .C(FIFO_CLK_c), .D(n6648));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3068_3069 (.Q(\REG.mem_31_18 ), .C(FIFO_CLK_c), .D(n6647));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3065_3066 (.Q(\REG.mem_31_17 ), .C(FIFO_CLK_c), .D(n6646));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3062_3063 (.Q(\REG.mem_31_16 ), .C(FIFO_CLK_c), .D(n6645));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3059_3060 (.Q(\REG.mem_31_15 ), .C(FIFO_CLK_c), .D(n6644));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3056_3057 (.Q(\REG.mem_31_14 ), .C(FIFO_CLK_c), .D(n6643));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3053_3054 (.Q(\REG.mem_31_13 ), .C(FIFO_CLK_c), .D(n6642));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3050_3051 (.Q(\REG.mem_31_12 ), .C(FIFO_CLK_c), .D(n6641));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3047_3048 (.Q(\REG.mem_31_11 ), .C(FIFO_CLK_c), .D(n6640));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3044_3045 (.Q(\REG.mem_31_10 ), .C(FIFO_CLK_c), .D(n6639));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3041_3042 (.Q(\REG.mem_31_9 ), .C(FIFO_CLK_c), .D(n6638));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3038_3039 (.Q(\REG.mem_31_8 ), .C(FIFO_CLK_c), .D(n6637));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3035_3036 (.Q(\REG.mem_31_7 ), .C(FIFO_CLK_c), .D(n6636));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3032_3033 (.Q(\REG.mem_31_6 ), .C(FIFO_CLK_c), .D(n6635));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3029_3030 (.Q(\REG.mem_31_5 ), .C(FIFO_CLK_c), .D(n6634));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3026_3027 (.Q(\REG.mem_31_4 ), .C(FIFO_CLK_c), .D(n6633));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3023_3024 (.Q(\REG.mem_31_3 ), .C(FIFO_CLK_c), .D(n6632));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3020_3021 (.Q(\REG.mem_31_2 ), .C(FIFO_CLK_c), .D(n6631));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3017_3018 (.Q(\REG.mem_31_1 ), .C(FIFO_CLK_c), .D(n6630));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3014_3015 (.Q(\REG.mem_31_0 ), .C(FIFO_CLK_c), .D(n6629));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3011_3012 (.Q(\REG.mem_30_31 ), .C(FIFO_CLK_c), .D(n6628));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3008_3009 (.Q(\REG.mem_30_30 ), .C(FIFO_CLK_c), .D(n6627));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3005_3006 (.Q(\REG.mem_30_29 ), .C(FIFO_CLK_c), .D(n6626));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3002_3003 (.Q(\REG.mem_30_28 ), .C(FIFO_CLK_c), .D(n6625));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2999_3000 (.Q(\REG.mem_30_27 ), .C(FIFO_CLK_c), .D(n6624));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2996_2997 (.Q(\REG.mem_30_26 ), .C(FIFO_CLK_c), .D(n6623));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2993_2994 (.Q(\REG.mem_30_25 ), .C(FIFO_CLK_c), .D(n6622));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2990_2991 (.Q(\REG.mem_30_24 ), .C(FIFO_CLK_c), .D(n6621));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2987_2988 (.Q(\REG.mem_30_23 ), .C(FIFO_CLK_c), .D(n6620));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2984_2985 (.Q(\REG.mem_30_22 ), .C(FIFO_CLK_c), .D(n6619));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2981_2982 (.Q(\REG.mem_30_21 ), .C(FIFO_CLK_c), .D(n6618));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2978_2979 (.Q(\REG.mem_30_20 ), .C(FIFO_CLK_c), .D(n6617));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2975_2976 (.Q(\REG.mem_30_19 ), .C(FIFO_CLK_c), .D(n6616));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2972_2973 (.Q(\REG.mem_30_18 ), .C(FIFO_CLK_c), .D(n6615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2969_2970 (.Q(\REG.mem_30_17 ), .C(FIFO_CLK_c), .D(n6614));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2966_2967 (.Q(\REG.mem_30_16 ), .C(FIFO_CLK_c), .D(n6613));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2963_2964 (.Q(\REG.mem_30_15 ), .C(FIFO_CLK_c), .D(n6612));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2960_2961 (.Q(\REG.mem_30_14 ), .C(FIFO_CLK_c), .D(n6611));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2957_2958 (.Q(\REG.mem_30_13 ), .C(FIFO_CLK_c), .D(n6610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2954_2955 (.Q(\REG.mem_30_12 ), .C(FIFO_CLK_c), .D(n6609));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2951_2952 (.Q(\REG.mem_30_11 ), .C(FIFO_CLK_c), .D(n6608));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2948_2949 (.Q(\REG.mem_30_10 ), .C(FIFO_CLK_c), .D(n6607));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2945_2946 (.Q(\REG.mem_30_9 ), .C(FIFO_CLK_c), .D(n6606));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2942_2943 (.Q(\REG.mem_30_8 ), .C(FIFO_CLK_c), .D(n6605));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2939_2940 (.Q(\REG.mem_30_7 ), .C(FIFO_CLK_c), .D(n6604));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2936_2937 (.Q(\REG.mem_30_6 ), .C(FIFO_CLK_c), .D(n6603));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2933_2934 (.Q(\REG.mem_30_5 ), .C(FIFO_CLK_c), .D(n6602));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2930_2931 (.Q(\REG.mem_30_4 ), .C(FIFO_CLK_c), .D(n6601));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2927_2928 (.Q(\REG.mem_30_3 ), .C(FIFO_CLK_c), .D(n6600));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2924_2925 (.Q(\REG.mem_30_2 ), .C(FIFO_CLK_c), .D(n6599));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2921_2922 (.Q(\REG.mem_30_1 ), .C(FIFO_CLK_c), .D(n6598));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2918_2919 (.Q(\REG.mem_30_0 ), .C(FIFO_CLK_c), .D(n6597));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2915_2916 (.Q(\REG.mem_29_31 ), .C(FIFO_CLK_c), .D(n6596));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2912_2913 (.Q(\REG.mem_29_30 ), .C(FIFO_CLK_c), .D(n6595));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2909_2910 (.Q(\REG.mem_29_29 ), .C(FIFO_CLK_c), .D(n6594));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2906_2907 (.Q(\REG.mem_29_28 ), .C(FIFO_CLK_c), .D(n6593));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2903_2904 (.Q(\REG.mem_29_27 ), .C(FIFO_CLK_c), .D(n6592));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2900_2901 (.Q(\REG.mem_29_26 ), .C(FIFO_CLK_c), .D(n6591));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2897_2898 (.Q(\REG.mem_29_25 ), .C(FIFO_CLK_c), .D(n6590));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2894_2895 (.Q(\REG.mem_29_24 ), .C(FIFO_CLK_c), .D(n6589));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2891_2892 (.Q(\REG.mem_29_23 ), .C(FIFO_CLK_c), .D(n6588));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2888_2889 (.Q(\REG.mem_29_22 ), .C(FIFO_CLK_c), .D(n6587));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2885_2886 (.Q(\REG.mem_29_21 ), .C(FIFO_CLK_c), .D(n6586));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2882_2883 (.Q(\REG.mem_29_20 ), .C(FIFO_CLK_c), .D(n6585));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2879_2880 (.Q(\REG.mem_29_19 ), .C(FIFO_CLK_c), .D(n6584));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2876_2877 (.Q(\REG.mem_29_18 ), .C(FIFO_CLK_c), .D(n6583));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2873_2874 (.Q(\REG.mem_29_17 ), .C(FIFO_CLK_c), .D(n6582));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2870_2871 (.Q(\REG.mem_29_16 ), .C(FIFO_CLK_c), .D(n6581));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2867_2868 (.Q(\REG.mem_29_15 ), .C(FIFO_CLK_c), .D(n6580));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2864_2865 (.Q(\REG.mem_29_14 ), .C(FIFO_CLK_c), .D(n6579));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2861_2862 (.Q(\REG.mem_29_13 ), .C(FIFO_CLK_c), .D(n6578));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2858_2859 (.Q(\REG.mem_29_12 ), .C(FIFO_CLK_c), .D(n6577));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2855_2856 (.Q(\REG.mem_29_11 ), .C(FIFO_CLK_c), .D(n6576));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2852_2853 (.Q(\REG.mem_29_10 ), .C(FIFO_CLK_c), .D(n6575));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2849_2850 (.Q(\REG.mem_29_9 ), .C(FIFO_CLK_c), .D(n6574));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2846_2847 (.Q(\REG.mem_29_8 ), .C(FIFO_CLK_c), .D(n6573));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2843_2844 (.Q(\REG.mem_29_7 ), .C(FIFO_CLK_c), .D(n6572));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2840_2841 (.Q(\REG.mem_29_6 ), .C(FIFO_CLK_c), .D(n6571));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2837_2838 (.Q(\REG.mem_29_5 ), .C(FIFO_CLK_c), .D(n6570));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2834_2835 (.Q(\REG.mem_29_4 ), .C(FIFO_CLK_c), .D(n6569));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2831_2832 (.Q(\REG.mem_29_3 ), .C(FIFO_CLK_c), .D(n6568));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2828_2829 (.Q(\REG.mem_29_2 ), .C(FIFO_CLK_c), .D(n6567));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2825_2826 (.Q(\REG.mem_29_1 ), .C(FIFO_CLK_c), .D(n6566));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2822_2823 (.Q(\REG.mem_29_0 ), .C(FIFO_CLK_c), .D(n6565));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2819_2820 (.Q(\REG.mem_28_31 ), .C(FIFO_CLK_c), .D(n6564));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2816_2817 (.Q(\REG.mem_28_30 ), .C(FIFO_CLK_c), .D(n6563));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2813_2814 (.Q(\REG.mem_28_29 ), .C(FIFO_CLK_c), .D(n6562));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2810_2811 (.Q(\REG.mem_28_28 ), .C(FIFO_CLK_c), .D(n6561));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2807_2808 (.Q(\REG.mem_28_27 ), .C(FIFO_CLK_c), .D(n6560));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2804_2805 (.Q(\REG.mem_28_26 ), .C(FIFO_CLK_c), .D(n6559));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2801_2802 (.Q(\REG.mem_28_25 ), .C(FIFO_CLK_c), .D(n6558));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2798_2799 (.Q(\REG.mem_28_24 ), .C(FIFO_CLK_c), .D(n6557));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2795_2796 (.Q(\REG.mem_28_23 ), .C(FIFO_CLK_c), .D(n6556));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2792_2793 (.Q(\REG.mem_28_22 ), .C(FIFO_CLK_c), .D(n6555));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2789_2790 (.Q(\REG.mem_28_21 ), .C(FIFO_CLK_c), .D(n6554));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2786_2787 (.Q(\REG.mem_28_20 ), .C(FIFO_CLK_c), .D(n6553));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2783_2784 (.Q(\REG.mem_28_19 ), .C(FIFO_CLK_c), .D(n6552));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2780_2781 (.Q(\REG.mem_28_18 ), .C(FIFO_CLK_c), .D(n6551));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2777_2778 (.Q(\REG.mem_28_17 ), .C(FIFO_CLK_c), .D(n6550));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2774_2775 (.Q(\REG.mem_28_16 ), .C(FIFO_CLK_c), .D(n6549));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2771_2772 (.Q(\REG.mem_28_15 ), .C(FIFO_CLK_c), .D(n6548));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2768_2769 (.Q(\REG.mem_28_14 ), .C(FIFO_CLK_c), .D(n6547));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2765_2766 (.Q(\REG.mem_28_13 ), .C(FIFO_CLK_c), .D(n6546));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2762_2763 (.Q(\REG.mem_28_12 ), .C(FIFO_CLK_c), .D(n6545));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2759_2760 (.Q(\REG.mem_28_11 ), .C(FIFO_CLK_c), .D(n6544));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2756_2757 (.Q(\REG.mem_28_10 ), .C(FIFO_CLK_c), .D(n6543));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2753_2754 (.Q(\REG.mem_28_9 ), .C(FIFO_CLK_c), .D(n6542));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2750_2751 (.Q(\REG.mem_28_8 ), .C(FIFO_CLK_c), .D(n6541));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2747_2748 (.Q(\REG.mem_28_7 ), .C(FIFO_CLK_c), .D(n6540));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2744_2745 (.Q(\REG.mem_28_6 ), .C(FIFO_CLK_c), .D(n6539));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2741_2742 (.Q(\REG.mem_28_5 ), .C(FIFO_CLK_c), .D(n6538));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2738_2739 (.Q(\REG.mem_28_4 ), .C(FIFO_CLK_c), .D(n6537));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2735_2736 (.Q(\REG.mem_28_3 ), .C(FIFO_CLK_c), .D(n6536));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2732_2733 (.Q(\REG.mem_28_2 ), .C(FIFO_CLK_c), .D(n6535));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2729_2730 (.Q(\REG.mem_28_1 ), .C(FIFO_CLK_c), .D(n6534));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2726_2727 (.Q(\REG.mem_28_0 ), .C(FIFO_CLK_c), .D(n6533));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2723_2724 (.Q(\REG.mem_27_31 ), .C(FIFO_CLK_c), .D(n6532));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2720_2721 (.Q(\REG.mem_27_30 ), .C(FIFO_CLK_c), .D(n6531));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2717_2718 (.Q(\REG.mem_27_29 ), .C(FIFO_CLK_c), .D(n6530));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2714_2715 (.Q(\REG.mem_27_28 ), .C(FIFO_CLK_c), .D(n6529));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2711_2712 (.Q(\REG.mem_27_27 ), .C(FIFO_CLK_c), .D(n6528));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2708_2709 (.Q(\REG.mem_27_26 ), .C(FIFO_CLK_c), .D(n6527));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2705_2706 (.Q(\REG.mem_27_25 ), .C(FIFO_CLK_c), .D(n6526));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2702_2703 (.Q(\REG.mem_27_24 ), .C(FIFO_CLK_c), .D(n6525));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2699_2700 (.Q(\REG.mem_27_23 ), .C(FIFO_CLK_c), .D(n6524));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2696_2697 (.Q(\REG.mem_27_22 ), .C(FIFO_CLK_c), .D(n6523));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2693_2694 (.Q(\REG.mem_27_21 ), .C(FIFO_CLK_c), .D(n6522));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2690_2691 (.Q(\REG.mem_27_20 ), .C(FIFO_CLK_c), .D(n6521));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2687_2688 (.Q(\REG.mem_27_19 ), .C(FIFO_CLK_c), .D(n6520));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2684_2685 (.Q(\REG.mem_27_18 ), .C(FIFO_CLK_c), .D(n6519));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2681_2682 (.Q(\REG.mem_27_17 ), .C(FIFO_CLK_c), .D(n6518));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2678_2679 (.Q(\REG.mem_27_16 ), .C(FIFO_CLK_c), .D(n6517));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2675_2676 (.Q(\REG.mem_27_15 ), .C(FIFO_CLK_c), .D(n6516));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2672_2673 (.Q(\REG.mem_27_14 ), .C(FIFO_CLK_c), .D(n6515));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2669_2670 (.Q(\REG.mem_27_13 ), .C(FIFO_CLK_c), .D(n6514));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2666_2667 (.Q(\REG.mem_27_12 ), .C(FIFO_CLK_c), .D(n6513));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2663_2664 (.Q(\REG.mem_27_11 ), .C(FIFO_CLK_c), .D(n6512));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2660_2661 (.Q(\REG.mem_27_10 ), .C(FIFO_CLK_c), .D(n6511));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2657_2658 (.Q(\REG.mem_27_9 ), .C(FIFO_CLK_c), .D(n6510));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2654_2655 (.Q(\REG.mem_27_8 ), .C(FIFO_CLK_c), .D(n6509));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2651_2652 (.Q(\REG.mem_27_7 ), .C(FIFO_CLK_c), .D(n6508));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2648_2649 (.Q(\REG.mem_27_6 ), .C(FIFO_CLK_c), .D(n6507));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2645_2646 (.Q(\REG.mem_27_5 ), .C(FIFO_CLK_c), .D(n6506));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2642_2643 (.Q(\REG.mem_27_4 ), .C(FIFO_CLK_c), .D(n6505));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2639_2640 (.Q(\REG.mem_27_3 ), .C(FIFO_CLK_c), .D(n6504));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2636_2637 (.Q(\REG.mem_27_2 ), .C(FIFO_CLK_c), .D(n6503));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2633_2634 (.Q(\REG.mem_27_1 ), .C(FIFO_CLK_c), .D(n6502));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2630_2631 (.Q(\REG.mem_27_0 ), .C(FIFO_CLK_c), .D(n6501));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2627_2628 (.Q(\REG.mem_26_31 ), .C(FIFO_CLK_c), .D(n6500));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2624_2625 (.Q(\REG.mem_26_30 ), .C(FIFO_CLK_c), .D(n6499));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2621_2622 (.Q(\REG.mem_26_29 ), .C(FIFO_CLK_c), .D(n6498));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2618_2619 (.Q(\REG.mem_26_28 ), .C(FIFO_CLK_c), .D(n6497));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2615_2616 (.Q(\REG.mem_26_27 ), .C(FIFO_CLK_c), .D(n6496));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2612_2613 (.Q(\REG.mem_26_26 ), .C(FIFO_CLK_c), .D(n6495));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2609_2610 (.Q(\REG.mem_26_25 ), .C(FIFO_CLK_c), .D(n6494));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2606_2607 (.Q(\REG.mem_26_24 ), .C(FIFO_CLK_c), .D(n6493));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2603_2604 (.Q(\REG.mem_26_23 ), .C(FIFO_CLK_c), .D(n6492));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2600_2601 (.Q(\REG.mem_26_22 ), .C(FIFO_CLK_c), .D(n6491));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2597_2598 (.Q(\REG.mem_26_21 ), .C(FIFO_CLK_c), .D(n6490));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2594_2595 (.Q(\REG.mem_26_20 ), .C(FIFO_CLK_c), .D(n6489));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2591_2592 (.Q(\REG.mem_26_19 ), .C(FIFO_CLK_c), .D(n6488));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2588_2589 (.Q(\REG.mem_26_18 ), .C(FIFO_CLK_c), .D(n6487));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2585_2586 (.Q(\REG.mem_26_17 ), .C(FIFO_CLK_c), .D(n6486));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2582_2583 (.Q(\REG.mem_26_16 ), .C(FIFO_CLK_c), .D(n6485));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2579_2580 (.Q(\REG.mem_26_15 ), .C(FIFO_CLK_c), .D(n6484));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2576_2577 (.Q(\REG.mem_26_14 ), .C(FIFO_CLK_c), .D(n6483));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2573_2574 (.Q(\REG.mem_26_13 ), .C(FIFO_CLK_c), .D(n6482));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2570_2571 (.Q(\REG.mem_26_12 ), .C(FIFO_CLK_c), .D(n6481));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2567_2568 (.Q(\REG.mem_26_11 ), .C(FIFO_CLK_c), .D(n6480));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2564_2565 (.Q(\REG.mem_26_10 ), .C(FIFO_CLK_c), .D(n6479));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2561_2562 (.Q(\REG.mem_26_9 ), .C(FIFO_CLK_c), .D(n6478));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2558_2559 (.Q(\REG.mem_26_8 ), .C(FIFO_CLK_c), .D(n6477));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2555_2556 (.Q(\REG.mem_26_7 ), .C(FIFO_CLK_c), .D(n6476));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2552_2553 (.Q(\REG.mem_26_6 ), .C(FIFO_CLK_c), .D(n6475));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2549_2550 (.Q(\REG.mem_26_5 ), .C(FIFO_CLK_c), .D(n6474));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2546_2547 (.Q(\REG.mem_26_4 ), .C(FIFO_CLK_c), .D(n6473));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2543_2544 (.Q(\REG.mem_26_3 ), .C(FIFO_CLK_c), .D(n6472));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2540_2541 (.Q(\REG.mem_26_2 ), .C(FIFO_CLK_c), .D(n6471));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2537_2538 (.Q(\REG.mem_26_1 ), .C(FIFO_CLK_c), .D(n6470));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2534_2535 (.Q(\REG.mem_26_0 ), .C(FIFO_CLK_c), .D(n6469));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2531_2532 (.Q(\REG.mem_25_31 ), .C(FIFO_CLK_c), .D(n6468));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2528_2529 (.Q(\REG.mem_25_30 ), .C(FIFO_CLK_c), .D(n6467));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2525_2526 (.Q(\REG.mem_25_29 ), .C(FIFO_CLK_c), .D(n6466));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2522_2523 (.Q(\REG.mem_25_28 ), .C(FIFO_CLK_c), .D(n6465));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2519_2520 (.Q(\REG.mem_25_27 ), .C(FIFO_CLK_c), .D(n6464));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2516_2517 (.Q(\REG.mem_25_26 ), .C(FIFO_CLK_c), .D(n6463));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2513_2514 (.Q(\REG.mem_25_25 ), .C(FIFO_CLK_c), .D(n6462));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2510_2511 (.Q(\REG.mem_25_24 ), .C(FIFO_CLK_c), .D(n6461));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2507_2508 (.Q(\REG.mem_25_23 ), .C(FIFO_CLK_c), .D(n6460));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2504_2505 (.Q(\REG.mem_25_22 ), .C(FIFO_CLK_c), .D(n6459));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2501_2502 (.Q(\REG.mem_25_21 ), .C(FIFO_CLK_c), .D(n6458));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2498_2499 (.Q(\REG.mem_25_20 ), .C(FIFO_CLK_c), .D(n6457));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2495_2496 (.Q(\REG.mem_25_19 ), .C(FIFO_CLK_c), .D(n6456));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2492_2493 (.Q(\REG.mem_25_18 ), .C(FIFO_CLK_c), .D(n6455));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2489_2490 (.Q(\REG.mem_25_17 ), .C(FIFO_CLK_c), .D(n6454));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2486_2487 (.Q(\REG.mem_25_16 ), .C(FIFO_CLK_c), .D(n6453));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2483_2484 (.Q(\REG.mem_25_15 ), .C(FIFO_CLK_c), .D(n6452));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2480_2481 (.Q(\REG.mem_25_14 ), .C(FIFO_CLK_c), .D(n6451));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2477_2478 (.Q(\REG.mem_25_13 ), .C(FIFO_CLK_c), .D(n6450));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2474_2475 (.Q(\REG.mem_25_12 ), .C(FIFO_CLK_c), .D(n6449));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2471_2472 (.Q(\REG.mem_25_11 ), .C(FIFO_CLK_c), .D(n6448));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2468_2469 (.Q(\REG.mem_25_10 ), .C(FIFO_CLK_c), .D(n6447));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2465_2466 (.Q(\REG.mem_25_9 ), .C(FIFO_CLK_c), .D(n6446));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2462_2463 (.Q(\REG.mem_25_8 ), .C(FIFO_CLK_c), .D(n6445));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2459_2460 (.Q(\REG.mem_25_7 ), .C(FIFO_CLK_c), .D(n6444));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2456_2457 (.Q(\REG.mem_25_6 ), .C(FIFO_CLK_c), .D(n6443));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2453_2454 (.Q(\REG.mem_25_5 ), .C(FIFO_CLK_c), .D(n6442));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2450_2451 (.Q(\REG.mem_25_4 ), .C(FIFO_CLK_c), .D(n6441));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2447_2448 (.Q(\REG.mem_25_3 ), .C(FIFO_CLK_c), .D(n6440));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2444_2445 (.Q(\REG.mem_25_2 ), .C(FIFO_CLK_c), .D(n6439));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2441_2442 (.Q(\REG.mem_25_1 ), .C(FIFO_CLK_c), .D(n6438));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2438_2439 (.Q(\REG.mem_25_0 ), .C(FIFO_CLK_c), .D(n6437));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2435_2436 (.Q(\REG.mem_24_31 ), .C(FIFO_CLK_c), .D(n6436));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2432_2433 (.Q(\REG.mem_24_30 ), .C(FIFO_CLK_c), .D(n6435));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2429_2430 (.Q(\REG.mem_24_29 ), .C(FIFO_CLK_c), .D(n6434));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2426_2427 (.Q(\REG.mem_24_28 ), .C(FIFO_CLK_c), .D(n6433));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2423_2424 (.Q(\REG.mem_24_27 ), .C(FIFO_CLK_c), .D(n6432));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2420_2421 (.Q(\REG.mem_24_26 ), .C(FIFO_CLK_c), .D(n6431));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2417_2418 (.Q(\REG.mem_24_25 ), .C(FIFO_CLK_c), .D(n6430));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2414_2415 (.Q(\REG.mem_24_24 ), .C(FIFO_CLK_c), .D(n6429));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2411_2412 (.Q(\REG.mem_24_23 ), .C(FIFO_CLK_c), .D(n6428));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2408_2409 (.Q(\REG.mem_24_22 ), .C(FIFO_CLK_c), .D(n6427));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2405_2406 (.Q(\REG.mem_24_21 ), .C(FIFO_CLK_c), .D(n6426));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2402_2403 (.Q(\REG.mem_24_20 ), .C(FIFO_CLK_c), .D(n6425));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2399_2400 (.Q(\REG.mem_24_19 ), .C(FIFO_CLK_c), .D(n6424));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2396_2397 (.Q(\REG.mem_24_18 ), .C(FIFO_CLK_c), .D(n6423));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2393_2394 (.Q(\REG.mem_24_17 ), .C(FIFO_CLK_c), .D(n6422));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2390_2391 (.Q(\REG.mem_24_16 ), .C(FIFO_CLK_c), .D(n6421));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2387_2388 (.Q(\REG.mem_24_15 ), .C(FIFO_CLK_c), .D(n6420));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2384_2385 (.Q(\REG.mem_24_14 ), .C(FIFO_CLK_c), .D(n6419));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2381_2382 (.Q(\REG.mem_24_13 ), .C(FIFO_CLK_c), .D(n6418));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2378_2379 (.Q(\REG.mem_24_12 ), .C(FIFO_CLK_c), .D(n6417));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2375_2376 (.Q(\REG.mem_24_11 ), .C(FIFO_CLK_c), .D(n6416));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2372_2373 (.Q(\REG.mem_24_10 ), .C(FIFO_CLK_c), .D(n6415));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2369_2370 (.Q(\REG.mem_24_9 ), .C(FIFO_CLK_c), .D(n6414));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2366_2367 (.Q(\REG.mem_24_8 ), .C(FIFO_CLK_c), .D(n6413));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2363_2364 (.Q(\REG.mem_24_7 ), .C(FIFO_CLK_c), .D(n6412));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2360_2361 (.Q(\REG.mem_24_6 ), .C(FIFO_CLK_c), .D(n6411));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2357_2358 (.Q(\REG.mem_24_5 ), .C(FIFO_CLK_c), .D(n6410));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2354_2355 (.Q(\REG.mem_24_4 ), .C(FIFO_CLK_c), .D(n6409));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2351_2352 (.Q(\REG.mem_24_3 ), .C(FIFO_CLK_c), .D(n6408));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2348_2349 (.Q(\REG.mem_24_2 ), .C(FIFO_CLK_c), .D(n6407));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2345_2346 (.Q(\REG.mem_24_1 ), .C(FIFO_CLK_c), .D(n6406));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2342_2343 (.Q(\REG.mem_24_0 ), .C(FIFO_CLK_c), .D(n6405));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2339_2340 (.Q(\REG.mem_23_31 ), .C(FIFO_CLK_c), .D(n6404));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2336_2337 (.Q(\REG.mem_23_30 ), .C(FIFO_CLK_c), .D(n6403));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2333_2334 (.Q(\REG.mem_23_29 ), .C(FIFO_CLK_c), .D(n6402));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2330_2331 (.Q(\REG.mem_23_28 ), .C(FIFO_CLK_c), .D(n6401));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2327_2328 (.Q(\REG.mem_23_27 ), .C(FIFO_CLK_c), .D(n6400));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2324_2325 (.Q(\REG.mem_23_26 ), .C(FIFO_CLK_c), .D(n6399));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2321_2322 (.Q(\REG.mem_23_25 ), .C(FIFO_CLK_c), .D(n6398));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2318_2319 (.Q(\REG.mem_23_24 ), .C(FIFO_CLK_c), .D(n6397));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2315_2316 (.Q(\REG.mem_23_23 ), .C(FIFO_CLK_c), .D(n6396));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2312_2313 (.Q(\REG.mem_23_22 ), .C(FIFO_CLK_c), .D(n6395));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2309_2310 (.Q(\REG.mem_23_21 ), .C(FIFO_CLK_c), .D(n6394));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2306_2307 (.Q(\REG.mem_23_20 ), .C(FIFO_CLK_c), .D(n6393));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2303_2304 (.Q(\REG.mem_23_19 ), .C(FIFO_CLK_c), .D(n6392));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2300_2301 (.Q(\REG.mem_23_18 ), .C(FIFO_CLK_c), .D(n6391));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2297_2298 (.Q(\REG.mem_23_17 ), .C(FIFO_CLK_c), .D(n6390));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2294_2295 (.Q(\REG.mem_23_16 ), .C(FIFO_CLK_c), .D(n6389));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2291_2292 (.Q(\REG.mem_23_15 ), .C(FIFO_CLK_c), .D(n6388));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2288_2289 (.Q(\REG.mem_23_14 ), .C(FIFO_CLK_c), .D(n6387));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2285_2286 (.Q(\REG.mem_23_13 ), .C(FIFO_CLK_c), .D(n6386));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2282_2283 (.Q(\REG.mem_23_12 ), .C(FIFO_CLK_c), .D(n6385));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2279_2280 (.Q(\REG.mem_23_11 ), .C(FIFO_CLK_c), .D(n6384));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2276_2277 (.Q(\REG.mem_23_10 ), .C(FIFO_CLK_c), .D(n6383));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2273_2274 (.Q(\REG.mem_23_9 ), .C(FIFO_CLK_c), .D(n6382));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2270_2271 (.Q(\REG.mem_23_8 ), .C(FIFO_CLK_c), .D(n6381));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2267_2268 (.Q(\REG.mem_23_7 ), .C(FIFO_CLK_c), .D(n6380));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2264_2265 (.Q(\REG.mem_23_6 ), .C(FIFO_CLK_c), .D(n6379));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2261_2262 (.Q(\REG.mem_23_5 ), .C(FIFO_CLK_c), .D(n6378));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2258_2259 (.Q(\REG.mem_23_4 ), .C(FIFO_CLK_c), .D(n6377));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2255_2256 (.Q(\REG.mem_23_3 ), .C(FIFO_CLK_c), .D(n6376));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2252_2253 (.Q(\REG.mem_23_2 ), .C(FIFO_CLK_c), .D(n6375));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2249_2250 (.Q(\REG.mem_23_1 ), .C(FIFO_CLK_c), .D(n6374));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2246_2247 (.Q(\REG.mem_23_0 ), .C(FIFO_CLK_c), .D(n6373));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2243_2244 (.Q(\REG.mem_22_31 ), .C(FIFO_CLK_c), .D(n6372));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2240_2241 (.Q(\REG.mem_22_30 ), .C(FIFO_CLK_c), .D(n6371));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2237_2238 (.Q(\REG.mem_22_29 ), .C(FIFO_CLK_c), .D(n6370));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2234_2235 (.Q(\REG.mem_22_28 ), .C(FIFO_CLK_c), .D(n6369));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2231_2232 (.Q(\REG.mem_22_27 ), .C(FIFO_CLK_c), .D(n6368));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2228_2229 (.Q(\REG.mem_22_26 ), .C(FIFO_CLK_c), .D(n6367));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2225_2226 (.Q(\REG.mem_22_25 ), .C(FIFO_CLK_c), .D(n6366));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2222_2223 (.Q(\REG.mem_22_24 ), .C(FIFO_CLK_c), .D(n6365));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2219_2220 (.Q(\REG.mem_22_23 ), .C(FIFO_CLK_c), .D(n6364));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2216_2217 (.Q(\REG.mem_22_22 ), .C(FIFO_CLK_c), .D(n6363));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2213_2214 (.Q(\REG.mem_22_21 ), .C(FIFO_CLK_c), .D(n6362));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2210_2211 (.Q(\REG.mem_22_20 ), .C(FIFO_CLK_c), .D(n6361));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2207_2208 (.Q(\REG.mem_22_19 ), .C(FIFO_CLK_c), .D(n6360));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2204_2205 (.Q(\REG.mem_22_18 ), .C(FIFO_CLK_c), .D(n6359));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2201_2202 (.Q(\REG.mem_22_17 ), .C(FIFO_CLK_c), .D(n6358));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2198_2199 (.Q(\REG.mem_22_16 ), .C(FIFO_CLK_c), .D(n6357));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2195_2196 (.Q(\REG.mem_22_15 ), .C(FIFO_CLK_c), .D(n6356));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2192_2193 (.Q(\REG.mem_22_14 ), .C(FIFO_CLK_c), .D(n6355));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2189_2190 (.Q(\REG.mem_22_13 ), .C(FIFO_CLK_c), .D(n6354));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2186_2187 (.Q(\REG.mem_22_12 ), .C(FIFO_CLK_c), .D(n6353));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2183_2184 (.Q(\REG.mem_22_11 ), .C(FIFO_CLK_c), .D(n6352));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2180_2181 (.Q(\REG.mem_22_10 ), .C(FIFO_CLK_c), .D(n6351));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2177_2178 (.Q(\REG.mem_22_9 ), .C(FIFO_CLK_c), .D(n6350));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2174_2175 (.Q(\REG.mem_22_8 ), .C(FIFO_CLK_c), .D(n6349));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2171_2172 (.Q(\REG.mem_22_7 ), .C(FIFO_CLK_c), .D(n6348));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2168_2169 (.Q(\REG.mem_22_6 ), .C(FIFO_CLK_c), .D(n6347));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2165_2166 (.Q(\REG.mem_22_5 ), .C(FIFO_CLK_c), .D(n6346));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2162_2163 (.Q(\REG.mem_22_4 ), .C(FIFO_CLK_c), .D(n6345));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2159_2160 (.Q(\REG.mem_22_3 ), .C(FIFO_CLK_c), .D(n6344));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2156_2157 (.Q(\REG.mem_22_2 ), .C(FIFO_CLK_c), .D(n6343));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2153_2154 (.Q(\REG.mem_22_1 ), .C(FIFO_CLK_c), .D(n6342));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2150_2151 (.Q(\REG.mem_22_0 ), .C(FIFO_CLK_c), .D(n6341));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2147_2148 (.Q(\REG.mem_21_31 ), .C(FIFO_CLK_c), .D(n6340));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2144_2145 (.Q(\REG.mem_21_30 ), .C(FIFO_CLK_c), .D(n6339));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2141_2142 (.Q(\REG.mem_21_29 ), .C(FIFO_CLK_c), .D(n6338));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2138_2139 (.Q(\REG.mem_21_28 ), .C(FIFO_CLK_c), .D(n6337));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2135_2136 (.Q(\REG.mem_21_27 ), .C(FIFO_CLK_c), .D(n6336));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2132_2133 (.Q(\REG.mem_21_26 ), .C(FIFO_CLK_c), .D(n6335));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2129_2130 (.Q(\REG.mem_21_25 ), .C(FIFO_CLK_c), .D(n6334));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2126_2127 (.Q(\REG.mem_21_24 ), .C(FIFO_CLK_c), .D(n6333));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2123_2124 (.Q(\REG.mem_21_23 ), .C(FIFO_CLK_c), .D(n6332));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2120_2121 (.Q(\REG.mem_21_22 ), .C(FIFO_CLK_c), .D(n6331));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2117_2118 (.Q(\REG.mem_21_21 ), .C(FIFO_CLK_c), .D(n6330));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2114_2115 (.Q(\REG.mem_21_20 ), .C(FIFO_CLK_c), .D(n6329));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2111_2112 (.Q(\REG.mem_21_19 ), .C(FIFO_CLK_c), .D(n6328));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2108_2109 (.Q(\REG.mem_21_18 ), .C(FIFO_CLK_c), .D(n6327));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2105_2106 (.Q(\REG.mem_21_17 ), .C(FIFO_CLK_c), .D(n6326));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2102_2103 (.Q(\REG.mem_21_16 ), .C(FIFO_CLK_c), .D(n6325));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2099_2100 (.Q(\REG.mem_21_15 ), .C(FIFO_CLK_c), .D(n6324));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2096_2097 (.Q(\REG.mem_21_14 ), .C(FIFO_CLK_c), .D(n6323));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2093_2094 (.Q(\REG.mem_21_13 ), .C(FIFO_CLK_c), .D(n6322));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2090_2091 (.Q(\REG.mem_21_12 ), .C(FIFO_CLK_c), .D(n6321));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2087_2088 (.Q(\REG.mem_21_11 ), .C(FIFO_CLK_c), .D(n6320));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2084_2085 (.Q(\REG.mem_21_10 ), .C(FIFO_CLK_c), .D(n6319));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2081_2082 (.Q(\REG.mem_21_9 ), .C(FIFO_CLK_c), .D(n6318));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2078_2079 (.Q(\REG.mem_21_8 ), .C(FIFO_CLK_c), .D(n6317));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2075_2076 (.Q(\REG.mem_21_7 ), .C(FIFO_CLK_c), .D(n6316));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2072_2073 (.Q(\REG.mem_21_6 ), .C(FIFO_CLK_c), .D(n6315));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2069_2070 (.Q(\REG.mem_21_5 ), .C(FIFO_CLK_c), .D(n6314));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2066_2067 (.Q(\REG.mem_21_4 ), .C(FIFO_CLK_c), .D(n6313));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2063_2064 (.Q(\REG.mem_21_3 ), .C(FIFO_CLK_c), .D(n6312));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2060_2061 (.Q(\REG.mem_21_2 ), .C(FIFO_CLK_c), .D(n6311));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2057_2058 (.Q(\REG.mem_21_1 ), .C(FIFO_CLK_c), .D(n6310));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2054_2055 (.Q(\REG.mem_21_0 ), .C(FIFO_CLK_c), .D(n6309));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2051_2052 (.Q(\REG.mem_20_31 ), .C(FIFO_CLK_c), .D(n6308));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2048_2049 (.Q(\REG.mem_20_30 ), .C(FIFO_CLK_c), .D(n6307));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2045_2046 (.Q(\REG.mem_20_29 ), .C(FIFO_CLK_c), .D(n6306));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2042_2043 (.Q(\REG.mem_20_28 ), .C(FIFO_CLK_c), .D(n6305));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2039_2040 (.Q(\REG.mem_20_27 ), .C(FIFO_CLK_c), .D(n6304));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2036_2037 (.Q(\REG.mem_20_26 ), .C(FIFO_CLK_c), .D(n6303));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2033_2034 (.Q(\REG.mem_20_25 ), .C(FIFO_CLK_c), .D(n6302));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2030_2031 (.Q(\REG.mem_20_24 ), .C(FIFO_CLK_c), .D(n6301));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2027_2028 (.Q(\REG.mem_20_23 ), .C(FIFO_CLK_c), .D(n6300));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2024_2025 (.Q(\REG.mem_20_22 ), .C(FIFO_CLK_c), .D(n6299));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2021_2022 (.Q(\REG.mem_20_21 ), .C(FIFO_CLK_c), .D(n6298));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2018_2019 (.Q(\REG.mem_20_20 ), .C(FIFO_CLK_c), .D(n6297));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2015_2016 (.Q(\REG.mem_20_19 ), .C(FIFO_CLK_c), .D(n6296));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2012_2013 (.Q(\REG.mem_20_18 ), .C(FIFO_CLK_c), .D(n6295));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2009_2010 (.Q(\REG.mem_20_17 ), .C(FIFO_CLK_c), .D(n6294));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2006_2007 (.Q(\REG.mem_20_16 ), .C(FIFO_CLK_c), .D(n6293));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2003_2004 (.Q(\REG.mem_20_15 ), .C(FIFO_CLK_c), .D(n6292));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2000_2001 (.Q(\REG.mem_20_14 ), .C(FIFO_CLK_c), .D(n6291));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1997_1998 (.Q(\REG.mem_20_13 ), .C(FIFO_CLK_c), .D(n6290));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1994_1995 (.Q(\REG.mem_20_12 ), .C(FIFO_CLK_c), .D(n6289));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1991_1992 (.Q(\REG.mem_20_11 ), .C(FIFO_CLK_c), .D(n6288));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1988_1989 (.Q(\REG.mem_20_10 ), .C(FIFO_CLK_c), .D(n6287));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1985_1986 (.Q(\REG.mem_20_9 ), .C(FIFO_CLK_c), .D(n6286));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1982_1983 (.Q(\REG.mem_20_8 ), .C(FIFO_CLK_c), .D(n6285));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1979_1980 (.Q(\REG.mem_20_7 ), .C(FIFO_CLK_c), .D(n6284));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1976_1977 (.Q(\REG.mem_20_6 ), .C(FIFO_CLK_c), .D(n6283));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1973_1974 (.Q(\REG.mem_20_5 ), .C(FIFO_CLK_c), .D(n6282));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1970_1971 (.Q(\REG.mem_20_4 ), .C(FIFO_CLK_c), .D(n6281));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1967_1968 (.Q(\REG.mem_20_3 ), .C(FIFO_CLK_c), .D(n6280));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1964_1965 (.Q(\REG.mem_20_2 ), .C(FIFO_CLK_c), .D(n6279));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1961_1962 (.Q(\REG.mem_20_1 ), .C(FIFO_CLK_c), .D(n6278));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1958_1959 (.Q(\REG.mem_20_0 ), .C(FIFO_CLK_c), .D(n6277));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1955_1956 (.Q(\REG.mem_19_31 ), .C(FIFO_CLK_c), .D(n6276));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1952_1953 (.Q(\REG.mem_19_30 ), .C(FIFO_CLK_c), .D(n6275));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1949_1950 (.Q(\REG.mem_19_29 ), .C(FIFO_CLK_c), .D(n6274));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1946_1947 (.Q(\REG.mem_19_28 ), .C(FIFO_CLK_c), .D(n6273));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1943_1944 (.Q(\REG.mem_19_27 ), .C(FIFO_CLK_c), .D(n6272));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1940_1941 (.Q(\REG.mem_19_26 ), .C(FIFO_CLK_c), .D(n6271));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1937_1938 (.Q(\REG.mem_19_25 ), .C(FIFO_CLK_c), .D(n6270));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1934_1935 (.Q(\REG.mem_19_24 ), .C(FIFO_CLK_c), .D(n6269));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1931_1932 (.Q(\REG.mem_19_23 ), .C(FIFO_CLK_c), .D(n6268));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1928_1929 (.Q(\REG.mem_19_22 ), .C(FIFO_CLK_c), .D(n6267));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1925_1926 (.Q(\REG.mem_19_21 ), .C(FIFO_CLK_c), .D(n6266));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1922_1923 (.Q(\REG.mem_19_20 ), .C(FIFO_CLK_c), .D(n6265));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1919_1920 (.Q(\REG.mem_19_19 ), .C(FIFO_CLK_c), .D(n6264));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1916_1917 (.Q(\REG.mem_19_18 ), .C(FIFO_CLK_c), .D(n6263));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1913_1914 (.Q(\REG.mem_19_17 ), .C(FIFO_CLK_c), .D(n6262));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1910_1911 (.Q(\REG.mem_19_16 ), .C(FIFO_CLK_c), .D(n6261));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1907_1908 (.Q(\REG.mem_19_15 ), .C(FIFO_CLK_c), .D(n6260));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1904_1905 (.Q(\REG.mem_19_14 ), .C(FIFO_CLK_c), .D(n6259));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1901_1902 (.Q(\REG.mem_19_13 ), .C(FIFO_CLK_c), .D(n6258));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1898_1899 (.Q(\REG.mem_19_12 ), .C(FIFO_CLK_c), .D(n6257));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1895_1896 (.Q(\REG.mem_19_11 ), .C(FIFO_CLK_c), .D(n6256));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1892_1893 (.Q(\REG.mem_19_10 ), .C(FIFO_CLK_c), .D(n6255));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1889_1890 (.Q(\REG.mem_19_9 ), .C(FIFO_CLK_c), .D(n6254));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1886_1887 (.Q(\REG.mem_19_8 ), .C(FIFO_CLK_c), .D(n6253));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1883_1884 (.Q(\REG.mem_19_7 ), .C(FIFO_CLK_c), .D(n6252));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1880_1881 (.Q(\REG.mem_19_6 ), .C(FIFO_CLK_c), .D(n6251));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1877_1878 (.Q(\REG.mem_19_5 ), .C(FIFO_CLK_c), .D(n6250));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1874_1875 (.Q(\REG.mem_19_4 ), .C(FIFO_CLK_c), .D(n6249));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1871_1872 (.Q(\REG.mem_19_3 ), .C(FIFO_CLK_c), .D(n6248));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1868_1869 (.Q(\REG.mem_19_2 ), .C(FIFO_CLK_c), .D(n6247));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1865_1866 (.Q(\REG.mem_19_1 ), .C(FIFO_CLK_c), .D(n6246));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1862_1863 (.Q(\REG.mem_19_0 ), .C(FIFO_CLK_c), .D(n6245));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1859_1860 (.Q(\REG.mem_18_31 ), .C(FIFO_CLK_c), .D(n6244));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1856_1857 (.Q(\REG.mem_18_30 ), .C(FIFO_CLK_c), .D(n6243));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1853_1854 (.Q(\REG.mem_18_29 ), .C(FIFO_CLK_c), .D(n6242));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1850_1851 (.Q(\REG.mem_18_28 ), .C(FIFO_CLK_c), .D(n6241));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1847_1848 (.Q(\REG.mem_18_27 ), .C(FIFO_CLK_c), .D(n6240));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1844_1845 (.Q(\REG.mem_18_26 ), .C(FIFO_CLK_c), .D(n6239));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1841_1842 (.Q(\REG.mem_18_25 ), .C(FIFO_CLK_c), .D(n6238));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1838_1839 (.Q(\REG.mem_18_24 ), .C(FIFO_CLK_c), .D(n6237));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1835_1836 (.Q(\REG.mem_18_23 ), .C(FIFO_CLK_c), .D(n6236));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1832_1833 (.Q(\REG.mem_18_22 ), .C(FIFO_CLK_c), .D(n6235));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1829_1830 (.Q(\REG.mem_18_21 ), .C(FIFO_CLK_c), .D(n6234));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1826_1827 (.Q(\REG.mem_18_20 ), .C(FIFO_CLK_c), .D(n6233));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1823_1824 (.Q(\REG.mem_18_19 ), .C(FIFO_CLK_c), .D(n6232));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1820_1821 (.Q(\REG.mem_18_18 ), .C(FIFO_CLK_c), .D(n6231));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1817_1818 (.Q(\REG.mem_18_17 ), .C(FIFO_CLK_c), .D(n6230));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1814_1815 (.Q(\REG.mem_18_16 ), .C(FIFO_CLK_c), .D(n6229));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1811_1812 (.Q(\REG.mem_18_15 ), .C(FIFO_CLK_c), .D(n6228));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1808_1809 (.Q(\REG.mem_18_14 ), .C(FIFO_CLK_c), .D(n6227));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1805_1806 (.Q(\REG.mem_18_13 ), .C(FIFO_CLK_c), .D(n6226));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1802_1803 (.Q(\REG.mem_18_12 ), .C(FIFO_CLK_c), .D(n6225));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1799_1800 (.Q(\REG.mem_18_11 ), .C(FIFO_CLK_c), .D(n6224));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1796_1797 (.Q(\REG.mem_18_10 ), .C(FIFO_CLK_c), .D(n6223));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1793_1794 (.Q(\REG.mem_18_9 ), .C(FIFO_CLK_c), .D(n6222));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1790_1791 (.Q(\REG.mem_18_8 ), .C(FIFO_CLK_c), .D(n6221));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1787_1788 (.Q(\REG.mem_18_7 ), .C(FIFO_CLK_c), .D(n6220));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1784_1785 (.Q(\REG.mem_18_6 ), .C(FIFO_CLK_c), .D(n6219));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1781_1782 (.Q(\REG.mem_18_5 ), .C(FIFO_CLK_c), .D(n6218));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1778_1779 (.Q(\REG.mem_18_4 ), .C(FIFO_CLK_c), .D(n6217));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1775_1776 (.Q(\REG.mem_18_3 ), .C(FIFO_CLK_c), .D(n6216));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1772_1773 (.Q(\REG.mem_18_2 ), .C(FIFO_CLK_c), .D(n6215));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1769_1770 (.Q(\REG.mem_18_1 ), .C(FIFO_CLK_c), .D(n6214));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1766_1767 (.Q(\REG.mem_18_0 ), .C(FIFO_CLK_c), .D(n6213));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1763_1764 (.Q(\REG.mem_17_31 ), .C(FIFO_CLK_c), .D(n6212));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1760_1761 (.Q(\REG.mem_17_30 ), .C(FIFO_CLK_c), .D(n6211));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1757_1758 (.Q(\REG.mem_17_29 ), .C(FIFO_CLK_c), .D(n6210));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1754_1755 (.Q(\REG.mem_17_28 ), .C(FIFO_CLK_c), .D(n6209));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1751_1752 (.Q(\REG.mem_17_27 ), .C(FIFO_CLK_c), .D(n6208));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1748_1749 (.Q(\REG.mem_17_26 ), .C(FIFO_CLK_c), .D(n6207));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1745_1746 (.Q(\REG.mem_17_25 ), .C(FIFO_CLK_c), .D(n6206));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1742_1743 (.Q(\REG.mem_17_24 ), .C(FIFO_CLK_c), .D(n6205));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1739_1740 (.Q(\REG.mem_17_23 ), .C(FIFO_CLK_c), .D(n6204));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1736_1737 (.Q(\REG.mem_17_22 ), .C(FIFO_CLK_c), .D(n6203));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1733_1734 (.Q(\REG.mem_17_21 ), .C(FIFO_CLK_c), .D(n6202));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1730_1731 (.Q(\REG.mem_17_20 ), .C(FIFO_CLK_c), .D(n6201));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1727_1728 (.Q(\REG.mem_17_19 ), .C(FIFO_CLK_c), .D(n6200));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1724_1725 (.Q(\REG.mem_17_18 ), .C(FIFO_CLK_c), .D(n6199));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1721_1722 (.Q(\REG.mem_17_17 ), .C(FIFO_CLK_c), .D(n6198));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1718_1719 (.Q(\REG.mem_17_16 ), .C(FIFO_CLK_c), .D(n6197));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1715_1716 (.Q(\REG.mem_17_15 ), .C(FIFO_CLK_c), .D(n6196));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1712_1713 (.Q(\REG.mem_17_14 ), .C(FIFO_CLK_c), .D(n6195));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1709_1710 (.Q(\REG.mem_17_13 ), .C(FIFO_CLK_c), .D(n6194));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1706_1707 (.Q(\REG.mem_17_12 ), .C(FIFO_CLK_c), .D(n6193));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1703_1704 (.Q(\REG.mem_17_11 ), .C(FIFO_CLK_c), .D(n6192));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1700_1701 (.Q(\REG.mem_17_10 ), .C(FIFO_CLK_c), .D(n6191));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1697_1698 (.Q(\REG.mem_17_9 ), .C(FIFO_CLK_c), .D(n6190));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1694_1695 (.Q(\REG.mem_17_8 ), .C(FIFO_CLK_c), .D(n6189));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1691_1692 (.Q(\REG.mem_17_7 ), .C(FIFO_CLK_c), .D(n6188));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1688_1689 (.Q(\REG.mem_17_6 ), .C(FIFO_CLK_c), .D(n6187));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1685_1686 (.Q(\REG.mem_17_5 ), .C(FIFO_CLK_c), .D(n6186));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1682_1683 (.Q(\REG.mem_17_4 ), .C(FIFO_CLK_c), .D(n6185));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1679_1680 (.Q(\REG.mem_17_3 ), .C(FIFO_CLK_c), .D(n6184));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1676_1677 (.Q(\REG.mem_17_2 ), .C(FIFO_CLK_c), .D(n6183));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1673_1674 (.Q(\REG.mem_17_1 ), .C(FIFO_CLK_c), .D(n6182));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1670_1671 (.Q(\REG.mem_17_0 ), .C(FIFO_CLK_c), .D(n6181));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1667_1668 (.Q(\REG.mem_16_31 ), .C(FIFO_CLK_c), .D(n6180));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1664_1665 (.Q(\REG.mem_16_30 ), .C(FIFO_CLK_c), .D(n6179));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1661_1662 (.Q(\REG.mem_16_29 ), .C(FIFO_CLK_c), .D(n6178));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1658_1659 (.Q(\REG.mem_16_28 ), .C(FIFO_CLK_c), .D(n6177));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1655_1656 (.Q(\REG.mem_16_27 ), .C(FIFO_CLK_c), .D(n6176));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1652_1653 (.Q(\REG.mem_16_26 ), .C(FIFO_CLK_c), .D(n6175));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1649_1650 (.Q(\REG.mem_16_25 ), .C(FIFO_CLK_c), .D(n6174));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1646_1647 (.Q(\REG.mem_16_24 ), .C(FIFO_CLK_c), .D(n6173));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1643_1644 (.Q(\REG.mem_16_23 ), .C(FIFO_CLK_c), .D(n6172));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1640_1641 (.Q(\REG.mem_16_22 ), .C(FIFO_CLK_c), .D(n6171));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1637_1638 (.Q(\REG.mem_16_21 ), .C(FIFO_CLK_c), .D(n6170));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1634_1635 (.Q(\REG.mem_16_20 ), .C(FIFO_CLK_c), .D(n6169));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1631_1632 (.Q(\REG.mem_16_19 ), .C(FIFO_CLK_c), .D(n6168));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1628_1629 (.Q(\REG.mem_16_18 ), .C(FIFO_CLK_c), .D(n6167));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1625_1626 (.Q(\REG.mem_16_17 ), .C(FIFO_CLK_c), .D(n6166));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1622_1623 (.Q(\REG.mem_16_16 ), .C(FIFO_CLK_c), .D(n6165));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1619_1620 (.Q(\REG.mem_16_15 ), .C(FIFO_CLK_c), .D(n6164));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1616_1617 (.Q(\REG.mem_16_14 ), .C(FIFO_CLK_c), .D(n6163));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1613_1614 (.Q(\REG.mem_16_13 ), .C(FIFO_CLK_c), .D(n6162));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1610_1611 (.Q(\REG.mem_16_12 ), .C(FIFO_CLK_c), .D(n6161));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1607_1608 (.Q(\REG.mem_16_11 ), .C(FIFO_CLK_c), .D(n6160));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1604_1605 (.Q(\REG.mem_16_10 ), .C(FIFO_CLK_c), .D(n6159));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1601_1602 (.Q(\REG.mem_16_9 ), .C(FIFO_CLK_c), .D(n6158));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1598_1599 (.Q(\REG.mem_16_8 ), .C(FIFO_CLK_c), .D(n6157));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1595_1596 (.Q(\REG.mem_16_7 ), .C(FIFO_CLK_c), .D(n6156));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1592_1593 (.Q(\REG.mem_16_6 ), .C(FIFO_CLK_c), .D(n6155));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1589_1590 (.Q(\REG.mem_16_5 ), .C(FIFO_CLK_c), .D(n6154));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1586_1587 (.Q(\REG.mem_16_4 ), .C(FIFO_CLK_c), .D(n6153));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1583_1584 (.Q(\REG.mem_16_3 ), .C(FIFO_CLK_c), .D(n6152));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1580_1581 (.Q(\REG.mem_16_2 ), .C(FIFO_CLK_c), .D(n6151));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1577_1578 (.Q(\REG.mem_16_1 ), .C(FIFO_CLK_c), .D(n6150));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1574_1575 (.Q(\REG.mem_16_0 ), .C(FIFO_CLK_c), .D(n6149));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1571_1572 (.Q(\REG.mem_15_31 ), .C(FIFO_CLK_c), .D(n6148));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1568_1569 (.Q(\REG.mem_15_30 ), .C(FIFO_CLK_c), .D(n6147));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1565_1566 (.Q(\REG.mem_15_29 ), .C(FIFO_CLK_c), .D(n6146));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1562_1563 (.Q(\REG.mem_15_28 ), .C(FIFO_CLK_c), .D(n6145));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1559_1560 (.Q(\REG.mem_15_27 ), .C(FIFO_CLK_c), .D(n6144));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1556_1557 (.Q(\REG.mem_15_26 ), .C(FIFO_CLK_c), .D(n6143));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1553_1554 (.Q(\REG.mem_15_25 ), .C(FIFO_CLK_c), .D(n6142));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n16983_bdd_4_lut (.I0(n16983), .I1(n15728), .I2(n15503), .I3(rd_addr_r[3]), 
            .O(n16986));
    defparam n16983_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5153_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_31_23 ), .O(n6652));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5153_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14214 (.I0(rd_addr_r[2]), .I1(n15239), 
            .I2(n15296), .I3(rd_addr_r[3]), .O(n16281));
    defparam rd_addr_r_2__bdd_4_lut_14214.LUT_INIT = 16'he4aa;
    SB_LUT4 i4598_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_14_12 ), .O(n6097));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4598_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5152_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_31_22 ), .O(n6651));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5152_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1550_1551 (.Q(\REG.mem_15_24 ), .C(FIFO_CLK_c), .D(n6141));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1547_1548 (.Q(\REG.mem_15_23 ), .C(FIFO_CLK_c), .D(n6140));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1544_1545 (.Q(\REG.mem_15_22 ), .C(FIFO_CLK_c), .D(n6139));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1541_1542 (.Q(\REG.mem_15_21 ), .C(FIFO_CLK_c), .D(n6138));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1538_1539 (.Q(\REG.mem_15_20 ), .C(FIFO_CLK_c), .D(n6137));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1535_1536 (.Q(\REG.mem_15_19 ), .C(FIFO_CLK_c), .D(n6136));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1532_1533 (.Q(\REG.mem_15_18 ), .C(FIFO_CLK_c), .D(n6135));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1529_1530 (.Q(\REG.mem_15_17 ), .C(FIFO_CLK_c), .D(n6134));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1526_1527 (.Q(\REG.mem_15_16 ), .C(FIFO_CLK_c), .D(n6133));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1523_1524 (.Q(\REG.mem_15_15 ), .C(FIFO_CLK_c), .D(n6132));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1520_1521 (.Q(\REG.mem_15_14 ), .C(FIFO_CLK_c), .D(n6131));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1517_1518 (.Q(\REG.mem_15_13 ), .C(FIFO_CLK_c), .D(n6130));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1514_1515 (.Q(\REG.mem_15_12 ), .C(FIFO_CLK_c), .D(n6129));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1511_1512 (.Q(\REG.mem_15_11 ), .C(FIFO_CLK_c), .D(n6128));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1508_1509 (.Q(\REG.mem_15_10 ), .C(FIFO_CLK_c), .D(n6127));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1505_1506 (.Q(\REG.mem_15_9 ), .C(FIFO_CLK_c), .D(n6126));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1502_1503 (.Q(\REG.mem_15_8 ), .C(FIFO_CLK_c), .D(n6125));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n16197_bdd_4_lut (.I0(n16197), .I1(\REG.mem_9_29 ), .I2(\REG.mem_8_29 ), 
            .I3(rd_addr_r[1]), .O(n16200));
    defparam n16197_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5151_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_31_21 ), .O(n6650));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5151_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5150_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_31_20 ), .O(n6649));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5150_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5149_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_31_19 ), .O(n6648));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5149_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15307 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_21 ), 
            .I2(\REG.mem_15_21 ), .I3(rd_addr_r[1]), .O(n17685));
    defparam rd_addr_r_0__bdd_4_lut_15307.LUT_INIT = 16'he4aa;
    SB_LUT4 n17685_bdd_4_lut (.I0(n17685), .I1(\REG.mem_13_21 ), .I2(\REG.mem_12_21 ), 
            .I3(rd_addr_r[1]), .O(n15134));
    defparam n17685_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13689_3_lut (.I0(\REG.mem_16_15 ), .I1(\REG.mem_17_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15813));
    defparam i13689_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1499_1500 (.Q(\REG.mem_15_7 ), .C(FIFO_CLK_c), .D(n6124));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1496_1497 (.Q(\REG.mem_15_6 ), .C(FIFO_CLK_c), .D(n6123));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i356_357 (.Q(\REG.mem_3_10 ), .C(FIFO_CLK_c), .D(n5743));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1493_1494 (.Q(\REG.mem_15_5 ), .C(FIFO_CLK_c), .D(n6122));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5148_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_31_18 ), .O(n6647));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5148_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5147_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_31_17 ), .O(n6646));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5147_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5146_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_31_16 ), .O(n6645));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5146_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i46_2_lut_3_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n12));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i46_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15332 (.I0(rd_addr_r[1]), .I1(n15006), 
            .I2(n15007), .I3(rd_addr_r[2]), .O(n17679));
    defparam rd_addr_r_1__bdd_4_lut_15332.LUT_INIT = 16'he4aa;
    SB_LUT4 i4597_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_14_11 ), .O(n6096));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4597_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1490_1491 (.Q(\REG.mem_15_4 ), .C(FIFO_CLK_c), .D(n6121));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1487_1488 (.Q(\REG.mem_15_3 ), .C(FIFO_CLK_c), .D(n6120));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1484_1485 (.Q(\REG.mem_15_2 ), .C(FIFO_CLK_c), .D(n6119));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1481_1482 (.Q(\REG.mem_15_1 ), .C(FIFO_CLK_c), .D(n6118));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1478_1479 (.Q(\REG.mem_15_0 ), .C(FIFO_CLK_c), .D(n6117));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1475_1476 (.Q(\REG.mem_14_31 ), .C(FIFO_CLK_c), .D(n6116));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1472_1473 (.Q(\REG.mem_14_30 ), .C(FIFO_CLK_c), .D(n6115));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1469_1470 (.Q(\REG.mem_14_29 ), .C(FIFO_CLK_c), .D(n6114));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i353_354 (.Q(\REG.mem_3_9 ), .C(FIFO_CLK_c), .D(n5742));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1466_1467 (.Q(\REG.mem_14_28 ), .C(FIFO_CLK_c), .D(n6113));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5145_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_31_15 ), .O(n6644));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5145_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5144_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_31_14 ), .O(n6643));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5144_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16281_bdd_4_lut (.I0(n16281), .I1(n15440), .I2(n15119), .I3(rd_addr_r[3]), 
            .O(n16284));
    defparam n16281_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5143_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_31_13 ), .O(n6642));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5143_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5142_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_31_12 ), .O(n6641));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5142_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5141_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_31_11 ), .O(n6640));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5141_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5140_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_31_10 ), .O(n6639));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5140_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4596_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_14_10 ), .O(n6095));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4596_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5139_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_31_9 ), .O(n6638));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5139_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4595_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_14_9 ), .O(n6094));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4595_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5138_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_31_8 ), .O(n6637));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5138_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5137_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_31_7 ), .O(n6636));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5137_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4594_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_14_8 ), .O(n6093));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4594_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4593_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_14_7 ), .O(n6092));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4593_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17679_bdd_4_lut (.I0(n17679), .I1(n15004), .I2(n15003), .I3(rd_addr_r[2]), 
            .O(n15139));
    defparam n17679_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1463_1464 (.Q(\REG.mem_14_27 ), .C(FIFO_CLK_c), .D(n6112));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5136_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_31_6 ), .O(n6635));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5136_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14723 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_15 ), 
            .I2(\REG.mem_27_15 ), .I3(rd_addr_r[1]), .O(n16971));
    defparam rd_addr_r_0__bdd_4_lut_14723.LUT_INIT = 16'he4aa;
    SB_DFF i1460_1461 (.Q(\REG.mem_14_26 ), .C(FIFO_CLK_c), .D(n6111));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5135_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_31_5 ), .O(n6634));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5135_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1457_1458 (.Q(\REG.mem_14_25 ), .C(FIFO_CLK_c), .D(n6110));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1454_1455 (.Q(\REG.mem_14_24 ), .C(FIFO_CLK_c), .D(n6109));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1451_1452 (.Q(\REG.mem_14_23 ), .C(FIFO_CLK_c), .D(n6108));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1448_1449 (.Q(\REG.mem_14_22 ), .C(FIFO_CLK_c), .D(n6107));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1445_1446 (.Q(\REG.mem_14_21 ), .C(FIFO_CLK_c), .D(n6106));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1442_1443 (.Q(\REG.mem_14_20 ), .C(FIFO_CLK_c), .D(n6105));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5134_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_31_4 ), .O(n6633));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5134_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5133_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_31_3 ), .O(n6632));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5133_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15302 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_23 ), 
            .I2(\REG.mem_3_23 ), .I3(rd_addr_r[1]), .O(n17673));
    defparam rd_addr_r_0__bdd_4_lut_15302.LUT_INIT = 16'he4aa;
    SB_LUT4 n17673_bdd_4_lut (.I0(n17673), .I1(\REG.mem_1_23 ), .I2(\REG.mem_0_23 ), 
            .I3(rd_addr_r[1]), .O(n15608));
    defparam n17673_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16971_bdd_4_lut (.I0(n16971), .I1(\REG.mem_25_15 ), .I2(\REG.mem_24_15 ), 
            .I3(rd_addr_r[1]), .O(n16974));
    defparam n16971_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4592_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_14_6 ), .O(n6091));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4592_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5132_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_31_2 ), .O(n6631));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5132_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4591_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_14_5 ), .O(n6090));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4591_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5131_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_31_1 ), .O(n6630));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5131_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1439_1440 (.Q(\REG.mem_14_19 ), .C(FIFO_CLK_c), .D(n6104));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14708 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_21 ), 
            .I2(\REG.mem_27_21 ), .I3(rd_addr_r[1]), .O(n16965));
    defparam rd_addr_r_0__bdd_4_lut_14708.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14139 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_17 ), 
            .I2(\REG.mem_27_17 ), .I3(rd_addr_r[1]), .O(n16275));
    defparam rd_addr_r_0__bdd_4_lut_14139.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15292 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_27 ), 
            .I2(\REG.mem_19_27 ), .I3(rd_addr_r[1]), .O(n17667));
    defparam rd_addr_r_0__bdd_4_lut_15292.LUT_INIT = 16'he4aa;
    SB_LUT4 n16275_bdd_4_lut (.I0(n16275), .I1(\REG.mem_25_17 ), .I2(\REG.mem_24_17 ), 
            .I3(rd_addr_r[1]), .O(n16278));
    defparam n16275_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5130_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_31_0 ), .O(n6629));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5130_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14134 (.I0(rd_addr_r[2]), .I1(n15314), 
            .I2(n15326), .I3(rd_addr_r[3]), .O(n16269));
    defparam rd_addr_r_2__bdd_4_lut_14134.LUT_INIT = 16'he4aa;
    SB_DFF i1436_1437 (.Q(\REG.mem_14_18 ), .C(FIFO_CLK_c), .D(n6103));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1433_1434 (.Q(\REG.mem_14_17 ), .C(FIFO_CLK_c), .D(n6102));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i50_2_lut_3_lut_4_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n10));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i50_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_DFF i1430_1431 (.Q(\REG.mem_14_16 ), .C(FIFO_CLK_c), .D(n6101));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1427_1428 (.Q(\REG.mem_14_15 ), .C(FIFO_CLK_c), .D(n6100));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1424_1425 (.Q(\REG.mem_14_14 ), .C(FIFO_CLK_c), .D(n6099));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1421_1422 (.Q(\REG.mem_14_13 ), .C(FIFO_CLK_c), .D(n6098));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1418_1419 (.Q(\REG.mem_14_12 ), .C(FIFO_CLK_c), .D(n6097));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1415_1416 (.Q(\REG.mem_14_11 ), .C(FIFO_CLK_c), .D(n6096));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i51_2_lut_3_lut_4_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n26));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i51_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_DFF i1412_1413 (.Q(\REG.mem_14_10 ), .C(FIFO_CLK_c), .D(n6095));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i350_351 (.Q(\REG.mem_3_8 ), .C(FIFO_CLK_c), .D(n5741));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4590_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_14_4 ), .O(n6089));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4590_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4589_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_14_3 ), .O(n6088));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4589_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4588_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_14_2 ), .O(n6087));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4588_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4587_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_14_1 ), .O(n6086));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4587_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17667_bdd_4_lut (.I0(n17667), .I1(\REG.mem_17_27 ), .I2(\REG.mem_16_27 ), 
            .I3(rd_addr_r[1]), .O(n15146));
    defparam n17667_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4586_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_14_0 ), .O(n6085));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4586_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i5_2_lut_4_lut (.I0(rd_grey_sync_r[5]), 
            .I1(rd_addr_p1_w[5]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_5__N_573[4] ), 
            .O(rd_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i5525_2_lut_4_lut (.I0(rd_grey_sync_r[5]), .I1(rd_addr_p1_w[5]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n7024));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i5525_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_DFF i1409_1410 (.Q(\REG.mem_14_9 ), .C(FIFO_CLK_c), .D(n6094));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4937_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_24_31 ), .O(n6436));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4937_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1406_1407 (.Q(\REG.mem_14_8 ), .C(FIFO_CLK_c), .D(n6093));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n16965_bdd_4_lut (.I0(n16965), .I1(\REG.mem_25_21 ), .I2(\REG.mem_24_21 ), 
            .I3(rd_addr_r[1]), .O(n15266));
    defparam n16965_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4936_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_24_30 ), .O(n6435));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4936_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1403_1404 (.Q(\REG.mem_14_7 ), .C(FIFO_CLK_c), .D(n6092));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1400_1401 (.Q(\REG.mem_14_6 ), .C(FIFO_CLK_c), .D(n6091));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1397_1398 (.Q(\REG.mem_14_5 ), .C(FIFO_CLK_c), .D(n6090));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4935_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_24_29 ), .O(n6434));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4935_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4745_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_18_31 ), .O(n6244));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4745_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4744_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_18_30 ), .O(n6243));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4744_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4743_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_18_29 ), .O(n6242));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4743_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4934_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_24_28 ), .O(n6433));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4934_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4933_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_24_27 ), .O(n6432));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4933_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4742_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_18_28 ), .O(n6241));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4742_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4741_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_18_27 ), .O(n6240));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4741_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4740_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_18_26 ), .O(n6239));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4740_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4739_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_18_25 ), .O(n6238));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4739_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4738_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_18_24 ), .O(n6237));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4738_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1394_1395 (.Q(\REG.mem_14_4 ), .C(FIFO_CLK_c), .D(n6089));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4737_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_18_23 ), .O(n6236));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4737_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4932_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_24_26 ), .O(n6431));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4932_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4736_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_18_22 ), .O(n6235));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4736_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4735_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_18_21 ), .O(n6234));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4735_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4734_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_18_20 ), .O(n6233));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4734_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4931_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_24_25 ), .O(n6430));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4931_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4930_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_24_24 ), .O(n6429));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4930_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4733_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_18_19 ), .O(n6232));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4733_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1391_1392 (.Q(\REG.mem_14_3 ), .C(FIFO_CLK_c), .D(n6088));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1388_1389 (.Q(\REG.mem_14_2 ), .C(FIFO_CLK_c), .D(n6087));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1385_1386 (.Q(\REG.mem_14_1 ), .C(FIFO_CLK_c), .D(n6086));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14703 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_22 ), 
            .I2(\REG.mem_7_22 ), .I3(rd_addr_r[1]), .O(n16959));
    defparam rd_addr_r_0__bdd_4_lut_14703.LUT_INIT = 16'he4aa;
    SB_LUT4 n16269_bdd_4_lut (.I0(n16269), .I1(n15428), .I2(n15260), .I3(rd_addr_r[3]), 
            .O(n16272));
    defparam n16269_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4929_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_24_23 ), .O(n6428));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4929_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13690_3_lut (.I0(\REG.mem_18_15 ), .I1(\REG.mem_19_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15814));
    defparam i13690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4732_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_18_18 ), .O(n6231));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4732_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4731_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_18_17 ), .O(n6230));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4731_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1382_1383 (.Q(\REG.mem_14_0 ), .C(FIFO_CLK_c), .D(n6085));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15287 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_23 ), 
            .I2(\REG.mem_7_23 ), .I3(rd_addr_r[1]), .O(n17661));
    defparam rd_addr_r_0__bdd_4_lut_15287.LUT_INIT = 16'he4aa;
    SB_LUT4 i4730_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_18_16 ), .O(n6229));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4730_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17661_bdd_4_lut (.I0(n17661), .I1(\REG.mem_5_23 ), .I2(\REG.mem_4_23 ), 
            .I3(rd_addr_r[1]), .O(n15614));
    defparam n17661_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14129 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_30 ), 
            .I2(\REG.mem_27_30 ), .I3(rd_addr_r[1]), .O(n16263));
    defparam rd_addr_r_0__bdd_4_lut_14129.LUT_INIT = 16'he4aa;
    SB_LUT4 i4729_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_18_15 ), .O(n6228));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4729_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4728_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_18_14 ), .O(n6227));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4728_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4928_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_24_22 ), .O(n6427));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4928_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4727_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_18_13 ), .O(n6226));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4727_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12819_3_lut (.I0(\REG.mem_16_24 ), .I1(\REG.mem_17_24 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14943));
    defparam i12819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4726_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_18_12 ), .O(n6225));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4726_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1379_1380 (.Q(\REG.mem_13_31 ), .C(FIFO_CLK_c), .D(n6084));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1376_1377 (.Q(\REG.mem_13_30 ), .C(FIFO_CLK_c), .D(n6083));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4725_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_18_11 ), .O(n6224));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4725_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1373_1374 (.Q(\REG.mem_13_29 ), .C(FIFO_CLK_c), .D(n6082));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4724_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_18_10 ), .O(n6223));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4724_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1370_1371 (.Q(\REG.mem_13_28 ), .C(FIFO_CLK_c), .D(n6081));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4723_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_18_9 ), .O(n6222));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4723_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16959_bdd_4_lut (.I0(n16959), .I1(\REG.mem_5_22 ), .I2(\REG.mem_4_22 ), 
            .I3(rd_addr_r[1]), .O(n16962));
    defparam n16959_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4722_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_18_8 ), .O(n6221));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4722_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12820_3_lut (.I0(\REG.mem_18_24 ), .I1(\REG.mem_19_24 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14944));
    defparam i12820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4721_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_18_7 ), .O(n6220));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4721_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12826_3_lut (.I0(\REG.mem_22_24 ), .I1(\REG.mem_23_24 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14950));
    defparam i12826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15282 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_23 ), 
            .I2(\REG.mem_11_23 ), .I3(rd_addr_r[1]), .O(n17655));
    defparam rd_addr_r_0__bdd_4_lut_15282.LUT_INIT = 16'he4aa;
    SB_LUT4 i4720_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_18_6 ), .O(n6219));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4720_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4719_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_18_5 ), .O(n6218));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4719_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1367_1368 (.Q(\REG.mem_13_27 ), .C(FIFO_CLK_c), .D(n6080));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1364_1365 (.Q(\REG.mem_13_26 ), .C(FIFO_CLK_c), .D(n6079));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i12825_3_lut (.I0(\REG.mem_20_24 ), .I1(\REG.mem_21_24 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14949));
    defparam i12825_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1361_1362 (.Q(\REG.mem_13_25 ), .C(FIFO_CLK_c), .D(n6078));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i347_348 (.Q(\REG.mem_3_7 ), .C(FIFO_CLK_c), .D(n5740));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4718_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_18_4 ), .O(n6217));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4718_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4927_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_24_21 ), .O(n6426));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4927_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1358_1359 (.Q(\REG.mem_13_24 ), .C(FIFO_CLK_c), .D(n6077));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4717_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_18_3 ), .O(n6216));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4717_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17655_bdd_4_lut (.I0(n17655), .I1(\REG.mem_9_23 ), .I2(\REG.mem_8_23 ), 
            .I3(rd_addr_r[1]), .O(n15617));
    defparam n17655_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4716_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_18_2 ), .O(n6215));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4716_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1355_1356 (.Q(\REG.mem_13_23 ), .C(FIFO_CLK_c), .D(n6076));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1352_1353 (.Q(\REG.mem_13_22 ), .C(FIFO_CLK_c), .D(n6075));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15277 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_20 ), 
            .I2(\REG.mem_19_20 ), .I3(rd_addr_r[1]), .O(n17649));
    defparam rd_addr_r_0__bdd_4_lut_15277.LUT_INIT = 16'he4aa;
    SB_DFF i1349_1350 (.Q(\REG.mem_13_21 ), .C(FIFO_CLK_c), .D(n6074));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n17649_bdd_4_lut (.I0(n17649), .I1(\REG.mem_17_20 ), .I2(\REG.mem_16_20 ), 
            .I3(rd_addr_r[1]), .O(n15149));
    defparam n17649_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16263_bdd_4_lut (.I0(n16263), .I1(\REG.mem_25_30 ), .I2(\REG.mem_24_30 ), 
            .I3(rd_addr_r[1]), .O(n16266));
    defparam n16263_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i344_345 (.Q(\REG.mem_3_6 ), .C(FIFO_CLK_c), .D(n5739));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4926_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_24_20 ), .O(n6425));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4926_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1346_1347 (.Q(\REG.mem_13_20 ), .C(FIFO_CLK_c), .D(n6073));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4715_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_18_1 ), .O(n6214));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4715_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1343_1344 (.Q(\REG.mem_13_19 ), .C(FIFO_CLK_c), .D(n6072));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4714_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_18_0 ), .O(n6213));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4714_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1340_1341 (.Q(\REG.mem_13_18 ), .C(FIFO_CLK_c), .D(n6071));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15297 (.I0(rd_addr_r[1]), .I1(n15570), 
            .I2(n15571), .I3(rd_addr_r[2]), .O(n17643));
    defparam rd_addr_r_1__bdd_4_lut_15297.LUT_INIT = 16'he4aa;
    SB_LUT4 i4925_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_24_19 ), .O(n6424));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4925_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4924_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_24_18 ), .O(n6423));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4924_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14698 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_1 ), 
            .I2(\REG.mem_27_1 ), .I3(rd_addr_r[1]), .O(n16953));
    defparam rd_addr_r_0__bdd_4_lut_14698.LUT_INIT = 16'he4aa;
    SB_DFF i341_342 (.Q(\REG.mem_3_5 ), .C(FIFO_CLK_c), .D(n5738));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5129_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_30_31 ), .O(n6628));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5129_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4923_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_24_17 ), .O(n6422));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4923_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5128_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_30_30 ), .O(n6627));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5128_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5127_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_30_29 ), .O(n6626));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5127_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5126_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_30_28 ), .O(n6625));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5126_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17643_bdd_4_lut (.I0(n17643), .I1(n15499), .I2(n15498), .I3(rd_addr_r[2]), 
            .O(n15885));
    defparam n17643_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16953_bdd_4_lut (.I0(n16953), .I1(\REG.mem_25_1 ), .I2(\REG.mem_24_1 ), 
            .I3(rd_addr_r[1]), .O(n15833));
    defparam n16953_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i338_339 (.Q(\REG.mem_3_4 ), .C(FIFO_CLK_c), .D(n5737));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5125_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_30_27 ), .O(n6624));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5125_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1337_1338 (.Q(\REG.mem_13_17 ), .C(FIFO_CLK_c), .D(n6070));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5124_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_30_26 ), .O(n6623));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5124_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5123_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_30_25 ), .O(n6622));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5123_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i335_336 (.Q(\REG.mem_3_3 ), .C(FIFO_CLK_c), .D(n5736));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i13699_3_lut (.I0(\REG.mem_22_15 ), .I1(\REG.mem_23_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15823));
    defparam i13699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5122_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_30_24 ), .O(n6621));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5122_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15272 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_18 ), 
            .I2(\REG.mem_11_18 ), .I3(rd_addr_r[1]), .O(n17631));
    defparam rd_addr_r_0__bdd_4_lut_15272.LUT_INIT = 16'he4aa;
    SB_LUT4 i4922_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_24_16 ), .O(n6421));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4922_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5121_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_30_23 ), .O(n6620));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5121_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13698_3_lut (.I0(\REG.mem_20_15 ), .I1(\REG.mem_21_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15822));
    defparam i13698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17631_bdd_4_lut (.I0(n17631), .I1(\REG.mem_9_18 ), .I2(\REG.mem_8_18 ), 
            .I3(rd_addr_r[1]), .O(n15623));
    defparam n17631_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5120_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_30_22 ), .O(n6619));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5120_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5119_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_30_21 ), .O(n6618));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5119_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5118_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_30_20 ), .O(n6617));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5118_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1334_1335 (.Q(\REG.mem_13_16 ), .C(FIFO_CLK_c), .D(n6069));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1331_1332 (.Q(\REG.mem_13_15 ), .C(FIFO_CLK_c), .D(n6068));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5117_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_30_19 ), .O(n6616));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5117_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15257 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_7 ), 
            .I2(\REG.mem_7_7 ), .I3(rd_addr_r[1]), .O(n17625));
    defparam rd_addr_r_0__bdd_4_lut_15257.LUT_INIT = 16'he4aa;
    SB_LUT4 i5116_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_30_18 ), .O(n6615));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5116_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1328_1329 (.Q(\REG.mem_13_14 ), .C(FIFO_CLK_c), .D(n6067));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14718 (.I0(rd_addr_r[2]), .I1(n15623), 
            .I2(n15650), .I3(rd_addr_r[3]), .O(n16947));
    defparam rd_addr_r_2__bdd_4_lut_14718.LUT_INIT = 16'he4aa;
    SB_DFF i1325_1326 (.Q(\REG.mem_13_13 ), .C(FIFO_CLK_c), .D(n6066));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i12879_3_lut (.I0(\REG.mem_24_13 ), .I1(\REG.mem_25_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15003));
    defparam i12879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5115_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_30_17 ), .O(n6614));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5115_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5114_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_30_16 ), .O(n6613));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5114_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17625_bdd_4_lut (.I0(n17625), .I1(\REG.mem_5_7 ), .I2(\REG.mem_4_7 ), 
            .I3(rd_addr_r[1]), .O(n17628));
    defparam n17625_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12880_3_lut (.I0(\REG.mem_26_13 ), .I1(\REG.mem_27_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15004));
    defparam i12880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13728_3_lut (.I0(\REG.mem_16_22 ), .I1(\REG.mem_17_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15852));
    defparam i13728_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1322_1323 (.Q(\REG.mem_13_12 ), .C(FIFO_CLK_c), .D(n6065));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1319_1320 (.Q(\REG.mem_13_11 ), .C(FIFO_CLK_c), .D(n6064));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i13729_3_lut (.I0(\REG.mem_18_22 ), .I1(\REG.mem_19_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15853));
    defparam i13729_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1316_1317 (.Q(\REG.mem_13_10 ), .C(FIFO_CLK_c), .D(n6063));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4921_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_24_15 ), .O(n6420));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4921_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5113_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_30_15 ), .O(n6612));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5113_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5112_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_30_14 ), .O(n6611));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5112_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5111_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_30_13 ), .O(n6610));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5111_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5110_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_30_12 ), .O(n6609));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5110_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4920_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_24_14 ), .O(n6419));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4920_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5109_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_30_11 ), .O(n6608));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5109_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15252 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_23 ), 
            .I2(\REG.mem_15_23 ), .I3(rd_addr_r[1]), .O(n17619));
    defparam rd_addr_r_0__bdd_4_lut_15252.LUT_INIT = 16'he4aa;
    SB_LUT4 i5108_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_30_10 ), .O(n6607));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5108_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5107_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_30_9 ), .O(n6606));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5107_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17619_bdd_4_lut (.I0(n17619), .I1(\REG.mem_13_23 ), .I2(\REG.mem_12_23 ), 
            .I3(rd_addr_r[1]), .O(n15626));
    defparam n17619_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5106_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_30_8 ), .O(n6605));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5106_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16947_bdd_4_lut (.I0(n16947), .I1(n16428), .I2(n15569), .I3(rd_addr_r[3]), 
            .O(n16950));
    defparam n16947_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4919_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_24_13 ), .O(n6418));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4919_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4918_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_24_12 ), .O(n6417));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4918_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1313_1314 (.Q(\REG.mem_13_9 ), .C(FIFO_CLK_c), .D(n6062));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5105_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_30_7 ), .O(n6604));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5105_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1310_1311 (.Q(\REG.mem_13_8 ), .C(FIFO_CLK_c), .D(n6061));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1307_1308 (.Q(\REG.mem_13_7 ), .C(FIFO_CLK_c), .D(n6060));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5104_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_30_6 ), .O(n6603));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5104_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14693 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_15 ), 
            .I2(\REG.mem_31_15 ), .I3(rd_addr_r[1]), .O(n16941));
    defparam rd_addr_r_0__bdd_4_lut_14693.LUT_INIT = 16'he4aa;
    SB_LUT4 i5103_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_30_5 ), .O(n6602));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5103_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1304_1305 (.Q(\REG.mem_13_6 ), .C(FIFO_CLK_c), .D(n6059));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15247 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_9 ), 
            .I2(\REG.mem_11_9 ), .I3(rd_addr_r[1]), .O(n17613));
    defparam rd_addr_r_0__bdd_4_lut_15247.LUT_INIT = 16'he4aa;
    SB_LUT4 n16941_bdd_4_lut (.I0(n16941), .I1(\REG.mem_29_15 ), .I2(\REG.mem_28_15 ), 
            .I3(rd_addr_r[1]), .O(n16944));
    defparam n16941_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5102_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_30_4 ), .O(n6601));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5102_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5101_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_30_3 ), .O(n6600));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5101_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17613_bdd_4_lut (.I0(n17613), .I1(\REG.mem_9_9 ), .I2(\REG.mem_8_9 ), 
            .I3(rd_addr_r[1]), .O(n14789));
    defparam n17613_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5100_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_30_2 ), .O(n6599));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5100_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5099_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_30_1 ), .O(n6598));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5099_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5098_3_lut_4_lut (.I0(n32), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_30_0 ), .O(n6597));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5098_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15267 (.I0(rd_addr_r[1]), .I1(n14718), 
            .I2(n14719), .I3(rd_addr_r[2]), .O(n17607));
    defparam rd_addr_r_1__bdd_4_lut_15267.LUT_INIT = 16'he4aa;
    SB_LUT4 n17607_bdd_4_lut (.I0(n17607), .I1(n14740), .I2(n14739), .I3(rd_addr_r[2]), 
            .O(n15660));
    defparam n17607_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14683 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_19 ), 
            .I2(\REG.mem_31_19 ), .I3(rd_addr_r[1]), .O(n16935));
    defparam rd_addr_r_0__bdd_4_lut_14683.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15242 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_19 ), 
            .I2(\REG.mem_19_19 ), .I3(rd_addr_r[1]), .O(n17601));
    defparam rd_addr_r_0__bdd_4_lut_15242.LUT_INIT = 16'he4aa;
    SB_LUT4 n16935_bdd_4_lut (.I0(n16935), .I1(\REG.mem_29_19 ), .I2(\REG.mem_28_19 ), 
            .I3(rd_addr_r[1]), .O(n16938));
    defparam n16935_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17601_bdd_4_lut (.I0(n17601), .I1(\REG.mem_17_19 ), .I2(\REG.mem_16_19 ), 
            .I3(rd_addr_r[1]), .O(n17604));
    defparam n17601_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14688 (.I0(rd_addr_r[2]), .I1(n15176), 
            .I2(n15200), .I3(rd_addr_r[3]), .O(n16929));
    defparam rd_addr_r_2__bdd_4_lut_14688.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i24_2_lut_3_lut_4_lut (.I0(n7_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n24));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i24_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_6_lut (.I0(n46), .I1(wp_sync_w[4]), 
            .I2(n1[4]), .I3(n13665), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_6_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 EnabledDecoder_2_i25_2_lut_3_lut_4_lut (.I0(n7_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n25_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i25_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15232 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_9 ), 
            .I2(\REG.mem_15_9 ), .I3(rd_addr_r[1]), .O(n17595));
    defparam rd_addr_r_0__bdd_4_lut_15232.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_5__I_0_i4_3_lut (.I0(rd_addr_r[3]), .I1(rd_addr_p1_w[3]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_5__N_573[3] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_5__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4142_2_lut_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_p1_w[0]), 
            .I2(rd_fifo_en_w), .I3(reset_per_frame), .O(n5641));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4142_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i1_2_lut_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_p1_w[0]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_5__N_573[1] ), .O(rd_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_5__I_0_138_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n16929_bdd_4_lut (.I0(n16929), .I1(n15122), .I2(n15098), .I3(rd_addr_r[3]), 
            .O(n16932));
    defparam n16929_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_5__I_0_i5_3_lut (.I0(rd_addr_r[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_5__N_573[4] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_5__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14678 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_1 ), 
            .I2(\REG.mem_31_1 ), .I3(rd_addr_r[1]), .O(n16923));
    defparam rd_addr_r_0__bdd_4_lut_14678.LUT_INIT = 16'he4aa;
    SB_LUT4 n16923_bdd_4_lut (.I0(n16923), .I1(\REG.mem_29_1 ), .I2(\REG.mem_28_1 ), 
            .I3(rd_addr_r[1]), .O(n15842));
    defparam n16923_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17595_bdd_4_lut (.I0(n17595), .I1(\REG.mem_13_9 ), .I2(\REG.mem_12_9 ), 
            .I3(rd_addr_r[1]), .O(n14798));
    defparam n17595_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i2_2_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(wr_fifo_en_w), .I3(\wr_addr_nxt_c[2] ), .O(wr_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_5__I_0_136_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14748 (.I0(rd_addr_r[1]), .I1(n14790), 
            .I2(n14791), .I3(rd_addr_r[2]), .O(n16917));
    defparam rd_addr_r_1__bdd_4_lut_14748.LUT_INIT = 16'he4aa;
    SB_DFF i1301_1302 (.Q(\REG.mem_13_5 ), .C(FIFO_CLK_c), .D(n6058));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5457_2_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(wr_fifo_en_w), .I3(reset_per_frame), .O(n6956));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i5457_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i1_2_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(wr_fifo_en_w), .I3(wr_addr_nxt_c[0]), .O(wr_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_5__I_0_136_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_15482 (.I0(rd_addr_r[2]), .I1(n15536), 
            .I2(n16368), .I3(rd_addr_r[3]), .O(n17589));
    defparam rd_addr_r_2__bdd_4_lut_15482.LUT_INIT = 16'he4aa;
    SB_LUT4 i5097_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_29_31 ), .O(n6596));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5097_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17589_bdd_4_lut (.I0(n17589), .I1(n15527), .I2(n16290), .I3(rd_addr_r[3]), 
            .O(n17592));
    defparam n17589_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16917_bdd_4_lut (.I0(n16917), .I1(n14785), .I2(n14784), .I3(rd_addr_r[2]), 
            .O(n14821));
    defparam n16917_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5096_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_29_30 ), .O(n6595));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5096_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4917_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_24_11 ), .O(n6416));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4917_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_6 (.CI(n13665), .I0(wp_sync_w[4]), 
            .I1(n1[4]), .CO(n13666));
    SB_LUT4 i5095_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_29_29 ), .O(n6594));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5095_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5094_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_29_28 ), .O(n6593));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5094_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14673 (.I0(rd_addr_r[2]), .I1(n15680), 
            .I2(n15692), .I3(rd_addr_r[3]), .O(n16911));
    defparam rd_addr_r_2__bdd_4_lut_14673.LUT_INIT = 16'he4aa;
    SB_LUT4 n16911_bdd_4_lut (.I0(n16911), .I1(n16596), .I2(n15665), .I3(rd_addr_r[3]), 
            .O(n16914));
    defparam n16911_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_5_lut (.I0(GND_net), .I1(wp_sync_w[3]), 
            .I2(n1[3]), .I3(n13664), .O(rd_sig_diff0_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5093_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_29_27 ), .O(n6592));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5093_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut (.I0(rd_addr_r[3]), .I1(n17400), .I2(n15520), 
            .I3(rd_addr_r[4]), .O(n17583));
    defparam rd_addr_r_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i12883_3_lut (.I0(\REG.mem_30_13 ), .I1(\REG.mem_31_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15007));
    defparam i12883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17583_bdd_4_lut (.I0(n17583), .I1(n15592), .I2(n17556), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[25]));
    defparam n17583_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12882_3_lut (.I0(\REG.mem_28_13 ), .I1(\REG.mem_29_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15006));
    defparam i12882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5092_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_29_26 ), .O(n6591));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5092_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5091_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_29_25 ), .O(n6590));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5091_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5090_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_29_24 ), .O(n6589));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5090_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5089_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_29_23 ), .O(n6588));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5089_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5088_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_29_22 ), .O(n6587));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5088_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5087_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_29_21 ), .O(n6586));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5087_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14658 (.I0(rd_addr_r[2]), .I1(n15800), 
            .I2(n15809), .I3(rd_addr_r[3]), .O(n16905));
    defparam rd_addr_r_2__bdd_4_lut_14658.LUT_INIT = 16'he4aa;
    SB_LUT4 i5086_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_29_20 ), .O(n6585));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5086_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16905_bdd_4_lut (.I0(n16905), .I1(n15794), .I2(n15254), .I3(rd_addr_r[3]), 
            .O(n16908));
    defparam n16905_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5085_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_29_19 ), .O(n6584));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5085_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14668 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_20 ), 
            .I2(\REG.mem_31_20 ), .I3(rd_addr_r[1]), .O(n16899));
    defparam rd_addr_r_0__bdd_4_lut_14668.LUT_INIT = 16'he4aa;
    SB_LUT4 n16899_bdd_4_lut (.I0(n16899), .I1(\REG.mem_29_20 ), .I2(\REG.mem_28_20 ), 
            .I3(rd_addr_r[1]), .O(n15278));
    defparam n16899_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4916_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_24_10 ), .O(n6415));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4916_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15227 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_20 ), 
            .I2(\REG.mem_23_20 ), .I3(rd_addr_r[1]), .O(n17571));
    defparam rd_addr_r_0__bdd_4_lut_15227.LUT_INIT = 16'he4aa;
    SB_LUT4 i5084_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_29_18 ), .O(n6583));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5084_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5083_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_29_17 ), .O(n6582));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5083_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5082_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_29_16 ), .O(n6581));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5082_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5081_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_29_15 ), .O(n6580));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5081_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5080_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_29_14 ), .O(n6579));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5080_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5079_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_29_13 ), .O(n6578));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5079_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17571_bdd_4_lut (.I0(n17571), .I1(\REG.mem_21_20 ), .I2(\REG.mem_20_20 ), 
            .I3(rd_addr_r[1]), .O(n15164));
    defparam n17571_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5078_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_29_12 ), .O(n6577));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5078_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5077_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_29_11 ), .O(n6576));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5077_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1298_1299 (.Q(\REG.mem_13_4 ), .C(FIFO_CLK_c), .D(n6057));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15207 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_23 ), 
            .I2(\REG.mem_19_23 ), .I3(rd_addr_r[1]), .O(n17565));
    defparam rd_addr_r_0__bdd_4_lut_15207.LUT_INIT = 16'he4aa;
    SB_LUT4 i4915_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_24_9 ), .O(n6414));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4915_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17565_bdd_4_lut (.I0(n17565), .I1(\REG.mem_17_23 ), .I2(\REG.mem_16_23 ), 
            .I3(rd_addr_r[1]), .O(n15635));
    defparam n17565_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4914_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_24_8 ), .O(n6413));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4914_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5076_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_29_10 ), .O(n6575));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5076_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5075_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_29_9 ), .O(n6574));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5075_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14648 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_27 ), 
            .I2(\REG.mem_23_27 ), .I3(rd_addr_r[1]), .O(n16893));
    defparam rd_addr_r_0__bdd_4_lut_14648.LUT_INIT = 16'he4aa;
    SB_LUT4 i4913_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_24_7 ), .O(n6412));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4913_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4912_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_24_6 ), .O(n6411));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4912_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16893_bdd_4_lut (.I0(n16893), .I1(\REG.mem_21_27 ), .I2(\REG.mem_20_27 ), 
            .I3(rd_addr_r[1]), .O(n15281));
    defparam n16893_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1295_1296 (.Q(\REG.mem_13_3 ), .C(FIFO_CLK_c), .D(n6056));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1292_1293 (.Q(\REG.mem_13_2 ), .C(FIFO_CLK_c), .D(n6055));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1289_1290 (.Q(\REG.mem_13_1 ), .C(FIFO_CLK_c), .D(n6054));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1286_1287 (.Q(\REG.mem_13_0 ), .C(FIFO_CLK_c), .D(n6053));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5074_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_29_8 ), .O(n6573));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5074_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5073_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_29_7 ), .O(n6572));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5073_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i332_333 (.Q(\REG.mem_3_2 ), .C(FIFO_CLK_c), .D(n5735));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i329_330 (.Q(\REG.mem_3_1 ), .C(FIFO_CLK_c), .D(n5734));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i326_327 (.Q(\REG.mem_3_0 ), .C(FIFO_CLK_c), .D(n5733));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15202 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_20 ), 
            .I2(\REG.mem_27_20 ), .I3(rd_addr_r[1]), .O(n17559));
    defparam rd_addr_r_0__bdd_4_lut_15202.LUT_INIT = 16'he4aa;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_5 (.CI(n13664), .I0(wp_sync_w[3]), 
            .I1(n1[3]), .CO(n13665));
    SB_LUT4 n17559_bdd_4_lut (.I0(n17559), .I1(\REG.mem_25_20 ), .I2(\REG.mem_24_20 ), 
            .I3(rd_addr_r[1]), .O(n15170));
    defparam n17559_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5072_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_29_6 ), .O(n6571));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5072_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5071_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_29_5 ), .O(n6570));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5071_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5070_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_29_4 ), .O(n6569));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5070_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5069_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_29_3 ), .O(n6568));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5069_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5068_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_29_2 ), .O(n6567));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5068_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5067_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_29_1 ), .O(n6566));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5067_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i323_324 (.Q(\REG.mem_2_31 ), .C(FIFO_CLK_c), .D(n5732));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14653 (.I0(rd_addr_r[2]), .I1(n15788), 
            .I2(n15797), .I3(rd_addr_r[3]), .O(n16887));
    defparam rd_addr_r_2__bdd_4_lut_14653.LUT_INIT = 16'he4aa;
    SB_LUT4 i5066_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_29_0 ), .O(n6565));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5066_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16887_bdd_4_lut (.I0(n16887), .I1(n15782), .I2(n15263), .I3(rd_addr_r[3]), 
            .O(n16890));
    defparam n16887_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15237 (.I0(rd_addr_r[1]), .I1(n15444), 
            .I2(n15445), .I3(rd_addr_r[2]), .O(n17553));
    defparam rd_addr_r_1__bdd_4_lut_15237.LUT_INIT = 16'he4aa;
    SB_LUT4 n17553_bdd_4_lut (.I0(n17553), .I1(n15412), .I2(n15411), .I3(rd_addr_r[2]), 
            .O(n17556));
    defparam n17553_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12609_3_lut (.I0(\REG.mem_0_28 ), .I1(\REG.mem_1_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14733));
    defparam i12609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12610_3_lut (.I0(\REG.mem_2_28 ), .I1(\REG.mem_3_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14734));
    defparam i12610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i22_2_lut_3_lut_4_lut (.I0(n6_adj_1378), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n22_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i22_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i12619_3_lut (.I0(\REG.mem_6_28 ), .I1(\REG.mem_7_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14743));
    defparam i12619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i23_2_lut_3_lut_4_lut (.I0(n6_adj_1378), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n23));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i23_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i12618_3_lut (.I0(\REG.mem_4_28 ), .I1(\REG.mem_5_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14742));
    defparam i12618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12642_3_lut (.I0(\REG.mem_24_28 ), .I1(\REG.mem_25_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14766));
    defparam i12642_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i320_321 (.Q(\REG.mem_2_30 ), .C(FIFO_CLK_c), .D(n5731));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i317_318 (.Q(\REG.mem_2_29 ), .C(FIFO_CLK_c), .D(n5730));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i314_315 (.Q(\REG.mem_2_28 ), .C(FIFO_CLK_c), .D(n5729));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i311_312 (.Q(\REG.mem_2_27 ), .C(FIFO_CLK_c), .D(n5728));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i308_309 (.Q(\REG.mem_2_26 ), .C(FIFO_CLK_c), .D(n5727));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14643 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_8 ), 
            .I2(\REG.mem_27_8 ), .I3(rd_addr_r[1]), .O(n16869));
    defparam rd_addr_r_0__bdd_4_lut_14643.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14144 (.I0(rd_addr_r[1]), .I1(n15864), 
            .I2(n15865), .I3(rd_addr_r[2]), .O(n16251));
    defparam rd_addr_r_1__bdd_4_lut_14144.LUT_INIT = 16'he4aa;
    SB_LUT4 i13048_3_lut (.I0(n16776), .I1(n17964), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15172));
    defparam i13048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n16869_bdd_4_lut (.I0(n16869), .I1(\REG.mem_25_8 ), .I2(\REG.mem_24_8 ), 
            .I3(rd_addr_r[1]), .O(n16872));
    defparam n16869_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14867 (.I0(rd_addr_r[3]), .I1(n16164), 
            .I2(n14722), .I3(rd_addr_r[4]), .O(n16863));
    defparam rd_addr_r_3__bdd_4_lut_14867.LUT_INIT = 16'he4aa;
    SB_LUT4 i12643_3_lut (.I0(\REG.mem_26_28 ), .I1(\REG.mem_27_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14767));
    defparam i12643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n16863_bdd_4_lut (.I0(n16863), .I1(n15241), .I2(n16860), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[10]));
    defparam n16863_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12646_3_lut (.I0(\REG.mem_30_28 ), .I1(\REG.mem_31_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14770));
    defparam i12646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12645_3_lut (.I0(\REG.mem_28_28 ), .I1(\REG.mem_29_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14769));
    defparam i12645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14663 (.I0(rd_addr_r[1]), .I1(n15195), 
            .I2(n15196), .I3(rd_addr_r[2]), .O(n16857));
    defparam rd_addr_r_1__bdd_4_lut_14663.LUT_INIT = 16'he4aa;
    SB_LUT4 n16857_bdd_4_lut (.I0(n16857), .I1(n15193), .I2(n15192), .I3(rd_addr_r[2]), 
            .O(n16860));
    defparam n16857_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_4_lut (.I0(n6_c), .I1(wp_sync_w[2]), 
            .I2(n1[2]), .I3(n13663), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_4_lut.LUT_INIT = 16'hebbe;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_4 (.CI(n13663), .I0(wp_sync_w[2]), 
            .I1(n1[2]), .CO(n13664));
    SB_LUT4 i12621_3_lut (.I0(\REG.mem_8_28 ), .I1(\REG.mem_9_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14745));
    defparam i12621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12622_3_lut (.I0(\REG.mem_10_28 ), .I1(\REG.mem_11_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14746));
    defparam i12622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_3_lut (.I0(n49), .I1(wp_sync_w[1]), 
            .I2(n1[1]), .I3(n13662), .O(n46)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_3 (.CI(n13662), .I0(wp_sync_w[1]), 
            .I1(n1[1]), .CO(n13663));
    SB_LUT4 i12628_3_lut (.I0(\REG.mem_14_28 ), .I1(\REG.mem_15_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14752));
    defparam i12628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_5__I_0_135_add_2_2_lut (.I0(n25), .I1(wp_sync_w[0]), 
            .I2(n1[0]), .I3(VCC_net), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_5__I_0_135_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i12627_3_lut (.I0(\REG.mem_12_28 ), .I1(\REG.mem_13_28 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14751));
    defparam i12627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4911_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_24_5 ), .O(n6410));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4911_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13335_3_lut (.I0(\REG.mem_8_25 ), .I1(\REG.mem_9_25 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15459));
    defparam i13335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15197 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_16 ), 
            .I2(\REG.mem_27_16 ), .I3(rd_addr_r[1]), .O(n17541));
    defparam rd_addr_r_0__bdd_4_lut_15197.LUT_INIT = 16'he4aa;
    SB_LUT4 i13336_3_lut (.I0(\REG.mem_10_25 ), .I1(\REG.mem_11_25 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15460));
    defparam i13336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17541_bdd_4_lut (.I0(n17541), .I1(\REG.mem_25_16 ), .I2(\REG.mem_24_16 ), 
            .I3(rd_addr_r[1]), .O(n15176));
    defparam n17541_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i6_1_lut (.I0(rd_grey_sync_r[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n1[5]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY wp_sync2_r_5__I_0_135_add_2_2 (.CI(VCC_net), .I0(wp_sync_w[0]), 
            .I1(n1[0]), .CO(n13662));
    SB_DFF i305_306 (.Q(\REG.mem_2_25 ), .C(FIFO_CLK_c), .D(n5726));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i302_303 (.Q(\REG.mem_2_24 ), .C(FIFO_CLK_c), .D(n5725));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i299_300 (.Q(\REG.mem_2_23 ), .C(FIFO_CLK_c), .D(n5724));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i296_297 (.Q(\REG.mem_2_22 ), .C(FIFO_CLK_c), .D(n5723));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i293_294 (.Q(\REG.mem_2_21 ), .C(FIFO_CLK_c), .D(n5722));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i290_291 (.Q(\REG.mem_2_20 ), .C(FIFO_CLK_c), .D(n5721));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i287_288 (.Q(\REG.mem_2_19 ), .C(FIFO_CLK_c), .D(n5720));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i284_285 (.Q(\REG.mem_2_18 ), .C(FIFO_CLK_c), .D(n5719));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i281_282 (.Q(\REG.mem_2_17 ), .C(FIFO_CLK_c), .D(n5718));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i13360_3_lut (.I0(\REG.mem_14_25 ), .I1(\REG.mem_15_25 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15484));
    defparam i13360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14623 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_22 ), 
            .I2(\REG.mem_27_22 ), .I3(rd_addr_r[1]), .O(n16845));
    defparam rd_addr_r_0__bdd_4_lut_14623.LUT_INIT = 16'he4aa;
    SB_DFF i1283_1284 (.Q(\REG.mem_12_31 ), .C(FIFO_CLK_c), .D(n6052));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n16251_bdd_4_lut (.I0(n16251), .I1(n15853), .I2(n15852), .I3(rd_addr_r[2]), 
            .O(n16254));
    defparam n16251_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16845_bdd_4_lut (.I0(n16845), .I1(\REG.mem_25_22 ), .I2(\REG.mem_24_22 ), 
            .I3(rd_addr_r[1]), .O(n16848));
    defparam n16845_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13359_3_lut (.I0(\REG.mem_12_25 ), .I1(\REG.mem_13_25 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15483));
    defparam i13359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15182 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_23 ), 
            .I2(\REG.mem_23_23 ), .I3(rd_addr_r[1]), .O(n17529));
    defparam rd_addr_r_0__bdd_4_lut_15182.LUT_INIT = 16'he4aa;
    SB_LUT4 i4910_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_24_4 ), .O(n6409));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4910_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14124 (.I0(rd_addr_r[2]), .I1(n15050), 
            .I2(n15083), .I3(rd_addr_r[3]), .O(n16245));
    defparam rd_addr_r_2__bdd_4_lut_14124.LUT_INIT = 16'he4aa;
    SB_LUT4 i4909_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_24_3 ), .O(n6408));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4909_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4908_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_24_2 ), .O(n6407));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4908_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14613 (.I0(rd_addr_r[1]), .I1(n15822), 
            .I2(n15823), .I3(rd_addr_r[2]), .O(n16839));
    defparam rd_addr_r_1__bdd_4_lut_14613.LUT_INIT = 16'he4aa;
    SB_LUT4 i4713_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_17_31 ), .O(n6212));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4713_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4712_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_17_30 ), .O(n6211));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4712_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17529_bdd_4_lut (.I0(n17529), .I1(\REG.mem_21_23 ), .I2(\REG.mem_20_23 ), 
            .I3(rd_addr_r[1]), .O(n15641));
    defparam n17529_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4907_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_24_1 ), .O(n6406));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4907_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4711_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_17_29 ), .O(n6210));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4711_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4710_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_17_28 ), .O(n6209));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4710_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16839_bdd_4_lut (.I0(n16839), .I1(n15814), .I2(n15813), .I3(rd_addr_r[2]), 
            .O(n16842));
    defparam n16839_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4709_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_17_27 ), .O(n6208));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4709_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4708_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_17_26 ), .O(n6207));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4708_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i278_279 (.Q(\REG.mem_2_16 ), .C(FIFO_CLK_c), .D(n5717));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i275_276 (.Q(\REG.mem_2_15 ), .C(FIFO_CLK_c), .D(n5716));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFE \REG.out_raw_i0_i1  (.Q(dc32_fifo_data_out[1]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[1]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_15222 (.I0(rd_addr_r[2]), .I1(n15590), 
            .I2(n15605), .I3(rd_addr_r[3]), .O(n17523));
    defparam rd_addr_r_2__bdd_4_lut_15222.LUT_INIT = 16'he4aa;
    SB_LUT4 n17523_bdd_4_lut (.I0(n17523), .I1(n16404), .I2(n15566), .I3(rd_addr_r[3]), 
            .O(n17526));
    defparam n17523_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15192 (.I0(rd_addr_r[1]), .I1(n15126), 
            .I2(n15127), .I3(rd_addr_r[2]), .O(n17517));
    defparam rd_addr_r_1__bdd_4_lut_15192.LUT_INIT = 16'he4aa;
    SB_DFFE \REG.out_raw_i0_i2  (.Q(dc32_fifo_data_out[2]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[2]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i3  (.Q(dc32_fifo_data_out[3]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[3]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i4  (.Q(dc32_fifo_data_out[4]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[4]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i5  (.Q(dc32_fifo_data_out[5]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[5]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i6  (.Q(dc32_fifo_data_out[6]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[6]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i7  (.Q(dc32_fifo_data_out[7]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[7]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i8  (.Q(dc32_fifo_data_out[8]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[8]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i9  (.Q(dc32_fifo_data_out[9]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[9]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i10  (.Q(dc32_fifo_data_out[10]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[10]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i11  (.Q(dc32_fifo_data_out[11]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[11]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i12  (.Q(dc32_fifo_data_out[12]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[12]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i13  (.Q(dc32_fifo_data_out[13]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[13]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i14  (.Q(dc32_fifo_data_out[14]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[14]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i15  (.Q(dc32_fifo_data_out[15]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[15]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i16  (.Q(dc32_fifo_data_out[16]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[16]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i17  (.Q(dc32_fifo_data_out[17]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[17]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i18  (.Q(dc32_fifo_data_out[18]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[18]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i19  (.Q(dc32_fifo_data_out[19]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[19]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i20  (.Q(dc32_fifo_data_out[20]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[20]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i21  (.Q(dc32_fifo_data_out[21]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[21]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i22  (.Q(dc32_fifo_data_out[22]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[22]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i23  (.Q(dc32_fifo_data_out[23]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[23]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i24  (.Q(dc32_fifo_data_out[24]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[24]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i25  (.Q(dc32_fifo_data_out[25]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[25]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i26  (.Q(dc32_fifo_data_out[26]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[26]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i27  (.Q(dc32_fifo_data_out[27]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[27]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i28  (.Q(dc32_fifo_data_out[28]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[28]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i29  (.Q(dc32_fifo_data_out[29]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[29]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i30  (.Q(dc32_fifo_data_out[30]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[30]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw_i0_i31  (.Q(dc32_fifo_data_out[31]), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(rd_data_o_31__N_598[31]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 n16245_bdd_4_lut (.I0(n16245), .I1(n15044), .I2(n15035), .I3(rd_addr_r[3]), 
            .O(n16248));
    defparam n16245_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14638 (.I0(rd_addr_r[2]), .I1(n15833), 
            .I2(n15842), .I3(rd_addr_r[3]), .O(n16833));
    defparam rd_addr_r_2__bdd_4_lut_14638.LUT_INIT = 16'he4aa;
    SB_LUT4 i4906_3_lut_4_lut (.I0(n20), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_24_0 ), .O(n6405));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4906_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4707_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_17_25 ), .O(n6206));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4707_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4706_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_17_24 ), .O(n6205));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4706_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16833_bdd_4_lut (.I0(n16833), .I1(n15818), .I2(n15806), .I3(rd_addr_r[3]), 
            .O(n16836));
    defparam n16833_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4705_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_17_23 ), .O(n6204));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4705_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i272_273 (.Q(\REG.mem_2_14 ), .C(FIFO_CLK_c), .D(n5715));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14598 (.I0(rd_addr_r[1]), .I1(n15456), 
            .I2(n15457), .I3(rd_addr_r[2]), .O(n16827));
    defparam rd_addr_r_1__bdd_4_lut_14598.LUT_INIT = 16'he4aa;
    SB_LUT4 i4704_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_17_22 ), .O(n6203));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4704_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1280_1281 (.Q(\REG.mem_12_30 ), .C(FIFO_CLK_c), .D(n6051));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1277_1278 (.Q(\REG.mem_12_29 ), .C(FIFO_CLK_c), .D(n6050));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14119 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_30 ), 
            .I2(\REG.mem_31_30 ), .I3(rd_addr_r[1]), .O(n16239));
    defparam rd_addr_r_0__bdd_4_lut_14119.LUT_INIT = 16'he4aa;
    SB_LUT4 n16827_bdd_4_lut (.I0(n16827), .I1(n15064), .I2(n15063), .I3(rd_addr_r[2]), 
            .O(n16830));
    defparam n16827_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16239_bdd_4_lut (.I0(n16239), .I1(\REG.mem_29_30 ), .I2(\REG.mem_28_30 ), 
            .I3(rd_addr_r[1]), .O(n16242));
    defparam n16239_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17517_bdd_4_lut (.I0(n17517), .I1(n15115), .I2(n15114), .I3(rd_addr_r[2]), 
            .O(n15181));
    defparam n17517_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15172 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_23 ), 
            .I2(\REG.mem_27_23 ), .I3(rd_addr_r[1]), .O(n17511));
    defparam rd_addr_r_0__bdd_4_lut_15172.LUT_INIT = 16'he4aa;
    SB_DFF i1274_1275 (.Q(\REG.mem_12_28 ), .C(FIFO_CLK_c), .D(n6049));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1271_1272 (.Q(\REG.mem_12_27 ), .C(FIFO_CLK_c), .D(n6048));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1268_1269 (.Q(\REG.mem_12_26 ), .C(FIFO_CLK_c), .D(n6047));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1265_1266 (.Q(\REG.mem_12_25 ), .C(FIFO_CLK_c), .D(n6046));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4703_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_17_21 ), .O(n6202));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4703_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4702_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_17_20 ), .O(n6201));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4702_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1262_1263 (.Q(\REG.mem_12_24 ), .C(FIFO_CLK_c), .D(n6045));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1259_1260 (.Q(\REG.mem_12_23 ), .C(FIFO_CLK_c), .D(n6044));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1256_1257 (.Q(\REG.mem_12_22 ), .C(FIFO_CLK_c), .D(n6043));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4701_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_17_19 ), .O(n6200));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4701_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14603 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_22 ), 
            .I2(\REG.mem_31_22 ), .I3(rd_addr_r[1]), .O(n16821));
    defparam rd_addr_r_0__bdd_4_lut_14603.LUT_INIT = 16'he4aa;
    SB_LUT4 n16821_bdd_4_lut (.I0(n16821), .I1(\REG.mem_29_22 ), .I2(\REG.mem_28_22 ), 
            .I3(rd_addr_r[1]), .O(n16824));
    defparam n16821_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1253_1254 (.Q(\REG.mem_12_21 ), .C(FIFO_CLK_c), .D(n6042));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n17511_bdd_4_lut (.I0(n17511), .I1(\REG.mem_25_23 ), .I2(\REG.mem_24_23 ), 
            .I3(rd_addr_r[1]), .O(n15647));
    defparam n17511_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4700_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_17_18 ), .O(n6199));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4700_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4699_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_17_17 ), .O(n6198));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4699_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4698_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_17_16 ), .O(n6197));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4698_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15157 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_18 ), 
            .I2(\REG.mem_15_18 ), .I3(rd_addr_r[1]), .O(n17505));
    defparam rd_addr_r_0__bdd_4_lut_15157.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i4_2_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(wr_fifo_en_w), .I3(\wr_addr_nxt_c[4] ), .O(wr_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_5__I_0_136_i4_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4697_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_17_15 ), .O(n6196));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4697_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i269_270 (.Q(\REG.mem_2_13 ), .C(FIFO_CLK_c), .D(n5714));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1250_1251 (.Q(\REG.mem_12_20 ), .C(FIFO_CLK_c), .D(n6041));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n17505_bdd_4_lut (.I0(n17505), .I1(\REG.mem_13_18 ), .I2(\REG.mem_12_18 ), 
            .I3(rd_addr_r[1]), .O(n15650));
    defparam n17505_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14593 (.I0(rd_addr_r[2]), .I1(n15101), 
            .I2(n15131), .I3(rd_addr_r[3]), .O(n16809));
    defparam rd_addr_r_2__bdd_4_lut_14593.LUT_INIT = 16'he4aa;
    SB_LUT4 n16809_bdd_4_lut (.I0(n16809), .I1(n15095), .I2(n15080), .I3(rd_addr_r[3]), 
            .O(n16812));
    defparam n16809_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15152 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_21 ), 
            .I2(\REG.mem_19_21 ), .I3(rd_addr_r[1]), .O(n17499));
    defparam rd_addr_r_0__bdd_4_lut_15152.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14618 (.I0(rd_addr_r[3]), .I1(n16386), 
            .I2(n14800), .I3(rd_addr_r[4]), .O(n16803));
    defparam rd_addr_r_3__bdd_4_lut_14618.LUT_INIT = 16'he4aa;
    SB_LUT4 n16803_bdd_4_lut (.I0(n16803), .I1(n15181), .I2(n16800), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[11]));
    defparam n16803_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1247_1248 (.Q(\REG.mem_12_19 ), .C(FIFO_CLK_c), .D(n6040));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1244_1245 (.Q(\REG.mem_12_18 ), .C(FIFO_CLK_c), .D(n6039));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1241_1242 (.Q(\REG.mem_12_17 ), .C(FIFO_CLK_c), .D(n6038));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1238_1239 (.Q(\REG.mem_12_16 ), .C(FIFO_CLK_c), .D(n6037));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n17499_bdd_4_lut (.I0(n17499), .I1(\REG.mem_17_21 ), .I2(\REG.mem_16_21 ), 
            .I3(rd_addr_r[1]), .O(n15185));
    defparam n17499_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_15167 (.I0(rd_addr_r[2]), .I1(n15617), 
            .I2(n15626), .I3(rd_addr_r[3]), .O(n17493));
    defparam rd_addr_r_2__bdd_4_lut_15167.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14588 (.I0(rd_addr_r[1]), .I1(n15108), 
            .I2(n15109), .I3(rd_addr_r[2]), .O(n16797));
    defparam rd_addr_r_1__bdd_4_lut_14588.LUT_INIT = 16'he4aa;
    SB_LUT4 n17493_bdd_4_lut (.I0(n17493), .I1(n15614), .I2(n15608), .I3(rd_addr_r[3]), 
            .O(n17496));
    defparam n17493_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4696_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_17_14 ), .O(n6195));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4696_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4695_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_17_13 ), .O(n6194));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4695_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16797_bdd_4_lut (.I0(n16797), .I1(n15091), .I2(n15090), .I3(rd_addr_r[2]), 
            .O(n16800));
    defparam n16797_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4694_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_17_12 ), .O(n6193));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4694_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i3_2_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(wr_fifo_en_w), .I3(\wr_addr_nxt_c[2] ), .O(wr_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_5__I_0_136_i3_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4693_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_17_11 ), .O(n6192));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4693_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1235_1236 (.Q(\REG.mem_12_15 ), .C(FIFO_CLK_c), .D(n6036));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1232_1233 (.Q(\REG.mem_12_14 ), .C(FIFO_CLK_c), .D(n6035));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4692_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_17_10 ), .O(n6191));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4692_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4691_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_17_9 ), .O(n6190));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4691_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4690_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_17_8 ), .O(n6189));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4690_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5455_2_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(wr_fifo_en_w), .I3(reset_per_frame), .O(n6954));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i5455_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_DFF i1229_1230 (.Q(\REG.mem_12_13 ), .C(FIFO_CLK_c), .D(n6034));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1226_1227 (.Q(\REG.mem_12_12 ), .C(FIFO_CLK_c), .D(n6033));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1223_1224 (.Q(\REG.mem_12_11 ), .C(FIFO_CLK_c), .D(n6032));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1220_1221 (.Q(\REG.mem_12_10 ), .C(FIFO_CLK_c), .D(n6031));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1217_1218 (.Q(\REG.mem_12_9 ), .C(FIFO_CLK_c), .D(n6030));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1214_1215 (.Q(\REG.mem_12_8 ), .C(FIFO_CLK_c), .D(n6029));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1211_1212 (.Q(\REG.mem_12_7 ), .C(FIFO_CLK_c), .D(n6028));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1208_1209 (.Q(\REG.mem_12_6 ), .C(FIFO_CLK_c), .D(n6027));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1205_1206 (.Q(\REG.mem_12_5 ), .C(FIFO_CLK_c), .D(n6026));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1202_1203 (.Q(\REG.mem_12_4 ), .C(FIFO_CLK_c), .D(n6025));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i13026_3_lut (.I0(\REG.mem_16_8 ), .I1(\REG.mem_17_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15150));
    defparam i13026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14563 (.I0(rd_addr_r[1]), .I1(n15651), 
            .I2(n15652), .I3(rd_addr_r[2]), .O(n16791));
    defparam rd_addr_r_1__bdd_4_lut_14563.LUT_INIT = 16'he4aa;
    SB_LUT4 i4689_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_17_7 ), .O(n6188));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4689_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13027_3_lut (.I0(\REG.mem_18_8 ), .I1(\REG.mem_19_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15151));
    defparam i13027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15162 (.I0(rd_addr_r[1]), .I1(n14763), 
            .I2(n14764), .I3(rd_addr_r[2]), .O(n17481));
    defparam rd_addr_r_1__bdd_4_lut_15162.LUT_INIT = 16'he4aa;
    SB_LUT4 n16791_bdd_4_lut (.I0(n16791), .I1(n15610), .I2(n15609), .I3(rd_addr_r[2]), 
            .O(n15886));
    defparam n16791_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14583 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_14 ), 
            .I2(\REG.mem_23_14 ), .I3(rd_addr_r[1]), .O(n16785));
    defparam rd_addr_r_0__bdd_4_lut_14583.LUT_INIT = 16'he4aa;
    SB_LUT4 n17481_bdd_4_lut (.I0(n17481), .I1(n14749), .I2(n14748), .I3(rd_addr_r[2]), 
            .O(n15190));
    defparam n17481_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i266_267 (.Q(\REG.mem_2_12 ), .C(FIFO_CLK_c), .D(n5713));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_nxt_c_5__I_0_136_i5_2_lut_4_lut (.I0(\wr_addr_r[5] ), 
            .I1(wr_addr_p1_w[5]), .I2(wr_fifo_en_w), .I3(\wr_addr_nxt_c[4] ), 
            .O(wr_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_5__I_0_136_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_DFF i263_264 (.Q(\REG.mem_2_11 ), .C(FIFO_CLK_c), .D(n5712));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5453_2_lut_4_lut (.I0(\wr_addr_r[5] ), .I1(wr_addr_p1_w[5]), 
            .I2(wr_fifo_en_w), .I3(reset_per_frame), .O(n6952));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i5453_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 n16785_bdd_4_lut (.I0(n16785), .I1(\REG.mem_21_14 ), .I2(\REG.mem_20_14 ), 
            .I3(rd_addr_r[1]), .O(n16788));
    defparam n16785_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15132 (.I0(rd_addr_r[1]), .I1(n15576), 
            .I2(n15577), .I3(rd_addr_r[2]), .O(n17475));
    defparam rd_addr_r_1__bdd_4_lut_15132.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14558 (.I0(rd_addr_r[1]), .I1(n15876), 
            .I2(n15877), .I3(rd_addr_r[2]), .O(n16779));
    defparam rd_addr_r_1__bdd_4_lut_14558.LUT_INIT = 16'he4aa;
    SB_LUT4 n16779_bdd_4_lut (.I0(n16779), .I1(n15859), .I2(n15858), .I3(rd_addr_r[2]), 
            .O(n16782));
    defparam n16779_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17475_bdd_4_lut (.I0(n17475), .I1(n14965), .I2(n14964), .I3(rd_addr_r[2]), 
            .O(n15552));
    defparam n17475_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR rd_grey_sync_r__i1 (.Q(rd_grey_sync_r[1]), .C(SLM_CLK_c), .D(rd_grey_w[1]), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i2 (.Q(rd_grey_sync_r[2]), .C(SLM_CLK_c), .D(rd_grey_w[2]), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i3 (.Q(rd_grey_sync_r[3]), .C(SLM_CLK_c), .D(rd_grey_w[3]), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i4 (.Q(rd_grey_sync_r[4]), .C(SLM_CLK_c), .D(rd_grey_w[4]), 
            .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR wr_grey_sync_r__i1 (.Q(\wr_grey_sync_r[1] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[1]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFSR wr_grey_sync_r__i2 (.Q(\wr_grey_sync_r[2] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[2]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_LUT4 i4688_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_17_6 ), .O(n6187));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4688_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4687_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_17_5 ), .O(n6186));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4687_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4686_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_17_4 ), .O(n6185));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4686_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14553 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_5 ), 
            .I2(\REG.mem_11_5 ), .I3(rd_addr_r[1]), .O(n16773));
    defparam rd_addr_r_0__bdd_4_lut_14553.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15147 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_2 ), 
            .I2(\REG.mem_3_2 ), .I3(rd_addr_r[1]), .O(n17463));
    defparam rd_addr_r_0__bdd_4_lut_15147.LUT_INIT = 16'he4aa;
    SB_LUT4 i4685_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_17_3 ), .O(n6184));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4685_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4684_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_17_2 ), .O(n6183));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4684_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFSR wr_grey_sync_r__i3 (.Q(\wr_grey_sync_r[3] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[3]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFSR wr_grey_sync_r__i4 (.Q(\wr_grey_sync_r[4] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[4]), .R(reset_per_frame));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_LUT4 i4683_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_17_1 ), .O(n6182));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4683_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4682_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_17_0 ), .O(n6181));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4682_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5065_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_28_31 ), .O(n6564));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5065_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5064_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_28_30 ), .O(n6563));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5064_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5063_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_28_29 ), .O(n6562));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5063_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5062_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_28_28 ), .O(n6561));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5062_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17463_bdd_4_lut (.I0(n17463), .I1(\REG.mem_1_2 ), .I2(\REG.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(n15665));
    defparam n17463_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16773_bdd_4_lut (.I0(n16773), .I1(\REG.mem_9_5 ), .I2(\REG.mem_8_5 ), 
            .I3(rd_addr_r[1]), .O(n16776));
    defparam n16773_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15117 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_18 ), 
            .I2(\REG.mem_19_18 ), .I3(rd_addr_r[1]), .O(n17457));
    defparam rd_addr_r_0__bdd_4_lut_15117.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14573 (.I0(rd_addr_r[2]), .I1(n15170), 
            .I2(n15278), .I3(rd_addr_r[3]), .O(n16767));
    defparam rd_addr_r_2__bdd_4_lut_14573.LUT_INIT = 16'he4aa;
    SB_LUT4 n16767_bdd_4_lut (.I0(n16767), .I1(n15164), .I2(n15149), .I3(rd_addr_r[3]), 
            .O(n16770));
    defparam n16767_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17457_bdd_4_lut (.I0(n17457), .I1(\REG.mem_17_18 ), .I2(\REG.mem_16_18 ), 
            .I3(rd_addr_r[1]), .O(n15668));
    defparam n17457_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1199_1200 (.Q(\REG.mem_12_3 ), .C(FIFO_CLK_c), .D(n6024));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1196_1197 (.Q(\REG.mem_12_2 ), .C(FIFO_CLK_c), .D(n6023));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14548 (.I0(rd_addr_r[1]), .I1(n15846), 
            .I2(n15847), .I3(rd_addr_r[2]), .O(n16761));
    defparam rd_addr_r_1__bdd_4_lut_14548.LUT_INIT = 16'he4aa;
    SB_LUT4 n16761_bdd_4_lut (.I0(n16761), .I1(n15475), .I2(n15474), .I3(rd_addr_r[2]), 
            .O(n15898));
    defparam n16761_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14543 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_9 ), 
            .I2(\REG.mem_27_9 ), .I3(rd_addr_r[1]), .O(n16755));
    defparam rd_addr_r_0__bdd_4_lut_14543.LUT_INIT = 16'he4aa;
    SB_LUT4 n16755_bdd_4_lut (.I0(n16755), .I1(\REG.mem_25_9 ), .I2(\REG.mem_24_9 ), 
            .I3(rd_addr_r[1]), .O(n16758));
    defparam n16755_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5061_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_28_27 ), .O(n6560));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5061_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5060_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_28_26 ), .O(n6559));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5060_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1193_1194 (.Q(\REG.mem_12_1 ), .C(FIFO_CLK_c), .D(n6022));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1190_1191 (.Q(\REG.mem_12_0 ), .C(FIFO_CLK_c), .D(n6021));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1187_1188 (.Q(\REG.mem_11_31 ), .C(FIFO_CLK_c), .D(n6020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1184_1185 (.Q(\REG.mem_11_30 ), .C(FIFO_CLK_c), .D(n6019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1181_1182 (.Q(\REG.mem_11_29 ), .C(FIFO_CLK_c), .D(n6018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1178_1179 (.Q(\REG.mem_11_28 ), .C(FIFO_CLK_c), .D(n6017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1175_1176 (.Q(\REG.mem_11_27 ), .C(FIFO_CLK_c), .D(n6016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1172_1173 (.Q(\REG.mem_11_26 ), .C(FIFO_CLK_c), .D(n6015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1169_1170 (.Q(\REG.mem_11_25 ), .C(FIFO_CLK_c), .D(n6014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1166_1167 (.Q(\REG.mem_11_24 ), .C(FIFO_CLK_c), .D(n6013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1163_1164 (.Q(\REG.mem_11_23 ), .C(FIFO_CLK_c), .D(n6012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1160_1161 (.Q(\REG.mem_11_22 ), .C(FIFO_CLK_c), .D(n6011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1157_1158 (.Q(\REG.mem_11_21 ), .C(FIFO_CLK_c), .D(n6010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1154_1155 (.Q(\REG.mem_11_20 ), .C(FIFO_CLK_c), .D(n6009));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1151_1152 (.Q(\REG.mem_11_19 ), .C(FIFO_CLK_c), .D(n6008));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1148_1149 (.Q(\REG.mem_11_18 ), .C(FIFO_CLK_c), .D(n6007));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15127 (.I0(rd_addr_r[1]), .I1(n15165), 
            .I2(n15166), .I3(rd_addr_r[2]), .O(n17451));
    defparam rd_addr_r_1__bdd_4_lut_15127.LUT_INIT = 16'he4aa;
    SB_LUT4 n17451_bdd_4_lut (.I0(n17451), .I1(n15160), .I2(n15159), .I3(rd_addr_r[2]), 
            .O(n14800));
    defparam n17451_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14528 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_21 ), 
            .I2(\REG.mem_31_21 ), .I3(rd_addr_r[1]), .O(n16749));
    defparam rd_addr_r_0__bdd_4_lut_14528.LUT_INIT = 16'he4aa;
    SB_LUT4 n16749_bdd_4_lut (.I0(n16749), .I1(\REG.mem_29_21 ), .I2(\REG.mem_28_21 ), 
            .I3(rd_addr_r[1]), .O(n15293));
    defparam n16749_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15112 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_6 ), 
            .I2(\REG.mem_11_6 ), .I3(rd_addr_r[1]), .O(n17445));
    defparam rd_addr_r_0__bdd_4_lut_15112.LUT_INIT = 16'he4aa;
    SB_LUT4 i5059_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_28_25 ), .O(n6558));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5059_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17445_bdd_4_lut (.I0(n17445), .I1(\REG.mem_9_6 ), .I2(\REG.mem_8_6 ), 
            .I3(rd_addr_r[1]), .O(n17448));
    defparam n17445_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5058_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_28_24 ), .O(n6557));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5058_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14523 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_17 ), 
            .I2(\REG.mem_15_17 ), .I3(rd_addr_r[1]), .O(n16743));
    defparam rd_addr_r_0__bdd_4_lut_14523.LUT_INIT = 16'he4aa;
    SB_LUT4 i5057_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_28_23 ), .O(n6556));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5057_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5056_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_28_22 ), .O(n6555));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5056_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5055_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_28_21 ), .O(n6554));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5055_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16743_bdd_4_lut (.I0(n16743), .I1(\REG.mem_13_17 ), .I2(\REG.mem_12_17 ), 
            .I3(rd_addr_r[1]), .O(n15296));
    defparam n16743_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5054_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_28_20 ), .O(n6553));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5054_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_15142 (.I0(rd_addr_r[2]), .I1(n15647), 
            .I2(n16536), .I3(rd_addr_r[3]), .O(n17439));
    defparam rd_addr_r_2__bdd_4_lut_15142.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14518 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_9 ), 
            .I2(\REG.mem_31_9 ), .I3(rd_addr_r[1]), .O(n16737));
    defparam rd_addr_r_0__bdd_4_lut_14518.LUT_INIT = 16'he4aa;
    SB_LUT4 n17439_bdd_4_lut (.I0(n17439), .I1(n15641), .I2(n15635), .I3(rd_addr_r[3]), 
            .O(n17442));
    defparam n17439_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5053_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_28_19 ), .O(n6552));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5053_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5052_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_28_18 ), .O(n6551));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5052_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1145_1146 (.Q(\REG.mem_11_17 ), .C(FIFO_CLK_c), .D(n6006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1142_1143 (.Q(\REG.mem_11_16 ), .C(FIFO_CLK_c), .D(n6005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1139_1140 (.Q(\REG.mem_11_15 ), .C(FIFO_CLK_c), .D(n6004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1136_1137 (.Q(\REG.mem_11_14 ), .C(FIFO_CLK_c), .D(n6003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1133_1134 (.Q(\REG.mem_11_13 ), .C(FIFO_CLK_c), .D(n6002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1130_1131 (.Q(\REG.mem_11_12 ), .C(FIFO_CLK_c), .D(n6001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1127_1128 (.Q(\REG.mem_11_11 ), .C(FIFO_CLK_c), .D(n6000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1124_1125 (.Q(\REG.mem_11_10 ), .C(FIFO_CLK_c), .D(n5999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1121_1122 (.Q(\REG.mem_11_9 ), .C(FIFO_CLK_c), .D(n5998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14105 (.I0(rd_addr_r[2]), .I1(n14909), 
            .I2(n14912), .I3(rd_addr_r[3]), .O(n16233));
    defparam rd_addr_r_2__bdd_4_lut_14105.LUT_INIT = 16'he4aa;
    SB_LUT4 i5051_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_28_17 ), .O(n6550));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5051_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16737_bdd_4_lut (.I0(n16737), .I1(\REG.mem_29_9 ), .I2(\REG.mem_28_9 ), 
            .I3(rd_addr_r[1]), .O(n16740));
    defparam n16737_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15102 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_16 ), 
            .I2(\REG.mem_31_16 ), .I3(rd_addr_r[1]), .O(n17433));
    defparam rd_addr_r_0__bdd_4_lut_15102.LUT_INIT = 16'he4aa;
    SB_LUT4 n17433_bdd_4_lut (.I0(n17433), .I1(\REG.mem_29_16 ), .I2(\REG.mem_28_16 ), 
            .I3(rd_addr_r[1]), .O(n15200));
    defparam n17433_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14533 (.I0(rd_addr_r[1]), .I1(n14997), 
            .I2(n14998), .I3(rd_addr_r[2]), .O(n16731));
    defparam rd_addr_r_1__bdd_4_lut_14533.LUT_INIT = 16'he4aa;
    SB_LUT4 n16731_bdd_4_lut (.I0(n16731), .I1(n14995), .I2(n14994), .I3(rd_addr_r[2]), 
            .O(n15138));
    defparam n16731_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_r_5__I_0_add_2_7_lut (.I0(n13844), .I1(\wr_addr_r[5] ), 
            .I2(n1_adj_1394[5]), .I3(n13702), .O(\afull_flag_impl.af_flag_nxt_w )) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 wr_addr_r_5__I_0_add_2_6_lut (.I0(n6_adj_1384), .I1(wr_addr_r[4]), 
            .I2(rp_sync_w[4]), .I3(n13701), .O(n8_adj_1383)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5050_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_28_16 ), .O(n6549));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5050_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY wr_addr_r_5__I_0_add_2_6 (.CI(n13701), .I0(wr_addr_r[4]), .I1(rp_sync_w[4]), 
            .CO(n13702));
    SB_LUT4 wr_addr_r_5__I_0_add_2_5_lut (.I0(wr_sig_diff0_w[1]), .I1(wr_addr_r[3]), 
            .I2(rp_sync_w[3]), .I3(n13700), .O(n6_adj_1384)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY wr_addr_r_5__I_0_add_2_5 (.CI(n13700), .I0(wr_addr_r[3]), .I1(rp_sync_w[3]), 
            .CO(n13701));
    SB_LUT4 wr_addr_r_5__I_0_add_2_4_lut (.I0(n14_adj_1386), .I1(wr_addr_r[2]), 
            .I2(rp_sync_w[2]), .I3(n13699), .O(n7_adj_1385)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY wr_addr_r_5__I_0_add_2_4 (.CI(n13699), .I0(wr_addr_r[2]), .I1(rp_sync_w[2]), 
            .CO(n13700));
    SB_LUT4 wr_addr_r_5__I_0_add_2_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), 
            .I2(rp_sync_w[1]), .I3(n13698), .O(wr_sig_diff0_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5049_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_28_15 ), .O(n6548));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5049_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14056 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_4 ), 
            .I2(\REG.mem_23_4 ), .I3(rd_addr_r[1]), .O(n16179));
    defparam rd_addr_r_0__bdd_4_lut_14056.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14513 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_2 ), 
            .I2(\REG.mem_31_2 ), .I3(rd_addr_r[1]), .O(n16719));
    defparam rd_addr_r_0__bdd_4_lut_14513.LUT_INIT = 16'he4aa;
    SB_LUT4 i5048_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_28_14 ), .O(n6547));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5048_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY wr_addr_r_5__I_0_add_2_3 (.CI(n13698), .I0(wr_addr_r[1]), .I1(rp_sync_w[1]), 
            .CO(n13699));
    SB_LUT4 n16719_bdd_4_lut (.I0(n16719), .I1(\REG.mem_29_2 ), .I2(\REG.mem_28_2 ), 
            .I3(rd_addr_r[1]), .O(n16722));
    defparam n16719_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_15217 (.I0(rd_addr_r[3]), .I1(n15579), 
            .I2(n15580), .I3(rd_addr_r[4]), .O(n17421));
    defparam rd_addr_r_3__bdd_4_lut_15217.LUT_INIT = 16'he4aa;
    SB_LUT4 n17421_bdd_4_lut (.I0(n17421), .I1(n15547), .I2(n15546), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[7]));
    defparam n17421_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_5__I_0_137_7_lut (.I0(GND_net), .I1(rd_grey_sync_r[5]), 
            .I2(GND_net), .I3(n13727), .O(rd_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wr_addr_r_5__I_0_add_2_2_lut (.I0(DEBUG_5_c), .I1(\wr_addr_r[0] ), 
            .I2(rp_sync_w[0]), .I3(VCC_net), .O(n14_adj_1386)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 rd_addr_r_5__I_0_137_6_lut (.I0(GND_net), .I1(rd_addr_r[4]), 
            .I2(GND_net), .I3(n13726), .O(rd_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_5__I_0_add_2_2 (.CI(VCC_net), .I0(\wr_addr_r[0] ), 
            .I1(rp_sync_w[0]), .CO(n13698));
    SB_CARRY rd_addr_r_5__I_0_137_6 (.CI(n13726), .I0(rd_addr_r[4]), .I1(GND_net), 
            .CO(n13727));
    SB_LUT4 i5047_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_28_13 ), .O(n6546));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5047_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_5__I_0_137_5_lut (.I0(GND_net), .I1(rd_addr_r[3]), 
            .I2(GND_net), .I3(n13725), .O(rd_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rd_addr_r_5__I_0_137_5 (.CI(n13725), .I0(rd_addr_r[3]), .I1(GND_net), 
            .CO(n13726));
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14498 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_27 ), 
            .I2(\REG.mem_3_27 ), .I3(rd_addr_r[1]), .O(n16707));
    defparam rd_addr_r_0__bdd_4_lut_14498.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_15097 (.I0(rd_addr_r[2]), .I1(n14960), 
            .I2(n15077), .I3(rd_addr_r[3]), .O(n17415));
    defparam rd_addr_r_2__bdd_4_lut_15097.LUT_INIT = 16'he4aa;
    SB_LUT4 i5046_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_28_12 ), .O(n6545));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5046_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16707_bdd_4_lut (.I0(n16707), .I1(\REG.mem_1_27 ), .I2(\REG.mem_0_27 ), 
            .I3(rd_addr_r[1]), .O(n16710));
    defparam n16707_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17415_bdd_4_lut (.I0(n17415), .I1(n14948), .I2(n16710), .I3(rd_addr_r[3]), 
            .O(n17418));
    defparam n17415_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_5__I_0_137_4_lut (.I0(GND_net), .I1(rd_addr_r[2]), 
            .I2(GND_net), .I3(n13724), .O(rd_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rd_addr_r_5__I_0_137_4 (.CI(n13724), .I0(rd_addr_r[2]), .I1(GND_net), 
            .CO(n13725));
    SB_LUT4 rd_addr_r_5__I_0_137_3_lut (.I0(GND_net), .I1(rd_addr_r[1]), 
            .I2(GND_net), .I3(n13723), .O(rd_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5045_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_28_11 ), .O(n6544));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5045_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY rd_addr_r_5__I_0_137_3 (.CI(n13723), .I0(rd_addr_r[1]), .I1(GND_net), 
            .CO(n13724));
    SB_LUT4 rd_addr_r_5__I_0_137_2_lut (.I0(GND_net), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(VCC_net), .O(rd_addr_p1_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_5__I_0_137_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15092 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_2 ), 
            .I2(\REG.mem_11_2 ), .I3(rd_addr_r[1]), .O(n17409));
    defparam rd_addr_r_0__bdd_4_lut_15092.LUT_INIT = 16'he4aa;
    SB_CARRY rd_addr_r_5__I_0_137_2 (.CI(VCC_net), .I0(rd_addr_r[0]), .I1(GND_net), 
            .CO(n13723));
    SB_LUT4 i5044_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_28_10 ), .O(n6543));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5044_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13054_3_lut (.I0(\REG.mem_22_8 ), .I1(\REG.mem_23_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15178));
    defparam i13054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5043_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_28_9 ), .O(n6542));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5043_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14488 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_2 ), 
            .I2(\REG.mem_19_2 ), .I3(rd_addr_r[1]), .O(n16695));
    defparam rd_addr_r_0__bdd_4_lut_14488.LUT_INIT = 16'he4aa;
    SB_LUT4 i13053_3_lut (.I0(\REG.mem_20_8 ), .I1(\REG.mem_21_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15177));
    defparam i13053_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1118_1119 (.Q(\REG.mem_11_8 ), .C(FIFO_CLK_c), .D(n5997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1115_1116 (.Q(\REG.mem_11_7 ), .C(FIFO_CLK_c), .D(n5996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1112_1113 (.Q(\REG.mem_11_6 ), .C(FIFO_CLK_c), .D(n5995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1109_1110 (.Q(\REG.mem_11_5 ), .C(FIFO_CLK_c), .D(n5994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i260_261 (.Q(\REG.mem_2_10 ), .C(FIFO_CLK_c), .D(n5711));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4297_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_4_31 ), .O(n5796));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4297_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i257_258 (.Q(\REG.mem_2_9 ), .C(FIFO_CLK_c), .D(n5710));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i254_255 (.Q(\REG.mem_2_8 ), .C(FIFO_CLK_c), .D(n5709));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i251_252 (.Q(\REG.mem_2_7 ), .C(FIFO_CLK_c), .D(n5708));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i248_249 (.Q(\REG.mem_2_6 ), .C(FIFO_CLK_c), .D(n5707));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i71_72 (.Q(\REG.mem_0_11 ), .C(FIFO_CLK_c), .D(n5706));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i74_75 (.Q(\REG.mem_0_12 ), .C(FIFO_CLK_c), .D(n5705));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i77_78 (.Q(\REG.mem_0_13 ), .C(FIFO_CLK_c), .D(n5704));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i80_81 (.Q(\REG.mem_0_14 ), .C(FIFO_CLK_c), .D(n5702));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4296_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_4_30 ), .O(n5795));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4296_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5042_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_28_8 ), .O(n6541));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5042_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17409_bdd_4_lut (.I0(n17409), .I1(\REG.mem_9_2 ), .I2(\REG.mem_8_2 ), 
            .I3(rd_addr_r[1]), .O(n15680));
    defparam n17409_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5041_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_28_7 ), .O(n6540));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5041_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5040_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_28_6 ), .O(n6539));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5040_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i30_2_lut (.I0(n14), .I1(wr_addr_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n30));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4295_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_4_29 ), .O(n5794));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4295_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16695_bdd_4_lut (.I0(n16695), .I1(\REG.mem_17_2 ), .I2(\REG.mem_16_2 ), 
            .I3(rd_addr_r[1]), .O(n16698));
    defparam n16695_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15072 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_6 ), 
            .I2(\REG.mem_15_6 ), .I3(rd_addr_r[1]), .O(n17403));
    defparam rd_addr_r_0__bdd_4_lut_15072.LUT_INIT = 16'he4aa;
    SB_DFF i83_84 (.Q(\REG.mem_0_15 ), .C(FIFO_CLK_c), .D(n5701));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i86_87 (.Q(\REG.mem_0_16 ), .C(FIFO_CLK_c), .D(n5700));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1106_1107 (.Q(\REG.mem_11_4 ), .C(FIFO_CLK_c), .D(n5993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i5039_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_28_5 ), .O(n6538));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5039_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17403_bdd_4_lut (.I0(n17403), .I1(\REG.mem_13_6 ), .I2(\REG.mem_12_6 ), 
            .I3(rd_addr_r[1]), .O(n17406));
    defparam n17403_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_r_5__I_0_123_i1_3_lut (.I0(\wr_addr_r[0] ), .I1(\wr_addr_p1_w[0] ), 
            .I2(wr_fifo_en_w), .I3(GND_net), .O(wr_addr_nxt_c[0]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_5__I_0_123_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15107 (.I0(rd_addr_r[1]), .I1(n15528), 
            .I2(n15529), .I3(rd_addr_r[2]), .O(n17397));
    defparam rd_addr_r_1__bdd_4_lut_15107.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14478 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_7 ), 
            .I2(\REG.mem_3_7 ), .I3(rd_addr_r[1]), .O(n16689));
    defparam rd_addr_r_0__bdd_4_lut_14478.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut (.I0(wp_sync2_r[5]), .I1(wp_sync2_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4962));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n16689_bdd_4_lut (.I0(n16689), .I1(\REG.mem_1_7 ), .I2(\REG.mem_0_7 ), 
            .I3(rd_addr_r[1]), .O(n16692));
    defparam n16689_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14473 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_18 ), 
            .I2(\REG.mem_23_18 ), .I3(rd_addr_r[1]), .O(n16683));
    defparam rd_addr_r_0__bdd_4_lut_14473.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_r_5__I_0_128_7_lut (.I0(GND_net), .I1(\wr_addr_r[5] ), 
            .I2(GND_net), .I3(n13722), .O(wr_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n16683_bdd_4_lut (.I0(n16683), .I1(\REG.mem_21_18 ), .I2(\REG.mem_20_18 ), 
            .I3(rd_addr_r[1]), .O(n16686));
    defparam n16683_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_88 (.I0(wp_sync2_r[2]), .I1(wp_sync_w[3]), .I2(GND_net), 
            .I3(GND_net), .O(wp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_88.LUT_INIT = 16'h6666;
    SB_LUT4 n17397_bdd_4_lut (.I0(n17397), .I1(n15514), .I2(n15513), .I3(rd_addr_r[2]), 
            .O(n17400));
    defparam n17397_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5038_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_28_4 ), .O(n6537));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5038_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_4_lut (.I0(wp_sync2_r[5]), .I1(rd_addr_p1_w[1]), .I2(rd_addr_p1_w[5]), 
            .I3(wp_sync_w[1]), .O(n8_adj_1387));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i5037_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_28_3 ), .O(n6536));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5037_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut (.I0(rd_addr_p1_w[2]), .I1(rd_addr_p1_w[0]), .I2(wp_sync_w[2]), 
            .I3(wp_sync_w[0]), .O(n7_adj_1388));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i1_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut (.I0(rd_addr_p1_w[3]), .I1(rd_addr_p1_w[4]), .I2(wp_sync_w[3]), 
            .I3(n4962), .O(n9));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 n16179_bdd_4_lut (.I0(n16179), .I1(\REG.mem_21_4 ), .I2(\REG.mem_20_4 ), 
            .I3(rd_addr_r[1]), .O(n16182));
    defparam n16179_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14076 (.I0(rd_addr_r[2]), .I1(n14789), 
            .I2(n14798), .I3(rd_addr_r[3]), .O(n16173));
    defparam rd_addr_r_2__bdd_4_lut_14076.LUT_INIT = 16'he4aa;
    SB_LUT4 i5036_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_28_2 ), .O(n6535));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5036_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5035_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_28_1 ), .O(n6534));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5035_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12505_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_r[2]), .I2(wp_sync_w[0]), 
            .I3(wp_sync_w[2]), .O(n14625));
    defparam i12505_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i5034_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_28_0 ), .O(n6533));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5034_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16173_bdd_4_lut (.I0(n16173), .I1(n14777), .I2(n15251), .I3(rd_addr_r[3]), 
            .O(n16176));
    defparam n16173_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12548_4_lut (.I0(rd_addr_r[3]), .I1(rd_addr_r[1]), .I2(wp_sync_w[3]), 
            .I3(wp_sync_w[1]), .O(n14670));
    defparam i12548_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14066 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_24 ), 
            .I2(\REG.mem_15_24 ), .I3(rd_addr_r[1]), .O(n16185));
    defparam rd_addr_r_0__bdd_4_lut_14066.LUT_INIT = 16'he4aa;
    SB_LUT4 i4294_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_4_28 ), .O(n5793));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4294_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_3_lut (.I0(n9), .I1(n7_adj_1388), .I2(n8_adj_1387), .I3(GND_net), 
            .O(n13865));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14568 (.I0(rd_addr_r[3]), .I1(n16656), 
            .I2(n15058), .I3(rd_addr_r[4]), .O(n16671));
    defparam rd_addr_r_3__bdd_4_lut_14568.LUT_INIT = 16'he4aa;
    SB_LUT4 i12583_4_lut (.I0(n14670), .I1(rd_addr_r[4]), .I2(n14625), 
            .I3(n4962), .O(n14706));
    defparam i12583_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 n16671_bdd_4_lut (.I0(n16671), .I1(n15886), .I2(n15885), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[26]));
    defparam n16671_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4293_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_4_27 ), .O(n5792));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4293_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i20_2_lut_3_lut_4_lut (.I0(n7_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n20));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i20_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i4292_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_4_26 ), .O(n5791));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4292_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1103_1104 (.Q(\REG.mem_11_3 ), .C(FIFO_CLK_c), .D(n5992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1100_1101 (.Q(\REG.mem_11_2 ), .C(FIFO_CLK_c), .D(n5991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1097_1098 (.Q(\REG.mem_11_1 ), .C(FIFO_CLK_c), .D(n5990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i13065_3_lut (.I0(n17370), .I1(n16788), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15189));
    defparam i13065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i21_2_lut_3_lut_4_lut (.I0(n7_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[2]), .O(n21));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i21_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 wr_addr_r_5__I_0_128_6_lut (.I0(GND_net), .I1(wr_addr_r[4]), 
            .I2(GND_net), .I3(n13721), .O(wr_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_5__I_0_128_6 (.CI(n13721), .I0(wr_addr_r[4]), .I1(GND_net), 
            .CO(n13722));
    SB_LUT4 i4681_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_16_31 ), .O(n6180));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4681_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14459 (.I0(rd_addr_r[3]), .I1(n16566), 
            .I2(n14968), .I3(rd_addr_r[4]), .O(n16665));
    defparam rd_addr_r_3__bdd_4_lut_14459.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_r_5__I_0_128_5_lut (.I0(GND_net), .I1(wr_addr_r[3]), 
            .I2(GND_net), .I3(n13720), .O(wr_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_5__I_0_128_5 (.CI(n13720), .I0(wr_addr_r[3]), .I1(GND_net), 
            .CO(n13721));
    SB_LUT4 i4680_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_16_30 ), .O(n6179));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4680_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4679_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_16_29 ), .O(n6178));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4679_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_r_5__I_0_128_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(GND_net), .I3(n13719), .O(wr_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_5__I_0_128_4 (.CI(n13719), .I0(wr_addr_r[2]), .I1(GND_net), 
            .CO(n13720));
    SB_LUT4 i2_3_lut (.I0(rp_sync2_r[3]), .I1(rp_sync2_r[4]), .I2(rp_sync2_r[5]), 
            .I3(GND_net), .O(rp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i2_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15062 (.I0(rd_addr_r[1]), .I1(n15087), 
            .I2(n15088), .I3(rd_addr_r[2]), .O(n17385));
    defparam rd_addr_r_1__bdd_4_lut_15062.LUT_INIT = 16'he4aa;
    SB_LUT4 i4678_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_16_28 ), .O(n6177));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4678_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_addr_r_5__I_0_128_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), 
            .I2(GND_net), .I3(n13718), .O(wr_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_89 (.I0(rp_sync2_r[2]), .I1(rp_sync_w[3]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_adj_89.LUT_INIT = 16'h6666;
    SB_LUT4 rp_sync2_r_5__I_0_124_i1_2_lut (.I0(rp_sync2_r[4]), .I1(rp_sync2_r[5]), 
            .I2(GND_net), .I3(GND_net), .O(rp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam rp_sync2_r_5__I_0_124_i1_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 n16665_bdd_4_lut (.I0(n16665), .I1(n14962), .I2(n16560), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[24]));
    defparam n16665_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17385_bdd_4_lut (.I0(n17385), .I1(n15073), .I2(n15072), .I3(rd_addr_r[2]), 
            .O(n15205));
    defparam n17385_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12527_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[4]), .I2(rp_sync_w[1]), 
            .I3(rp_sync_w[4]), .O(n14649));
    defparam i12527_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14454 (.I0(rd_addr_r[3]), .I1(n16650), 
            .I2(n15055), .I3(rd_addr_r[4]), .O(n16659));
    defparam rd_addr_r_3__bdd_4_lut_14454.LUT_INIT = 16'he4aa;
    SB_LUT4 i4677_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_16_27 ), .O(n6176));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4677_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4676_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_16_26 ), .O(n6175));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4676_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12541_4_lut (.I0(wr_addr_r[3]), .I1(\wr_addr_r[0] ), .I2(rp_sync_w[3]), 
            .I3(rp_sync_w[0]), .O(n14663));
    defparam i12541_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i2_4_lut_adj_90 (.I0(wr_addr_p1_w[2]), .I1(wr_addr_p1_w[5]), 
            .I2(rp_sync_w[2]), .I3(rp_sync2_r[5]), .O(n8_adj_1389));
    defparam i2_4_lut_adj_90.LUT_INIT = 16'h1248;
    SB_LUT4 n16659_bdd_4_lut (.I0(n16659), .I1(n15052), .I2(n16644), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[12]));
    defparam n16659_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12473_4_lut (.I0(wr_addr_p1_w[3]), .I1(\wr_addr_p1_w[0] ), 
            .I2(rp_sync_w[3]), .I3(rp_sync_w[0]), .O(n14593));
    defparam i12473_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14508 (.I0(rd_addr_r[1]), .I1(n15492), 
            .I2(n15493), .I3(rd_addr_r[2]), .O(n16653));
    defparam rd_addr_r_1__bdd_4_lut_14508.LUT_INIT = 16'he4aa;
    SB_LUT4 n16233_bdd_4_lut (.I0(n16233), .I1(n14906), .I2(n14903), .I3(rd_addr_r[3]), 
            .O(n16236));
    defparam n16233_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16653_bdd_4_lut (.I0(n16653), .I1(n15697), .I2(n15696), .I3(rd_addr_r[2]), 
            .O(n16656));
    defparam n16653_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12493_4_lut (.I0(wr_addr_p1_w[4]), .I1(wr_addr_p1_w[1]), .I2(rp_sync_w[4]), 
            .I3(rp_sync_w[1]), .O(n14613));
    defparam i12493_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i12581_4_lut (.I0(n14663), .I1(wr_addr_r[2]), .I2(n14649), 
            .I3(rp_sync_w[2]), .O(n14704));
    defparam i12581_4_lut.LUT_INIT = 16'hfefb;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14444 (.I0(rd_addr_r[1]), .I1(n15036), 
            .I2(n15037), .I3(rd_addr_r[2]), .O(n16647));
    defparam rd_addr_r_1__bdd_4_lut_14444.LUT_INIT = 16'he4aa;
    SB_LUT4 i13909_3_lut (.I0(n14613), .I1(n14593), .I2(n8_adj_1389), 
            .I3(GND_net), .O(n15904));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam i13909_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 full_nxt_c_I_10_4_lut (.I0(n15904), .I1(n14704), .I2(dc32_fifo_full), 
            .I3(DEBUG_5_c), .O(full_nxt_c_N_633));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam full_nxt_c_I_10_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 rd_addr_r_5__I_0_i2_3_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1_w[1]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_5__N_573[1] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_5__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n16647_bdd_4_lut (.I0(n16647), .I1(n15031), .I2(n15030), .I3(rd_addr_r[2]), 
            .O(n16650));
    defparam n16647_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i32_2_lut (.I0(n16), .I1(wr_addr_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4291_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_4_25 ), .O(n5790));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4291_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14439 (.I0(rd_addr_r[1]), .I1(n15024), 
            .I2(n15025), .I3(rd_addr_r[2]), .O(n16641));
    defparam rd_addr_r_1__bdd_4_lut_14439.LUT_INIT = 16'he4aa;
    SB_LUT4 n16641_bdd_4_lut (.I0(n16641), .I1(n15019), .I2(n15018), .I3(rd_addr_r[2]), 
            .O(n16644));
    defparam n16641_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14449 (.I0(rd_addr_r[3]), .I1(n16632), 
            .I2(n15022), .I3(rd_addr_r[4]), .O(n16635));
    defparam rd_addr_r_3__bdd_4_lut_14449.LUT_INIT = 16'he4aa;
    SB_LUT4 i4675_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_16_25 ), .O(n6174));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4675_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4674_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_16_24 ), .O(n6173));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4674_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4673_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_16_23 ), .O(n6172));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4673_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4672_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_16_22 ), .O(n6171));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4672_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4290_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_4_24 ), .O(n5789));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4290_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4671_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_16_21 ), .O(n6170));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4671_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4289_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_4_23 ), .O(n5788));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4289_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16635_bdd_4_lut (.I0(n16635), .I1(n15016), .I2(n16620), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[0]));
    defparam n16635_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4670_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_16_20 ), .O(n6169));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4670_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14110 (.I0(rd_addr_r[1]), .I1(n14931), 
            .I2(n14932), .I3(rd_addr_r[2]), .O(n16191));
    defparam rd_addr_r_1__bdd_4_lut_14110.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14434 (.I0(rd_addr_r[1]), .I1(n14991), 
            .I2(n14992), .I3(rd_addr_r[2]), .O(n16629));
    defparam rd_addr_r_1__bdd_4_lut_14434.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14071 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_29 ), 
            .I2(\REG.mem_11_29 ), .I3(rd_addr_r[1]), .O(n16197));
    defparam rd_addr_r_0__bdd_4_lut_14071.LUT_INIT = 16'he4aa;
    SB_LUT4 n16629_bdd_4_lut (.I0(n16629), .I1(n14983), .I2(n14982), .I3(rd_addr_r[2]), 
            .O(n16632));
    defparam n16629_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4669_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_16_19 ), .O(n6168));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4669_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4668_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_16_18 ), .O(n6167));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4668_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15067 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_14 ), 
            .I2(\REG.mem_19_14 ), .I3(rd_addr_r[1]), .O(n17367));
    defparam rd_addr_r_0__bdd_4_lut_15067.LUT_INIT = 16'he4aa;
    SB_LUT4 i4667_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_16_17 ), .O(n6166));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4667_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14429 (.I0(rd_addr_r[3]), .I1(n15138), 
            .I2(n15139), .I3(rd_addr_r[4]), .O(n16623));
    defparam rd_addr_r_3__bdd_4_lut_14429.LUT_INIT = 16'he4aa;
    SB_LUT4 i4666_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_16_16 ), .O(n6165));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4666_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4288_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_4_22 ), .O(n5787));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4288_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4287_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_4_21 ), .O(n5786));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4287_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13308_3_lut (.I0(\REG.mem_24_7 ), .I1(\REG.mem_25_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15432));
    defparam i13308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4233_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_2_31 ), .O(n5732));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4233_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13309_3_lut (.I0(\REG.mem_26_7 ), .I1(\REG.mem_27_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15433));
    defparam i13309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4232_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_2_30 ), .O(n5731));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4232_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4665_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_16_15 ), .O(n6164));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4665_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13348_3_lut (.I0(\REG.mem_30_7 ), .I1(\REG.mem_31_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15472));
    defparam i13348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13347_3_lut (.I0(\REG.mem_28_7 ), .I1(\REG.mem_29_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15471));
    defparam i13347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_91 (.I0(dc32_fifo_empty), .I1(FT_OE_N_496), .I2(GND_net), 
            .I3(GND_net), .O(n12_adj_3));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i1_2_lut_adj_91.LUT_INIT = 16'hdddd;
    SB_LUT4 i4231_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_2_29 ), .O(n5730));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4231_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4286_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_4_20 ), .O(n5785));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4286_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4664_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_16_14 ), .O(n6163));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4664_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4230_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_2_28 ), .O(n5729));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4230_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4229_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_2_27 ), .O(n5728));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4229_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4663_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_16_13 ), .O(n6162));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4663_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4228_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_2_26 ), .O(n5727));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4228_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4227_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_2_25 ), .O(n5726));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4227_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4226_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_2_24 ), .O(n5725));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4226_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4662_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_16_12 ), .O(n6161));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4662_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4225_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_2_23 ), .O(n5724));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4225_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4224_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_2_22 ), .O(n5723));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4224_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4223_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_2_21 ), .O(n5722));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4223_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4285_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_4_19 ), .O(n5784));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4285_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4661_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_16_11 ), .O(n6160));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4661_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4284_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_4_18 ), .O(n5783));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4284_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4222_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_2_20 ), .O(n5721));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4222_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4660_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_16_10 ), .O(n6159));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4660_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4221_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_2_19 ), .O(n5720));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4221_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4220_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_2_18 ), .O(n5719));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4220_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4219_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_2_17 ), .O(n5718));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4219_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17367_bdd_4_lut (.I0(n17367), .I1(\REG.mem_17_14 ), .I2(\REG.mem_16_14 ), 
            .I3(rd_addr_r[1]), .O(n17370));
    defparam n17367_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4659_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_16_9 ), .O(n6158));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4659_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4218_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_2_16 ), .O(n5717));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4218_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15037 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_2 ), 
            .I2(\REG.mem_15_2 ), .I3(rd_addr_r[1]), .O(n17361));
    defparam rd_addr_r_0__bdd_4_lut_15037.LUT_INIT = 16'he4aa;
    SB_LUT4 i4217_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_2_15 ), .O(n5716));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4217_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4283_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_4_17 ), .O(n5782));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4283_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4658_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_16_8 ), .O(n6157));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4658_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4657_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_16_7 ), .O(n6156));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4657_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4216_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_2_14 ), .O(n5715));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4216_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4656_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_16_6 ), .O(n6155));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4656_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4655_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_16_5 ), .O(n6154));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4655_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4215_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_2_13 ), .O(n5714));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4215_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4654_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_16_4 ), .O(n6153));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4654_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4214_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_2_12 ), .O(n5713));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4214_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4653_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_16_3 ), .O(n6152));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4653_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4282_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_4_16 ), .O(n5781));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4282_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4213_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_2_11 ), .O(n5712));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4213_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4212_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_2_10 ), .O(n5711));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4212_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4211_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_2_9 ), .O(n5710));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4211_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4210_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_2_8 ), .O(n5709));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4210_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4652_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_16_2 ), .O(n6151));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4652_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16623_bdd_4_lut (.I0(n16623), .I1(n15013), .I2(n16614), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[13]));
    defparam n16623_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4208_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_2_6 ), .O(n5707));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4208_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4186_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_2_4 ), .O(n5685));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4186_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17361_bdd_4_lut (.I0(n17361), .I1(\REG.mem_13_2 ), .I2(\REG.mem_12_2 ), 
            .I3(rd_addr_r[1]), .O(n15692));
    defparam n17361_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4188_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_2_0 ), .O(n5687));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4188_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4281_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_4_15 ), .O(n5780));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4281_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14424 (.I0(rd_addr_r[1]), .I1(n14802), 
            .I2(n14803), .I3(rd_addr_r[2]), .O(n16617));
    defparam rd_addr_r_1__bdd_4_lut_14424.LUT_INIT = 16'he4aa;
    SB_LUT4 n16617_bdd_4_lut (.I0(n16617), .I1(n15895), .I2(n15894), .I3(rd_addr_r[2]), 
            .O(n16620));
    defparam n16617_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4209_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_2_7 ), .O(n5708));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4209_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15052 (.I0(rd_addr_r[1]), .I1(n15507), 
            .I2(n15508), .I3(rd_addr_r[2]), .O(n17355));
    defparam rd_addr_r_1__bdd_4_lut_15052.LUT_INIT = 16'he4aa;
    SB_LUT4 n17355_bdd_4_lut (.I0(n17355), .I1(n15628), .I2(n15627), .I3(rd_addr_r[2]), 
            .O(n17358));
    defparam n17355_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4182_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_2_5 ), .O(n5681));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4182_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4100_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_2_3 ), .O(n5599));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4100_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4124_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_2_1 ), .O(n5623));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4124_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_92 (.I0(dc32_fifo_empty), .I1(dc32_fifo_read_enable), 
            .I2(GND_net), .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i1_2_lut_adj_92.LUT_INIT = 16'h4444;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14414 (.I0(rd_addr_r[1]), .I1(n14979), 
            .I2(n14980), .I3(rd_addr_r[2]), .O(n16611));
    defparam rd_addr_r_1__bdd_4_lut_14414.LUT_INIT = 16'he4aa;
    SB_LUT4 i4651_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_16_1 ), .O(n6150));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4651_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4104_3_lut_4_lut (.I0(n25_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_2_2 ), .O(n5603));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4104_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4650_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_16_0 ), .O(n6149));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4650_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4280_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_4_14 ), .O(n5779));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4280_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16611_bdd_4_lut (.I0(n16611), .I1(n14977), .I2(n14976), .I3(rd_addr_r[2]), 
            .O(n16614));
    defparam n16611_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4279_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_4_13 ), .O(n5778));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4279_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4553_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_12_31 ), .O(n6052));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4553_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4278_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_4_12 ), .O(n5777));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4278_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4277_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_4_11 ), .O(n5776));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4277_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4552_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_12_30 ), .O(n6051));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4552_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4551_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_12_29 ), .O(n6050));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4551_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4550_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_12_28 ), .O(n6049));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4550_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1094_1095 (.Q(\REG.mem_11_0 ), .C(FIFO_CLK_c), .D(n5989));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14061 (.I0(rd_addr_r[1]), .I1(n15222), 
            .I2(n15223), .I3(rd_addr_r[2]), .O(n16161));
    defparam rd_addr_r_1__bdd_4_lut_14061.LUT_INIT = 16'he4aa;
    SB_DFF i1091_1092 (.Q(\REG.mem_10_31 ), .C(FIFO_CLK_c), .D(n5988));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1088_1089 (.Q(\REG.mem_10_30 ), .C(FIFO_CLK_c), .D(n5987));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1085_1086 (.Q(\REG.mem_10_29 ), .C(FIFO_CLK_c), .D(n5986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1082_1083 (.Q(\REG.mem_10_28 ), .C(FIFO_CLK_c), .D(n5985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1079_1080 (.Q(\REG.mem_10_27 ), .C(FIFO_CLK_c), .D(n5984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1076_1077 (.Q(\REG.mem_10_26 ), .C(FIFO_CLK_c), .D(n5983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1073_1074 (.Q(\REG.mem_10_25 ), .C(FIFO_CLK_c), .D(n5982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1070_1071 (.Q(\REG.mem_10_24 ), .C(FIFO_CLK_c), .D(n5981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1067_1068 (.Q(\REG.mem_10_23 ), .C(FIFO_CLK_c), .D(n5980));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1064_1065 (.Q(\REG.mem_10_22 ), .C(FIFO_CLK_c), .D(n5979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1061_1062 (.Q(\REG.mem_10_21 ), .C(FIFO_CLK_c), .D(n5978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1058_1059 (.Q(\REG.mem_10_20 ), .C(FIFO_CLK_c), .D(n5977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1055_1056 (.Q(\REG.mem_10_19 ), .C(FIFO_CLK_c), .D(n5976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1052_1053 (.Q(\REG.mem_10_18 ), .C(FIFO_CLK_c), .D(n5975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1049_1050 (.Q(\REG.mem_10_17 ), .C(FIFO_CLK_c), .D(n5974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1046_1047 (.Q(\REG.mem_10_16 ), .C(FIFO_CLK_c), .D(n5973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1043_1044 (.Q(\REG.mem_10_15 ), .C(FIFO_CLK_c), .D(n5972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1040_1041 (.Q(\REG.mem_10_14 ), .C(FIFO_CLK_c), .D(n5971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1037_1038 (.Q(\REG.mem_10_13 ), .C(FIFO_CLK_c), .D(n5970));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1034_1035 (.Q(\REG.mem_10_12 ), .C(FIFO_CLK_c), .D(n5969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1031_1032 (.Q(\REG.mem_10_11 ), .C(FIFO_CLK_c), .D(n5968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1028_1029 (.Q(\REG.mem_10_10 ), .C(FIFO_CLK_c), .D(n5967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1025_1026 (.Q(\REG.mem_10_9 ), .C(FIFO_CLK_c), .D(n5966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1022_1023 (.Q(\REG.mem_10_8 ), .C(FIFO_CLK_c), .D(n5965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1019_1020 (.Q(\REG.mem_10_7 ), .C(FIFO_CLK_c), .D(n5964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1016_1017 (.Q(\REG.mem_10_6 ), .C(FIFO_CLK_c), .D(n5963));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1013_1014 (.Q(\REG.mem_10_5 ), .C(FIFO_CLK_c), .D(n5962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1010_1011 (.Q(\REG.mem_10_4 ), .C(FIFO_CLK_c), .D(n5961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1007_1008 (.Q(\REG.mem_10_3 ), .C(FIFO_CLK_c), .D(n5960));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1004_1005 (.Q(\REG.mem_10_2 ), .C(FIFO_CLK_c), .D(n5959));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1001_1002 (.Q(\REG.mem_10_1 ), .C(FIFO_CLK_c), .D(n5958));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i998_999 (.Q(\REG.mem_10_0 ), .C(FIFO_CLK_c), .D(n5957));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i995_996 (.Q(\REG.mem_9_31 ), .C(FIFO_CLK_c), .D(n5956));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i992_993 (.Q(\REG.mem_9_30 ), .C(FIFO_CLK_c), .D(n5955));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i989_990 (.Q(\REG.mem_9_29 ), .C(FIFO_CLK_c), .D(n5954));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i986_987 (.Q(\REG.mem_9_28 ), .C(FIFO_CLK_c), .D(n5953));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i983_984 (.Q(\REG.mem_9_27 ), .C(FIFO_CLK_c), .D(n5952));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i980_981 (.Q(\REG.mem_9_26 ), .C(FIFO_CLK_c), .D(n5951));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i977_978 (.Q(\REG.mem_9_25 ), .C(FIFO_CLK_c), .D(n5950));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i974_975 (.Q(\REG.mem_9_24 ), .C(FIFO_CLK_c), .D(n5949));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i971_972 (.Q(\REG.mem_9_23 ), .C(FIFO_CLK_c), .D(n5948));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i968_969 (.Q(\REG.mem_9_22 ), .C(FIFO_CLK_c), .D(n5947));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i965_966 (.Q(\REG.mem_9_21 ), .C(FIFO_CLK_c), .D(n5946));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i962_963 (.Q(\REG.mem_9_20 ), .C(FIFO_CLK_c), .D(n5945));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i959_960 (.Q(\REG.mem_9_19 ), .C(FIFO_CLK_c), .D(n5944));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i956_957 (.Q(\REG.mem_9_18 ), .C(FIFO_CLK_c), .D(n5943));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i953_954 (.Q(\REG.mem_9_17 ), .C(FIFO_CLK_c), .D(n5942));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i950_951 (.Q(\REG.mem_9_16 ), .C(FIFO_CLK_c), .D(n5941));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i947_948 (.Q(\REG.mem_9_15 ), .C(FIFO_CLK_c), .D(n5940));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i944_945 (.Q(\REG.mem_9_14 ), .C(FIFO_CLK_c), .D(n5939));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i941_942 (.Q(\REG.mem_9_13 ), .C(FIFO_CLK_c), .D(n5938));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i938_939 (.Q(\REG.mem_9_12 ), .C(FIFO_CLK_c), .D(n5937));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i935_936 (.Q(\REG.mem_9_11 ), .C(FIFO_CLK_c), .D(n5936));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i932_933 (.Q(\REG.mem_9_10 ), .C(FIFO_CLK_c), .D(n5935));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i929_930 (.Q(\REG.mem_9_9 ), .C(FIFO_CLK_c), .D(n5934));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i926_927 (.Q(\REG.mem_9_8 ), .C(FIFO_CLK_c), .D(n5933));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i923_924 (.Q(\REG.mem_9_7 ), .C(FIFO_CLK_c), .D(n5932));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i920_921 (.Q(\REG.mem_9_6 ), .C(FIFO_CLK_c), .D(n5931));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i917_918 (.Q(\REG.mem_9_5 ), .C(FIFO_CLK_c), .D(n5930));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i914_915 (.Q(\REG.mem_9_4 ), .C(FIFO_CLK_c), .D(n5929));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i911_912 (.Q(\REG.mem_9_3 ), .C(FIFO_CLK_c), .D(n5928));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i908_909 (.Q(\REG.mem_9_2 ), .C(FIFO_CLK_c), .D(n5927));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i905_906 (.Q(\REG.mem_9_1 ), .C(FIFO_CLK_c), .D(n5926));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i902_903 (.Q(\REG.mem_9_0 ), .C(FIFO_CLK_c), .D(n5925));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i899_900 (.Q(\REG.mem_8_31 ), .C(FIFO_CLK_c), .D(n5924));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i896_897 (.Q(\REG.mem_8_30 ), .C(FIFO_CLK_c), .D(n5923));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i893_894 (.Q(\REG.mem_8_29 ), .C(FIFO_CLK_c), .D(n5922));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i890_891 (.Q(\REG.mem_8_28 ), .C(FIFO_CLK_c), .D(n5921));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i887_888 (.Q(\REG.mem_8_27 ), .C(FIFO_CLK_c), .D(n5920));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i884_885 (.Q(\REG.mem_8_26 ), .C(FIFO_CLK_c), .D(n5919));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i881_882 (.Q(\REG.mem_8_25 ), .C(FIFO_CLK_c), .D(n5918));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i878_879 (.Q(\REG.mem_8_24 ), .C(FIFO_CLK_c), .D(n5917));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i875_876 (.Q(\REG.mem_8_23 ), .C(FIFO_CLK_c), .D(n5916));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i872_873 (.Q(\REG.mem_8_22 ), .C(FIFO_CLK_c), .D(n5915));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i869_870 (.Q(\REG.mem_8_21 ), .C(FIFO_CLK_c), .D(n5914));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i866_867 (.Q(\REG.mem_8_20 ), .C(FIFO_CLK_c), .D(n5913));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i863_864 (.Q(\REG.mem_8_19 ), .C(FIFO_CLK_c), .D(n5912));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i860_861 (.Q(\REG.mem_8_18 ), .C(FIFO_CLK_c), .D(n5911));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i857_858 (.Q(\REG.mem_8_17 ), .C(FIFO_CLK_c), .D(n5910));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i854_855 (.Q(\REG.mem_8_16 ), .C(FIFO_CLK_c), .D(n5909));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i851_852 (.Q(\REG.mem_8_15 ), .C(FIFO_CLK_c), .D(n5908));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i848_849 (.Q(\REG.mem_8_14 ), .C(FIFO_CLK_c), .D(n5907));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i845_846 (.Q(\REG.mem_8_13 ), .C(FIFO_CLK_c), .D(n5906));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i842_843 (.Q(\REG.mem_8_12 ), .C(FIFO_CLK_c), .D(n5905));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i839_840 (.Q(\REG.mem_8_11 ), .C(FIFO_CLK_c), .D(n5904));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i836_837 (.Q(\REG.mem_8_10 ), .C(FIFO_CLK_c), .D(n5903));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i833_834 (.Q(\REG.mem_8_9 ), .C(FIFO_CLK_c), .D(n5902));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i830_831 (.Q(\REG.mem_8_8 ), .C(FIFO_CLK_c), .D(n5901));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i827_828 (.Q(\REG.mem_8_7 ), .C(FIFO_CLK_c), .D(n5900));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i824_825 (.Q(\REG.mem_8_6 ), .C(FIFO_CLK_c), .D(n5899));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i821_822 (.Q(\REG.mem_8_5 ), .C(FIFO_CLK_c), .D(n5898));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i818_819 (.Q(\REG.mem_8_4 ), .C(FIFO_CLK_c), .D(n5897));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i815_816 (.Q(\REG.mem_8_3 ), .C(FIFO_CLK_c), .D(n5896));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i812_813 (.Q(\REG.mem_8_2 ), .C(FIFO_CLK_c), .D(n5895));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i809_810 (.Q(\REG.mem_8_1 ), .C(FIFO_CLK_c), .D(n5894));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i806_807 (.Q(\REG.mem_8_0 ), .C(FIFO_CLK_c), .D(n5893));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i803_804 (.Q(\REG.mem_7_31 ), .C(FIFO_CLK_c), .D(n5892));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i800_801 (.Q(\REG.mem_7_30 ), .C(FIFO_CLK_c), .D(n5891));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i797_798 (.Q(\REG.mem_7_29 ), .C(FIFO_CLK_c), .D(n5890));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i794_795 (.Q(\REG.mem_7_28 ), .C(FIFO_CLK_c), .D(n5889));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i791_792 (.Q(\REG.mem_7_27 ), .C(FIFO_CLK_c), .D(n5888));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i788_789 (.Q(\REG.mem_7_26 ), .C(FIFO_CLK_c), .D(n5887));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i785_786 (.Q(\REG.mem_7_25 ), .C(FIFO_CLK_c), .D(n5886));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i782_783 (.Q(\REG.mem_7_24 ), .C(FIFO_CLK_c), .D(n5885));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i779_780 (.Q(\REG.mem_7_23 ), .C(FIFO_CLK_c), .D(n5884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i776_777 (.Q(\REG.mem_7_22 ), .C(FIFO_CLK_c), .D(n5883));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i773_774 (.Q(\REG.mem_7_21 ), .C(FIFO_CLK_c), .D(n5882));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i770_771 (.Q(\REG.mem_7_20 ), .C(FIFO_CLK_c), .D(n5881));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i767_768 (.Q(\REG.mem_7_19 ), .C(FIFO_CLK_c), .D(n5880));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i764_765 (.Q(\REG.mem_7_18 ), .C(FIFO_CLK_c), .D(n5879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i761_762 (.Q(\REG.mem_7_17 ), .C(FIFO_CLK_c), .D(n5878));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i758_759 (.Q(\REG.mem_7_16 ), .C(FIFO_CLK_c), .D(n5877));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i755_756 (.Q(\REG.mem_7_15 ), .C(FIFO_CLK_c), .D(n5876));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i752_753 (.Q(\REG.mem_7_14 ), .C(FIFO_CLK_c), .D(n5875));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i749_750 (.Q(\REG.mem_7_13 ), .C(FIFO_CLK_c), .D(n5874));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i746_747 (.Q(\REG.mem_7_12 ), .C(FIFO_CLK_c), .D(n5873));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i743_744 (.Q(\REG.mem_7_11 ), .C(FIFO_CLK_c), .D(n5872));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i740_741 (.Q(\REG.mem_7_10 ), .C(FIFO_CLK_c), .D(n5871));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i737_738 (.Q(\REG.mem_7_9 ), .C(FIFO_CLK_c), .D(n5870));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i734_735 (.Q(\REG.mem_7_8 ), .C(FIFO_CLK_c), .D(n5869));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i731_732 (.Q(\REG.mem_7_7 ), .C(FIFO_CLK_c), .D(n5868));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i728_729 (.Q(\REG.mem_7_6 ), .C(FIFO_CLK_c), .D(n5867));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i725_726 (.Q(\REG.mem_7_5 ), .C(FIFO_CLK_c), .D(n5866));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i722_723 (.Q(\REG.mem_7_4 ), .C(FIFO_CLK_c), .D(n5865));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i719_720 (.Q(\REG.mem_7_3 ), .C(FIFO_CLK_c), .D(n5864));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i716_717 (.Q(\REG.mem_7_2 ), .C(FIFO_CLK_c), .D(n5863));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i713_714 (.Q(\REG.mem_7_1 ), .C(FIFO_CLK_c), .D(n5862));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i710_711 (.Q(\REG.mem_7_0 ), .C(FIFO_CLK_c), .D(n5861));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i707_708 (.Q(\REG.mem_6_31 ), .C(FIFO_CLK_c), .D(n5860));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i704_705 (.Q(\REG.mem_6_30 ), .C(FIFO_CLK_c), .D(n5859));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i701_702 (.Q(\REG.mem_6_29 ), .C(FIFO_CLK_c), .D(n5858));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i698_699 (.Q(\REG.mem_6_28 ), .C(FIFO_CLK_c), .D(n5857));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i695_696 (.Q(\REG.mem_6_27 ), .C(FIFO_CLK_c), .D(n5856));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i692_693 (.Q(\REG.mem_6_26 ), .C(FIFO_CLK_c), .D(n5855));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i689_690 (.Q(\REG.mem_6_25 ), .C(FIFO_CLK_c), .D(n5854));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i686_687 (.Q(\REG.mem_6_24 ), .C(FIFO_CLK_c), .D(n5853));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i683_684 (.Q(\REG.mem_6_23 ), .C(FIFO_CLK_c), .D(n5852));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i680_681 (.Q(\REG.mem_6_22 ), .C(FIFO_CLK_c), .D(n5851));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4549_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_12_27 ), .O(n6048));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4549_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_3_lut (.I0(dc32_fifo_almost_empty), .I1(\state[3] ), .I2(n4843), 
            .I3(GND_net), .O(n1224));   // src/fifo_dc_32_lut_gen.v(669[37] 672[40])
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i4548_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_12_26 ), .O(n6047));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4548_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4276_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_4_10 ), .O(n5775));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4276_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14419 (.I0(rd_addr_r[3]), .I1(n15189), 
            .I2(n15190), .I3(rd_addr_r[4]), .O(n16605));
    defparam rd_addr_r_3__bdd_4_lut_14419.LUT_INIT = 16'he4aa;
    SB_DFF i677_678 (.Q(\REG.mem_6_21 ), .C(FIFO_CLK_c), .D(n5850));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i674_675 (.Q(\REG.mem_6_20 ), .C(FIFO_CLK_c), .D(n5849));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i671_672 (.Q(\REG.mem_6_19 ), .C(FIFO_CLK_c), .D(n5848));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i668_669 (.Q(\REG.mem_6_18 ), .C(FIFO_CLK_c), .D(n5847));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i665_666 (.Q(\REG.mem_6_17 ), .C(FIFO_CLK_c), .D(n5846));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i662_663 (.Q(\REG.mem_6_16 ), .C(FIFO_CLK_c), .D(n5845));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i659_660 (.Q(\REG.mem_6_15 ), .C(FIFO_CLK_c), .D(n5844));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i656_657 (.Q(\REG.mem_6_14 ), .C(FIFO_CLK_c), .D(n5843));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i89_90 (.Q(\REG.mem_0_17 ), .C(FIFO_CLK_c), .D(n5699));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i92_93 (.Q(\REG.mem_0_18 ), .C(FIFO_CLK_c), .D(n5695));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i95_96 (.Q(\REG.mem_0_19 ), .C(FIFO_CLK_c), .D(n5694));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i98_99 (.Q(\REG.mem_0_20 ), .C(FIFO_CLK_c), .D(n5693));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4547_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_12_25 ), .O(n6046));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4547_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16605_bdd_4_lut (.I0(n16605), .I1(n16542), .I2(n16482), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[14]));
    defparam n16605_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i653_654 (.Q(\REG.mem_6_13 ), .C(FIFO_CLK_c), .D(n5842));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i650_651 (.Q(\REG.mem_6_12 ), .C(FIFO_CLK_c), .D(n5841));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i647_648 (.Q(\REG.mem_6_11 ), .C(FIFO_CLK_c), .D(n5840));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i644_645 (.Q(\REG.mem_6_10 ), .C(FIFO_CLK_c), .D(n5839));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i641_642 (.Q(\REG.mem_6_9 ), .C(FIFO_CLK_c), .D(n5838));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i638_639 (.Q(\REG.mem_6_8 ), .C(FIFO_CLK_c), .D(n5837));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i635_636 (.Q(\REG.mem_6_7 ), .C(FIFO_CLK_c), .D(n5836));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i632_633 (.Q(\REG.mem_6_6 ), .C(FIFO_CLK_c), .D(n5835));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i629_630 (.Q(\REG.mem_6_5 ), .C(FIFO_CLK_c), .D(n5834));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i101_102 (.Q(\REG.mem_0_21 ), .C(FIFO_CLK_c), .D(n5689));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i104_105 (.Q(\REG.mem_0_22 ), .C(FIFO_CLK_c), .D(n5688));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i230_231 (.Q(\REG.mem_2_0 ), .C(FIFO_CLK_c), .D(n5687));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i107_108 (.Q(\REG.mem_0_23 ), .C(FIFO_CLK_c), .D(n5686));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i242_243 (.Q(\REG.mem_2_4 ), .C(FIFO_CLK_c), .D(n5685));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i110_111 (.Q(\REG.mem_0_24 ), .C(FIFO_CLK_c), .D(n5684));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i113_114 (.Q(\REG.mem_0_25 ), .C(FIFO_CLK_c), .D(n5683));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i116_117 (.Q(\REG.mem_0_26 ), .C(FIFO_CLK_c), .D(n5682));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i626_627 (.Q(\REG.mem_6_4 ), .C(FIFO_CLK_c), .D(n5833));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4546_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_12_24 ), .O(n6045));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4546_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4545_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_12_23 ), .O(n6044));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4545_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4275_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_4_9 ), .O(n5774));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4275_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4274_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_4_8 ), .O(n5773));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4274_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4273_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_4_7 ), .O(n5772));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4273_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4544_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_12_22 ), .O(n6043));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4544_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4272_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_4_6 ), .O(n5771));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4272_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i245_246 (.Q(\REG.mem_2_5 ), .C(FIFO_CLK_c), .D(n5681));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4207_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_0_11 ), .O(n5706));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4207_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4543_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_12_21 ), .O(n6042));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4543_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4177_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_0_0 ), .O(n5676));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4177_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4180_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_0_28 ), .O(n5679));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4180_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14468 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_4 ), 
            .I2(\REG.mem_11_4 ), .I3(rd_addr_r[1]), .O(n16599));
    defparam rd_addr_r_0__bdd_4_lut_14468.LUT_INIT = 16'he4aa;
    SB_LUT4 n16599_bdd_4_lut (.I0(n16599), .I1(\REG.mem_9_4 ), .I2(\REG.mem_8_4 ), 
            .I3(rd_addr_r[1]), .O(n15314));
    defparam n16599_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4542_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_12_20 ), .O(n6041));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4542_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4181_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_0_27 ), .O(n5680));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4181_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4271_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_4_5 ), .O(n5770));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4271_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4541_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_12_19 ), .O(n6040));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4541_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4183_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_0_26 ), .O(n5682));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4183_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4184_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_0_25 ), .O(n5683));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4184_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4540_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_12_18 ), .O(n6039));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4540_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4185_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_0_24 ), .O(n5684));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4185_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i119_120 (.Q(\REG.mem_0_27 ), .C(FIFO_CLK_c), .D(n5680));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4539_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_12_17 ), .O(n6038));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4539_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4270_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_4_4 ), .O(n5769));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4270_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4187_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_0_23 ), .O(n5686));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4187_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4189_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_0_22 ), .O(n5688));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4189_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4190_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_0_21 ), .O(n5689));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4190_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4194_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_0_20 ), .O(n5693));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4194_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4195_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_0_19 ), .O(n5694));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4195_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14399 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_2 ), 
            .I2(\REG.mem_7_2 ), .I3(rd_addr_r[1]), .O(n16593));
    defparam rd_addr_r_0__bdd_4_lut_14399.LUT_INIT = 16'he4aa;
    SB_LUT4 i4538_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_12_16 ), .O(n6037));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4538_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4196_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_0_18 ), .O(n5695));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4196_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4200_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_0_17 ), .O(n5699));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4200_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4537_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_12_15 ), .O(n6036));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4537_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i623_624 (.Q(\REG.mem_6_3 ), .C(FIFO_CLK_c), .D(n5832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i620_621 (.Q(\REG.mem_6_2 ), .C(FIFO_CLK_c), .D(n5831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n16593_bdd_4_lut (.I0(n16593), .I1(\REG.mem_5_2 ), .I2(\REG.mem_4_2 ), 
            .I3(rd_addr_r[1]), .O(n16596));
    defparam n16593_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4201_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_0_16 ), .O(n5700));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4201_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4269_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_4_3 ), .O(n5768));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4269_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4536_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_12_14 ), .O(n6035));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4536_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4535_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_12_13 ), .O(n6034));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4535_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4534_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_12_12 ), .O(n6033));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4534_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i617_618 (.Q(\REG.mem_6_1 ), .C(FIFO_CLK_c), .D(n5830));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_15082 (.I0(rd_addr_r[3]), .I1(n16830), 
            .I2(n15205), .I3(rd_addr_r[4]), .O(n17319));
    defparam rd_addr_r_3__bdd_4_lut_15082.LUT_INIT = 16'he4aa;
    SB_LUT4 i4533_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_12_11 ), .O(n6032));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4533_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4202_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_0_15 ), .O(n5701));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4202_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i614_615 (.Q(\REG.mem_6_0 ), .C(FIFO_CLK_c), .D(n5829));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4268_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_4_2 ), .O(n5767));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4268_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4267_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_4_1 ), .O(n5766));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4267_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4532_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_12_10 ), .O(n6031));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4532_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4203_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_0_14 ), .O(n5702));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4203_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4205_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_0_13 ), .O(n5704));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4205_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14394 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_7 ), 
            .I2(\REG.mem_15_7 ), .I3(rd_addr_r[1]), .O(n16587));
    defparam rd_addr_r_0__bdd_4_lut_14394.LUT_INIT = 16'he4aa;
    SB_DFF i611_612 (.Q(\REG.mem_5_31 ), .C(FIFO_CLK_c), .D(n5828));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4531_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_12_9 ), .O(n6030));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4531_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4530_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_12_8 ), .O(n6029));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4530_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4529_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_12_7 ), .O(n6028));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4529_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4206_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_0_12 ), .O(n5705));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4206_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4122_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_0_10 ), .O(n5621));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4122_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4123_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_0_9 ), .O(n5622));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4123_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4127_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_0_8 ), .O(n5626));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4127_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16587_bdd_4_lut (.I0(n16587), .I1(\REG.mem_13_7 ), .I2(\REG.mem_12_7 ), 
            .I3(rd_addr_r[1]), .O(n16590));
    defparam n16587_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4528_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_12_6 ), .O(n6027));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4528_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i122_123 (.Q(\REG.mem_0_28 ), .C(FIFO_CLK_c), .D(n5679));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4128_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_0_7 ), .O(n5627));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4128_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4527_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_12_5 ), .O(n6026));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4527_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4133_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_0_6 ), .O(n5632));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4133_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i608_609 (.Q(\REG.mem_5_30 ), .C(FIFO_CLK_c), .D(n5827));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4526_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_12_4 ), .O(n6025));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4526_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i125_126 (.Q(\REG.mem_0_29 ), .C(FIFO_CLK_c), .D(n5678));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4134_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_0_5 ), .O(n5633));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4134_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4164_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_0_4 ), .O(n5663));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4164_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4170_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_0_3 ), .O(n5669));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4170_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4266_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_4_0 ), .O(n5765));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4266_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4172_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_0_31 ), .O(n5671));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4172_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4525_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_12_3 ), .O(n6024));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4525_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4173_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_0_2 ), .O(n5672));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4173_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4176_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_0_1 ), .O(n5675));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4176_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i605_606 (.Q(\REG.mem_5_29 ), .C(FIFO_CLK_c), .D(n5826));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14389 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_24 ), 
            .I2(\REG.mem_11_24 ), .I3(rd_addr_r[1]), .O(n16581));
    defparam rd_addr_r_0__bdd_4_lut_14389.LUT_INIT = 16'he4aa;
    SB_DFF i128_129 (.Q(\REG.mem_0_30 ), .C(FIFO_CLK_c), .D(n5677));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4178_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_0_30 ), .O(n5677));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4178_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4179_3_lut_4_lut (.I0(n21), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_0_29 ), .O(n5678));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4179_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i602_603 (.Q(\REG.mem_5_28 ), .C(FIFO_CLK_c), .D(n5825));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4524_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_12_2 ), .O(n6023));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4524_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17319_bdd_4_lut (.I0(n17319), .I1(n15172), .I2(n16782), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[5]));
    defparam n17319_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4523_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_12_1 ), .O(n6022));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4523_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i38_39 (.Q(\REG.mem_0_0 ), .C(FIFO_CLK_c), .D(n5676));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i41_42 (.Q(\REG.mem_0_1 ), .C(FIFO_CLK_c), .D(n5675));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i599_600 (.Q(\REG.mem_5_27 ), .C(FIFO_CLK_c), .D(n5824));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4522_3_lut_4_lut (.I0(n28_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_12_0 ), .O(n6021));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4522_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i596_597 (.Q(\REG.mem_5_26 ), .C(FIFO_CLK_c), .D(n5823));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4649_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_15_31 ), .O(n6148));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4649_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i593_594 (.Q(\REG.mem_5_25 ), .C(FIFO_CLK_c), .D(n5822));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i44_45 (.Q(\REG.mem_0_2 ), .C(FIFO_CLK_c), .D(n5672));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i590_591 (.Q(\REG.mem_5_24 ), .C(FIFO_CLK_c), .D(n5821));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i131_132 (.Q(\REG.mem_0_31 ), .C(FIFO_CLK_c), .D(n5671));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4648_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_15_30 ), .O(n6147));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4648_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i587_588 (.Q(\REG.mem_5_23 ), .C(FIFO_CLK_c), .D(n5820));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n16581_bdd_4_lut (.I0(n16581), .I1(\REG.mem_9_24 ), .I2(\REG.mem_8_24 ), 
            .I3(rd_addr_r[1]), .O(n16584));
    defparam n16581_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4647_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_15_29 ), .O(n6146));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4647_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4585_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_13_31 ), .O(n6084));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4585_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i134_135 (.Q(\REG.mem_1_0 ), .C(FIFO_CLK_c), .D(n5670));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4646_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_15_28 ), .O(n6145));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4646_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i47_48 (.Q(\REG.mem_0_3 ), .C(FIFO_CLK_c), .D(n5669));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i584_585 (.Q(\REG.mem_5_22 ), .C(FIFO_CLK_c), .D(n5819));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i581_582 (.Q(\REG.mem_5_21 ), .C(FIFO_CLK_c), .D(n5818));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i137_138 (.Q(\REG.mem_1_1 ), .C(FIFO_CLK_c), .D(n5668));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4584_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_13_30 ), .O(n6083));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4584_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i140_141 (.Q(\REG.mem_1_2 ), .C(FIFO_CLK_c), .D(n5667));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4583_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_13_29 ), .O(n6082));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4583_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4582_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_13_28 ), .O(n6081));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4582_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i578_579 (.Q(\REG.mem_5_20 ), .C(FIFO_CLK_c), .D(n5817));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i143_144 (.Q(\REG.mem_1_3 ), .C(FIFO_CLK_c), .D(n5666));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i575_576 (.Q(\REG.mem_5_19 ), .C(FIFO_CLK_c), .D(n5816));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i146_147 (.Q(\REG.mem_1_4 ), .C(FIFO_CLK_c), .D(n5665));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i572_573 (.Q(\REG.mem_5_18 ), .C(FIFO_CLK_c), .D(n5815));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4645_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_15_27 ), .O(n6144));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4645_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i50_51 (.Q(\REG.mem_0_4 ), .C(FIFO_CLK_c), .D(n5663));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i569_570 (.Q(\REG.mem_5_17 ), .C(FIFO_CLK_c), .D(n5814));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i566_567 (.Q(\REG.mem_5_16 ), .C(FIFO_CLK_c), .D(n5813));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4581_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_13_27 ), .O(n6080));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4581_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i206_207 (.Q(\REG.mem_1_24 ), .C(FIFO_CLK_c), .D(n5662));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i563_564 (.Q(\REG.mem_5_15 ), .C(FIFO_CLK_c), .D(n5812));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i10_2_lut (.I0(n6_adj_1378), .I1(wr_addr_r[1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i10_2_lut.LUT_INIT = 16'h8888;
    SB_DFF i194_195 (.Q(\REG.mem_1_20 ), .C(FIFO_CLK_c), .D(n5660));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i227_228 (.Q(\REG.mem_1_31 ), .C(FIFO_CLK_c), .D(n5659));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i560_561 (.Q(\REG.mem_5_14 ), .C(FIFO_CLK_c), .D(n5811));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i557_558 (.Q(\REG.mem_5_13 ), .C(FIFO_CLK_c), .D(n5810));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14384 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_29 ), 
            .I2(\REG.mem_15_29 ), .I3(rd_addr_r[1]), .O(n16575));
    defparam rd_addr_r_0__bdd_4_lut_14384.LUT_INIT = 16'he4aa;
    SB_DFF i554_555 (.Q(\REG.mem_5_12 ), .C(FIFO_CLK_c), .D(n5809));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4644_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_15_26 ), .O(n6143));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4644_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16575_bdd_4_lut (.I0(n16575), .I1(\REG.mem_13_29 ), .I2(\REG.mem_12_29 ), 
            .I3(rd_addr_r[1]), .O(n16578));
    defparam n16575_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i551_552 (.Q(\REG.mem_5_11 ), .C(FIFO_CLK_c), .D(n5808));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4643_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_15_25 ), .O(n6142));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4643_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY wr_addr_r_5__I_0_128_3 (.CI(n13718), .I0(wr_addr_r[1]), .I1(GND_net), 
            .CO(n13719));
    SB_LUT4 i4642_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_15_24 ), .O(n6141));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4642_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i548_549 (.Q(\REG.mem_5_10 ), .C(FIFO_CLK_c), .D(n5807));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4641_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_15_23 ), .O(n6140));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4641_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i545_546 (.Q(\REG.mem_5_9 ), .C(FIFO_CLK_c), .D(n5806));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i221_222 (.Q(\REG.mem_1_29 ), .C(FIFO_CLK_c), .D(n5655));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4640_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_15_22 ), .O(n6139));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4640_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4639_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_15_21 ), .O(n6138));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4639_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4638_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_15_20 ), .O(n6137));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4638_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i542_543 (.Q(\REG.mem_5_8 ), .C(FIFO_CLK_c), .D(n5805));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i539_540 (.Q(\REG.mem_5_7 ), .C(FIFO_CLK_c), .D(n5804));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15032 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_18 ), 
            .I2(\REG.mem_27_18 ), .I3(rd_addr_r[1]), .O(n17307));
    defparam rd_addr_r_0__bdd_4_lut_15032.LUT_INIT = 16'he4aa;
    SB_LUT4 i4637_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_15_19 ), .O(n6136));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4637_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4636_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_15_18 ), .O(n6135));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4636_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i149_150 (.Q(\REG.mem_1_5 ), .C(FIFO_CLK_c), .D(n5654));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4635_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_15_17 ), .O(n6134));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4635_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14379 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_31 ), 
            .I2(\REG.mem_7_31 ), .I3(rd_addr_r[1]), .O(n16569));
    defparam rd_addr_r_0__bdd_4_lut_14379.LUT_INIT = 16'he4aa;
    SB_LUT4 n16569_bdd_4_lut (.I0(n16569), .I1(\REG.mem_5_31 ), .I2(\REG.mem_4_31 ), 
            .I3(rd_addr_r[1]), .O(n14879));
    defparam n16569_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4634_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_15_16 ), .O(n6133));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4634_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i152_153 (.Q(\REG.mem_1_6 ), .C(FIFO_CLK_c), .D(n5653));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4633_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_15_15 ), .O(n6132));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4633_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14409 (.I0(rd_addr_r[1]), .I1(n14949), 
            .I2(n14950), .I3(rd_addr_r[2]), .O(n16563));
    defparam rd_addr_r_1__bdd_4_lut_14409.LUT_INIT = 16'he4aa;
    SB_LUT4 i4632_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_15_14 ), .O(n6131));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4632_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4631_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_15_13 ), .O(n6130));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4631_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i155_156 (.Q(\REG.mem_1_7 ), .C(FIFO_CLK_c), .D(n5652));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n16563_bdd_4_lut (.I0(n16563), .I1(n14944), .I2(n14943), .I3(rd_addr_r[2]), 
            .O(n16566));
    defparam n16563_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14100 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_31 ), 
            .I2(\REG.mem_3_31 ), .I3(rd_addr_r[1]), .O(n16221));
    defparam rd_addr_r_0__bdd_4_lut_14100.LUT_INIT = 16'he4aa;
    SB_DFF i158_159 (.Q(\REG.mem_1_8 ), .C(FIFO_CLK_c), .D(n5651));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i161_162 (.Q(\REG.mem_1_9 ), .C(FIFO_CLK_c), .D(n5650));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4580_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_13_26 ), .O(n6079));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4580_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4630_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_15_12 ), .O(n6129));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4630_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4579_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_13_25 ), .O(n6078));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4579_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17307_bdd_4_lut (.I0(n17307), .I1(\REG.mem_25_18 ), .I2(\REG.mem_24_18 ), 
            .I3(rd_addr_r[1]), .O(n15707));
    defparam n17307_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4629_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_15_11 ), .O(n6128));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4629_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i536_537 (.Q(\REG.mem_5_6 ), .C(FIFO_CLK_c), .D(n5803));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4628_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_15_10 ), .O(n6127));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4628_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i533_534 (.Q(\REG.mem_5_5 ), .C(FIFO_CLK_c), .D(n5802));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i164_165 (.Q(\REG.mem_1_10 ), .C(FIFO_CLK_c), .D(n5649));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wp_sync2_r__i0 (.Q(wp_sync2_r[0]), .C(SLM_CLK_c), .D(n5648));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 n16221_bdd_4_lut (.I0(n16221), .I1(\REG.mem_1_31 ), .I2(\REG.mem_0_31 ), 
            .I3(rd_addr_r[1]), .O(n16224));
    defparam n16221_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4627_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_15_9 ), .O(n6126));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4627_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_r_5__I_0_128_2_lut (.I0(GND_net), .I1(\wr_addr_r[0] ), 
            .I2(GND_net), .I3(VCC_net), .O(\wr_addr_p1_w[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_5__I_0_128_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF i530_531 (.Q(\REG.mem_5_4 ), .C(FIFO_CLK_c), .D(n5801));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4578_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_13_24 ), .O(n6077));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4578_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4626_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_15_8 ), .O(n6125));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4626_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4625_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_15_7 ), .O(n6124));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4625_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4624_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_15_6 ), .O(n6123));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4624_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4623_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_15_5 ), .O(n6122));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4623_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4577_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_13_23 ), .O(n6076));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4577_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4576_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_13_22 ), .O(n6075));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4576_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4575_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_13_21 ), .O(n6074));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4575_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4622_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_15_4 ), .O(n6121));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4622_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i527_528 (.Q(\REG.mem_5_3 ), .C(FIFO_CLK_c), .D(n5800));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4574_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_13_20 ), .O(n6073));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4574_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4621_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_15_3 ), .O(n6120));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4621_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY wr_addr_r_5__I_0_128_2 (.CI(VCC_net), .I0(\wr_addr_r[0] ), 
            .I1(GND_net), .CO(n13718));
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14369 (.I0(rd_addr_r[1]), .I1(n14838), 
            .I2(n14839), .I3(rd_addr_r[2]), .O(n16557));
    defparam rd_addr_r_1__bdd_4_lut_14369.LUT_INIT = 16'he4aa;
    SB_LUT4 i4573_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_13_19 ), .O(n6072));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4573_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4572_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_13_18 ), .O(n6071));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4572_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16557_bdd_4_lut (.I0(n16557), .I1(n14830), .I2(n14829), .I3(rd_addr_r[2]), 
            .O(n16560));
    defparam n16557_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4571_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_13_17 ), .O(n6070));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4571_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i224_225 (.Q(\REG.mem_1_30 ), .C(FIFO_CLK_c), .D(n5644));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4570_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_13_16 ), .O(n6069));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4570_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i209_210 (.Q(\REG.mem_1_25 ), .C(FIFO_CLK_c), .D(n5643));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14987 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_2 ), 
            .I2(\REG.mem_23_2 ), .I3(rd_addr_r[1]), .O(n17295));
    defparam rd_addr_r_0__bdd_4_lut_14987.LUT_INIT = 16'he4aa;
    SB_DFF wp_sync1_r__i0 (.Q(wp_sync1_r[0]), .C(SLM_CLK_c), .D(n5642));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n5641));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_LUT4 i4620_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_15_2 ), .O(n6119));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4620_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16161_bdd_4_lut (.I0(n16161), .I1(n15220), .I2(n15219), .I3(rd_addr_r[2]), 
            .O(n16164));
    defparam n16161_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i197_198 (.Q(\REG.mem_1_21 ), .C(FIFO_CLK_c), .D(n5640));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync2_r__i0 (.Q(rp_sync2_r[0]), .C(FIFO_CLK_c), .D(n5639));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_LUT4 n16191_bdd_4_lut (.I0(n16191), .I1(n14929), .I2(n14928), .I3(rd_addr_r[2]), 
            .O(n16194));
    defparam n16191_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4569_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_13_15 ), .O(n6068));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4569_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF rp_sync1_r__i0 (.Q(rp_sync1_r[0]), .C(FIFO_CLK_c), .D(n5638));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i167_168 (.Q(\REG.mem_1_11 ), .C(FIFO_CLK_c), .D(n5637));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i170_171 (.Q(\REG.mem_1_12 ), .C(FIFO_CLK_c), .D(n5635));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i173_174 (.Q(\REG.mem_1_13 ), .C(FIFO_CLK_c), .D(n5634));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i53_54 (.Q(\REG.mem_0_5 ), .C(FIFO_CLK_c), .D(n5633));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14259 (.I0(rd_addr_r[3]), .I1(n15660), 
            .I2(n15661), .I3(rd_addr_r[4]), .O(n16215));
    defparam rd_addr_r_3__bdd_4_lut_14259.LUT_INIT = 16'he4aa;
    SB_DFF i56_57 (.Q(\REG.mem_0_6 ), .C(FIFO_CLK_c), .D(n5632));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n17295_bdd_4_lut (.I0(n17295), .I1(\REG.mem_21_2 ), .I2(\REG.mem_20_2 ), 
            .I3(rd_addr_r[1]), .O(n15713));
    defparam n17295_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i176_177 (.Q(\REG.mem_1_14 ), .C(FIFO_CLK_c), .D(n5630));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i524_525 (.Q(\REG.mem_5_2 ), .C(FIFO_CLK_c), .D(n5799));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4619_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_15_1 ), .O(n6118));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4619_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i59_60 (.Q(\REG.mem_0_7 ), .C(FIFO_CLK_c), .D(n5627));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i521_522 (.Q(\REG.mem_5_1 ), .C(FIFO_CLK_c), .D(n5798));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i62_63 (.Q(\REG.mem_0_8 ), .C(FIFO_CLK_c), .D(n5626));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4618_3_lut_4_lut (.I0(n34), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_15_0 ), .O(n6117));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4618_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5001_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_26_31 ), .O(n6500));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5001_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5000_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_26_30 ), .O(n6499));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i5000_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4568_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_13_14 ), .O(n6067));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4568_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i518_519 (.Q(\REG.mem_5_0 ), .C(FIFO_CLK_c), .D(n5797));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i233_234 (.Q(\REG.mem_2_1 ), .C(FIFO_CLK_c), .D(n5623));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4999_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_26_29 ), .O(n6498));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4999_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14374 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_31 ), 
            .I2(\REG.mem_11_31 ), .I3(rd_addr_r[1]), .O(n16551));
    defparam rd_addr_r_0__bdd_4_lut_14374.LUT_INIT = 16'he4aa;
    SB_DFF i515_516 (.Q(\REG.mem_4_31 ), .C(FIFO_CLK_c), .D(n5796));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i65_66 (.Q(\REG.mem_0_9 ), .C(FIFO_CLK_c), .D(n5622));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4998_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_26_28 ), .O(n6497));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4998_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i68_69 (.Q(\REG.mem_0_10 ), .C(FIFO_CLK_c), .D(n5621));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i512_513 (.Q(\REG.mem_4_30 ), .C(FIFO_CLK_c), .D(n5795));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i212_213 (.Q(\REG.mem_1_26 ), .C(FIFO_CLK_c), .D(n5619));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i179_180 (.Q(\REG.mem_1_15 ), .C(FIFO_CLK_c), .D(n5616));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14977 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_21 ), 
            .I2(\REG.mem_23_21 ), .I3(rd_addr_r[1]), .O(n17289));
    defparam rd_addr_r_0__bdd_4_lut_14977.LUT_INIT = 16'he4aa;
    SB_LUT4 i4567_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_13_13 ), .O(n6066));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4567_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i182_183 (.Q(\REG.mem_1_16 ), .C(FIFO_CLK_c), .D(n5615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4997_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_26_27 ), .O(n6496));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4997_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17289_bdd_4_lut (.I0(n17289), .I1(\REG.mem_21_21 ), .I2(\REG.mem_20_21 ), 
            .I3(rd_addr_r[1]), .O(n15230));
    defparam n17289_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16551_bdd_4_lut (.I0(n16551), .I1(\REG.mem_9_31 ), .I2(\REG.mem_8_31 ), 
            .I3(rd_addr_r[1]), .O(n14882));
    defparam n16551_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i509_510 (.Q(\REG.mem_4_29 ), .C(FIFO_CLK_c), .D(n5794));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i506_507 (.Q(\REG.mem_4_28 ), .C(FIFO_CLK_c), .D(n5793));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14364 (.I0(rd_addr_r[1]), .I1(n15600), 
            .I2(n15601), .I3(rd_addr_r[2]), .O(n16545));
    defparam rd_addr_r_1__bdd_4_lut_14364.LUT_INIT = 16'he4aa;
    SB_LUT4 i4996_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_26_26 ), .O(n6495));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4996_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4566_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_13_12 ), .O(n6065));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4566_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4995_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_26_25 ), .O(n6494));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4995_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4994_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_26_24 ), .O(n6493));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4994_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4993_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_26_23 ), .O(n6492));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4993_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4992_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_26_22 ), .O(n6491));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4992_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i503_504 (.Q(\REG.mem_4_27 ), .C(FIFO_CLK_c), .D(n5792));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4991_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_26_21 ), .O(n6490));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4991_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4990_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_26_20 ), .O(n6489));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4990_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4989_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_26_19 ), .O(n6488));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4989_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16545_bdd_4_lut (.I0(n16545), .I1(n14815), .I2(n14814), .I3(rd_addr_r[2]), 
            .O(n16548));
    defparam n16545_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4988_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_26_18 ), .O(n6487));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4988_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14354 (.I0(rd_addr_r[1]), .I1(n15879), 
            .I2(n15880), .I3(rd_addr_r[2]), .O(n16539));
    defparam rd_addr_r_1__bdd_4_lut_14354.LUT_INIT = 16'he4aa;
    SB_DFF i500_501 (.Q(\REG.mem_4_26 ), .C(FIFO_CLK_c), .D(n5791));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i497_498 (.Q(\REG.mem_4_25 ), .C(FIFO_CLK_c), .D(n5790));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i494_495 (.Q(\REG.mem_4_24 ), .C(FIFO_CLK_c), .D(n5789));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i491_492 (.Q(\REG.mem_4_23 ), .C(FIFO_CLK_c), .D(n5788));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i488_489 (.Q(\REG.mem_4_22 ), .C(FIFO_CLK_c), .D(n5787));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i485_486 (.Q(\REG.mem_4_21 ), .C(FIFO_CLK_c), .D(n5786));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i482_483 (.Q(\REG.mem_4_20 ), .C(FIFO_CLK_c), .D(n5785));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i479_480 (.Q(\REG.mem_4_19 ), .C(FIFO_CLK_c), .D(n5784));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i476_477 (.Q(\REG.mem_4_18 ), .C(FIFO_CLK_c), .D(n5783));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i185_186 (.Q(\REG.mem_1_17 ), .C(FIFO_CLK_c), .D(n5610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i188_189 (.Q(\REG.mem_1_18 ), .C(FIFO_CLK_c), .D(n5607));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i200_201 (.Q(\REG.mem_1_22 ), .C(FIFO_CLK_c), .D(n5606));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wr_addr_r__i0 (.Q(\wr_addr_r[0] ), .C(FIFO_CLK_c), .D(n5605));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i236_237 (.Q(\REG.mem_2_2 ), .C(FIFO_CLK_c), .D(n5603));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i215_216 (.Q(\REG.mem_1_27 ), .C(FIFO_CLK_c), .D(n5602));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i473_474 (.Q(\REG.mem_4_17 ), .C(FIFO_CLK_c), .D(n5782));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4987_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_26_17 ), .O(n6486));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4987_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i470_471 (.Q(\REG.mem_4_16 ), .C(FIFO_CLK_c), .D(n5781));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i467_468 (.Q(\REG.mem_4_15 ), .C(FIFO_CLK_c), .D(n5780));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i464_465 (.Q(\REG.mem_4_14 ), .C(FIFO_CLK_c), .D(n5779));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i461_462 (.Q(\REG.mem_4_13 ), .C(FIFO_CLK_c), .D(n5778));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i203_204 (.Q(\REG.mem_1_23 ), .C(FIFO_CLK_c), .D(n5601));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i191_192 (.Q(\REG.mem_1_19 ), .C(FIFO_CLK_c), .D(n5600));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i239_240 (.Q(\REG.mem_2_3 ), .C(FIFO_CLK_c), .D(n5599));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i218_219 (.Q(\REG.mem_1_28 ), .C(FIFO_CLK_c), .D(n5598));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i458_459 (.Q(\REG.mem_4_12 ), .C(FIFO_CLK_c), .D(n5777));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4565_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_13_11 ), .O(n6064));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4565_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16539_bdd_4_lut (.I0(n16539), .I1(n15868), .I2(n15867), .I3(rd_addr_r[2]), 
            .O(n16542));
    defparam n16539_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4986_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_26_16 ), .O(n6485));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4986_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i1_1_lut (.I0(rd_addr_r[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i2_1_lut (.I0(rd_addr_r[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14359 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_23 ), 
            .I2(\REG.mem_31_23 ), .I3(rd_addr_r[1]), .O(n16533));
    defparam rd_addr_r_0__bdd_4_lut_14359.LUT_INIT = 16'he4aa;
    SB_LUT4 i4985_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_26_15 ), .O(n6484));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4985_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4984_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_26_14 ), .O(n6483));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4984_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16533_bdd_4_lut (.I0(n16533), .I1(\REG.mem_29_23 ), .I2(\REG.mem_28_23 ), 
            .I3(rd_addr_r[1]), .O(n16536));
    defparam n16533_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4983_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_26_13 ), .O(n6482));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4983_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_15077 (.I0(rd_addr_r[2]), .I1(n16266), 
            .I2(n16242), .I3(rd_addr_r[3]), .O(n17277));
    defparam rd_addr_r_2__bdd_4_lut_15077.LUT_INIT = 16'he4aa;
    SB_LUT4 n17277_bdd_4_lut (.I0(n17277), .I1(n16326), .I2(n16344), .I3(rd_addr_r[3]), 
            .O(n17280));
    defparam n17277_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4489_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_10_31 ), .O(n5988));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4489_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14344 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_31 ), 
            .I2(\REG.mem_15_31 ), .I3(rd_addr_r[1]), .O(n16527));
    defparam rd_addr_r_0__bdd_4_lut_14344.LUT_INIT = 16'he4aa;
    SB_LUT4 i4982_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_26_12 ), .O(n6481));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4982_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i3_1_lut (.I0(rd_addr_r[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n16527_bdd_4_lut (.I0(n16527), .I1(\REG.mem_13_31 ), .I2(\REG.mem_12_31 ), 
            .I3(rd_addr_r[1]), .O(n14885));
    defparam n16527_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4488_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_10_30 ), .O(n5987));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4488_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4487_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_10_29 ), .O(n5986));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4487_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i29_2_lut (.I0(n12_adj_1391), .I1(wr_addr_r[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i29_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4486_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_10_28 ), .O(n5985));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4486_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4485_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_10_27 ), .O(n5984));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4485_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13068_3_lut (.I0(\REG.mem_0_10 ), .I1(\REG.mem_1_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15192));
    defparam i13068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4484_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_10_26 ), .O(n5983));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4484_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14972 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_2 ), 
            .I2(\REG.mem_27_2 ), .I3(rd_addr_r[1]), .O(n17271));
    defparam rd_addr_r_0__bdd_4_lut_14972.LUT_INIT = 16'he4aa;
    SB_LUT4 i4981_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_26_11 ), .O(n6480));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4981_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4483_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_10_25 ), .O(n5982));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4483_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14339 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_31 ), 
            .I2(\REG.mem_19_31 ), .I3(rd_addr_r[1]), .O(n16521));
    defparam rd_addr_r_0__bdd_4_lut_14339.LUT_INIT = 16'he4aa;
    SB_LUT4 i4482_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_10_24 ), .O(n5981));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4482_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4980_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_26_10 ), .O(n6479));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4980_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4481_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_10_23 ), .O(n5980));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4481_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13069_3_lut (.I0(\REG.mem_2_10 ), .I1(\REG.mem_3_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15193));
    defparam i13069_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i455_456 (.Q(\REG.mem_4_11 ), .C(FIFO_CLK_c), .D(n5776));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i452_453 (.Q(\REG.mem_4_10 ), .C(FIFO_CLK_c), .D(n5775));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i449_450 (.Q(\REG.mem_4_9 ), .C(FIFO_CLK_c), .D(n5774));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i446_447 (.Q(\REG.mem_4_8 ), .C(FIFO_CLK_c), .D(n5773));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4979_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_26_9 ), .O(n6478));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4979_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i443_444 (.Q(\REG.mem_4_7 ), .C(FIFO_CLK_c), .D(n5772));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i440_441 (.Q(\REG.mem_4_6 ), .C(FIFO_CLK_c), .D(n5771));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4480_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_10_22 ), .O(n5979));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4480_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i437_438 (.Q(\REG.mem_4_5 ), .C(FIFO_CLK_c), .D(n5770));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i434_435 (.Q(\REG.mem_4_4 ), .C(FIFO_CLK_c), .D(n5769));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i13072_3_lut (.I0(\REG.mem_6_10 ), .I1(\REG.mem_7_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15196));
    defparam i13072_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i431_432 (.Q(\REG.mem_4_3 ), .C(FIFO_CLK_c), .D(n5768));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i428_429 (.Q(\REG.mem_4_2 ), .C(FIFO_CLK_c), .D(n5767));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n17271_bdd_4_lut (.I0(n17271), .I1(\REG.mem_25_2 ), .I2(\REG.mem_24_2 ), 
            .I3(rd_addr_r[1]), .O(n15722));
    defparam n17271_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i425_426 (.Q(\REG.mem_4_1 ), .C(FIFO_CLK_c), .D(n5766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i422_423 (.Q(\REG.mem_4_0 ), .C(FIFO_CLK_c), .D(n5765));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i419_420 (.Q(\REG.mem_3_31 ), .C(FIFO_CLK_c), .D(n5764));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i416_417 (.Q(\REG.mem_3_30 ), .C(FIFO_CLK_c), .D(n5763));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4978_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_26_8 ), .O(n6477));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4978_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4977_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_26_7 ), .O(n6476));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4977_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4564_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_13_10 ), .O(n6063));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4564_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16521_bdd_4_lut (.I0(n16521), .I1(\REG.mem_17_31 ), .I2(\REG.mem_16_31 ), 
            .I3(rd_addr_r[1]), .O(n16524));
    defparam n16521_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4479_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_10_21 ), .O(n5978));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4479_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i413_414 (.Q(\REG.mem_3_29 ), .C(FIFO_CLK_c), .D(n5762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4478_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_10_20 ), .O(n5977));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4478_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4477_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_10_19 ), .O(n5976));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4477_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i410_411 (.Q(\REG.mem_3_28 ), .C(FIFO_CLK_c), .D(n5761));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\REG.mem_26_27 ), 
            .I2(\REG.mem_27_27 ), .I3(rd_addr_r[1]), .O(n18027));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF i407_408 (.Q(\REG.mem_3_27 ), .C(FIFO_CLK_c), .D(n5760));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n18027_bdd_4_lut (.I0(n18027), .I1(\REG.mem_25_27 ), .I2(\REG.mem_24_27 ), 
            .I3(rd_addr_r[1]), .O(n15392));
    defparam n18027_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14334 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_31 ), 
            .I2(\REG.mem_23_31 ), .I3(rd_addr_r[1]), .O(n16515));
    defparam rd_addr_r_0__bdd_4_lut_14334.LUT_INIT = 16'he4aa;
    SB_LUT4 i13071_3_lut (.I0(\REG.mem_4_10 ), .I1(\REG.mem_5_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15195));
    defparam i13071_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i404_405 (.Q(\REG.mem_3_26 ), .C(FIFO_CLK_c), .D(n5759));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n16515_bdd_4_lut (.I0(n16515), .I1(\REG.mem_21_31 ), .I2(\REG.mem_20_31 ), 
            .I3(rd_addr_r[1]), .O(n16518));
    defparam n16515_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4476_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_10_18 ), .O(n5975));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4476_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4475_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_10_17 ), .O(n5974));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4475_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i401_402 (.Q(\REG.mem_3_25 ), .C(FIFO_CLK_c), .D(n5758));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i398_399 (.Q(\REG.mem_3_24 ), .C(FIFO_CLK_c), .D(n5757));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14329 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_31 ), 
            .I2(\REG.mem_27_31 ), .I3(rd_addr_r[1]), .O(n16503));
    defparam rd_addr_r_0__bdd_4_lut_14329.LUT_INIT = 16'he4aa;
    SB_DFF i395_396 (.Q(\REG.mem_3_23 ), .C(FIFO_CLK_c), .D(n5756));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4474_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_10_16 ), .O(n5973));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4474_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4976_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_26_6 ), .O(n6475));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4976_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15587 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_27 ), 
            .I2(\REG.mem_7_27 ), .I3(rd_addr_r[1]), .O(n18021));
    defparam rd_addr_r_0__bdd_4_lut_15587.LUT_INIT = 16'he4aa;
    SB_DFF i392_393 (.Q(\REG.mem_3_22 ), .C(FIFO_CLK_c), .D(n5755));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n16215_bdd_4_lut (.I0(n16215), .I1(n14731), .I2(n16194), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[29]));
    defparam n16215_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i389_390 (.Q(\REG.mem_3_21 ), .C(FIFO_CLK_c), .D(n5754));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n18021_bdd_4_lut (.I0(n18021), .I1(\REG.mem_5_27 ), .I2(\REG.mem_4_27 ), 
            .I3(rd_addr_r[1]), .O(n14948));
    defparam n18021_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4975_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_26_5 ), .O(n6474));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4975_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16503_bdd_4_lut (.I0(n16503), .I1(\REG.mem_25_31 ), .I2(\REG.mem_24_31 ), 
            .I3(rd_addr_r[1]), .O(n16506));
    defparam n16503_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4974_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_26_4 ), .O(n6473));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4974_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4473_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_10_15 ), .O(n5972));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4473_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4472_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_10_14 ), .O(n5971));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4472_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4471_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_10_13 ), .O(n5970));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4471_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4973_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_26_3 ), .O(n6472));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4973_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4563_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_13_9 ), .O(n6062));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4563_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4470_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_10_12 ), .O(n5969));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4470_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4562_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_13_8 ), .O(n6061));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4562_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14957 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_6 ), 
            .I2(\REG.mem_23_6 ), .I3(rd_addr_r[1]), .O(n17259));
    defparam rd_addr_r_0__bdd_4_lut_14957.LUT_INIT = 16'he4aa;
    SB_LUT4 i4469_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_10_11 ), .O(n5968));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4469_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17259_bdd_4_lut (.I0(n17259), .I1(\REG.mem_21_6 ), .I2(\REG.mem_20_6 ), 
            .I3(rd_addr_r[1]), .O(n15728));
    defparam n17259_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4468_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_10_10 ), .O(n5967));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4468_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4972_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_26_2 ), .O(n6471));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4972_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15582 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_27 ), 
            .I2(\REG.mem_31_27 ), .I3(rd_addr_r[1]), .O(n18015));
    defparam rd_addr_r_0__bdd_4_lut_15582.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14319 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_4 ), 
            .I2(\REG.mem_15_4 ), .I3(rd_addr_r[1]), .O(n16497));
    defparam rd_addr_r_0__bdd_4_lut_14319.LUT_INIT = 16'he4aa;
    SB_LUT4 n16497_bdd_4_lut (.I0(n16497), .I1(\REG.mem_13_4 ), .I2(\REG.mem_12_4 ), 
            .I3(rd_addr_r[1]), .O(n15326));
    defparam n16497_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4971_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_26_1 ), .O(n6470));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4971_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12598_3_lut (.I0(n17256), .I1(n17214), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n14722));
    defparam i12598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4467_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_10_9 ), .O(n5966));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4467_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n18015_bdd_4_lut (.I0(n18015), .I1(\REG.mem_29_27 ), .I2(\REG.mem_28_27 ), 
            .I3(rd_addr_r[1]), .O(n15401));
    defparam n18015_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4466_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_10_8 ), .O(n5965));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4466_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4465_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_10_7 ), .O(n5964));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4465_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4464_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_10_6 ), .O(n5963));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4464_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13741_3_lut (.I0(\REG.mem_22_22 ), .I1(\REG.mem_23_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15865));
    defparam i13741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14947 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_10 ), 
            .I2(\REG.mem_27_10 ), .I3(rd_addr_r[1]), .O(n17253));
    defparam rd_addr_r_0__bdd_4_lut_14947.LUT_INIT = 16'he4aa;
    SB_LUT4 n17253_bdd_4_lut (.I0(n17253), .I1(\REG.mem_25_10 ), .I2(\REG.mem_24_10 ), 
            .I3(rd_addr_r[1]), .O(n17256));
    defparam n17253_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15577 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_4 ), 
            .I2(\REG.mem_27_4 ), .I3(rd_addr_r[1]), .O(n18009));
    defparam rd_addr_r_0__bdd_4_lut_15577.LUT_INIT = 16'he4aa;
    SB_LUT4 n18009_bdd_4_lut (.I0(n18009), .I1(\REG.mem_25_4 ), .I2(\REG.mem_24_4 ), 
            .I3(rd_addr_r[1]), .O(n15407));
    defparam n18009_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13740_3_lut (.I0(\REG.mem_20_22 ), .I1(\REG.mem_21_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15864));
    defparam i13740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14942 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_18 ), 
            .I2(\REG.mem_31_18 ), .I3(rd_addr_r[1]), .O(n17247));
    defparam rd_addr_r_0__bdd_4_lut_14942.LUT_INIT = 16'he4aa;
    SB_LUT4 n17247_bdd_4_lut (.I0(n17247), .I1(\REG.mem_29_18 ), .I2(\REG.mem_28_18 ), 
            .I3(rd_addr_r[1]), .O(n15731));
    defparam n17247_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4970_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_26_0 ), .O(n6469));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4970_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15572 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_24 ), 
            .I2(\REG.mem_27_24 ), .I3(rd_addr_r[1]), .O(n18003));
    defparam rd_addr_r_0__bdd_4_lut_15572.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14349 (.I0(rd_addr_r[1]), .I1(n15861), 
            .I2(n15862), .I3(rd_addr_r[2]), .O(n16479));
    defparam rd_addr_r_1__bdd_4_lut_14349.LUT_INIT = 16'he4aa;
    SB_LUT4 i4463_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_10_5 ), .O(n5962));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4463_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16479_bdd_4_lut (.I0(n16479), .I1(n15850), .I2(n15849), .I3(rd_addr_r[2]), 
            .O(n16482));
    defparam n16479_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n18003_bdd_4_lut (.I0(n18003), .I1(\REG.mem_25_24 ), .I2(\REG.mem_24_24 ), 
            .I3(rd_addr_r[1]), .O(n18006));
    defparam n18003_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14404 (.I0(rd_addr_r[3]), .I1(n16254), 
            .I2(n14755), .I3(rd_addr_r[4]), .O(n16473));
    defparam rd_addr_r_3__bdd_4_lut_14404.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15567 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_4 ), 
            .I2(\REG.mem_19_4 ), .I3(rd_addr_r[1]), .O(n17997));
    defparam rd_addr_r_0__bdd_4_lut_15567.LUT_INIT = 16'he4aa;
    SB_LUT4 i4462_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_10_4 ), .O(n5961));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4462_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16473_bdd_4_lut (.I0(n16473), .I1(n15898), .I2(n15897), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[22]));
    defparam n16473_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17997_bdd_4_lut (.I0(n17997), .I1(\REG.mem_17_4 ), .I2(\REG.mem_16_4 ), 
            .I3(rd_addr_r[1]), .O(n15419));
    defparam n17997_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13099_3_lut (.I0(\REG.mem_22_10 ), .I1(\REG.mem_23_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15223));
    defparam i13099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13098_3_lut (.I0(\REG.mem_20_10 ), .I1(\REG.mem_21_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15222));
    defparam i13098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12852_3_lut (.I0(\REG.mem_0_13 ), .I1(\REG.mem_1_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14976));
    defparam i12852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12853_3_lut (.I0(\REG.mem_2_13 ), .I1(\REG.mem_3_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14977));
    defparam i12853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12856_3_lut (.I0(\REG.mem_6_13 ), .I1(\REG.mem_7_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14980));
    defparam i12856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12855_3_lut (.I0(\REG.mem_4_13 ), .I1(\REG.mem_5_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14979));
    defparam i12855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13503_3_lut (.I0(\REG.mem_0_6 ), .I1(\REG.mem_1_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15627));
    defparam i13503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13504_3_lut (.I0(\REG.mem_2_6 ), .I1(\REG.mem_3_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15628));
    defparam i13504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13384_3_lut (.I0(\REG.mem_6_6 ), .I1(\REG.mem_7_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15508));
    defparam i13384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13383_3_lut (.I0(\REG.mem_4_6 ), .I1(\REG.mem_5_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15507));
    defparam i13383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13770_3_lut (.I0(\REG.mem_0_0 ), .I1(\REG.mem_1_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15894));
    defparam i13770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13771_3_lut (.I0(\REG.mem_2_0 ), .I1(\REG.mem_3_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15895));
    defparam i13771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12679_3_lut (.I0(\REG.mem_6_0 ), .I1(\REG.mem_7_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14803));
    defparam i12679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12678_3_lut (.I0(\REG.mem_4_0 ), .I1(\REG.mem_5_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14802));
    defparam i12678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12858_3_lut (.I0(\REG.mem_16_0 ), .I1(\REG.mem_17_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14982));
    defparam i12858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12859_3_lut (.I0(\REG.mem_18_0 ), .I1(\REG.mem_19_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14983));
    defparam i12859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12868_3_lut (.I0(\REG.mem_22_0 ), .I1(\REG.mem_23_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14992));
    defparam i12868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12867_3_lut (.I0(\REG.mem_20_0 ), .I1(\REG.mem_21_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14991));
    defparam i12867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12808_3_lut (.I0(\REG.mem_6_29 ), .I1(\REG.mem_7_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14932));
    defparam i12808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12807_3_lut (.I0(\REG.mem_4_29 ), .I1(\REG.mem_5_29 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14931));
    defparam i12807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12894_3_lut (.I0(\REG.mem_0_12 ), .I1(\REG.mem_1_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15018));
    defparam i12894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12895_3_lut (.I0(\REG.mem_2_12 ), .I1(\REG.mem_3_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15019));
    defparam i12895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12901_3_lut (.I0(\REG.mem_6_12 ), .I1(\REG.mem_7_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15025));
    defparam i12901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12900_3_lut (.I0(\REG.mem_4_12 ), .I1(\REG.mem_5_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15024));
    defparam i12900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4461_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_10_3 ), .O(n5960));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4461_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15562 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_27 ), 
            .I2(\REG.mem_11_27 ), .I3(rd_addr_r[1]), .O(n17991));
    defparam rd_addr_r_0__bdd_4_lut_15562.LUT_INIT = 16'he4aa;
    SB_LUT4 i12906_3_lut (.I0(\REG.mem_16_12 ), .I1(\REG.mem_17_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15030));
    defparam i12906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4460_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_10_2 ), .O(n5959));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4460_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4459_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_10_1 ), .O(n5958));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4459_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17991_bdd_4_lut (.I0(n17991), .I1(\REG.mem_9_27 ), .I2(\REG.mem_8_27 ), 
            .I3(rd_addr_r[1]), .O(n14960));
    defparam n17991_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14538 (.I0(rd_addr_r[2]), .I1(n15392), 
            .I2(n15401), .I3(rd_addr_r[3]), .O(n16455));
    defparam rd_addr_r_2__bdd_4_lut_14538.LUT_INIT = 16'he4aa;
    SB_LUT4 n16455_bdd_4_lut (.I0(n16455), .I1(n15281), .I2(n15146), .I3(rd_addr_r[3]), 
            .O(n16458));
    defparam n16455_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14294 (.I0(rd_addr_r[3]), .I1(n15594), 
            .I2(n15595), .I3(rd_addr_r[4]), .O(n16449));
    defparam rd_addr_r_3__bdd_4_lut_14294.LUT_INIT = 16'he4aa;
    SB_LUT4 i12907_3_lut (.I0(\REG.mem_18_12 ), .I1(\REG.mem_19_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15031));
    defparam i12907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12913_3_lut (.I0(\REG.mem_22_12 ), .I1(\REG.mem_23_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15037));
    defparam i12913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12912_3_lut (.I0(\REG.mem_20_12 ), .I1(\REG.mem_21_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15036));
    defparam i12912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13572_3_lut (.I0(\REG.mem_16_26 ), .I1(\REG.mem_17_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15696));
    defparam i13572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13573_3_lut (.I0(\REG.mem_18_26 ), .I1(\REG.mem_19_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15697));
    defparam i13573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15557 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_17 ), 
            .I2(\REG.mem_31_17 ), .I3(rd_addr_r[1]), .O(n17979));
    defparam rd_addr_r_0__bdd_4_lut_15557.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14937 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_6 ), 
            .I2(\REG.mem_27_6 ), .I3(rd_addr_r[1]), .O(n17217));
    defparam rd_addr_r_0__bdd_4_lut_14937.LUT_INIT = 16'he4aa;
    SB_LUT4 n17217_bdd_4_lut (.I0(n17217), .I1(\REG.mem_25_6 ), .I2(\REG.mem_24_6 ), 
            .I3(rd_addr_r[1]), .O(n15746));
    defparam n17217_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17979_bdd_4_lut (.I0(n17979), .I1(\REG.mem_29_17 ), .I2(\REG.mem_28_17 ), 
            .I3(rd_addr_r[1]), .O(n15425));
    defparam n17979_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14912 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_10 ), 
            .I2(\REG.mem_31_10 ), .I3(rd_addr_r[1]), .O(n17211));
    defparam rd_addr_r_0__bdd_4_lut_14912.LUT_INIT = 16'he4aa;
    SB_LUT4 n16449_bdd_4_lut (.I0(n16449), .I1(n14821), .I2(n16422), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[19]));
    defparam n16449_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15547 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_4 ), 
            .I2(\REG.mem_7_4 ), .I3(rd_addr_r[1]), .O(n17973));
    defparam rd_addr_r_0__bdd_4_lut_15547.LUT_INIT = 16'he4aa;
    SB_LUT4 i4458_3_lut_4_lut (.I0(n24), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_10_0 ), .O(n5957));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4458_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13369_3_lut (.I0(\REG.mem_22_26 ), .I1(\REG.mem_23_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15493));
    defparam i13369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13368_3_lut (.I0(\REG.mem_20_26 ), .I1(\REG.mem_21_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15492));
    defparam i13368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12928_3_lut (.I0(n17706), .I1(n17928), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15052));
    defparam i12928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12948_3_lut (.I0(\REG.mem_24_5 ), .I1(\REG.mem_25_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15072));
    defparam i12948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12949_3_lut (.I0(\REG.mem_26_5 ), .I1(\REG.mem_27_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15073));
    defparam i12949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12838_3_lut (.I0(n16584), .I1(n16188), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n14962));
    defparam i12838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12964_3_lut (.I0(\REG.mem_30_5 ), .I1(\REG.mem_31_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15088));
    defparam i12964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12963_3_lut (.I0(\REG.mem_28_5 ), .I1(\REG.mem_29_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15087));
    defparam i12963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12844_3_lut (.I0(n18006), .I1(n17772), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n14968));
    defparam i12844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12934_3_lut (.I0(n17148), .I1(n17082), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15058));
    defparam i12934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13389_3_lut (.I0(\REG.mem_16_25 ), .I1(\REG.mem_17_25 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15513));
    defparam i13389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13390_3_lut (.I0(\REG.mem_18_25 ), .I1(\REG.mem_19_25 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15514));
    defparam i13390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17973_bdd_4_lut (.I0(n17973), .I1(\REG.mem_5_4 ), .I2(\REG.mem_4_4 ), 
            .I3(rd_addr_r[1]), .O(n15428));
    defparam n17973_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17211_bdd_4_lut (.I0(n17211), .I1(\REG.mem_29_10 ), .I2(\REG.mem_28_10 ), 
            .I3(rd_addr_r[1]), .O(n17214));
    defparam n17211_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4809_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_20_31 ), .O(n6308));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4809_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15542 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_17 ), 
            .I2(\REG.mem_7_17 ), .I3(rd_addr_r[1]), .O(n17967));
    defparam rd_addr_r_0__bdd_4_lut_15542.LUT_INIT = 16'he4aa;
    SB_LUT4 i4808_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_20_30 ), .O(n6307));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4808_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17967_bdd_4_lut (.I0(n17967), .I1(\REG.mem_5_17 ), .I2(\REG.mem_4_17 ), 
            .I3(rd_addr_r[1]), .O(n15440));
    defparam n17967_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14314 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_31 ), 
            .I2(\REG.mem_31_31 ), .I3(rd_addr_r[1]), .O(n16437));
    defparam rd_addr_r_0__bdd_4_lut_14314.LUT_INIT = 16'he4aa;
    SB_LUT4 n16437_bdd_4_lut (.I0(n16437), .I1(\REG.mem_29_31 ), .I2(\REG.mem_28_31 ), 
            .I3(rd_addr_r[1]), .O(n16440));
    defparam n16437_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14962 (.I0(rd_addr_r[2]), .I1(n15722), 
            .I2(n16722), .I3(rd_addr_r[3]), .O(n17205));
    defparam rd_addr_r_2__bdd_4_lut_14962.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15537 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_5 ), 
            .I2(\REG.mem_15_5 ), .I3(rd_addr_r[1]), .O(n17961));
    defparam rd_addr_r_0__bdd_4_lut_15537.LUT_INIT = 16'he4aa;
    SB_LUT4 n17961_bdd_4_lut (.I0(n17961), .I1(\REG.mem_13_5 ), .I2(\REG.mem_12_5 ), 
            .I3(rd_addr_r[1]), .O(n17964));
    defparam n17961_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4807_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_20_29 ), .O(n6306));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4807_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4806_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_20_28 ), .O(n6305));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4806_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4805_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_20_27 ), .O(n6304));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4805_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17205_bdd_4_lut (.I0(n17205), .I1(n15713), .I2(n16698), .I3(rd_addr_r[3]), 
            .O(n17208));
    defparam n17205_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14274 (.I0(rd_addr_r[3]), .I1(n16410), 
            .I2(n14809), .I3(rd_addr_r[4]), .O(n16431));
    defparam rd_addr_r_3__bdd_4_lut_14274.LUT_INIT = 16'he4aa;
    SB_LUT4 n16431_bdd_4_lut (.I0(n16431), .I1(n14782), .I2(n16296), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[28]));
    defparam n16431_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4804_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_20_26 ), .O(n6303));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4804_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14264 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_18 ), 
            .I2(\REG.mem_7_18 ), .I3(rd_addr_r[1]), .O(n16425));
    defparam rd_addr_r_0__bdd_4_lut_14264.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut (.I0(rd_addr_r[1]), .I1(n14988), .I2(n14989), 
            .I3(rd_addr_r[2]), .O(n17955));
    defparam rd_addr_r_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n17955_bdd_4_lut (.I0(n17955), .I1(n14986), .I2(n14985), .I3(rd_addr_r[2]), 
            .O(n15013));
    defparam n17955_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15527 (.I0(rd_addr_r[1]), .I1(n14973), 
            .I2(n14974), .I3(rd_addr_r[2]), .O(n17949));
    defparam rd_addr_r_1__bdd_4_lut_15527.LUT_INIT = 16'he4aa;
    SB_LUT4 i4561_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_13_7 ), .O(n6060));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4561_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13287_3_lut (.I0(\REG.mem_0_25 ), .I1(\REG.mem_1_25 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15411));
    defparam i13287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17949_bdd_4_lut (.I0(n17949), .I1(n14971), .I2(n14970), .I3(rd_addr_r[2]), 
            .O(n15016));
    defparam n17949_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16425_bdd_4_lut (.I0(n16425), .I1(\REG.mem_5_18 ), .I2(\REG.mem_4_18 ), 
            .I3(rd_addr_r[1]), .O(n16428));
    defparam n16425_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13288_3_lut (.I0(\REG.mem_2_25 ), .I1(\REG.mem_3_25 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15412));
    defparam i13288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4803_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_20_25 ), .O(n6302));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4803_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4802_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_20_24 ), .O(n6301));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4802_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4801_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_20_23 ), .O(n6300));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4801_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13405_3_lut (.I0(\REG.mem_22_25 ), .I1(\REG.mem_23_25 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15529));
    defparam i13405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13404_3_lut (.I0(\REG.mem_20_25 ), .I1(\REG.mem_21_25 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15528));
    defparam i13404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14299 (.I0(rd_addr_r[1]), .I1(n14778), 
            .I2(n14779), .I3(rd_addr_r[2]), .O(n16419));
    defparam rd_addr_r_1__bdd_4_lut_14299.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut (.I0(rd_addr_r[2]), .I1(n15407), .I2(n16206), 
            .I3(rd_addr_r[3]), .O(n17943));
    defparam rd_addr_r_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n17943_bdd_4_lut (.I0(n17943), .I1(n16182), .I2(n15419), .I3(rd_addr_r[3]), 
            .O(n17946));
    defparam n17943_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4560_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_13_6 ), .O(n6059));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4560_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16419_bdd_4_lut (.I0(n16419), .I1(n14773), .I2(n14772), .I3(rd_addr_r[2]), 
            .O(n16422));
    defparam n16419_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4800_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_20_22 ), .O(n6299));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4800_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15522 (.I0(rd_addr_r[1]), .I1(n15009), 
            .I2(n15010), .I3(rd_addr_r[2]), .O(n17937));
    defparam rd_addr_r_1__bdd_4_lut_15522.LUT_INIT = 16'he4aa;
    SB_LUT4 i4799_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_20_21 ), .O(n6298));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4799_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4798_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_20_20 ), .O(n6297));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4798_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14254 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_17 ), 
            .I2(\REG.mem_19_17 ), .I3(rd_addr_r[1]), .O(n16413));
    defparam rd_addr_r_0__bdd_4_lut_14254.LUT_INIT = 16'he4aa;
    SB_LUT4 n16413_bdd_4_lut (.I0(n16413), .I1(\REG.mem_17_17 ), .I2(\REG.mem_16_17 ), 
            .I3(rd_addr_r[1]), .O(n16416));
    defparam n16413_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4797_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_20_19 ), .O(n6296));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4797_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4171_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_1_0 ), .O(n5670));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4171_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17937_bdd_4_lut (.I0(n17937), .I1(n15001), .I2(n15000), .I3(rd_addr_r[2]), 
            .O(n15022));
    defparam n17937_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4145_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_1_30 ), .O(n5644));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4145_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15532 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_6 ), 
            .I2(\REG.mem_31_6 ), .I3(rd_addr_r[1]), .O(n17931));
    defparam rd_addr_r_0__bdd_4_lut_15532.LUT_INIT = 16'he4aa;
    SB_LUT4 n17931_bdd_4_lut (.I0(n17931), .I1(\REG.mem_29_6 ), .I2(\REG.mem_28_6 ), 
            .I3(rd_addr_r[1]), .O(n15488));
    defparam n17931_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14907 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_17 ), 
            .I2(\REG.mem_11_17 ), .I3(rd_addr_r[1]), .O(n17181));
    defparam rd_addr_r_0__bdd_4_lut_14907.LUT_INIT = 16'he4aa;
    SB_LUT4 n17181_bdd_4_lut (.I0(n17181), .I1(\REG.mem_9_17 ), .I2(\REG.mem_8_17 ), 
            .I3(rd_addr_r[1]), .O(n15239));
    defparam n17181_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15507 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_12 ), 
            .I2(\REG.mem_15_12 ), .I3(rd_addr_r[1]), .O(n17925));
    defparam rd_addr_r_0__bdd_4_lut_15507.LUT_INIT = 16'he4aa;
    SB_LUT4 i4796_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_20_18 ), .O(n6295));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4796_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4795_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_20_17 ), .O(n6294));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4795_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4160_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_1_31 ), .O(n5659));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4160_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14249 (.I0(rd_addr_r[1]), .I1(n14760), 
            .I2(n14761), .I3(rd_addr_r[2]), .O(n16407));
    defparam rd_addr_r_1__bdd_4_lut_14249.LUT_INIT = 16'he4aa;
    SB_LUT4 i4559_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_13_5 ), .O(n6058));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4559_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4794_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_20_16 ), .O(n6293));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4794_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4558_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_13_4 ), .O(n6057));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4558_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4101_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_1_19 ), .O(n5600));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4101_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17925_bdd_4_lut (.I0(n17925), .I1(\REG.mem_13_12 ), .I2(\REG.mem_12_12 ), 
            .I3(rd_addr_r[1]), .O(n17928));
    defparam n17925_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4793_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_20_15 ), .O(n6292));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4793_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16407_bdd_4_lut (.I0(n16407), .I1(n14758), .I2(n14757), .I3(rd_addr_r[2]), 
            .O(n16410));
    defparam n16407_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4792_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_20_14 ), .O(n6291));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4792_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4791_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_20_13 ), .O(n6290));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4791_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4790_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_20_12 ), .O(n6289));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4790_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4789_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_20_11 ), .O(n6288));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4789_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4557_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_13_3 ), .O(n6056));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4557_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4788_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_20_10 ), .O(n6287));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4788_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4787_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_20_9 ), .O(n6286));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4787_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14244 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_3 ), 
            .I2(\REG.mem_23_3 ), .I3(rd_addr_r[1]), .O(n16401));
    defparam rd_addr_r_0__bdd_4_lut_14244.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15502 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_6 ), 
            .I2(\REG.mem_19_6 ), .I3(rd_addr_r[1]), .O(n17919));
    defparam rd_addr_r_0__bdd_4_lut_15502.LUT_INIT = 16'he4aa;
    SB_LUT4 i4786_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_20_8 ), .O(n6285));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4786_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4785_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_20_7 ), .O(n6284));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4785_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4784_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_20_6 ), .O(n6283));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4784_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n16401_bdd_4_lut (.I0(n16401), .I1(\REG.mem_21_3 ), .I2(\REG.mem_20_3 ), 
            .I3(rd_addr_r[1]), .O(n16404));
    defparam n16401_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4783_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_20_5 ), .O(n6282));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4783_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4556_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_13_2 ), .O(n6055));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4556_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4782_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_20_4 ), .O(n6281));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4782_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4781_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_20_3 ), .O(n6280));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4781_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4107_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_1_22 ), .O(n5606));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4107_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4141_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_1_21 ), .O(n5640));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4141_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17919_bdd_4_lut (.I0(n17919), .I1(\REG.mem_17_6 ), .I2(\REG.mem_16_6 ), 
            .I3(rd_addr_r[1]), .O(n15503));
    defparam n17919_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4555_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_13_1 ), .O(n6054));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4555_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4780_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_20_2 ), .O(n6279));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4780_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4779_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_20_1 ), .O(n6278));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4779_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4778_3_lut_4_lut (.I0(n29), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_20_0 ), .O(n6277));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4778_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4155_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_1_5 ), .O(n5654));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4155_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4099_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_1_28 ), .O(n5598));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4099_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14095 (.I0(rd_addr_r[2]), .I1(n15266), 
            .I2(n15293), .I3(rd_addr_r[3]), .O(n16209));
    defparam rd_addr_r_2__bdd_4_lut_14095.LUT_INIT = 16'he4aa;
    SB_LUT4 i4103_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_1_27 ), .O(n5602));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4103_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4554_3_lut_4_lut (.I0(n30), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_13_0 ), .O(n6053));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4554_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4120_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_1_26 ), .O(n5619));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4120_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4144_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_1_25 ), .O(n5643));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4144_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14279 (.I0(rd_addr_r[2]), .I1(n14882), 
            .I2(n14885), .I3(rd_addr_r[3]), .O(n16395));
    defparam rd_addr_r_2__bdd_4_lut_14279.LUT_INIT = 16'he4aa;
    SB_LUT4 i4156_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_1_29 ), .O(n5655));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4156_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4102_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_1_23 ), .O(n5601));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4102_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4108_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_1_18 ), .O(n5607));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4108_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4111_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_1_17 ), .O(n5610));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4111_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16395_bdd_4_lut (.I0(n16395), .I1(n14879), .I2(n16224), .I3(rd_addr_r[3]), 
            .O(n16398));
    defparam n16395_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15027 (.I0(rd_addr_r[1]), .I1(n15213), 
            .I2(n15214), .I3(rd_addr_r[2]), .O(n17169));
    defparam rd_addr_r_1__bdd_4_lut_15027.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15497 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_16 ), 
            .I2(\REG.mem_3_16 ), .I3(rd_addr_r[1]), .O(n17907));
    defparam rd_addr_r_0__bdd_4_lut_15497.LUT_INIT = 16'he4aa;
    SB_LUT4 n17169_bdd_4_lut (.I0(n17169), .I1(n15208), .I2(n15207), .I3(rd_addr_r[2]), 
            .O(n15241));
    defparam n17169_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17907_bdd_4_lut (.I0(n17907), .I1(\REG.mem_1_16 ), .I2(\REG.mem_0_16 ), 
            .I3(rd_addr_r[1]), .O(n15035));
    defparam n17907_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_14239 (.I0(rd_addr_r[1]), .I1(n15141), 
            .I2(n15142), .I3(rd_addr_r[2]), .O(n16383));
    defparam rd_addr_r_1__bdd_4_lut_14239.LUT_INIT = 16'he4aa;
    SB_LUT4 n16383_bdd_4_lut (.I0(n16383), .I1(n15136), .I2(n15135), .I3(rd_addr_r[2]), 
            .O(n16386));
    defparam n16383_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4116_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_1_16 ), .O(n5615));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4116_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_15517 (.I0(rd_addr_r[2]), .I1(n16278), 
            .I2(n15425), .I3(rd_addr_r[3]), .O(n17901));
    defparam rd_addr_r_2__bdd_4_lut_15517.LUT_INIT = 16'he4aa;
    SB_LUT4 n17901_bdd_4_lut (.I0(n17901), .I1(n16320), .I2(n16416), .I3(rd_addr_r[3]), 
            .O(n17904));
    defparam n17901_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13321_3_lut (.I0(\REG.mem_6_25 ), .I1(\REG.mem_7_25 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15445));
    defparam i13321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_14997 (.I0(rd_addr_r[3]), .I1(n17052), 
            .I2(n15415), .I3(rd_addr_r[4]), .O(n17163));
    defparam rd_addr_r_3__bdd_4_lut_14997.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15487 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_21 ), 
            .I2(\REG.mem_3_21 ), .I3(rd_addr_r[1]), .O(n17895));
    defparam rd_addr_r_0__bdd_4_lut_15487.LUT_INIT = 16'he4aa;
    SB_LUT4 n17895_bdd_4_lut (.I0(n17895), .I1(\REG.mem_1_21 ), .I2(\REG.mem_0_21 ), 
            .I3(rd_addr_r[1]), .O(n15518));
    defparam n17895_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17163_bdd_4_lut (.I0(n17163), .I1(n15553), .I2(n15552), .I3(rd_addr_r[4]), 
            .O(rd_data_o_31__N_598[8]));
    defparam n17163_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14229 (.I0(rd_addr_r[2]), .I1(n15104), 
            .I2(n15134), .I3(rd_addr_r[3]), .O(n16377));
    defparam rd_addr_r_2__bdd_4_lut_14229.LUT_INIT = 16'he4aa;
    SB_LUT4 i13320_3_lut (.I0(\REG.mem_4_25 ), .I1(\REG.mem_5_25 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15444));
    defparam i13320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n16377_bdd_4_lut (.I0(n16377), .I1(n15542), .I2(n15518), .I3(rd_addr_r[3]), 
            .O(n16380));
    defparam n16377_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14234 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_30 ), 
            .I2(\REG.mem_3_30 ), .I3(rd_addr_r[1]), .O(n16371));
    defparam rd_addr_r_0__bdd_4_lut_14234.LUT_INIT = 16'he4aa;
    SB_LUT4 n16371_bdd_4_lut (.I0(n16371), .I1(\REG.mem_1_30 ), .I2(\REG.mem_0_30 ), 
            .I3(rd_addr_r[1]), .O(n14903));
    defparam n16371_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4117_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_1_15 ), .O(n5616));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4117_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13422_3_lut (.I0(n16692), .I1(n17628), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15546));
    defparam i13422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13423_3_lut (.I0(n17154), .I1(n16590), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15547));
    defparam i13423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14902 (.I0(rd_addr_r[2]), .I1(n15707), 
            .I2(n15731), .I3(rd_addr_r[3]), .O(n17157));
    defparam rd_addr_r_2__bdd_4_lut_14902.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15477 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_3 ), 
            .I2(\REG.mem_7_3 ), .I3(rd_addr_r[1]), .O(n17883));
    defparam rd_addr_r_0__bdd_4_lut_15477.LUT_INIT = 16'he4aa;
    SB_LUT4 n17157_bdd_4_lut (.I0(n17157), .I1(n16686), .I2(n15668), .I3(rd_addr_r[3]), 
            .O(n17160));
    defparam n17157_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13455_3_lut (.I0(n16302), .I1(n17880), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15579));
    defparam i13455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17883_bdd_4_lut (.I0(n17883), .I1(\REG.mem_5_3 ), .I2(\REG.mem_4_3 ), 
            .I3(rd_addr_r[1]), .O(n15527));
    defparam n17883_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_2_lut (.I0(n7_adj_1385), .I1(n8_adj_1383), .I2(GND_net), 
            .I3(GND_net), .O(n13844));   // src/top.v(119[12:19])
    defparam i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 wr_addr_r_5__I_0_inv_0_i6_1_lut (.I0(rp_sync2_r[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1394[5]));   // src/fifo_dc_32_lut_gen.v(212[47:78])
    defparam wr_addr_r_5__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12870_3_lut (.I0(\REG.mem_16_13 ), .I1(\REG.mem_17_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14994));
    defparam i12870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12871_3_lut (.I0(\REG.mem_18_13 ), .I1(\REG.mem_19_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14995));
    defparam i12871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12874_3_lut (.I0(\REG.mem_22_13 ), .I1(\REG.mem_23_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14998));
    defparam i12874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12873_3_lut (.I0(\REG.mem_20_13 ), .I1(\REG.mem_21_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14997));
    defparam i12873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4131_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_1_14 ), .O(n5630));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4131_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4135_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_1_13 ), .O(n5634));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4135_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4457_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_9_31 ), .O(n5956));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4457_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4456_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_9_30 ), .O(n5955));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4456_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4455_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_9_29 ), .O(n5954));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4455_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14882 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_7 ), 
            .I2(\REG.mem_11_7 ), .I3(rd_addr_r[1]), .O(n17151));
    defparam rd_addr_r_0__bdd_4_lut_14882.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15467 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_7 ), 
            .I2(\REG.mem_23_7 ), .I3(rd_addr_r[1]), .O(n17877));
    defparam rd_addr_r_0__bdd_4_lut_15467.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14209 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_3 ), 
            .I2(\REG.mem_15_3 ), .I3(rd_addr_r[1]), .O(n16365));
    defparam rd_addr_r_0__bdd_4_lut_14209.LUT_INIT = 16'he4aa;
    SB_LUT4 n17151_bdd_4_lut (.I0(n17151), .I1(\REG.mem_9_7 ), .I2(\REG.mem_8_7 ), 
            .I3(rd_addr_r[1]), .O(n17154));
    defparam n17151_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17877_bdd_4_lut (.I0(n17877), .I1(\REG.mem_21_7 ), .I2(\REG.mem_20_7 ), 
            .I3(rd_addr_r[1]), .O(n17880));
    defparam n17877_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4454_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_9_28 ), .O(n5953));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4454_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4136_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_1_12 ), .O(n5635));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4136_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4138_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_1_11 ), .O(n5637));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4138_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4150_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_1_10 ), .O(n5649));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4150_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13035_3_lut (.I0(\REG.mem_24_11 ), .I1(\REG.mem_25_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15159));
    defparam i13035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13036_3_lut (.I0(\REG.mem_26_11 ), .I1(\REG.mem_27_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15160));
    defparam i13036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13042_3_lut (.I0(\REG.mem_30_11 ), .I1(\REG.mem_31_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15166));
    defparam i13042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13041_3_lut (.I0(\REG.mem_28_11 ), .I1(\REG.mem_29_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15165));
    defparam i13041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4151_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_1_9 ), .O(n5650));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4151_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14857 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_26 ), 
            .I2(\REG.mem_27_26 ), .I3(rd_addr_r[1]), .O(n17145));
    defparam rd_addr_r_0__bdd_4_lut_14857.LUT_INIT = 16'he4aa;
    SB_LUT4 n17145_bdd_4_lut (.I0(n17145), .I1(\REG.mem_25_26 ), .I2(\REG.mem_24_26 ), 
            .I3(rd_addr_r[1]), .O(n17148));
    defparam n17145_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4453_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_9_27 ), .O(n5952));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4453_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16365_bdd_4_lut (.I0(n16365), .I1(\REG.mem_13_3 ), .I2(\REG.mem_12_3 ), 
            .I3(rd_addr_r[1]), .O(n16368));
    defparam n16365_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4152_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_1_8 ), .O(n5651));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4152_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4153_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_1_7 ), .O(n5652));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4153_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14204 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_30 ), 
            .I2(\REG.mem_7_30 ), .I3(rd_addr_r[1]), .O(n16359));
    defparam rd_addr_r_0__bdd_4_lut_14204.LUT_INIT = 16'he4aa;
    SB_LUT4 i4154_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_1_6 ), .O(n5653));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4154_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(wp_sync2_r[0]), .I1(wp_sync2_r[1]), 
            .I2(wp_sync2_r[2]), .I3(wp_sync_w[3]), .O(wp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_93 (.I0(rp_sync2_r[0]), .I1(rp_sync2_r[2]), 
            .I2(rp_sync_w[3]), .I3(rp_sync2_r[1]), .O(rp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_3_lut_4_lut_adj_93.LUT_INIT = 16'h6996;
    SB_LUT4 i4452_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_9_26 ), .O(n5951));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4452_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4451_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_9_25 ), .O(n5950));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4451_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15462 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_3 ), 
            .I2(\REG.mem_11_3 ), .I3(rd_addr_r[1]), .O(n17871));
    defparam rd_addr_r_0__bdd_4_lut_15462.LUT_INIT = 16'he4aa;
    SB_LUT4 i13350_3_lut (.I0(\REG.mem_8_22 ), .I1(\REG.mem_9_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15474));
    defparam i13350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13351_3_lut (.I0(\REG.mem_10_22 ), .I1(\REG.mem_11_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15475));
    defparam i13351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13723_3_lut (.I0(\REG.mem_14_22 ), .I1(\REG.mem_15_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15847));
    defparam i13723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13722_3_lut (.I0(\REG.mem_12_22 ), .I1(\REG.mem_13_22 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15846));
    defparam i13722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4450_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_9_24 ), .O(n5949));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4450_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4161_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_1_20 ), .O(n5660));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4161_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16359_bdd_4_lut (.I0(n16359), .I1(\REG.mem_5_30 ), .I2(\REG.mem_4_30 ), 
            .I3(rd_addr_r[1]), .O(n14906));
    defparam n16359_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17871_bdd_4_lut (.I0(n17871), .I1(\REG.mem_9_3 ), .I2(\REG.mem_8_3 ), 
            .I3(rd_addr_r[1]), .O(n15536));
    defparam n17871_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4163_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_1_24 ), .O(n5662));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4163_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15457 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_16 ), 
            .I2(\REG.mem_7_16 ), .I3(rd_addr_r[1]), .O(n17865));
    defparam rd_addr_r_0__bdd_4_lut_15457.LUT_INIT = 16'he4aa;
    SB_LUT4 n17865_bdd_4_lut (.I0(n17865), .I1(\REG.mem_5_16 ), .I2(\REG.mem_4_16 ), 
            .I3(rd_addr_r[1]), .O(n15044));
    defparam n17865_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_14862 (.I0(rd_addr_r[2]), .I1(n16506), 
            .I2(n16440), .I3(rd_addr_r[3]), .O(n17139));
    defparam rd_addr_r_2__bdd_4_lut_14862.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14199 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_30 ), 
            .I2(\REG.mem_11_30 ), .I3(rd_addr_r[1]), .O(n16353));
    defparam rd_addr_r_0__bdd_4_lut_14199.LUT_INIT = 16'he4aa;
    SB_LUT4 i4166_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_1_4 ), .O(n5665));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4166_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4167_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_1_3 ), .O(n5666));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4167_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4168_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_1_2 ), .O(n5667));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4168_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4169_3_lut_4_lut (.I0(n23), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_1_1 ), .O(n5668));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4169_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16353_bdd_4_lut (.I0(n16353), .I1(\REG.mem_9_30 ), .I2(\REG.mem_8_30 ), 
            .I3(rd_addr_r[1]), .O(n14909));
    defparam n16353_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15452 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_25 ), 
            .I2(\REG.mem_27_25 ), .I3(rd_addr_r[1]), .O(n17859));
    defparam rd_addr_r_0__bdd_4_lut_15452.LUT_INIT = 16'he4aa;
    SB_LUT4 n17139_bdd_4_lut (.I0(n17139), .I1(n16518), .I2(n16524), .I3(rd_addr_r[3]), 
            .O(n17142));
    defparam n17139_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17859_bdd_4_lut (.I0(n17859), .I1(\REG.mem_25_25 ), .I2(\REG.mem_24_25 ), 
            .I3(rd_addr_r[1]), .O(n17862));
    defparam n17859_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14194 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_30 ), 
            .I2(\REG.mem_15_30 ), .I3(rd_addr_r[1]), .O(n16347));
    defparam rd_addr_r_0__bdd_4_lut_14194.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15447 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_16 ), 
            .I2(\REG.mem_11_16 ), .I3(rd_addr_r[1]), .O(n17853));
    defparam rd_addr_r_0__bdd_4_lut_15447.LUT_INIT = 16'he4aa;
    SB_LUT4 n16347_bdd_4_lut (.I0(n16347), .I1(\REG.mem_13_30 ), .I2(\REG.mem_12_30 ), 
            .I3(rd_addr_r[1]), .O(n14912));
    defparam n16347_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17853_bdd_4_lut (.I0(n17853), .I1(\REG.mem_9_16 ), .I2(\REG.mem_8_16 ), 
            .I3(rd_addr_r[1]), .O(n15050));
    defparam n17853_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14189 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_30 ), 
            .I2(\REG.mem_19_30 ), .I3(rd_addr_r[1]), .O(n16341));
    defparam rd_addr_r_0__bdd_4_lut_14189.LUT_INIT = 16'he4aa;
    SB_LUT4 n16341_bdd_4_lut (.I0(n16341), .I1(\REG.mem_17_30 ), .I2(\REG.mem_16_30 ), 
            .I3(rd_addr_r[1]), .O(n16344));
    defparam n16341_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i6_2_lut_3_lut (.I0(DEBUG_5_c), .I1(dc32_fifo_full), 
            .I2(\wr_addr_r[0] ), .I3(GND_net), .O(n6_adj_1378));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i6_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_15512 (.I0(rd_addr_r[1]), .I1(n15045), 
            .I2(n15046), .I3(rd_addr_r[2]), .O(n17847));
    defparam rd_addr_r_1__bdd_4_lut_15512.LUT_INIT = 16'he4aa;
    SB_LUT4 i4449_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_9_23 ), .O(n5948));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4449_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4448_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_9_22 ), .O(n5947));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4448_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14852 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_1 ), 
            .I2(\REG.mem_7_1 ), .I3(rd_addr_r[1]), .O(n17127));
    defparam rd_addr_r_0__bdd_4_lut_14852.LUT_INIT = 16'he4aa;
    SB_LUT4 i4969_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[31]), 
            .I3(\REG.mem_25_31 ), .O(n6468));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4969_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4968_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[30]), 
            .I3(\REG.mem_25_30 ), .O(n6467));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4968_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4967_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[29]), 
            .I3(\REG.mem_25_29 ), .O(n6466));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4967_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i7_2_lut_3_lut (.I0(DEBUG_5_c), .I1(dc32_fifo_full), 
            .I2(\wr_addr_r[0] ), .I3(GND_net), .O(n7_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i7_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut (.I0(rp_sync2_r[2]), .I1(rp_sync_w[3]), .I2(rp_sync2_r[1]), 
            .I3(GND_net), .O(rp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 rd_addr_nxt_c_5__I_0_138_i4_2_lut (.I0(\rd_addr_nxt_c_5__N_573[3] ), 
            .I1(\rd_addr_nxt_c_5__N_573[4] ), .I2(GND_net), .I3(GND_net), 
            .O(rd_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(504[28:66])
    defparam rd_addr_nxt_c_5__I_0_138_i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 EnabledDecoder_2_i12_2_lut_3_lut_4_lut (.I0(wr_fifo_en_w), .I1(\wr_addr_r[0] ), 
            .I2(wr_addr_r[1]), .I3(wr_addr_r[2]), .O(n12_adj_1391));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i12_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_adj_94 (.I0(wp_sync2_r[1]), .I1(wp_sync2_r[2]), 
            .I2(wp_sync_w[3]), .I3(GND_net), .O(wp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_94.LUT_INIT = 16'h9696;
    SB_LUT4 i12840_3_lut (.I0(\REG.mem_0_8 ), .I1(\REG.mem_1_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14964));
    defparam i12840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12841_3_lut (.I0(\REG.mem_2_8 ), .I1(\REG.mem_3_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14965));
    defparam i12841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13734_3_lut (.I0(\REG.mem_0_5 ), .I1(\REG.mem_1_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15858));
    defparam i13734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13735_3_lut (.I0(\REG.mem_2_5 ), .I1(\REG.mem_3_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15859));
    defparam i13735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13753_3_lut (.I0(\REG.mem_6_5 ), .I1(\REG.mem_7_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15877));
    defparam i13753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13752_3_lut (.I0(\REG.mem_4_5 ), .I1(\REG.mem_5_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15876));
    defparam i13752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13453_3_lut (.I0(\REG.mem_6_8 ), .I1(\REG.mem_7_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15577));
    defparam i13453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13452_3_lut (.I0(\REG.mem_4_8 ), .I1(\REG.mem_5_8 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15576));
    defparam i13452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_95 (.I0(wp_sync2_r[3]), .I1(wp_sync2_r[5]), 
            .I2(wp_sync2_r[4]), .I3(GND_net), .O(wp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_95.LUT_INIT = 16'h9696;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14184 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_30 ), 
            .I2(\REG.mem_23_30 ), .I3(rd_addr_r[1]), .O(n16323));
    defparam rd_addr_r_0__bdd_4_lut_14184.LUT_INIT = 16'he4aa;
    SB_LUT4 n17847_bdd_4_lut (.I0(n17847), .I1(n15040), .I2(n15039), .I3(rd_addr_r[2]), 
            .O(n15055));
    defparam n17847_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16323_bdd_4_lut (.I0(n16323), .I1(\REG.mem_21_30 ), .I2(\REG.mem_20_30 ), 
            .I3(rd_addr_r[1]), .O(n16326));
    defparam n16323_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4966_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[28]), 
            .I3(\REG.mem_25_28 ), .O(n6465));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4966_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15442 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_21 ), 
            .I2(\REG.mem_7_21 ), .I3(rd_addr_r[1]), .O(n17841));
    defparam rd_addr_r_0__bdd_4_lut_15442.LUT_INIT = 16'he4aa;
    SB_LUT4 i4447_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_9_21 ), .O(n5946));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4447_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4965_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[27]), 
            .I3(\REG.mem_25_27 ), .O(n6464));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4965_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4446_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_9_20 ), .O(n5945));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4446_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17841_bdd_4_lut (.I0(n17841), .I1(\REG.mem_5_21 ), .I2(\REG.mem_4_21 ), 
            .I3(rd_addr_r[1]), .O(n15542));
    defparam n17841_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12624_3_lut (.I0(\REG.mem_24_14 ), .I1(\REG.mem_25_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14748));
    defparam i12624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12625_3_lut (.I0(\REG.mem_26_14 ), .I1(\REG.mem_27_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14749));
    defparam i12625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4964_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[26]), 
            .I3(\REG.mem_25_26 ), .O(n6463));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4964_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4445_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_9_19 ), .O(n5944));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4445_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4963_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[25]), 
            .I3(\REG.mem_25_25 ), .O(n6462));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4963_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13485_3_lut (.I0(\REG.mem_8_26 ), .I1(\REG.mem_9_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15609));
    defparam i13485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13486_3_lut (.I0(\REG.mem_10_26 ), .I1(\REG.mem_11_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15610));
    defparam i13486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12640_3_lut (.I0(\REG.mem_30_14 ), .I1(\REG.mem_31_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14764));
    defparam i12640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12639_3_lut (.I0(\REG.mem_28_14 ), .I1(\REG.mem_29_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14763));
    defparam i12639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13528_3_lut (.I0(\REG.mem_14_26 ), .I1(\REG.mem_15_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15652));
    defparam i13528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13527_3_lut (.I0(\REG.mem_12_26 ), .I1(\REG.mem_13_26 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15651));
    defparam i13527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4444_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_9_18 ), .O(n5943));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4444_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4443_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_9_17 ), .O(n5942));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4443_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4442_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_9_16 ), .O(n5941));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4442_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i28_2_lut_4_lut (.I0(n7_c), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n28_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i28_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i4962_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[24]), 
            .I3(\REG.mem_25_24 ), .O(n6461));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4962_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4961_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[23]), 
            .I3(\REG.mem_25_23 ), .O(n6460));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4961_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4441_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_9_15 ), .O(n5940));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4441_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4440_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_9_14 ), .O(n5939));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4440_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4960_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[22]), 
            .I3(\REG.mem_25_22 ), .O(n6459));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4960_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4959_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[21]), 
            .I3(\REG.mem_25_21 ), .O(n6458));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4959_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4958_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[20]), 
            .I3(\REG.mem_25_20 ), .O(n6457));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4958_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4439_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_9_13 ), .O(n5938));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4439_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17127_bdd_4_lut (.I0(n17127), .I1(\REG.mem_5_1 ), .I2(\REG.mem_4_1 ), 
            .I3(rd_addr_r[1]), .O(n15782));
    defparam n17127_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14837 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_9 ), 
            .I2(\REG.mem_3_9 ), .I3(rd_addr_r[1]), .O(n17121));
    defparam rd_addr_r_0__bdd_4_lut_14837.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14169 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_17 ), 
            .I2(\REG.mem_23_17 ), .I3(rd_addr_r[1]), .O(n16317));
    defparam rd_addr_r_0__bdd_4_lut_14169.LUT_INIT = 16'he4aa;
    SB_LUT4 i4438_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_9_12 ), .O(n5937));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4438_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16317_bdd_4_lut (.I0(n16317), .I1(\REG.mem_21_17 ), .I2(\REG.mem_20_17 ), 
            .I3(rd_addr_r[1]), .O(n16320));
    defparam n16317_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17121_bdd_4_lut (.I0(n17121), .I1(\REG.mem_1_9 ), .I2(\REG.mem_0_9 ), 
            .I3(rd_addr_r[1]), .O(n15251));
    defparam n17121_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4957_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[19]), 
            .I3(\REG.mem_25_19 ), .O(n6456));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4957_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15432 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_25 ), 
            .I2(\REG.mem_31_25 ), .I3(rd_addr_r[1]), .O(n17829));
    defparam rd_addr_r_0__bdd_4_lut_15432.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i14_2_lut_3_lut_4_lut (.I0(wr_fifo_en_w), .I1(\wr_addr_r[0] ), 
            .I2(wr_addr_r[1]), .I3(wr_addr_r[2]), .O(n14));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i14_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i4956_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[18]), 
            .I3(\REG.mem_25_18 ), .O(n6455));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4956_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14832 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_1 ), 
            .I2(\REG.mem_11_1 ), .I3(rd_addr_r[1]), .O(n17109));
    defparam rd_addr_r_0__bdd_4_lut_14832.LUT_INIT = 16'he4aa;
    SB_LUT4 i4437_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[11]), 
            .I3(\REG.mem_9_11 ), .O(n5936));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4437_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n16209_bdd_4_lut (.I0(n16209), .I1(n15230), .I2(n15185), .I3(rd_addr_r[3]), 
            .O(n16212));
    defparam n16209_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n17109_bdd_4_lut (.I0(n17109), .I1(\REG.mem_9_1 ), .I2(\REG.mem_8_1 ), 
            .I3(rd_addr_r[1]), .O(n15788));
    defparam n17109_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4955_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[17]), 
            .I3(\REG.mem_25_17 ), .O(n6454));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4955_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4436_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[10]), 
            .I3(\REG.mem_9_10 ), .O(n5935));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4436_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4954_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[16]), 
            .I3(\REG.mem_25_16 ), .O(n6453));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4954_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i16_2_lut_3_lut_4_lut (.I0(wr_fifo_en_w), .I1(\wr_addr_r[0] ), 
            .I2(wr_addr_r[1]), .I3(wr_addr_r[2]), .O(n16));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i16_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i34_2_lut_3_lut_4_lut (.I0(n6_adj_1378), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n34));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i34_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4435_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[9]), 
            .I3(\REG.mem_9_9 ), .O(n5934));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4435_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13396_3_lut (.I0(n17862), .I1(n17832), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n15520));
    defparam i13396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n17829_bdd_4_lut (.I0(n17829), .I1(\REG.mem_29_25 ), .I2(\REG.mem_28_25 ), 
            .I3(rd_addr_r[1]), .O(n17832));
    defparam n17829_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_5__I_0_135_inv_0_i4_1_lut (.I0(rd_addr_r[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_5__I_0_135_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 EnabledDecoder_2_i49_2_lut_3_lut (.I0(n16), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n27));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i49_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i4434_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[8]), 
            .I3(\REG.mem_9_8 ), .O(n5933));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4434_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12660_3_lut (.I0(\REG.mem_8_19 ), .I1(\REG.mem_9_19 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14784));
    defparam i12660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12661_3_lut (.I0(\REG.mem_10_19 ), .I1(\REG.mem_11_19 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14785));
    defparam i12661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12667_3_lut (.I0(\REG.mem_14_19 ), .I1(\REG.mem_15_19 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14791));
    defparam i12667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4953_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[15]), 
            .I3(\REG.mem_25_15 ), .O(n6452));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4953_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12666_3_lut (.I0(\REG.mem_12_19 ), .I1(\REG.mem_13_19 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n14790));
    defparam i12666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14085 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_4 ), 
            .I2(\REG.mem_31_4 ), .I3(rd_addr_r[1]), .O(n16203));
    defparam rd_addr_r_0__bdd_4_lut_14085.LUT_INIT = 16'he4aa;
    SB_LUT4 i4433_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[7]), 
            .I3(\REG.mem_9_7 ), .O(n5932));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4433_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4432_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[6]), 
            .I3(\REG.mem_9_6 ), .O(n5931));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4432_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15422 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_8 ), 
            .I2(\REG.mem_31_8 ), .I3(rd_addr_r[1]), .O(n17823));
    defparam rd_addr_r_0__bdd_4_lut_15422.LUT_INIT = 16'he4aa;
    SB_LUT4 i4431_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[5]), 
            .I3(\REG.mem_9_5 ), .O(n5930));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4431_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4430_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[4]), 
            .I3(\REG.mem_9_4 ), .O(n5929));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4430_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4429_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[3]), 
            .I3(\REG.mem_9_3 ), .O(n5928));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4429_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n17823_bdd_4_lut (.I0(n17823), .I1(\REG.mem_29_8 ), .I2(\REG.mem_28_8 ), 
            .I3(rd_addr_r[1]), .O(n17826));
    defparam n17823_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4428_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[2]), 
            .I3(\REG.mem_9_2 ), .O(n5927));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4428_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4427_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[1]), 
            .I3(\REG.mem_9_1 ), .O(n5926));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4427_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4952_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[14]), 
            .I3(\REG.mem_25_14 ), .O(n6451));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4952_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12966_3_lut (.I0(\REG.mem_0_11 ), .I1(\REG.mem_1_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15090));
    defparam i12966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12967_3_lut (.I0(\REG.mem_2_11 ), .I1(\REG.mem_3_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15091));
    defparam i12967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12985_3_lut (.I0(\REG.mem_6_11 ), .I1(\REG.mem_7_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15109));
    defparam i12985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12984_3_lut (.I0(\REG.mem_4_11 ), .I1(\REG.mem_5_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n15108));
    defparam i12984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i27_2_lut_3_lut_4_lut (.I0(n6_adj_1378), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[3]), .O(n27_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i27_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i4951_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[13]), 
            .I3(\REG.mem_25_13 ), .O(n6450));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4951_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15417 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_27 ), 
            .I2(\REG.mem_15_27 ), .I3(rd_addr_r[1]), .O(n17817));
    defparam rd_addr_r_0__bdd_4_lut_15417.LUT_INIT = 16'he4aa;
    SB_LUT4 n17817_bdd_4_lut (.I0(n17817), .I1(\REG.mem_13_27 ), .I2(\REG.mem_12_27 ), 
            .I3(rd_addr_r[1]), .O(n15077));
    defparam n17817_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n16203_bdd_4_lut (.I0(n16203), .I1(\REG.mem_29_4 ), .I2(\REG.mem_28_4 ), 
            .I3(rd_addr_r[1]), .O(n16206));
    defparam n16203_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i48_2_lut_3_lut (.I0(n16), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n11));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i48_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i47_2_lut_3_lut (.I0(n14), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n28));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i47_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_14822 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_15 ), 
            .I2(\REG.mem_7_15 ), .I3(rd_addr_r[1]), .O(n17097));
    defparam rd_addr_r_0__bdd_4_lut_14822.LUT_INIT = 16'he4aa;
    SB_LUT4 i4426_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[0]), 
            .I3(\REG.mem_9_0 ), .O(n5925));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4426_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_15412 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_20 ), 
            .I2(\REG.mem_3_20 ), .I3(rd_addr_r[1]), .O(n17811));
    defparam rd_addr_r_0__bdd_4_lut_15412.LUT_INIT = 16'he4aa;
    SB_LUT4 i4950_3_lut_4_lut (.I0(n22_c), .I1(wr_addr_r[4]), .I2(dc32_fifo_data_in[12]), 
            .I3(\REG.mem_25_12 ), .O(n6449));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4950_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n17097_bdd_4_lut (.I0(n17097), .I1(\REG.mem_5_15 ), .I2(\REG.mem_4_15 ), 
            .I3(rd_addr_r[1]), .O(n15794));
    defparam n17097_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module clock
//

module clock (GND_net, VCC_net, ICE_SYSCLK_c, pll_clk_unbuf) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    input ICE_SYSCLK_c;
    output pll_clk_unbuf;
    
    
    SB_PLL40_CORE pll_config (.REFERENCECLK(ICE_SYSCLK_c), .PLLOUTGLOBAL(pll_clk_unbuf), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=15, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/top.v(222[7] 228[3])
    defparam pll_config.FEEDBACK_PATH = "SIMPLE";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll_config.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll_config.FDA_FEEDBACK = 0;
    defparam pll_config.FDA_RELATIVE = 0;
    defparam pll_config.PLLOUT_SELECT = "GENCLK";
    defparam pll_config.DIVR = 4'b0001;
    defparam pll_config.DIVF = 7'b1010010;
    defparam pll_config.DIVQ = 3'b100;
    defparam pll_config.FILTER_RANGE = 3'b001;
    defparam pll_config.ENABLE_ICEGATE = 1'b0;
    defparam pll_config.TEST_MODE = 1'b0;
    defparam pll_config.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module spi
//

module spi (SLM_CLK_c, SOUT_c, n5025, \rx_shift_reg[0] , n4999, SDAT_c_15, 
            n7013, rx_buf_byte, n7012, n7011, n7010, n7009, n7008, 
            n7007, n7006, \rx_shift_reg[7] , n7005, \rx_shift_reg[6] , 
            n7004, \rx_shift_reg[5] , n7003, \rx_shift_reg[4] , n7002, 
            \rx_shift_reg[3] , n7001, \rx_shift_reg[2] , n7000, \rx_shift_reg[1] , 
            n14116, VCC_net, \tx_shift_reg[0] , multi_byte_spi_trans_flag_r, 
            GND_net, n2555, spi_start_transfer_r, tx_addr_byte, SEN_c_1, 
            spi_rx_byte_ready, SCK_c_0, n5636, \tx_data_byte[7] , \tx_data_byte[6] , 
            \tx_data_byte[5] , \tx_data_byte[4] , \tx_data_byte[3] , \tx_data_byte[2] , 
            \tx_data_byte[1] , n4086) /* synthesis syn_module_defined=1 */ ;
    input SLM_CLK_c;
    input SOUT_c;
    output n5025;
    output \rx_shift_reg[0] ;
    output n4999;
    output SDAT_c_15;
    input n7013;
    output [7:0]rx_buf_byte;
    input n7012;
    input n7011;
    input n7010;
    input n7009;
    input n7008;
    input n7007;
    input n7006;
    output \rx_shift_reg[7] ;
    input n7005;
    output \rx_shift_reg[6] ;
    input n7004;
    output \rx_shift_reg[5] ;
    input n7003;
    output \rx_shift_reg[4] ;
    input n7002;
    output \rx_shift_reg[3] ;
    input n7001;
    output \rx_shift_reg[2] ;
    input n7000;
    output \rx_shift_reg[1] ;
    input n14116;
    input VCC_net;
    output \tx_shift_reg[0] ;
    input multi_byte_spi_trans_flag_r;
    input GND_net;
    output n2555;
    input spi_start_transfer_r;
    input [7:0]tx_addr_byte;
    output SEN_c_1;
    output spi_rx_byte_ready;
    output SCK_c_0;
    input n5636;
    input \tx_data_byte[7] ;
    input \tx_data_byte[6] ;
    input \tx_data_byte[5] ;
    input \tx_data_byte[4] ;
    input \tx_data_byte[3] ;
    input \tx_data_byte[2] ;
    input \tx_data_byte[1] ;
    output n4086;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [7:0]n315;
    
    wire n5157;
    wire [7:0]multi_byte_counter;   // src/spi.v(68[11:29])
    
    wire n5428;
    wire [3:0]state_3__N_1123;
    
    wire n18032;
    wire [3:0]state;   // src/spi.v(71[11:16])
    wire [9:0]n45;
    
    wire n5059;
    wire [9:0]counter;   // src/spi.v(69[11:18])
    
    wire n5583;
    wire [15:0]n2556;
    
    wire n3, CS_N_1193, n3_adj_1367, n13785, n13784, n13783, n13782;
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    
    wire n13781, n13780, n13779, n13778, n13777, n4, n34;
    wire [7:0]n2634;
    
    wire n13734, n24, n35, n16, n14, n10, n14_adj_1368, n15909, 
        n15976, n34_adj_1369;
    wire [2:0]n1116;
    
    wire n37, n4919, n4922, n14527, n14526, n19, n13733, n13732, 
        n13731, n13730, n13729, n13728, n5381, n14659, n5189, 
        n5038, n6, n3787, n4657, n4_adj_1370, n31, n14708, n14674, 
        n15910, n7, n12, n15951, n15952, n24_adj_1371, n15969, 
        n14678, n21, n7_adj_1372, n22, n14525, n3_adj_1373, n10087, 
        n15962;
    
    SB_DFFESR multi_byte_counter_i6 (.Q(multi_byte_counter[6]), .C(SLM_CLK_c), 
            .E(n5157), .D(n315[6]), .R(n5428));   // src/spi.v(76[8] 221[4])
    SB_DFFESS multi_byte_counter_i5 (.Q(multi_byte_counter[5]), .C(SLM_CLK_c), 
            .E(n5157), .D(n315[5]), .S(n5428));   // src/spi.v(76[8] 221[4])
    SB_DFFE rx_shift_reg_i0 (.Q(\rx_shift_reg[0] ), .C(SLM_CLK_c), .E(n5025), 
            .D(SOUT_c));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n18032), .D(state_3__N_1123[0]));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_1469__i9 (.Q(counter[9]), .C(SLM_CLK_c), .E(n5059), 
            .D(n45[9]), .R(n5583));   // src/spi.v(183[28:41])
    SB_DFFESS counter_1469__i8 (.Q(counter[8]), .C(SLM_CLK_c), .E(n5059), 
            .D(n45[8]), .S(n5583));   // src/spi.v(183[28:41])
    SB_DFFE tx_shift_reg_i0_i15 (.Q(SDAT_c_15), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[15]));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_1469__i7 (.Q(counter[7]), .C(SLM_CLK_c), .E(n5059), 
            .D(n45[7]), .R(n5583));   // src/spi.v(183[28:41])
    SB_DFF Rx_Recv_Byte_i7 (.Q(rx_buf_byte[7]), .C(SLM_CLK_c), .D(n7013));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i6 (.Q(rx_buf_byte[6]), .C(SLM_CLK_c), .D(n7012));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i5 (.Q(rx_buf_byte[5]), .C(SLM_CLK_c), .D(n7011));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i4 (.Q(rx_buf_byte[4]), .C(SLM_CLK_c), .D(n7010));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i3 (.Q(rx_buf_byte[3]), .C(SLM_CLK_c), .D(n7009));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i2 (.Q(rx_buf_byte[2]), .C(SLM_CLK_c), .D(n7008));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i1 (.Q(rx_buf_byte[1]), .C(SLM_CLK_c), .D(n7007));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i7 (.Q(\rx_shift_reg[7] ), .C(SLM_CLK_c), .D(n7006));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i6 (.Q(\rx_shift_reg[6] ), .C(SLM_CLK_c), .D(n7005));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i5 (.Q(\rx_shift_reg[5] ), .C(SLM_CLK_c), .D(n7004));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i4 (.Q(\rx_shift_reg[4] ), .C(SLM_CLK_c), .D(n7003));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i3 (.Q(\rx_shift_reg[3] ), .C(SLM_CLK_c), .D(n7002));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i2 (.Q(\rx_shift_reg[2] ), .C(SLM_CLK_c), .D(n7001));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i1 (.Q(\rx_shift_reg[1] ), .C(SLM_CLK_c), .D(n7000));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i0 (.Q(\tx_shift_reg[0] ), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n14116));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_1469__i6 (.Q(counter[6]), .C(SLM_CLK_c), .E(n5059), 
            .D(n45[6]), .R(n5583));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1469__i5 (.Q(counter[5]), .C(SLM_CLK_c), .E(n5059), 
            .D(n45[5]), .R(n5583));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1469__i4 (.Q(counter[4]), .C(SLM_CLK_c), .E(n5059), 
            .D(n45[4]), .R(n5583));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1469__i3 (.Q(counter[3]), .C(SLM_CLK_c), .E(n5059), 
            .D(n45[3]), .R(n5583));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1469__i2 (.Q(counter[2]), .C(SLM_CLK_c), .E(n5059), 
            .D(n45[2]), .R(n5583));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1469__i0 (.Q(counter[0]), .C(SLM_CLK_c), .E(n5059), 
            .D(n45[0]), .R(n5583));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1469__i1 (.Q(counter[1]), .C(SLM_CLK_c), .E(n5059), 
            .D(n45[1]), .R(n5583));   // src/spi.v(183[28:41])
    SB_DFFESR multi_byte_counter_i0 (.Q(multi_byte_counter[0]), .C(SLM_CLK_c), 
            .E(n5157), .D(n315[0]), .R(n5428));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_56_Mux_1_i3_3_lut_3_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(GND_net), .O(n3));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i3_3_lut_3_lut.LUT_INIT = 16'h3e3e;
    SB_LUT4 mux_56_Mux_0_i3_4_lut_4_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(CS_N_1193), .O(n3_adj_1367));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_0_i3_4_lut_4_lut.LUT_INIT = 16'h31c1;
    SB_LUT4 counter_1469_add_4_11_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[9]), 
            .I3(n13785), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1469_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1469_add_4_10_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[8]), 
            .I3(n13784), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1469_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1469_add_4_10 (.CI(n13784), .I0(VCC_net), .I1(counter[8]), 
            .CO(n13785));
    SB_LUT4 counter_1469_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[7]), 
            .I3(n13783), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1469_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1469_add_4_9 (.CI(n13783), .I0(VCC_net), .I1(counter[7]), 
            .CO(n13784));
    SB_LUT4 counter_1469_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[6]), 
            .I3(n13782), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1469_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFE tx_shift_reg_i0_i1 (.Q(tx_shift_reg[1]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[1]));   // src/spi.v(76[8] 221[4])
    SB_CARRY counter_1469_add_4_8 (.CI(n13782), .I0(VCC_net), .I1(counter[6]), 
            .CO(n13783));
    SB_LUT4 counter_1469_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[5]), 
            .I3(n13781), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1469_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1469_add_4_7 (.CI(n13781), .I0(VCC_net), .I1(counter[5]), 
            .CO(n13782));
    SB_LUT4 counter_1469_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[4]), 
            .I3(n13780), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1469_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFE tx_shift_reg_i0_i2 (.Q(tx_shift_reg[2]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i3 (.Q(tx_shift_reg[3]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[3]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i4 (.Q(tx_shift_reg[4]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[4]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i5 (.Q(tx_shift_reg[5]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[5]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i6 (.Q(tx_shift_reg[6]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[6]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i7 (.Q(tx_shift_reg[7]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[7]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i8 (.Q(tx_shift_reg[8]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[8]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i9 (.Q(tx_shift_reg[9]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[9]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i10 (.Q(tx_shift_reg[10]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[10]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i11 (.Q(tx_shift_reg[11]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[11]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i12 (.Q(tx_shift_reg[12]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[12]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i13 (.Q(tx_shift_reg[13]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[13]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i14 (.Q(tx_shift_reg[14]), .C(SLM_CLK_c), .E(n4999), 
            .D(n2556[14]));   // src/spi.v(76[8] 221[4])
    SB_CARRY counter_1469_add_4_6 (.CI(n13780), .I0(VCC_net), .I1(counter[4]), 
            .CO(n13781));
    SB_LUT4 counter_1469_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[3]), 
            .I3(n13779), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1469_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1469_add_4_5 (.CI(n13779), .I0(VCC_net), .I1(counter[3]), 
            .CO(n13780));
    SB_LUT4 counter_1469_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[2]), 
            .I3(n13778), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1469_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1469_add_4_4 (.CI(n13778), .I0(VCC_net), .I1(counter[2]), 
            .CO(n13779));
    SB_LUT4 counter_1469_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[1]), 
            .I3(n13777), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1469_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1469_add_4_3 (.CI(n13777), .I0(VCC_net), .I1(counter[1]), 
            .CO(n13778));
    SB_LUT4 counter_1469_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1469_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1469_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n13777));
    SB_LUT4 i1_4_lut (.I0(counter[3]), .I1(n4), .I2(counter[4]), .I3(n34), 
            .O(n2555));
    defparam i1_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 add_1300_9_lut (.I0(GND_net), .I1(multi_byte_counter[7]), .I2(n2634[6]), 
            .I3(n13734), .O(n315[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1300_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR multi_byte_counter_i4 (.Q(multi_byte_counter[4]), .C(SLM_CLK_c), 
            .E(n5157), .D(n315[4]), .R(n5428));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i3 (.Q(multi_byte_counter[3]), .C(SLM_CLK_c), 
            .E(n5157), .D(n315[3]), .R(n5428));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i30_4_lut (.I0(spi_start_transfer_r), .I1(state[3]), .I2(state[1]), 
            .I3(state[0]), .O(n24));   // src/spi.v(88[9] 219[16])
    defparam i30_4_lut.LUT_INIT = 16'hcfc1;
    SB_LUT4 i1_4_lut_adj_74 (.I0(n35), .I1(state[3]), .I2(counter[4]), 
            .I3(state[1]), .O(n16));   // src/spi.v(88[9] 219[16])
    defparam i1_4_lut_adj_74.LUT_INIT = 16'hf5c4;
    SB_DFFESR multi_byte_counter_i2 (.Q(multi_byte_counter[2]), .C(SLM_CLK_c), 
            .E(n5157), .D(n315[2]), .R(n5428));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_1276_i16_3_lut (.I0(tx_addr_byte[7]), .I1(tx_shift_reg[14]), 
            .I2(n2555), .I3(GND_net), .O(n2556[15]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), .I3(GND_net), 
            .O(n14));   // src/spi.v(88[9] 219[16])
    defparam i1_3_lut.LUT_INIT = 16'hcdcd;
    SB_LUT4 i2_2_lut (.I0(multi_byte_counter[2]), .I1(multi_byte_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // src/spi.v(208[21:52])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(multi_byte_counter[3]), .I1(multi_byte_counter[1]), 
            .I2(multi_byte_counter[5]), .I3(multi_byte_counter[7]), .O(n14_adj_1368));   // src/spi.v(208[21:52])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(multi_byte_counter[0]), .I1(n14_adj_1368), .I2(n10), 
            .I3(multi_byte_counter[6]), .O(n2634[6]));   // src/spi.v(208[21:52])
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_DFFESR multi_byte_counter_i1 (.Q(multi_byte_counter[1]), .C(SLM_CLK_c), 
            .E(n5157), .D(n315[1]), .R(n5428));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i13864_3_lut (.I0(state[0]), .I1(state[2]), .I2(CS_N_1193), 
            .I3(GND_net), .O(n15909));
    defparam i13864_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i13929_3_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), 
            .I3(GND_net), .O(n15976));
    defparam i13929_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i65_3_lut (.I0(n14), .I1(n15909), .I2(state[1]), .I3(GND_net), 
            .O(n34_adj_1369));
    defparam i65_3_lut.LUT_INIT = 16'hc5c5;
    SB_DFF byte_recv_92_i2 (.Q(SEN_c_1), .C(SLM_CLK_c), .D(n1116[1]));   // src/spi.v(88[9] 219[16])
    SB_LUT4 i66_4_lut (.I0(n15976), .I1(n2634[6]), .I2(state[1]), .I3(state[3]), 
            .O(n37));
    defparam i66_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut_adj_75 (.I0(state[3]), .I1(n37), .I2(n34_adj_1369), 
            .I3(n4919), .O(n5583));
    defparam i1_4_lut_adj_75.LUT_INIT = 16'h50dc;
    SB_LUT4 i13995_4_lut (.I0(state[3]), .I1(state[1]), .I2(n4922), .I3(n14), 
            .O(n5059));   // src/spi.v(88[9] 219[16])
    defparam i13995_4_lut.LUT_INIT = 16'h4c5f;
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n14527), .D(state_3__N_1123[1]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n14526), .D(state_3__N_1123[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(n19), .D(state_3__N_1123[3]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 add_1300_8_lut (.I0(GND_net), .I1(multi_byte_counter[6]), .I2(n2634[6]), 
            .I3(n13733), .O(n315[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1300_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF byte_recv_92_i3 (.Q(spi_rx_byte_ready), .C(SLM_CLK_c), .D(n1116[2]));   // src/spi.v(88[9] 219[16])
    SB_DFF byte_recv_92_i1 (.Q(SCK_c_0), .C(SLM_CLK_c), .D(n1116[0]));   // src/spi.v(88[9] 219[16])
    SB_CARRY add_1300_8 (.CI(n13733), .I0(multi_byte_counter[6]), .I1(n2634[6]), 
            .CO(n13734));
    SB_LUT4 add_1300_7_lut (.I0(GND_net), .I1(multi_byte_counter[5]), .I2(n2634[6]), 
            .I3(n13732), .O(n315[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1300_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1300_7 (.CI(n13732), .I0(multi_byte_counter[5]), .I1(n2634[6]), 
            .CO(n13733));
    SB_LUT4 add_1300_6_lut (.I0(GND_net), .I1(multi_byte_counter[4]), .I2(n2634[6]), 
            .I3(n13731), .O(n315[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1300_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1300_6 (.CI(n13731), .I0(multi_byte_counter[4]), .I1(n2634[6]), 
            .CO(n13732));
    SB_LUT4 add_1300_5_lut (.I0(GND_net), .I1(multi_byte_counter[3]), .I2(n2634[6]), 
            .I3(n13730), .O(n315[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1300_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1300_5 (.CI(n13730), .I0(multi_byte_counter[3]), .I1(n2634[6]), 
            .CO(n13731));
    SB_LUT4 add_1300_4_lut (.I0(GND_net), .I1(multi_byte_counter[2]), .I2(n2634[6]), 
            .I3(n13729), .O(n315[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1300_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1300_4 (.CI(n13729), .I0(multi_byte_counter[2]), .I1(n2634[6]), 
            .CO(n13730));
    SB_LUT4 add_1300_3_lut (.I0(GND_net), .I1(multi_byte_counter[1]), .I2(n2634[6]), 
            .I3(n13728), .O(n315[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1300_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1300_3 (.CI(n13728), .I0(multi_byte_counter[1]), .I1(n2634[6]), 
            .CO(n13729));
    SB_LUT4 add_1300_2_lut (.I0(GND_net), .I1(multi_byte_counter[0]), .I2(n2634[6]), 
            .I3(GND_net), .O(n315[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1300_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1300_2 (.CI(GND_net), .I0(multi_byte_counter[0]), .I1(n2634[6]), 
            .CO(n13728));
    SB_LUT4 i12491_2_lut (.I0(state[3]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5381));
    defparam i12491_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12537_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n14659));
    defparam i12537_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(CS_N_1193), .I1(state[3]), .I2(state[2]), .I3(n14659), 
            .O(n5189));
    defparam i3_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i3_4_lut_adj_76 (.I0(spi_start_transfer_r), .I1(state[1]), .I2(state[0]), 
            .I3(n5381), .O(n5038));
    defparam i3_4_lut_adj_76.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(state[3]), .I1(n5038), .I2(CS_N_1193), .I3(state[0]), 
            .O(n6));
    defparam i2_4_lut.LUT_INIT = 16'hccc4;
    SB_LUT4 i2302_2_lut (.I0(state[1]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n3787));   // src/spi.v(88[9] 219[16])
    defparam i2302_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_77 (.I0(n3787), .I1(n6), .I2(n5189), .I3(state[3]), 
            .O(n18032));
    defparam i3_4_lut_adj_77.LUT_INIT = 16'h40c0;
    SB_LUT4 i3883_3_lut (.I0(n3_adj_1367), .I1(state[0]), .I2(n5381), 
            .I3(GND_net), .O(state_3__N_1123[0]));   // src/spi.v(88[9] 219[16])
    defparam i3883_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i2_3_lut (.I0(counter[2]), .I1(counter[1]), .I2(counter[0]), 
            .I3(GND_net), .O(n34));   // src/spi.v(183[28:41])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut (.I0(state[0]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n4919));   // src/spi.v(88[9] 219[16])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13997_3_lut (.I0(counter[4]), .I1(n35), .I2(n4657), .I3(GND_net), 
            .O(n5025));   // src/spi.v(88[9] 219[16])
    defparam i13997_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_adj_78 (.I0(state[3]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_1370));
    defparam i1_2_lut_adj_78.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_79 (.I0(counter[3]), .I1(counter[1]), .I2(counter[2]), 
            .I3(GND_net), .O(n31));
    defparam i2_3_lut_adj_79.LUT_INIT = 16'hfefe;
    SB_LUT4 i12585_4_lut (.I0(n31), .I1(counter[8]), .I2(counter[7]), 
            .I3(counter[9]), .O(n14708));
    defparam i12585_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12552_2_lut (.I0(counter[5]), .I1(counter[6]), .I2(GND_net), 
            .I3(GND_net), .O(n14674));
    defparam i12552_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_80 (.I0(n14674), .I1(counter[0]), .I2(n14708), 
            .I3(counter[4]), .O(CS_N_1193));
    defparam i2_4_lut_adj_80.LUT_INIT = 16'h0004;
    SB_LUT4 i3929_2_lut (.I0(n5157), .I1(state[3]), .I2(GND_net), .I3(GND_net), 
            .O(n5428));   // src/spi.v(76[8] 221[4])
    defparam i3929_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13873_3_lut (.I0(state[3]), .I1(CS_N_1193), .I2(state[2]), 
            .I3(GND_net), .O(n15910));
    defparam i13873_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_4_lut_adj_81 (.I0(state[1]), .I1(n4_adj_1370), .I2(n15910), 
            .I3(state[0]), .O(n5157));
    defparam i1_4_lut_adj_81.LUT_INIT = 16'ha088;
    SB_DFF Rx_Recv_Byte_i0 (.Q(rx_buf_byte[0]), .C(SLM_CLK_c), .D(n5636));   // src/spi.v(76[8] 221[4])
    SB_DFFESS multi_byte_counter_i7 (.Q(multi_byte_counter[7]), .C(SLM_CLK_c), 
            .E(n5157), .D(n315[7]), .S(n5428));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_1276_i15_3_lut (.I0(tx_addr_byte[6]), .I1(tx_shift_reg[13]), 
            .I2(n2555), .I3(GND_net), .O(n2556[14]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1276_i14_3_lut (.I0(tx_addr_byte[5]), .I1(tx_shift_reg[12]), 
            .I2(n2555), .I3(GND_net), .O(n2556[13]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1276_i13_3_lut (.I0(tx_addr_byte[4]), .I1(tx_shift_reg[11]), 
            .I2(n2555), .I3(GND_net), .O(n2556[12]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1276_i12_3_lut (.I0(tx_addr_byte[3]), .I1(tx_shift_reg[10]), 
            .I2(n2555), .I3(GND_net), .O(n2556[11]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1276_i11_3_lut (.I0(tx_addr_byte[2]), .I1(tx_shift_reg[9]), 
            .I2(n2555), .I3(GND_net), .O(n2556[10]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1276_i10_3_lut (.I0(tx_addr_byte[1]), .I1(tx_shift_reg[8]), 
            .I2(n2555), .I3(GND_net), .O(n2556[9]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1276_i9_3_lut (.I0(tx_addr_byte[0]), .I1(tx_shift_reg[7]), 
            .I2(n2555), .I3(GND_net), .O(n2556[8]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1276_i8_3_lut (.I0(\tx_data_byte[7] ), .I1(tx_shift_reg[6]), 
            .I2(n2555), .I3(GND_net), .O(n2556[7]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1276_i7_3_lut (.I0(\tx_data_byte[6] ), .I1(tx_shift_reg[5]), 
            .I2(n2555), .I3(GND_net), .O(n2556[6]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1276_i6_3_lut (.I0(\tx_data_byte[5] ), .I1(tx_shift_reg[4]), 
            .I2(n2555), .I3(GND_net), .O(n2556[5]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1276_i5_3_lut (.I0(\tx_data_byte[4] ), .I1(tx_shift_reg[3]), 
            .I2(n2555), .I3(GND_net), .O(n2556[4]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1276_i4_3_lut (.I0(\tx_data_byte[3] ), .I1(tx_shift_reg[2]), 
            .I2(n2555), .I3(GND_net), .O(n2556[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1276_i3_3_lut (.I0(\tx_data_byte[2] ), .I1(tx_shift_reg[1]), 
            .I2(n2555), .I3(GND_net), .O(n2556[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_373_Mux_1_i7_4_lut_4_lut (.I0(state[0]), .I1(state[2]), 
            .I2(CS_N_1193), .I3(state[1]), .O(n7));   // src/spi.v(88[9] 219[16])
    defparam mux_373_Mux_1_i7_4_lut_4_lut.LUT_INIT = 16'h20dd;
    SB_LUT4 i13894_4_lut (.I0(n12), .I1(state[1]), .I2(state[0]), .I3(state[2]), 
            .O(n15951));   // src/spi.v(88[9] 219[16])
    defparam i13894_4_lut.LUT_INIT = 16'hc08c;
    SB_LUT4 i1_4_lut_adj_82 (.I0(counter[4]), .I1(n15951), .I2(n15952), 
            .I3(state[3]), .O(n1116[0]));   // src/spi.v(88[9] 219[16])
    defparam i1_4_lut_adj_82.LUT_INIT = 16'ha088;
    SB_LUT4 mux_1276_i2_3_lut (.I0(\tx_data_byte[1] ), .I1(\tx_shift_reg[0] ), 
            .I2(n2555), .I3(GND_net), .O(n2556[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_1276_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n24_adj_1371));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i13861_2_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n15969));   // src/spi.v(88[9] 219[16])
    defparam i13861_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i12556_3_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(spi_start_transfer_r), 
            .I3(state[1]), .O(n14678));
    defparam i12556_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i43_4_lut_4_lut (.I0(state[0]), .I1(state[3]), .I2(state[2]), 
            .I3(state[1]), .O(n21));
    defparam i43_4_lut_4_lut.LUT_INIT = 16'hab44;
    SB_LUT4 mux_373_Mux_2_i15_4_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[2]), .I3(state[3]), .O(n1116[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_373_Mux_2_i15_4_lut_4_lut.LUT_INIT = 16'h0420;
    SB_LUT4 mux_56_Mux_1_i15_3_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[3]), .I3(n7_adj_1372), .O(state_3__N_1123[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i15_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i1_2_lut_4_lut (.I0(counter[0]), .I1(counter[3]), .I2(counter[1]), 
            .I3(counter[2]), .O(n12));   // src/spi.v(88[9] 219[16])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_83 (.I0(counter[2]), .I1(counter[1]), .I2(counter[0]), 
            .I3(counter[3]), .O(n35));
    defparam i1_2_lut_4_lut_adj_83.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_84 (.I0(CS_N_1193), .I1(n21), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i1_2_lut_adj_84.LUT_INIT = 16'h4444;
    SB_LUT4 i14003_4_lut (.I0(n22), .I1(n14678), .I2(n24_adj_1371), .I3(state[3]), 
            .O(n19));
    defparam i14003_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 mux_56_Mux_3_i15_4_lut (.I0(n15969), .I1(state[1]), .I2(state[3]), 
            .I3(n2634[6]), .O(state_3__N_1123[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_3_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i1_2_lut_adj_85 (.I0(n5189), .I1(n14525), .I2(GND_net), .I3(GND_net), 
            .O(n14526));
    defparam i1_2_lut_adj_85.LUT_INIT = 16'h8888;
    SB_LUT4 mux_56_Mux_2_i3_3_lut (.I0(multi_byte_spi_trans_flag_r), .I1(state[0]), 
            .I2(state[1]), .I3(GND_net), .O(n3_adj_1373));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i3_3_lut.LUT_INIT = 16'hc2c2;
    SB_LUT4 mux_56_Mux_2_i15_4_lut (.I0(n3_adj_1373), .I1(state[2]), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_1123[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 i1_4_lut_adj_86 (.I0(n5038), .I1(n5381), .I2(CS_N_1193), .I3(state[1]), 
            .O(n14525));
    defparam i1_4_lut_adj_86.LUT_INIT = 16'ha8aa;
    SB_LUT4 i1_3_lut_adj_87 (.I0(state[3]), .I1(n14525), .I2(n24_adj_1371), 
            .I3(GND_net), .O(n14527));
    defparam i1_3_lut_adj_87.LUT_INIT = 16'h4c4c;
    SB_LUT4 mux_56_Mux_1_i7_4_lut (.I0(n3), .I1(n10087), .I2(state[2]), 
            .I3(state[1]), .O(n7_adj_1372));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i7_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_3_lut_4_lut (.I0(n2634[6]), .I1(state[0]), .I2(state[2]), 
            .I3(state[1]), .O(n4922));   // src/spi.v(88[9] 219[16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i14020_3_lut_4_lut (.I0(state[2]), .I1(state[0]), .I2(n16), 
            .I3(n24), .O(n4999));   // src/spi.v(88[9] 219[16])
    defparam i14020_3_lut_4_lut.LUT_INIT = 16'h000d;
    SB_LUT4 i1_4_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(state[1]), 
            .I3(state[3]), .O(n4));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h01b0;
    SB_LUT4 i3161_4_lut_4_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(state[3]), .O(n4657));   // src/spi.v(88[9] 219[16])
    defparam i3161_4_lut_4_lut_4_lut.LUT_INIT = 16'hfe75;
    SB_LUT4 i13889_2_lut_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(n12), .O(n15952));   // src/spi.v(88[9] 219[16])
    defparam i13889_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i2600_4_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(state[1]), 
            .I3(state[3]), .O(n4086));   // src/spi.v(88[9] 219[16])
    defparam i2600_4_lut_4_lut.LUT_INIT = 16'hfdfb;
    SB_LUT4 i8600_2_lut (.I0(CS_N_1193), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n10087));
    defparam i8600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13919_3_lut (.I0(n2634[6]), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n15962));   // src/spi.v(88[9] 219[16])
    defparam i13919_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 mux_373_Mux_1_i15_4_lut (.I0(n7), .I1(n15962), .I2(state[3]), 
            .I3(state[2]), .O(n1116[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_373_Mux_1_i15_4_lut.LUT_INIT = 16'hfaca;
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=20) 
//

module \uart_rx(CLKS_PER_BIT=20)  (n14672, SLM_CLK_c, n14688, r_Rx_Data, 
            DEBUG_2_c_c, n4935, GND_net, n4, n4_adj_1, \r_Bit_Index[0] , 
            n4942, n4938, n4_adj_2, n6981, pc_data_rx, VCC_net, 
            debug_led3, n6977, n5624, n5620, n5613, n5612, n5611, 
            n5609, n5608) /* synthesis syn_module_defined=1 */ ;
    output n14672;
    input SLM_CLK_c;
    output n14688;
    output r_Rx_Data;
    input DEBUG_2_c_c;
    output n4935;
    input GND_net;
    output n4;
    output n4_adj_1;
    output \r_Bit_Index[0] ;
    output n4942;
    output n4938;
    output n4_adj_2;
    input n6981;
    output [7:0]pc_data_rx;
    input VCC_net;
    output debug_led3;
    input n6977;
    input n5624;
    input n5620;
    input n5613;
    input n5612;
    input n5611;
    input n5609;
    input n5608;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [2:0]n340;
    wire [2:0]r_Bit_Index;   // src/uart_rx.v(33[17:28])
    wire [9:0]n45;
    
    wire n5058;
    wire [9:0]r_Clock_Count;   // src/uart_rx.v(32[17:30])
    
    wire n5440, n3;
    wire [2:0]r_SM_Main;   // src/uart_rx.v(36[17:26])
    
    wire r_Rx_Data_R;
    wire [2:0]r_SM_Main_2__N_950;
    
    wire n14523, n4_c, n10099, n4848, n14032, n5011, n13743, n13742, 
        n13741, n13740, n13739, n13738, n13737, n13736, n13735, 
        n10031, n10081;
    wire [2:0]r_SM_Main_2__N_956;
    
    wire n1, n4846, n8, n14694, n6, n6_adj_1365, n4_adj_1366;
    
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(SLM_CLK_c), .E(n14672), 
            .D(n340[2]), .R(n14688));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1472__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n5058), .D(n45[3]), .R(n5440));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(SLM_CLK_c), .E(n14672), 
            .D(n340[1]), .R(n14688));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1472__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n5058), .D(n45[2]), .R(n5440));   // src/uart_rx.v(120[34:51])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n3), .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(SLM_CLK_c), .D(r_Rx_Data_R));   // src/uart_rx.v(41[10] 45[8])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(r_SM_Main_2__N_950[2]), 
            .R(n14523));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1472__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n5058), .D(n45[1]), .R(n5440));   // src/uart_rx.v(120[34:51])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(SLM_CLK_c), .D(DEBUG_2_c_c));   // src/uart_rx.v(41[10] 45[8])
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_950[2]), 
            .I2(r_SM_Main[1]), .I3(n4_c), .O(n10099));   // src/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h707a;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[2]), .I1(n4848), .I2(r_Bit_Index[1]), 
            .I3(GND_net), .O(n4935));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 equal_144_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // src/uart_rx.v(97[17:39])
    defparam equal_144_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_147_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // src/uart_rx.v(97[17:39])
    defparam equal_147_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut (.I0(n4848), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n4942));   // src/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main_2__N_950[2]), .O(n4848));   // src/uart_rx.v(52[7] 143[14])
    defparam i2_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_adj_71 (.I0(\r_Bit_Index[0] ), .I1(n4848), .I2(GND_net), 
            .I3(GND_net), .O(n4938));   // src/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_71.LUT_INIT = 16'heeee;
    SB_LUT4 equal_149_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // src/uart_rx.v(97[17:39])
    defparam equal_149_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFF r_Rx_Byte_i0 (.Q(pc_data_rx[0]), .C(SLM_CLK_c), .D(n6981));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Rx_DV_52 (.Q(debug_led3), .C(SLM_CLK_c), .E(VCC_net), .D(n14032));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n6977));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_950[2]), 
            .I3(r_SM_Main[0]), .O(n5011));   // src/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n5011), 
            .I3(debug_led3), .O(n14032));   // src/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i14006_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n14523));   // src/uart_rx.v(52[7] 143[14])
    defparam i14006_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFFESR r_Clock_Count_1472__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n5058), .D(n45[0]), .R(n5440));   // src/uart_rx.v(120[34:51])
    SB_LUT4 r_Clock_Count_1472_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n13743), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1472_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1472_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n13742), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1472_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1472_add_4_10 (.CI(n13742), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n13743));
    SB_LUT4 r_Clock_Count_1472_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n13741), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1472_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1472_add_4_9 (.CI(n13741), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n13742));
    SB_LUT4 r_Clock_Count_1472_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n13740), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1472_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1472_add_4_8 (.CI(n13740), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n13741));
    SB_LUT4 r_Clock_Count_1472_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n13739), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1472_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1472_add_4_7 (.CI(n13739), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n13740));
    SB_LUT4 r_Clock_Count_1472_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n13738), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1472_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1472_add_4_6 (.CI(n13738), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n13739));
    SB_LUT4 r_Clock_Count_1472_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n13737), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1472_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1472_add_4_5 (.CI(n13737), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n13738));
    SB_LUT4 r_Clock_Count_1472_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n13736), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1472_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1472_add_4_4 (.CI(n13736), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n13737));
    SB_LUT4 r_Clock_Count_1472_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n13735), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1472_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1472_add_4_3 (.CI(n13735), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n13736));
    SB_LUT4 r_Clock_Count_1472_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1472_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1472_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n13735));
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n10099), 
            .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1472__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n5058), .D(n45[9]), .R(n5440));   // src/uart_rx.v(120[34:51])
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n10031));   // src/uart_rx.v(102[36:51])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1643_2_lut_3_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n340[2]));   // src/uart_rx.v(102[36:51])
    defparam i1643_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n10031), .I1(r_SM_Main_2__N_950[2]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n10081));   // src/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_956[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // src/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n10081), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // src/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFESR r_Clock_Count_1472__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n5058), .D(n45[8]), .R(n5440));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1472__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n5058), .D(n45[7]), .R(n5440));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1472__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n5058), .D(n45[6]), .R(n5440));   // src/uart_rx.v(120[34:51])
    SB_LUT4 i1636_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n340[1]));   // src/uart_rx.v(102[36:51])
    defparam i1636_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Byte_i1 (.Q(pc_data_rx[1]), .C(SLM_CLK_c), .D(n5624));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(pc_data_rx[2]), .C(SLM_CLK_c), .D(n5620));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(pc_data_rx[3]), .C(SLM_CLK_c), .D(n5613));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(pc_data_rx[4]), .C(SLM_CLK_c), .D(n5612));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(pc_data_rx[5]), .C(SLM_CLK_c), .D(n5611));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1472__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n5058), .D(n45[5]), .R(n5440));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1472__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n5058), .D(n45[4]), .R(n5440));   // src/uart_rx.v(120[34:51])
    SB_DFF r_Rx_Byte_i6 (.Q(pc_data_rx[6]), .C(SLM_CLK_c), .D(n5609));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(pc_data_rx[7]), .C(SLM_CLK_c), .D(n5608));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[4]), .I2(r_Clock_Count[3]), 
            .I3(n4846), .O(n8));   // src/uart_rx.v(68[17:52])
    defparam i3_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i4_3_lut (.I0(r_Clock_Count[1]), .I1(n8), .I2(r_Clock_Count[2]), 
            .I3(GND_net), .O(r_SM_Main_2__N_956[0]));   // src/uart_rx.v(68[17:52])
    defparam i4_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_72 (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_956[0]), 
            .I2(GND_net), .I3(GND_net), .O(n4_c));
    defparam i1_2_lut_adj_72.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n14694), .I2(r_SM_Main_2__N_950[2]), 
            .I3(r_SM_Main[1]), .O(n5440));
    defparam i1_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i2_2_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_956[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13992_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6), 
            .I3(r_SM_Main[0]), .O(n5058));   // src/uart_rx.v(52[7] 143[14])
    defparam i13992_4_lut.LUT_INIT = 16'h4555;
    SB_LUT4 i1_2_lut_adj_73 (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[9]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_1365));   // src/uart_rx.v(68[17:52])
    defparam i1_2_lut_adj_73.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[5]), 
            .I3(n6_adj_1365), .O(n4846));   // src/uart_rx.v(68[17:52])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n4_adj_1366));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i8591_4_lut (.I0(r_Clock_Count[3]), .I1(n4846), .I2(r_Clock_Count[4]), 
            .I3(n4_adj_1366), .O(r_SM_Main_2__N_950[2]));
    defparam i8591_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i12572_2_lut_3_lut (.I0(r_SM_Main[0]), .I1(r_Rx_Data), .I2(r_SM_Main_2__N_956[0]), 
            .I3(GND_net), .O(n14694));
    defparam i12572_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i14012_3_lut (.I0(n14672), .I1(n10031), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n14688));
    defparam i14012_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i14034_4_lut (.I0(r_SM_Main_2__N_950[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n14672));
    defparam i14034_4_lut.LUT_INIT = 16'h0023;
    
endmodule
//
// Verilog Description of module \uart_tx(CLKS_PER_BIT=20) 
//

module \uart_tx(CLKS_PER_BIT=20)  (n14684, SLM_CLK_c, n14690, DEBUG_1_c, 
            r_SM_Main, \r_SM_Main_2__N_1026[1] , \r_SM_Main_2__N_1029[0] , 
            n14508, \r_Bit_Index[0] , r_Tx_Data, GND_net, n18034, 
            n6999, n6998, n6997, n6996, n6995, n6994, n6993, n6974, 
            VCC_net, n4435, n5629, n5628, tx_uart_active_flag) /* synthesis syn_module_defined=1 */ ;
    output n14684;
    input SLM_CLK_c;
    output n14690;
    output DEBUG_1_c;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_1026[1] ;
    input \r_SM_Main_2__N_1029[0] ;
    output n14508;
    output \r_Bit_Index[0] ;
    output [7:0]r_Tx_Data;
    input GND_net;
    input n18034;
    input n6999;
    input n6998;
    input n6997;
    input n6996;
    input n6995;
    input n6994;
    input n6993;
    input n6974;
    input VCC_net;
    output n4435;
    input n5629;
    input n5628;
    output tx_uart_active_flag;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [2:0]n312;
    wire [2:0]r_Bit_Index;   // src/uart_tx.v(33[16:27])
    
    wire n3, n1, n3775, n17043, n17046, n5442;
    wire [9:0]n45;
    wire [9:0]r_Clock_Count;   // src/uart_tx.v(32[16:29])
    
    wire n13750, n10035, n13751, n13749, n13748, n13747, n13746, 
        n13745, n13744, n3_adj_1361, n4, n8, n7, n3774, n17136, 
        o_Tx_Serial_N_1058, n13752, n17133;
    
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(SLM_CLK_c), .E(n14684), 
            .D(n312[1]), .R(n14690));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFE o_Tx_Serial_44 (.Q(DEBUG_1_c), .C(SLM_CLK_c), .E(n1), .D(n3));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n3775), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i13938_4_lut_4_lut (.I0(\r_SM_Main_2__N_1026[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_1029[0] ), .O(n14508));
    defparam i13938_4_lut_4_lut.LUT_INIT = 16'h8380;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_14842 (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n17043));
    defparam r_Bit_Index_0__bdd_4_lut_14842.LUT_INIT = 16'he4aa;
    SB_LUT4 n17043_bdd_4_lut (.I0(n17043), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n17046));
    defparam n17043_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13986_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_1026[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n5442));
    defparam i13986_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 r_Clock_Count_1474_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n13750), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1474_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(n18034));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(SLM_CLK_c), .D(n6999));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(SLM_CLK_c), .D(n6998));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(SLM_CLK_c), .D(n6997));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(SLM_CLK_c), .D(n6996));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(SLM_CLK_c), .D(n6995));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(SLM_CLK_c), .D(n6994));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(SLM_CLK_c), .D(n6993));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n6974));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i1665_2_lut_3_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n312[2]));   // src/uart_tx.v(96[36:51])
    defparam i1665_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n10035));   // src/uart_tx.v(96[36:51])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFFESR r_Clock_Count_1474__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[0]), .R(n5442));   // src/uart_tx.v(116[34:51])
    SB_CARRY r_Clock_Count_1474_add_4_9 (.CI(n13750), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n13751));
    SB_LUT4 r_Clock_Count_1474_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n13749), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1474_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1474_add_4_8 (.CI(n13749), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n13750));
    SB_LUT4 r_Clock_Count_1474_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n13748), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1474_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1474_add_4_7 (.CI(n13748), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n13749));
    SB_LUT4 r_Clock_Count_1474_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n13747), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1474_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1474_add_4_6 (.CI(n13747), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n13748));
    SB_LUT4 r_Clock_Count_1474_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n13746), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1474_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1474_add_4_5 (.CI(n13746), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n13747));
    SB_LUT4 r_Clock_Count_1474_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n13745), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1474_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1474_add_4_4 (.CI(n13745), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n13746));
    SB_LUT4 r_Clock_Count_1474_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n13744), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1474_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1474_add_4_3 (.CI(n13744), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n13745));
    SB_LUT4 r_Clock_Count_1474_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1474_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Clock_Count_1474__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[9]), .R(n5442));   // src/uart_tx.v(116[34:51])
    SB_CARRY r_Clock_Count_1474_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n13744));
    SB_DFFESR r_Clock_Count_1474__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[8]), .R(n5442));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1474__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[7]), .R(n5442));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1474__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[6]), .R(n5442));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1474__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[5]), .R(n5442));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1474__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[4]), .R(n5442));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1474__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[3]), .R(n5442));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1474__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[2]), .R(n5442));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1474__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[1]), .R(n5442));   // src/uart_tx.v(116[34:51])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_1029[0] ), .O(n4435));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i13964_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_1026[1] ), .O(n14684));
    defparam i13964_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n3_adj_1361), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n4));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[9]), .I2(GND_net), 
            .I3(GND_net), .O(n8));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[4]), 
            .I3(n4), .O(n7));
    defparam i1_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i5_4_lut (.I0(r_Clock_Count[5]), .I1(n7), .I2(r_Clock_Count[8]), 
            .I3(n8), .O(\r_SM_Main_2__N_1026[1] ));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2289_4_lut (.I0(\r_SM_Main_2__N_1029[0] ), .I1(n10035), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_1026[1] ), .O(n3774));   // src/uart_tx.v(41[7] 140[14])
    defparam i2289_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i2290_3_lut (.I0(n3774), .I1(\r_SM_Main_2__N_1026[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n3775));   // src/uart_tx.v(41[7] 140[14])
    defparam i2290_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9052256_i1_3_lut (.I0(n17136), .I1(n17046), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_1058));
    defparam i9052256_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_55_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_1058), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // src/uart_tx.v(41[7] 140[14])
    defparam r_SM_Main_2__I_0_55_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i2849_2_lut_3_lut (.I0(\r_SM_Main_2__N_1026[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_1361));
    defparam i2849_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(SLM_CLK_c), .D(n5629));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Active_46 (.Q(tx_uart_active_flag), .C(SLM_CLK_c), .D(n5628));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(SLM_CLK_c), .E(n14684), 
            .D(n312[2]), .R(n14690));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 r_Clock_Count_1474_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n13752), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1474_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1474_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n13751), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1474_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1474_add_4_10 (.CI(n13751), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n13752));
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n17133));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n17133_bdd_4_lut (.I0(n17133), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n17136));
    defparam n17133_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14015_3_lut (.I0(n14684), .I1(n10035), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n14690));
    defparam i14015_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1658_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n312[1]));   // src/uart_tx.v(96[36:51])
    defparam i1658_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module usb3_if
//

module usb3_if (FIFO_CLK_c, reset_per_frame, SLM_CLK_c, dc32_fifo_empty, 
            VCC_net, FT_RD_c, dc32_fifo_data_in, DEBUG_5_c, buffer_switch_done, 
            buffer_switch_done_latched, FT_OE_N_496, GND_net, FIFO_D0_c_31, 
            FIFO_D1_c_30, FIFO_D2_c_29, DEBUG_9_c_c, FIFO_D3_c_28, FIFO_D4_c_27, 
            FIFO_D5_c_26, FIFO_D6_c_25, FIFO_D7_c_24, FIFO_D8_c_23, 
            FIFO_D9_c_22, FIFO_D10_c_21, FIFO_D31_c_0, FIFO_D11_c_20, 
            FIFO_D12_c_19, FIFO_D13_c_18, FIFO_D14_c_17, FIFO_D15_c_16, 
            FIFO_D16_c_15, FIFO_D17_c_14, FIFO_D18_c_13, FIFO_D19_c_12, 
            FIFO_D20_c_11, FIFO_D21_c_10, FIFO_D22_c_9, FT_OE_c, FIFO_D23_c_8, 
            FIFO_D24_c_7, FIFO_D25_c_6, FIFO_D26_c_5, FIFO_D27_c_4, 
            n12, FIFO_D28_c_3, n14706, n13865, rd_fifo_en_w, empty_nxt_c_N_636, 
            dc32_fifo_almost_full, FIFO_D29_c_2, dc32_fifo_full, wr_fifo_en_w, 
            FIFO_D30_c_1) /* synthesis syn_module_defined=1 */ ;
    input FIFO_CLK_c;
    input reset_per_frame;
    input SLM_CLK_c;
    input dc32_fifo_empty;
    input VCC_net;
    output FT_RD_c;
    output [31:0]dc32_fifo_data_in;
    output DEBUG_5_c;
    input buffer_switch_done;
    output buffer_switch_done_latched;
    output FT_OE_N_496;
    input GND_net;
    input FIFO_D0_c_31;
    input FIFO_D1_c_30;
    input FIFO_D2_c_29;
    input DEBUG_9_c_c;
    input FIFO_D3_c_28;
    input FIFO_D4_c_27;
    input FIFO_D5_c_26;
    input FIFO_D6_c_25;
    input FIFO_D7_c_24;
    input FIFO_D8_c_23;
    input FIFO_D9_c_22;
    input FIFO_D10_c_21;
    input FIFO_D31_c_0;
    input FIFO_D11_c_20;
    input FIFO_D12_c_19;
    input FIFO_D13_c_18;
    input FIFO_D14_c_17;
    input FIFO_D15_c_16;
    input FIFO_D16_c_15;
    input FIFO_D17_c_14;
    input FIFO_D18_c_13;
    input FIFO_D19_c_12;
    input FIFO_D20_c_11;
    input FIFO_D21_c_10;
    input FIFO_D22_c_9;
    output FT_OE_c;
    input FIFO_D23_c_8;
    input FIFO_D24_c_7;
    input FIFO_D25_c_6;
    input FIFO_D26_c_5;
    input FIFO_D27_c_4;
    input n12;
    input FIFO_D28_c_3;
    input n14706;
    input n13865;
    input rd_fifo_en_w;
    output empty_nxt_c_N_636;
    input dc32_fifo_almost_full;
    input FIFO_D29_c_2;
    input dc32_fifo_full;
    output wr_fifo_en_w;
    input FIFO_D30_c_1;
    
    wire FIFO_CLK_c /* synthesis SET_AS_NETWORK=FIFO_CLK_c, is_clock=1 */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n14517, n4990;
    wire [4:0]state_timeout_counter;   // src/usb3_if.v(64[11:32])
    
    wire reset_per_frame_latched, dc32_fifo_empty_latched, FT_RD_N_501;
    wire [31:0]dc32_fifo_data_in_latched;   // src/usb3_if.v(66[12:37])
    
    wire write_to_dc32_fifo_latched;
    wire [5:0]n29;
    
    wire n8362;
    wire [5:0]num_words_curr_line;   // src/usb3_if.v(60[11:30])
    
    wire n8360;
    wire [15:0]n650;
    
    wire n1236, n4393, n10, n3525;
    wire [10:0]num_lines_clocked_out_10__N_441;
    
    wire n5098;
    wire [10:0]num_lines_clocked_out;   // src/usb3_if.v(63[12:33])
    
    wire n5217, n5432, write_to_dc32_fifo_latched_N_503, n15981, n609, 
        FT_OE_N_495, FT_OE_N_490, n7039, n15965, n14577, n13888, 
        FT_OE_N_491, n9, n32_adj_1353, n13790, n13712, n13789, n13788, 
        n13787, n13786;
    wire [4:0]n2034;
    
    wire n10053, n13711, n13710, n13709, n13708, n13707, n13706, 
        n13705, n15955, n1, n13704, n703, n859, n18, n16, n20, 
        n8464, n4, n14479, n696, n3510, n3506, n706, n709, n13703, 
        n6, n2118, n15945, n13825, n16_adj_1354, n8, n7, n15, 
        n4923, n894, n9698, n688, n7_adj_1355, n6_adj_1356, n2, 
        n8_adj_1357, n7_adj_1358, n8_adj_1359, n62;
    wire [4:0]n2024;
    
    wire n4578, n18_adj_1360, n614, n15944, n2122, n2120, n16067;
    
    SB_DFFE state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(FIFO_CLK_c), 
            .E(n4990), .D(n14517));   // src/usb3_if.v(86[8] 201[4])
    SB_DFF reset_per_frame_latched_111 (.Q(reset_per_frame_latched), .C(SLM_CLK_c), 
           .D(reset_per_frame));   // src/usb3_if.v(70[8] 83[4])
    SB_DFF dc32_fifo_empty_latched_112 (.Q(dc32_fifo_empty_latched), .C(SLM_CLK_c), 
           .D(dc32_fifo_empty));   // src/usb3_if.v(70[8] 83[4])
    SB_DFFESS FT_RD_114 (.Q(FT_RD_c), .C(FIFO_CLK_c), .E(VCC_net), .D(FT_RD_N_501), 
            .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFN dc32_fifo_data_in_i0 (.Q(dc32_fifo_data_in[0]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[0]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN write_to_dc32_fifo_122 (.Q(DEBUG_5_c), .C(FIFO_CLK_c), .D(write_to_dc32_fifo_latched));   // src/usb3_if.v(204[8] 207[4])
    SB_DFF buffer_switch_done_latched_110 (.Q(buffer_switch_done_latched), 
           .C(SLM_CLK_c), .D(buffer_switch_done));   // src/usb3_if.v(70[8] 83[4])
    SB_DFFESS num_words_curr_line_1470__i5 (.Q(num_words_curr_line[5]), .C(FIFO_CLK_c), 
            .E(n8362), .D(n29[5]), .S(n8360));   // src/usb3_if.v(148[44:69])
    SB_DFFESR num_words_curr_line_1470__i4 (.Q(num_words_curr_line[4]), .C(FIFO_CLK_c), 
            .E(n8362), .D(n29[4]), .R(n8360));   // src/usb3_if.v(148[44:69])
    SB_DFFESS num_words_curr_line_1470__i3 (.Q(num_words_curr_line[3]), .C(FIFO_CLK_c), 
            .E(n8362), .D(n29[3]), .S(n8360));   // src/usb3_if.v(148[44:69])
    SB_LUT4 i2_3_lut_4_lut (.I0(dc32_fifo_empty), .I1(n650[2]), .I2(FT_OE_N_496), 
            .I3(n1236), .O(n4393));   // src/usb3_if.v(97[9] 199[16])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_3_lut (.I0(dc32_fifo_empty), .I1(n650[2]), .I2(state_timeout_counter[0]), 
            .I3(GND_net), .O(n10));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFFSS state_FSM_i1 (.Q(n650[0]), .C(FIFO_CLK_c), .D(n3525), .S(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFESR num_words_curr_line_1470__i2 (.Q(num_words_curr_line[2]), .C(FIFO_CLK_c), 
            .E(n8362), .D(n29[2]), .R(n8360));   // src/usb3_if.v(148[44:69])
    SB_DFFESS num_lines_clocked_out_i10 (.Q(num_lines_clocked_out[10]), .C(FIFO_CLK_c), 
            .E(n5098), .D(num_lines_clocked_out_10__N_441[10]), .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_words_curr_line_1470__i1 (.Q(num_words_curr_line[1]), .C(FIFO_CLK_c), 
            .E(n8362), .D(n29[1]), .R(n8360));   // src/usb3_if.v(148[44:69])
    SB_DFFESR dc32_fifo_data_in_latched__i31 (.Q(dc32_fifo_data_in_latched[31]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D0_c_31), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i30 (.Q(dc32_fifo_data_in_latched[30]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D1_c_30), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i9 (.Q(num_lines_clocked_out[9]), .C(FIFO_CLK_c), 
            .E(n5098), .D(num_lines_clocked_out_10__N_441[9]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESS num_lines_clocked_out_i8 (.Q(num_lines_clocked_out[8]), .C(FIFO_CLK_c), 
            .E(n5098), .D(num_lines_clocked_out_10__N_441[8]), .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i7 (.Q(num_lines_clocked_out[7]), .C(FIFO_CLK_c), 
            .E(n5098), .D(num_lines_clocked_out_10__N_441[7]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i6 (.Q(num_lines_clocked_out[6]), .C(FIFO_CLK_c), 
            .E(n5098), .D(num_lines_clocked_out_10__N_441[6]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i5 (.Q(num_lines_clocked_out[5]), .C(FIFO_CLK_c), 
            .E(n5098), .D(num_lines_clocked_out_10__N_441[5]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i4 (.Q(num_lines_clocked_out[4]), .C(FIFO_CLK_c), 
            .E(n5098), .D(num_lines_clocked_out_10__N_441[4]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i3 (.Q(num_lines_clocked_out[3]), .C(FIFO_CLK_c), 
            .E(n5098), .D(num_lines_clocked_out_10__N_441[3]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i2 (.Q(num_lines_clocked_out[2]), .C(FIFO_CLK_c), 
            .E(n5098), .D(num_lines_clocked_out_10__N_441[2]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i1 (.Q(num_lines_clocked_out[1]), .C(FIFO_CLK_c), 
            .E(n5098), .D(num_lines_clocked_out_10__N_441[1]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFSR write_to_dc32_fifo_latched_116 (.Q(write_to_dc32_fifo_latched), 
            .C(FIFO_CLK_c), .D(write_to_dc32_fifo_latched_N_503), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i1_4_lut (.I0(n15981), .I1(n609), .I2(FT_OE_N_495), .I3(n650[2]), 
            .O(FT_OE_N_490));
    defparam i1_4_lut.LUT_INIT = 16'hcfaa;
    SB_DFF state_FSM_i5 (.Q(n650[4]), .C(FIFO_CLK_c), .D(n7039));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFESR dc32_fifo_data_in_latched__i29 (.Q(dc32_fifo_data_in_latched[29]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D2_c_29), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i1_4_lut_4_lut (.I0(n650[5]), .I1(FT_OE_N_496), .I2(DEBUG_9_c_c), 
            .I3(n15965), .O(FT_RD_N_501));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hf7a2;
    SB_DFFESR num_words_curr_line_1470__i0 (.Q(num_words_curr_line[0]), .C(FIFO_CLK_c), 
            .E(n8362), .D(n29[0]), .R(n8360));   // src/usb3_if.v(148[44:69])
    SB_LUT4 i2_3_lut_4_lut_adj_36 (.I0(n650[5]), .I1(FT_OE_N_496), .I2(n14577), 
            .I3(n650[2]), .O(n13888));   // src/usb3_if.v(97[9] 199[16])
    defparam i2_3_lut_4_lut_adj_36.LUT_INIT = 16'hf222;
    SB_LUT4 i1_3_lut_4_lut (.I0(n650[5]), .I1(FT_OE_N_491), .I2(n9), .I3(reset_per_frame_latched), 
            .O(n8362));   // src/usb3_if.v(96[10] 200[8])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hff70;
    SB_LUT4 i13930_3_lut_4_lut (.I0(n650[5]), .I1(FT_OE_N_491), .I2(n650[0]), 
            .I3(n32_adj_1353), .O(n15981));   // src/usb3_if.v(96[10] 200[8])
    defparam i13930_3_lut_4_lut.LUT_INIT = 16'hfff8;
    SB_DFFESR dc32_fifo_data_in_latched__i28 (.Q(dc32_fifo_data_in_latched[28]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D3_c_28), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i27 (.Q(dc32_fifo_data_in_latched[27]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D4_c_27), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i26 (.Q(dc32_fifo_data_in_latched[26]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D5_c_26), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i25 (.Q(dc32_fifo_data_in_latched[25]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D6_c_25), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i24 (.Q(dc32_fifo_data_in_latched[24]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D7_c_24), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i23 (.Q(dc32_fifo_data_in_latched[23]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D8_c_23), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i22 (.Q(dc32_fifo_data_in_latched[22]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D9_c_22), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i21 (.Q(dc32_fifo_data_in_latched[21]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D10_c_21), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i0 (.Q(dc32_fifo_data_in_latched[0]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D31_c_0), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i20 (.Q(dc32_fifo_data_in_latched[20]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D11_c_20), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i19 (.Q(dc32_fifo_data_in_latched[19]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D12_c_19), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR num_lines_clocked_out_i0 (.Q(num_lines_clocked_out[0]), .C(FIFO_CLK_c), 
            .E(n5098), .D(num_lines_clocked_out_10__N_441[0]), .R(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 num_words_curr_line_1470_add_4_7_lut (.I0(GND_net), .I1(VCC_net), 
            .I2(num_words_curr_line[5]), .I3(n13790), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam num_words_curr_line_1470_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_116_add_2_12_lut (.I0(GND_net), .I1(num_lines_clocked_out[10]), 
            .I2(VCC_net), .I3(n13712), .O(num_lines_clocked_out_10__N_441[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 num_words_curr_line_1470_add_4_6_lut (.I0(GND_net), .I1(VCC_net), 
            .I2(num_words_curr_line[4]), .I3(n13789), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam num_words_curr_line_1470_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY num_words_curr_line_1470_add_4_6 (.CI(n13789), .I0(VCC_net), 
            .I1(num_words_curr_line[4]), .CO(n13790));
    SB_LUT4 num_words_curr_line_1470_add_4_5_lut (.I0(GND_net), .I1(VCC_net), 
            .I2(num_words_curr_line[3]), .I3(n13788), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam num_words_curr_line_1470_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY num_words_curr_line_1470_add_4_5 (.CI(n13788), .I0(VCC_net), 
            .I1(num_words_curr_line[3]), .CO(n13789));
    SB_LUT4 num_words_curr_line_1470_add_4_4_lut (.I0(GND_net), .I1(VCC_net), 
            .I2(num_words_curr_line[2]), .I3(n13787), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam num_words_curr_line_1470_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut (.I0(reset_per_frame_latched), .I1(n650[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7039));   // src/usb3_if.v(70[8] 83[4])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY num_words_curr_line_1470_add_4_4 (.CI(n13787), .I0(VCC_net), 
            .I1(num_words_curr_line[2]), .CO(n13788));
    SB_LUT4 num_words_curr_line_1470_add_4_3_lut (.I0(GND_net), .I1(VCC_net), 
            .I2(num_words_curr_line[1]), .I3(n13786), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam num_words_curr_line_1470_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY num_words_curr_line_1470_add_4_3 (.CI(n13786), .I0(VCC_net), 
            .I1(num_words_curr_line[1]), .CO(n13787));
    SB_LUT4 num_words_curr_line_1470_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(num_words_curr_line[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam num_words_curr_line_1470_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFE state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(FIFO_CLK_c), 
            .E(n4990), .D(n2034[4]));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFE state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(FIFO_CLK_c), 
            .E(n4990), .D(n2034[3]));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFE state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(FIFO_CLK_c), 
            .E(n4990), .D(n2034[2]));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFE state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(FIFO_CLK_c), 
            .E(n4990), .D(n10053));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 sub_116_add_2_11_lut (.I0(GND_net), .I1(num_lines_clocked_out[9]), 
            .I2(VCC_net), .I3(n13711), .O(num_lines_clocked_out_10__N_441[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY num_words_curr_line_1470_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(num_words_curr_line[0]), .CO(n13786));
    SB_DFFESR dc32_fifo_data_in_latched__i18 (.Q(dc32_fifo_data_in_latched[18]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D13_c_18), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i17 (.Q(dc32_fifo_data_in_latched[17]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D14_c_17), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_CARRY sub_116_add_2_11 (.CI(n13711), .I0(num_lines_clocked_out[9]), 
            .I1(VCC_net), .CO(n13712));
    SB_LUT4 sub_116_add_2_10_lut (.I0(GND_net), .I1(num_lines_clocked_out[8]), 
            .I2(VCC_net), .I3(n13710), .O(num_lines_clocked_out_10__N_441[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_10 (.CI(n13710), .I0(num_lines_clocked_out[8]), 
            .I1(VCC_net), .CO(n13711));
    SB_LUT4 sub_116_add_2_9_lut (.I0(GND_net), .I1(num_lines_clocked_out[7]), 
            .I2(VCC_net), .I3(n13709), .O(num_lines_clocked_out_10__N_441[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_9 (.CI(n13709), .I0(num_lines_clocked_out[7]), 
            .I1(VCC_net), .CO(n13710));
    SB_LUT4 sub_116_add_2_8_lut (.I0(GND_net), .I1(num_lines_clocked_out[6]), 
            .I2(VCC_net), .I3(n13708), .O(num_lines_clocked_out_10__N_441[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_8 (.CI(n13708), .I0(num_lines_clocked_out[6]), 
            .I1(VCC_net), .CO(n13709));
    SB_LUT4 sub_116_add_2_7_lut (.I0(GND_net), .I1(num_lines_clocked_out[5]), 
            .I2(VCC_net), .I3(n13707), .O(num_lines_clocked_out_10__N_441[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_7 (.CI(n13707), .I0(num_lines_clocked_out[5]), 
            .I1(VCC_net), .CO(n13708));
    SB_LUT4 sub_116_add_2_6_lut (.I0(GND_net), .I1(num_lines_clocked_out[4]), 
            .I2(VCC_net), .I3(n13706), .O(num_lines_clocked_out_10__N_441[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_6 (.CI(n13706), .I0(num_lines_clocked_out[4]), 
            .I1(VCC_net), .CO(n13707));
    SB_LUT4 sub_116_add_2_5_lut (.I0(GND_net), .I1(num_lines_clocked_out[3]), 
            .I2(VCC_net), .I3(n13705), .O(num_lines_clocked_out_10__N_441[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_4_lut (.I0(n15955), .I1(n1), .I2(n650[5]), .I3(n609), 
            .O(write_to_dc32_fifo_latched_N_503));   // src/usb3_if.v(97[9] 199[16])
    defparam i13_4_lut.LUT_INIT = 16'h303a;
    SB_CARRY sub_116_add_2_5 (.CI(n13705), .I0(num_lines_clocked_out[3]), 
            .I1(VCC_net), .CO(n13706));
    SB_DFFN dc32_fifo_data_in_i1 (.Q(dc32_fifo_data_in[1]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[1]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i2 (.Q(dc32_fifo_data_in[2]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[2]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i3 (.Q(dc32_fifo_data_in[3]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[3]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i4 (.Q(dc32_fifo_data_in[4]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[4]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i5 (.Q(dc32_fifo_data_in[5]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[5]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i6 (.Q(dc32_fifo_data_in[6]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[6]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i7 (.Q(dc32_fifo_data_in[7]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[7]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i8 (.Q(dc32_fifo_data_in[8]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[8]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i9 (.Q(dc32_fifo_data_in[9]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[9]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i10 (.Q(dc32_fifo_data_in[10]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[10]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i11 (.Q(dc32_fifo_data_in[11]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[11]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i12 (.Q(dc32_fifo_data_in[12]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[12]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i13 (.Q(dc32_fifo_data_in[13]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[13]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i14 (.Q(dc32_fifo_data_in[14]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[14]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i15 (.Q(dc32_fifo_data_in[15]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[15]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i16 (.Q(dc32_fifo_data_in[16]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[16]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i17 (.Q(dc32_fifo_data_in[17]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[17]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i18 (.Q(dc32_fifo_data_in[18]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[18]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i19 (.Q(dc32_fifo_data_in[19]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[19]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i20 (.Q(dc32_fifo_data_in[20]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[20]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i21 (.Q(dc32_fifo_data_in[21]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[21]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i22 (.Q(dc32_fifo_data_in[22]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[22]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i23 (.Q(dc32_fifo_data_in[23]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[23]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i24 (.Q(dc32_fifo_data_in[24]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[24]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i25 (.Q(dc32_fifo_data_in[25]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[25]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i26 (.Q(dc32_fifo_data_in[26]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[26]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i27 (.Q(dc32_fifo_data_in[27]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[27]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i28 (.Q(dc32_fifo_data_in[28]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[28]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i29 (.Q(dc32_fifo_data_in[29]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[29]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i30 (.Q(dc32_fifo_data_in[30]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[30]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFN dc32_fifo_data_in_i31 (.Q(dc32_fifo_data_in[31]), .C(FIFO_CLK_c), 
            .D(dc32_fifo_data_in_latched[31]));   // src/usb3_if.v(204[8] 207[4])
    SB_DFFESR dc32_fifo_data_in_latched__i16 (.Q(dc32_fifo_data_in_latched[16]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D15_c_16), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i15 (.Q(dc32_fifo_data_in_latched[15]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D16_c_15), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i14 (.Q(dc32_fifo_data_in_latched[14]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D17_c_14), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i13 (.Q(dc32_fifo_data_in_latched[13]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D18_c_13), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i12 (.Q(dc32_fifo_data_in_latched[12]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D19_c_12), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i11 (.Q(dc32_fifo_data_in_latched[11]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D20_c_11), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i10 (.Q(dc32_fifo_data_in_latched[10]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D21_c_10), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i9 (.Q(dc32_fifo_data_in_latched[9]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D22_c_9), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESS FT_OE_113 (.Q(FT_OE_c), .C(FIFO_CLK_c), .E(VCC_net), .D(FT_OE_N_490), 
            .S(reset_per_frame_latched));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i8 (.Q(dc32_fifo_data_in_latched[8]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D23_c_8), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 sub_116_add_2_4_lut (.I0(GND_net), .I1(num_lines_clocked_out[2]), 
            .I2(VCC_net), .I3(n13704), .O(num_lines_clocked_out_10__N_441[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR dc32_fifo_data_in_latched__i7 (.Q(dc32_fifo_data_in_latched[7]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D24_c_7), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i6 (.Q(dc32_fifo_data_in_latched[6]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D25_c_6), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_DFFESR dc32_fifo_data_in_latched__i5 (.Q(dc32_fifo_data_in_latched[5]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D26_c_5), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i1_2_lut_adj_37 (.I0(DEBUG_9_c_c), .I1(FT_OE_N_496), .I2(GND_net), 
            .I3(GND_net), .O(n1));
    defparam i1_2_lut_adj_37.LUT_INIT = 16'h8888;
    SB_LUT4 i2201_4_lut (.I0(n650[2]), .I1(reset_per_frame_latched), .I2(n703), 
            .I3(n859), .O(n5432));   // src/usb3_if.v(86[8] 201[4])
    defparam i2201_4_lut.LUT_INIT = 16'hfcdd;
    SB_DFFESR dc32_fifo_data_in_latched__i4 (.Q(dc32_fifo_data_in_latched[4]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D27_c_4), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i7_4_lut (.I0(num_lines_clocked_out[3]), .I1(num_lines_clocked_out[1]), 
            .I2(num_lines_clocked_out[8]), .I3(num_lines_clocked_out[4]), 
            .O(n18));   // src/usb3_if.v(86[8] 201[4])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(num_lines_clocked_out[6]), .I1(num_lines_clocked_out[7]), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // src/usb3_if.v(86[8] 201[4])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut (.I0(num_lines_clocked_out[5]), .I1(n18), .I2(num_lines_clocked_out[2]), 
            .I3(num_lines_clocked_out[10]), .O(n20));   // src/usb3_if.v(86[8] 201[4])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(num_lines_clocked_out[0]), .I1(n20), .I2(n16), 
            .I3(num_lines_clocked_out[9]), .O(n8464));   // src/usb3_if.v(86[8] 201[4])
    defparam i10_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i2047_3_lut (.I0(n4), .I1(n4393), .I2(n8464), .I3(GND_net), 
            .O(n3525));   // src/usb3_if.v(97[9] 199[16])
    defparam i2047_3_lut.LUT_INIT = 16'haeae;
    SB_DFFSR state_FSM_i2 (.Q(n650[1]), .C(FIFO_CLK_c), .D(n14479), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i3 (.Q(n650[2]), .C(FIFO_CLK_c), .D(n13888), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i4 (.Q(n650[3]), .C(FIFO_CLK_c), .D(n696), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i6 (.Q(n650[5]), .C(FIFO_CLK_c), .D(n3510), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i7 (.Q(n650[6]), .C(FIFO_CLK_c), .D(n3506), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i8 (.Q(n650[7]), .C(FIFO_CLK_c), .D(n706), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_DFFSR state_FSM_i9 (.Q(n650[8]), .C(FIFO_CLK_c), .D(n709), .R(reset_per_frame_latched));   // src/usb3_if.v(97[9] 199[16])
    SB_CARRY sub_116_add_2_4 (.CI(n13704), .I0(num_lines_clocked_out[2]), 
            .I1(VCC_net), .CO(n13705));
    SB_LUT4 sub_116_add_2_3_lut (.I0(GND_net), .I1(num_lines_clocked_out[1]), 
            .I2(VCC_net), .I3(n13703), .O(num_lines_clocked_out_10__N_441[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_3 (.CI(n13703), .I0(num_lines_clocked_out[1]), 
            .I1(VCC_net), .CO(n13704));
    SB_LUT4 sub_116_add_2_2_lut (.I0(GND_net), .I1(num_lines_clocked_out[0]), 
            .I2(n12), .I3(VCC_net), .O(num_lines_clocked_out_10__N_441[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_2 (.CI(VCC_net), .I0(num_lines_clocked_out[0]), 
            .I1(n12), .CO(n13703));
    SB_DFFESR dc32_fifo_data_in_latched__i3 (.Q(dc32_fifo_data_in_latched[3]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D28_c_3), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i6658_4_lut (.I0(n14706), .I1(n13865), .I2(rd_fifo_en_w), 
            .I3(dc32_fifo_empty), .O(empty_nxt_c_N_636));   // src/fifo_dc_32_lut_gen.v(241[14:26])
    defparam i6658_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1601_2_lut_3_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(state_timeout_counter[2]), .I3(GND_net), .O(n6));   // src/usb3_if.v(180[42:69])
    defparam i1601_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i13870_3_lut_4_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(n2118), .I3(state_timeout_counter[2]), .O(n15945));   // src/usb3_if.v(180[42:69])
    defparam i13870_3_lut_4_lut.LUT_INIT = 16'he010;
    SB_LUT4 i1_2_lut_adj_38 (.I0(n650[4]), .I1(n650[5]), .I2(GND_net), 
            .I3(GND_net), .O(n859));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_adj_38.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(FT_OE_N_496), .I1(state_timeout_counter[1]), .I2(dc32_fifo_almost_full), 
            .I3(num_words_curr_line[5]), .O(n13825));   // src/usb3_if.v(97[9] 199[16])
    defparam i2_4_lut.LUT_INIT = 16'h0031;
    SB_LUT4 i7_4_lut_adj_39 (.I0(state_timeout_counter[2]), .I1(state_timeout_counter[4]), 
            .I2(num_words_curr_line[2]), .I3(n10), .O(n16_adj_1354));
    defparam i7_4_lut_adj_39.LUT_INIT = 16'h0100;
    SB_LUT4 i6_4_lut (.I0(state_timeout_counter[3]), .I1(n8), .I2(n7), 
            .I3(n13825), .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_40 (.I0(n8362), .I1(n15), .I2(n4923), .I3(n16_adj_1354), 
            .O(n8360));   // src/usb3_if.v(59[5:28])
    defparam i1_4_lut_adj_40.LUT_INIT = 16'ha8a0;
    SB_LUT4 i22_4_lut (.I0(n650[3]), .I1(n14577), .I2(n650[2]), .I3(n859), 
            .O(n9));   // src/usb3_if.v(70[8] 83[4])
    defparam i22_4_lut.LUT_INIT = 16'h3f3a;
    SB_LUT4 i1_2_lut_adj_41 (.I0(n650[4]), .I1(n650[8]), .I2(GND_net), 
            .I3(GND_net), .O(n894));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_adj_41.LUT_INIT = 16'heeee;
    SB_LUT4 i13936_4_lut (.I0(n650[2]), .I1(n894), .I2(FT_OE_N_495), .I3(n609), 
            .O(n15965));   // src/usb3_if.v(97[9] 199[16])
    defparam i13936_4_lut.LUT_INIT = 16'h3313;
    SB_DFFESR dc32_fifo_data_in_latched__i2 (.Q(dc32_fifo_data_in_latched[2]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D29_c_2), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i1_2_lut_adj_42 (.I0(DEBUG_5_c), .I1(dc32_fifo_full), .I2(GND_net), 
            .I3(GND_net), .O(wr_fifo_en_w));   // src/usb3_if.v(204[8] 207[4])
    defparam i1_2_lut_adj_42.LUT_INIT = 16'h2222;
    SB_DFFESR dc32_fifo_data_in_latched__i1 (.Q(dc32_fifo_data_in_latched[1]), 
            .C(FIFO_CLK_c), .E(n5217), .D(FIFO_D30_c_1), .R(n5432));   // src/usb3_if.v(86[8] 201[4])
    SB_LUT4 i1_4_lut_adj_43 (.I0(n9698), .I1(n688), .I2(n650[1]), .I3(n609), 
            .O(n7_adj_1355));   // src/usb3_if.v(154[17] 177[20])
    defparam i1_4_lut_adj_43.LUT_INIT = 16'hccec;
    SB_LUT4 FT_OE_I_8_2_lut (.I0(FT_OE_N_496), .I1(dc32_fifo_almost_full), 
            .I2(GND_net), .I3(GND_net), .O(FT_OE_N_495));   // src/usb3_if.v(155[25:87])
    defparam FT_OE_I_8_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i8217_2_lut (.I0(DEBUG_9_c_c), .I1(dc32_fifo_almost_full), .I2(GND_net), 
            .I3(GND_net), .O(n9698));
    defparam i8217_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_44 (.I0(n650[1]), .I1(n650[6]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_1353));
    defparam i1_2_lut_adj_44.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_45 (.I0(state_timeout_counter[4]), .I1(state_timeout_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_1356));   // src/usb3_if.v(86[8] 201[4])
    defparam i1_2_lut_adj_45.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(state_timeout_counter[0]), .I1(state_timeout_counter[2]), 
            .I2(state_timeout_counter[3]), .I3(n6_adj_1356), .O(n609));   // src/usb3_if.v(86[8] 201[4])
    defparam i4_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_4_lut_adj_46 (.I0(n2), .I1(n609), .I2(n32_adj_1353), .I3(n9698), 
            .O(n8_adj_1357));
    defparam i1_4_lut_adj_46.LUT_INIT = 16'heafa;
    SB_LUT4 i1_2_lut_adj_47 (.I0(num_words_curr_line[1]), .I1(num_words_curr_line[4]), 
            .I2(GND_net), .I3(GND_net), .O(n8));
    defparam i1_2_lut_adj_47.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_48 (.I0(num_words_curr_line[3]), .I1(num_words_curr_line[0]), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // src/usb3_if.v(148[44:69])
    defparam i1_2_lut_adj_48.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(num_words_curr_line[5]), .I1(num_words_curr_line[2]), 
            .I2(n7), .I3(n8), .O(FT_OE_N_496));   // src/usb3_if.v(133[21:47])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_49 (.I0(DEBUG_9_c_c), .I1(FT_OE_N_496), .I2(GND_net), 
            .I3(GND_net), .O(FT_OE_N_491));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam i1_2_lut_adj_49.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_50 (.I0(reset_per_frame_latched), .I1(n650[3]), 
            .I2(GND_net), .I3(GND_net), .O(n4923));   // src/usb3_if.v(70[8] 83[4])
    defparam i1_2_lut_adj_50.LUT_INIT = 16'heeee;
    SB_LUT4 i14023_4_lut (.I0(n4), .I1(n7_adj_1358), .I2(n650[4]), .I3(n8_adj_1359), 
            .O(n4990));   // src/usb3_if.v(96[10] 200[8])
    defparam i14023_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_adj_51 (.I0(state_timeout_counter[0]), .I1(n8_adj_1357), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // src/usb3_if.v(64[11:32])
    defparam i1_2_lut_adj_51.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_52 (.I0(reset_per_frame_latched), .I1(n7_adj_1355), 
            .I2(n62), .I3(n4393), .O(n14517));   // src/usb3_if.v(70[8] 83[4])
    defparam i1_4_lut_adj_52.LUT_INIT = 16'h1110;
    SB_LUT4 i1_3_lut_4_lut_adj_53 (.I0(dc32_fifo_empty_latched), .I1(buffer_switch_done_latched), 
            .I2(DEBUG_9_c_c), .I3(n650[0]), .O(n4));   // src/usb3_if.v(70[8] 83[4])
    defparam i1_3_lut_4_lut_adj_53.LUT_INIT = 16'hf700;
    SB_LUT4 i2_3_lut_4_lut_adj_54 (.I0(dc32_fifo_empty_latched), .I1(buffer_switch_done_latched), 
            .I2(DEBUG_9_c_c), .I3(n650[0]), .O(n688));   // src/usb3_if.v(70[8] 83[4])
    defparam i2_3_lut_4_lut_adj_54.LUT_INIT = 16'h0800;
    SB_LUT4 i1_4_lut_adj_55 (.I0(n650[2]), .I1(n650[7]), .I2(FT_OE_N_495), 
            .I3(n609), .O(n709));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_4_lut_adj_55.LUT_INIT = 16'hccec;
    SB_LUT4 i1_4_lut_adj_56 (.I0(DEBUG_9_c_c), .I1(n894), .I2(FT_OE_N_496), 
            .I3(n650[5]), .O(n3510));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_4_lut_adj_56.LUT_INIT = 16'hdccc;
    SB_LUT4 i1_2_lut_3_lut_adj_57 (.I0(reset_per_frame_latched), .I1(n7_adj_1355), 
            .I2(n8464), .I3(GND_net), .O(n2024[3]));
    defparam i1_2_lut_3_lut_adj_57.LUT_INIT = 16'hb0b0;
    SB_LUT4 i1_2_lut_4_lut (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[0]), .I3(state_timeout_counter[2]), 
            .O(n4578));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h5556;
    SB_LUT4 i1_2_lut_adj_58 (.I0(n4393), .I1(n8464), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_1360));
    defparam i1_2_lut_adj_58.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_59 (.I0(n688), .I1(n650[1]), .I2(n18_adj_1360), 
            .I3(n614), .O(n14479));
    defparam i1_4_lut_adj_59.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n650[6]), .I1(n609), .I2(DEBUG_9_c_c), 
            .I3(dc32_fifo_almost_full), .O(n706));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_60 (.I0(n650[1]), .I1(n609), .I2(DEBUG_9_c_c), 
            .I3(dc32_fifo_almost_full), .O(n696));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_3_lut_4_lut_adj_60.LUT_INIT = 16'h0002;
    SB_LUT4 i164_2_lut_3_lut (.I0(n609), .I1(DEBUG_9_c_c), .I2(dc32_fifo_almost_full), 
            .I3(GND_net), .O(n614));   // src/usb3_if.v(115[26] 117[24])
    defparam i164_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2028_3_lut_4_lut (.I0(n650[6]), .I1(n703), .I2(n609), .I3(n9698), 
            .O(n3506));   // src/usb3_if.v(97[9] 199[16])
    defparam i2028_3_lut_4_lut.LUT_INIT = 16'heeec;
    SB_LUT4 i13878_2_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n15944));   // src/usb3_if.v(96[10] 200[8])
    defparam i13878_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1013_i2_4_lut (.I0(n15944), .I1(n7_adj_1355), .I2(n2122), 
            .I3(n2118), .O(n10053));   // src/usb3_if.v(96[10] 200[8])
    defparam mux_1013_i2_4_lut.LUT_INIT = 16'h353f;
    SB_LUT4 i1_2_lut_3_lut_adj_61 (.I0(n650[8]), .I1(reset_per_frame_latched), 
            .I2(n650[3]), .I3(GND_net), .O(n7_adj_1358));   // src/usb3_if.v(96[10] 200[8])
    defparam i1_2_lut_3_lut_adj_61.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_62 (.I0(n650[5]), .I1(n650[7]), .I2(DEBUG_9_c_c), 
            .I3(FT_OE_N_496), .O(n8_adj_1359));   // src/usb3_if.v(96[10] 200[8])
    defparam i2_3_lut_4_lut_adj_62.LUT_INIT = 16'hcecc;
    SB_LUT4 i1_2_lut_3_lut_adj_63 (.I0(FT_OE_N_496), .I1(dc32_fifo_almost_full), 
            .I2(n609), .I3(GND_net), .O(n1236));   // src/usb3_if.v(86[8] 201[4])
    defparam i1_2_lut_3_lut_adj_63.LUT_INIT = 16'hf2f2;
    SB_LUT4 mux_1013_i3_4_lut (.I0(n15945), .I1(n2120), .I2(n2122), .I3(n8464), 
            .O(n2034[2]));   // src/usb3_if.v(96[10] 200[8])
    defparam mux_1013_i3_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 mux_1013_i4_4_lut (.I0(n4578), .I1(n2024[3]), .I2(n2122), 
            .I3(n2118), .O(n2034[3]));   // src/usb3_if.v(96[10] 200[8])
    defparam mux_1013_i4_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i1_3_lut_4_lut_adj_64 (.I0(FT_OE_N_496), .I1(dc32_fifo_almost_full), 
            .I2(n609), .I3(dc32_fifo_empty), .O(n14577));
    defparam i1_3_lut_4_lut_adj_64.LUT_INIT = 16'hf8fd;
    SB_LUT4 i1_2_lut_adj_65 (.I0(reset_per_frame_latched), .I1(n7_adj_1355), 
            .I2(GND_net), .I3(GND_net), .O(n2120));   // src/usb3_if.v(70[8] 83[4])
    defparam i1_2_lut_adj_65.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_66 (.I0(reset_per_frame_latched), .I1(n8_adj_1357), 
            .I2(GND_net), .I3(GND_net), .O(n2118));   // src/usb3_if.v(70[8] 83[4])
    defparam i1_2_lut_adj_66.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut (.I0(reset_per_frame_latched), .I1(n4393), .I2(n7_adj_1355), 
            .I3(GND_net), .O(n2122));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_3_lut_4_lut_adj_67 (.I0(FT_OE_N_495), .I1(n609), .I2(reset_per_frame_latched), 
            .I3(n650[2]), .O(n5098));
    defparam i1_3_lut_4_lut_adj_67.LUT_INIT = 16'hf1f0;
    SB_LUT4 i1_3_lut_4_lut_adj_68 (.I0(n650[4]), .I1(n650[5]), .I2(n5432), 
            .I3(n703), .O(n5217));
    defparam i1_3_lut_4_lut_adj_68.LUT_INIT = 16'hf0fe;
    SB_LUT4 i1_2_lut_3_lut_adj_69 (.I0(n650[5]), .I1(DEBUG_9_c_c), .I2(FT_OE_N_496), 
            .I3(GND_net), .O(n703));
    defparam i1_2_lut_3_lut_adj_69.LUT_INIT = 16'h8080;
    SB_LUT4 i13943_3_lut (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[4]), 
            .I2(n6), .I3(GND_net), .O(n16067));   // src/usb3_if.v(96[10] 200[8])
    defparam i13943_3_lut.LUT_INIT = 16'h3636;
    SB_LUT4 mux_1013_i5_4_lut (.I0(n16067), .I1(n2024[3]), .I2(n2122), 
            .I3(n2118), .O(n2034[4]));   // src/usb3_if.v(96[10] 200[8])
    defparam mux_1013_i5_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i13928_2_lut_3_lut (.I0(FT_OE_N_496), .I1(dc32_fifo_almost_full), 
            .I2(n650[2]), .I3(GND_net), .O(n15955));   // src/usb3_if.v(97[9] 199[16])
    defparam i13928_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_4_lut_adj_70 (.I0(n650[2]), .I1(FT_OE_N_496), .I2(dc32_fifo_almost_full), 
            .I3(n609), .O(n2));   // src/usb3_if.v(97[9] 199[16])
    defparam i1_2_lut_4_lut_adj_70.LUT_INIT = 16'haa08;
    
endmodule

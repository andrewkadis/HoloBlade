-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Jan 31 2020 15:13:18

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    SOUT : in std_logic;
    SCK : out std_logic;
    FIFO_D31 : out std_logic;
    FIFO_D20 : out std_logic;
    FIFO_D13 : out std_logic;
    FIFO_D1 : out std_logic;
    FIFO_CLK : out std_logic;
    FIFO_BE2 : out std_logic;
    DATA15 : out std_logic;
    DATA4 : out std_logic;
    DATA23 : out std_logic;
    RST : out std_logic;
    FIFO_D4 : out std_logic;
    FIFO_D14 : out std_logic;
    UART_TX : out std_logic;
    DATA10 : out std_logic;
    DATA28 : out std_logic;
    DATA19 : out std_logic;
    SDAT : out std_logic;
    FT_SIWU : out std_logic;
    DATA0 : out std_logic;
    FT_WR : out std_logic;
    FIFO_D27 : out std_logic;
    FIFO_D10 : out std_logic;
    FIFO_D0 : out std_logic;
    FIFO_BE3 : out std_logic;
    DEBUG_0 : out std_logic;
    FIFO_D9 : out std_logic;
    DATA14 : out std_logic;
    UPDATE : out std_logic;
    RESET : out std_logic;
    FIFO_D21 : out std_logic;
    FIFO_D12 : out std_logic;
    FIFO_BE1 : out std_logic;
    DEBUG_6 : out std_logic;
    DATA5 : out std_logic;
    DATA24 : out std_logic;
    SEN : out std_logic;
    FIFO_D7 : out std_logic;
    FIFO_D15 : out std_logic;
    ICE_CREST : out std_logic;
    FIFO_D23 : out std_logic;
    DATA3 : out std_logic;
    DATA22 : out std_logic;
    DATA13 : out std_logic;
    INVERT : out std_logic;
    FT_RD : out std_logic;
    FIFO_D5 : out std_logic;
    FIFO_D24 : out std_logic;
    FIFO_D17 : out std_logic;
    DSR : out std_logic;
    DEBUG_3 : out std_logic;
    DATA29 : out std_logic;
    DATA18 : out std_logic;
    ICE_SYSCLK : in std_logic;
    ICE_CLK : out std_logic;
    DATA20 : out std_logic;
    DATA11 : out std_logic;
    DATA1 : out std_logic;
    VALID : out std_logic;
    SYNC : out std_logic;
    FIFO_D3 : out std_logic;
    FIFO_D26 : out std_logic;
    FIFO_D11 : out std_logic;
    DEBUG_1 : out std_logic;
    DATA8 : out std_logic;
    DATA31 : out std_logic;
    DATA27 : out std_logic;
    CTS : out std_logic;
    FIFO_D8 : out std_logic;
    FIFO_D18 : out std_logic;
    DEBUG_8 : out std_logic;
    DCD : out std_logic;
    DATA17 : out std_logic;
    SLM_CLK : out std_logic;
    DATA6 : out std_logic;
    DATA25 : out std_logic;
    ICE_CDONE : out std_logic;
    FIFO_D6 : out std_logic;
    FIFO_D29 : out std_logic;
    UART_RX : in std_logic;
    FIFO_D22 : out std_logic;
    FIFO_BE0 : out std_logic;
    DEBUG_5 : out std_logic;
    DATA12 : out std_logic;
    DTR : out std_logic;
    DATA21 : out std_logic;
    DATA2 : out std_logic;
    FIFO_D25 : out std_logic;
    FIFO_D2 : out std_logic;
    FIFO_D16 : out std_logic;
    DEBUG_2 : out std_logic;
    DATA9 : out std_logic;
    DATA30 : out std_logic;
    FT_TXE : out std_logic;
    FR_RXF : out std_logic;
    FIFO_D19 : out std_logic;
    DEBUG_9 : out std_logic;
    DATA16 : out std_logic;
    FT_OE : out std_logic;
    DATA7 : out std_logic;
    DATA26 : out std_logic;
    FIFO_D30 : out std_logic;
    FIFO_D28 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__13369\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \ICE_SYSCLK_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \RESET_c\ : std_logic;
signal pll_clk_unbuf : std_logic;
signal \GB_BUFFER_pll_clk_unbuf_THRU_CO\ : std_logic;
signal \reset_all_w_N_61_cascade_\ : std_logic;
signal \n2_adj_493_cascade_\ : std_logic;
signal reset_clk_counter_3 : std_logic;
signal reset_clk_counter_0 : std_logic;
signal reset_clk_counter_1 : std_logic;
signal \reset_all_w_N_61\ : std_logic;
signal reset_clk_counter_2 : std_logic;
signal fifo_temp_output_5 : std_logic;
signal \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r\ : std_logic;
signal \mem_LUT_data_raw_r_7\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal fifo_temp_output_4 : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal fifo_temp_output_3 : std_logic;
signal fifo_temp_output_7 : std_logic;
signal fifo_temp_output_6 : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_7\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_4\ : std_logic;
signal fifo_temp_output_2 : std_logic;
signal \n32_cascade_\ : std_logic;
signal n4_adj_500 : std_logic;
signal \n24_adj_499_cascade_\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_2\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3534_cascade_\ : std_logic;
signal \mem_LUT_data_raw_r_2\ : std_logic;
signal n1827 : std_logic;
signal fifo_temp_output_1 : std_logic;
signal \mem_LUT_data_raw_r_0\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_1\ : std_logic;
signal \mem_LUT_data_raw_r_1\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3570\ : std_logic;
signal \mem_LUT_data_raw_r_4\ : std_logic;
signal \mem_LUT_data_raw_r_5\ : std_logic;
signal \rd_addr_p1_w_2_cascade_\ : std_logic;
signal n3428 : std_logic;
signal rd_addr_p1_w_2 : std_logic;
signal \tx_fifo.lscc_fifo_inst.rd_fifo_en_w_cascade_\ : std_logic;
signal \n1_cascade_\ : std_logic;
signal rd_addr_p1_w_1 : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_1\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3528\ : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal \pc_tx.n3461_cascade_\ : std_logic;
signal \pc_tx.n3462\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0\ : std_logic;
signal \pc_tx.r_Bit_Index_2\ : std_logic;
signal \pc_tx.n3456\ : std_logic;
signal \pc_tx.n3455\ : std_logic;
signal \pc_tx.r_Bit_Index_1\ : std_logic;
signal \pc_tx.n3522\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_5\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_5\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3558\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.rd_addr_r_2\ : std_logic;
signal n1 : std_logic;
signal \n3110_cascade_\ : std_logic;
signal wr_addr_p1_w_2 : std_logic;
signal \wr_addr_p1_w_2_cascade_\ : std_logic;
signal wr_addr_r_2 : std_logic;
signal \tx_fifo.lscc_fifo_inst.n2\ : std_logic;
signal n3414 : std_logic;
signal n15_adj_498 : std_logic;
signal wr_fifo_en_w : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3546\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_6\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6\ : std_logic;
signal \mem_LUT_data_raw_r_6\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3540\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_3\ : std_logic;
signal \mem_LUT_data_raw_r_3\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.rd_fifo_en_w\ : std_logic;
signal \bfn_14_3_0_\ : std_logic;
signal \pc_rx.n3060\ : std_logic;
signal \pc_rx.n3061\ : std_logic;
signal \pc_rx.n3062\ : std_logic;
signal \pc_rx.n3063\ : std_logic;
signal \pc_rx.n3064\ : std_logic;
signal \pc_rx.n3065\ : std_logic;
signal \pc_rx.n3066\ : std_logic;
signal \pc_rx.n3067\ : std_logic;
signal \bfn_14_4_0_\ : std_logic;
signal \pc_rx.n3068\ : std_logic;
signal fifo_temp_output_0 : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_0\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3564\ : std_logic;
signal rd_addr_r_1 : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3552\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_4\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_0\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_7\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3_cascade_\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_2\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_6\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n4_cascade_\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n4\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3\ : std_logic;
signal wr_addr_r_1 : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_3\ : std_logic;
signal \pc_rx.n6\ : std_logic;
signal \pc_rx.n3399_cascade_\ : std_logic;
signal \pc_rx.n3430\ : std_logic;
signal \pc_rx.r_Clock_Count_0\ : std_logic;
signal \pc_rx.r_Clock_Count_3\ : std_logic;
signal \pc_rx.r_Clock_Count_2\ : std_logic;
signal \pc_rx.r_Clock_Count_1\ : std_logic;
signal \pc_rx.r_Clock_Count_5\ : std_logic;
signal \pc_rx.r_Clock_Count_6\ : std_logic;
signal \pc_rx.n3400_cascade_\ : std_logic;
signal \pc_rx.r_Clock_Count_4\ : std_logic;
signal \pc_rx.r_Clock_Count_8\ : std_logic;
signal \pc_rx.r_Clock_Count_9\ : std_logic;
signal \pc_rx.n2605_cascade_\ : std_logic;
signal \pc_rx.r_Clock_Count_7\ : std_logic;
signal \r_Bit_Index_0_adj_489\ : std_logic;
signal \pc_tx.o_Tx_Serial_N_212\ : std_logic;
signal \pc_tx.n3\ : std_logic;
signal n1851 : std_logic;
signal \pc_tx.n2597\ : std_logic;
signal \n1851_cascade_\ : std_logic;
signal n1934 : std_logic;
signal pc_data_rx_4 : std_logic;
signal n1697 : std_logic;
signal \n3381_cascade_\ : std_logic;
signal pc_data_rx_0 : std_logic;
signal pc_data_rx_6 : std_logic;
signal spi_busy_falling_edge : std_logic;
signal tx_uart_active_flag : std_logic;
signal \r_SM_Main_2_N_183_0\ : std_logic;
signal spi_busy_prev : std_logic;
signal tx_data_byte_6 : std_logic;
signal tx_addr_byte_5 : std_logic;
signal tx_shift_reg_12 : std_logic;
signal tx_addr_byte_6 : std_logic;
signal tx_shift_reg_13 : std_logic;
signal tx_shift_reg_2 : std_logic;
signal tx_data_byte_5 : std_logic;
signal tx_shift_reg_5 : std_logic;
signal tx_shift_reg_3 : std_logic;
signal tx_shift_reg_4 : std_logic;
signal \INVspi0.tx_shift_reg_i6C_net\ : std_logic;
signal tx_shift_reg_14 : std_logic;
signal tx_addr_byte_7 : std_logic;
signal \DEBUG_8_c\ : std_logic;
signal \INVspi0.tx_shift_reg_i15C_net\ : std_logic;
signal tx_data_byte_4 : std_logic;
signal tx_addr_byte_4 : std_logic;
signal \pc_rx.n3412_cascade_\ : std_logic;
signal \pc_rx.n1946\ : std_logic;
signal \pc_rx.n6_adj_487_cascade_\ : std_logic;
signal \pc_rx.n1849\ : std_logic;
signal \n6_cascade_\ : std_logic;
signal \pc_tx.n1518\ : std_logic;
signal n1782 : std_logic;
signal tx_data_byte_3 : std_logic;
signal pc_data_rx_3 : std_logic;
signal pc_data_rx_2 : std_logic;
signal tx_data_byte_2 : std_logic;
signal pc_data_rx_5 : std_logic;
signal tx_data_byte_0 : std_logic;
signal \INVspi0.tx_shift_reg_i0C_net\ : std_logic;
signal tx_shift_reg_6 : std_logic;
signal \n1763_cascade_\ : std_logic;
signal tx_shift_reg_0 : std_logic;
signal tx_shift_reg_1 : std_logic;
signal tx_addr_byte_3 : std_logic;
signal tx_shift_reg_11 : std_logic;
signal tx_addr_byte_2 : std_logic;
signal tx_shift_reg_9 : std_logic;
signal \n3418_cascade_\ : std_logic;
signal tx_shift_reg_10 : std_logic;
signal n1763 : std_logic;
signal tx_shift_reg_7 : std_logic;
signal tx_addr_byte_0 : std_logic;
signal tx_shift_reg_8 : std_logic;
signal \INVspi0.tx_shift_reg_i7C_net\ : std_logic;
signal \spi0.n3467\ : std_logic;
signal \spi0.n3467_cascade_\ : std_logic;
signal \spi0.state_next_2_cascade_\ : std_logic;
signal \spi0.n500\ : std_logic;
signal \spi0.n4_cascade_\ : std_logic;
signal \spi0.n492\ : std_logic;
signal \spi0.state_next_1_cascade_\ : std_logic;
signal \spi0.n493\ : std_logic;
signal \spi0.n494\ : std_logic;
signal \spi0.n495\ : std_logic;
signal \spi0.n496\ : std_logic;
signal \spi0.n497\ : std_logic;
signal \pc_rx.r_SM_Main_2_N_107_0_cascade_\ : std_logic;
signal \n1801_cascade_\ : std_logic;
signal n6 : std_logic;
signal \pc_rx.r_SM_Main_2_N_107_0\ : std_logic;
signal \pc_rx.n2615\ : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal \pc_rx.n3432\ : std_logic;
signal n3191 : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal n4_adj_495 : std_logic;
signal n4_adj_494 : std_logic;
signal n2527 : std_logic;
signal \n2527_cascade_\ : std_logic;
signal \pc_rx.r_Bit_Index_1\ : std_logic;
signal \pc_rx.r_Bit_Index_2\ : std_logic;
signal pc_data_rx_7 : std_logic;
signal tx_data_byte_7 : std_logic;
signal \rx_shift_reg_15__N_315_cascade_\ : std_logic;
signal rx_buf_byte_7 : std_logic;
signal rx_shift_reg_8 : std_logic;
signal rx_buf_byte_5 : std_logic;
signal rx_shift_reg_7 : std_logic;
signal rx_buf_byte_6 : std_logic;
signal rx_buf_byte_4 : std_logic;
signal spi_busy : std_logic;
signal is_tx_fifo_full_flag : std_logic;
signal fifo_write_cmd : std_logic;
signal wr_addr_r_0 : std_logic;
signal fifo_read_cmd : std_logic;
signal is_fifo_empty_flag : std_logic;
signal rd_addr_r_0 : std_logic;
signal \spi0.n895\ : std_logic;
signal \n888_cascade_\ : std_logic;
signal \spi0.n507\ : std_logic;
signal \spi0.state_next_2__N_307\ : std_logic;
signal \spi0.n3476_cascade_\ : std_logic;
signal \spi0.n25\ : std_logic;
signal \spi0.n13\ : std_logic;
signal n888 : std_logic;
signal \spi0.n1458\ : std_logic;
signal \spi0.n13_cascade_\ : std_logic;
signal \spi0.state_next_0\ : std_logic;
signal \spi0.n499\ : std_logic;
signal \spi0.n498\ : std_logic;
signal \spi0.n502\ : std_logic;
signal \state_next_2__N_308\ : std_logic;
signal \spi0.n911\ : std_logic;
signal \spi0.n503\ : std_logic;
signal \spi0.state_next_2__N_306\ : std_logic;
signal \spi0.state_next_1\ : std_logic;
signal \spi0.n4\ : std_logic;
signal \spi0.n504\ : std_logic;
signal \pc_rx.n1\ : std_logic;
signal \pc_rx.r_SM_Main_2_N_110_0\ : std_logic;
signal \pc_rx.n4\ : std_logic;
signal \pc_rx.n1798\ : std_logic;
signal \pc_rx.r_SM_Main_1\ : std_logic;
signal \pc_rx.r_SM_Main_2_N_104_2\ : std_logic;
signal \pc_rx.r_SM_Main_0\ : std_logic;
signal \pc_rx.r_SM_Main_2\ : std_logic;
signal n1787 : std_logic;
signal \r_Rx_Data\ : std_logic;
signal n4 : std_logic;
signal pc_data_rx_1 : std_logic;
signal reset_all_w : std_logic;
signal rx_shift_reg_6 : std_logic;
signal rx_buf_byte_2 : std_logic;
signal rx_buf_byte_3 : std_logic;
signal rx_buf_byte_1 : std_logic;
signal \rx_shift_reg_15__N_315\ : std_logic;
signal rx_buf_byte_0 : std_logic;
signal rx_shift_reg_4 : std_logic;
signal rx_shift_reg_5 : std_logic;
signal \DEBUG_5_c_c\ : std_logic;
signal rx_shift_reg_0 : std_logic;
signal rx_shift_reg_3 : std_logic;
signal rx_shift_reg_1 : std_logic;
signal n3418 : std_logic;
signal rx_shift_reg_2 : std_logic;
signal \spi0.CS_w\ : std_logic;
signal tx_data_byte_1 : std_logic;
signal tx_addr_byte_1 : std_logic;
signal \DEBUG_9_c\ : std_logic;
signal \DEBUG_6_c\ : std_logic;
signal \pc_tx.n3125_cascade_\ : std_logic;
signal \pc_tx.n29_cascade_\ : std_logic;
signal \r_SM_Main_2_N_180_1\ : std_logic;
signal \pc_tx.r_Clock_Count_0\ : std_logic;
signal \bfn_19_7_0_\ : std_logic;
signal \pc_tx.r_Clock_Count_1\ : std_logic;
signal \pc_tx.n3069\ : std_logic;
signal \pc_tx.r_Clock_Count_2\ : std_logic;
signal \pc_tx.n3070\ : std_logic;
signal \pc_tx.r_Clock_Count_3\ : std_logic;
signal \pc_tx.n3071\ : std_logic;
signal \pc_tx.r_Clock_Count_4\ : std_logic;
signal \pc_tx.n3072\ : std_logic;
signal \pc_tx.r_Clock_Count_5\ : std_logic;
signal \pc_tx.n3073\ : std_logic;
signal \pc_tx.r_Clock_Count_6\ : std_logic;
signal \pc_tx.n3074\ : std_logic;
signal \pc_tx.r_Clock_Count_7\ : std_logic;
signal \pc_tx.n3075\ : std_logic;
signal \pc_tx.n3076\ : std_logic;
signal \pc_tx.r_Clock_Count_8\ : std_logic;
signal \bfn_19_8_0_\ : std_logic;
signal \pc_tx.n3077\ : std_logic;
signal \pc_tx.r_Clock_Count_9\ : std_logic;
signal \pc_tx.n1\ : std_logic;
signal \pc_tx.n1930\ : std_logic;
signal \spi0.n10_cascade_\ : std_logic;
signal \spi0.n1931_cascade_\ : std_logic;
signal \spi0.spi_clk\ : std_logic;
signal state_reg_2 : std_logic;
signal state_reg_0 : std_logic;
signal state_reg_1 : std_logic;
signal \spi0.spi_clk_counter_0\ : std_logic;
signal \bfn_19_10_0_\ : std_logic;
signal \spi0.spi_clk_counter_1\ : std_logic;
signal \spi0.n3055\ : std_logic;
signal \spi0.spi_clk_counter_2\ : std_logic;
signal \spi0.n3056\ : std_logic;
signal \spi0.spi_clk_counter_3\ : std_logic;
signal \spi0.n3057\ : std_logic;
signal \spi0.spi_clk_counter_4\ : std_logic;
signal \spi0.n3058\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \spi0.n3059\ : std_logic;
signal \spi0.spi_clk_counter_5\ : std_logic;
signal \spi0.n1931\ : std_logic;
signal start_transfer_prev : std_logic;
signal n5_adj_496 : std_logic;
signal start_transfer_edge : std_logic;
signal \UART_RX_c\ : std_logic;
signal \pc_rx.r_Rx_Data_R\ : std_logic;
signal \DEBUG_1_c\ : std_logic;
signal uart_rx_complete_prev : std_logic;
signal \DEBUG_2_c\ : std_logic;
signal uart_rx_complete_rising_edge : std_logic;
signal even_byte_flag : std_logic;
signal n25 : std_logic;
signal \bfn_24_8_0_\ : std_logic;
signal n24 : std_logic;
signal n3078 : std_logic;
signal n23 : std_logic;
signal n3079 : std_logic;
signal n22 : std_logic;
signal n3080 : std_logic;
signal n21 : std_logic;
signal n3081 : std_logic;
signal n20 : std_logic;
signal n3082 : std_logic;
signal n19 : std_logic;
signal n3083 : std_logic;
signal n18 : std_logic;
signal n3084 : std_logic;
signal n3085 : std_logic;
signal n17 : std_logic;
signal \bfn_24_9_0_\ : std_logic;
signal n16 : std_logic;
signal n3086 : std_logic;
signal n15 : std_logic;
signal n3087 : std_logic;
signal n14 : std_logic;
signal n3088 : std_logic;
signal n13 : std_logic;
signal n3089 : std_logic;
signal n12 : std_logic;
signal n3090 : std_logic;
signal n11 : std_logic;
signal n3091 : std_logic;
signal n10 : std_logic;
signal n3092 : std_logic;
signal n3093 : std_logic;
signal n9 : std_logic;
signal \bfn_24_10_0_\ : std_logic;
signal n8_adj_490 : std_logic;
signal n3094 : std_logic;
signal n7 : std_logic;
signal n3095 : std_logic;
signal n6_adj_491 : std_logic;
signal n3096 : std_logic;
signal n5 : std_logic;
signal n3097 : std_logic;
signal n4_adj_492 : std_logic;
signal n3098 : std_logic;
signal n3 : std_logic;
signal n3099 : std_logic;
signal n2 : std_logic;
signal n3100 : std_logic;
signal n3101 : std_logic;
signal \bfn_24_11_0_\ : std_logic;
signal \DEBUG_0_c_24\ : std_logic;
signal \SLM_CLK_c\ : std_logic;
signal \GB_BUFFER_SLM_CLK_c_THRU_CO\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \FIFO_BE1_wire\ : std_logic;
signal \VALID_wire\ : std_logic;
signal \FIFO_D14_wire\ : std_logic;
signal \FIFO_CLK_wire\ : std_logic;
signal \DATA30_wire\ : std_logic;
signal \DEBUG_9_wire\ : std_logic;
signal \FIFO_D8_wire\ : std_logic;
signal \DATA7_wire\ : std_logic;
signal \DEBUG_1_wire\ : std_logic;
signal \DATA4_wire\ : std_logic;
signal \FIFO_D26_wire\ : std_logic;
signal \DATA24_wire\ : std_logic;
signal \DTR_wire\ : std_logic;
signal \DATA29_wire\ : std_logic;
signal \FIFO_D16_wire\ : std_logic;
signal \FT_SIWU_wire\ : std_logic;
signal \DEBUG_6_wire\ : std_logic;
signal \DATA17_wire\ : std_logic;
signal \DATA21_wire\ : std_logic;
signal \SYNC_wire\ : std_logic;
signal \SCK_wire\ : std_logic;
signal \UPDATE_wire\ : std_logic;
signal \DATA3_wire\ : std_logic;
signal \DATA18_wire\ : std_logic;
signal \DATA25_wire\ : std_logic;
signal \DEBUG_5_wire\ : std_logic;
signal \RESET_wire\ : std_logic;
signal \DATA22_wire\ : std_logic;
signal \DSR_wire\ : std_logic;
signal \FT_WR_wire\ : std_logic;
signal \FIFO_D0_wire\ : std_logic;
signal \DATA12_wire\ : std_logic;
signal \FIFO_D31_wire\ : std_logic;
signal \DATA11_wire\ : std_logic;
signal \DATA26_wire\ : std_logic;
signal \FT_RD_wire\ : std_logic;
signal \DATA1_wire\ : std_logic;
signal \DATA31_wire\ : std_logic;
signal \FIFO_D10_wire\ : std_logic;
signal \DATA5_wire\ : std_logic;
signal \INVERT_wire\ : std_logic;
signal \FIFO_D13_wire\ : std_logic;
signal \ICE_CREST_wire\ : std_logic;
signal \DEBUG_3_wire\ : std_logic;
signal \FIFO_D17_wire\ : std_logic;
signal \DATA8_wire\ : std_logic;
signal \FIFO_D27_wire\ : std_logic;
signal \FIFO_D1_wire\ : std_logic;
signal \DATA15_wire\ : std_logic;
signal \DATA20_wire\ : std_logic;
signal \SOUT_wire\ : std_logic;
signal \DATA16_wire\ : std_logic;
signal \DATA28_wire\ : std_logic;
signal \FIFO_D23_wire\ : std_logic;
signal \ICE_CLK_wire\ : std_logic;
signal \CTS_wire\ : std_logic;
signal \SLM_CLK_wire\ : std_logic;
signal \FIFO_D20_wire\ : std_logic;
signal \FT_OE_wire\ : std_logic;
signal \FT_TXE_wire\ : std_logic;
signal \FIFO_BE3_wire\ : std_logic;
signal \FIFO_D19_wire\ : std_logic;
signal \FIFO_D7_wire\ : std_logic;
signal \UART_RX_wire\ : std_logic;
signal \FIFO_D6_wire\ : std_logic;
signal \SDAT_wire\ : std_logic;
signal \FIFO_BE0_wire\ : std_logic;
signal \DATA19_wire\ : std_logic;
signal \FIFO_D28_wire\ : std_logic;
signal \DATA14_wire\ : std_logic;
signal \DATA10_wire\ : std_logic;
signal \DATA6_wire\ : std_logic;
signal \FIFO_BE2_wire\ : std_logic;
signal \FIFO_D11_wire\ : std_logic;
signal \FIFO_D3_wire\ : std_logic;
signal \RST_wire\ : std_logic;
signal \FIFO_D25_wire\ : std_logic;
signal \ICE_CDONE_wire\ : std_logic;
signal \SEN_wire\ : std_logic;
signal \DCD_wire\ : std_logic;
signal \FIFO_D9_wire\ : std_logic;
signal \DATA9_wire\ : std_logic;
signal \FIFO_D12_wire\ : std_logic;
signal \DATA27_wire\ : std_logic;
signal \DEBUG_0_wire\ : std_logic;
signal \DATA2_wire\ : std_logic;
signal \FIFO_D24_wire\ : std_logic;
signal \FIFO_D2_wire\ : std_logic;
signal \FIFO_D22_wire\ : std_logic;
signal \UART_TX_wire\ : std_logic;
signal \FIFO_D29_wire\ : std_logic;
signal \FIFO_D21_wire\ : std_logic;
signal \FR_RXF_wire\ : std_logic;
signal \DEBUG_8_wire\ : std_logic;
signal \FIFO_D15_wire\ : std_logic;
signal \DEBUG_2_wire\ : std_logic;
signal \DATA13_wire\ : std_logic;
signal \FIFO_D5_wire\ : std_logic;
signal \FIFO_D4_wire\ : std_logic;
signal \FIFO_D18_wire\ : std_logic;
signal \DATA23_wire\ : std_logic;
signal \ICE_SYSCLK_wire\ : std_logic;
signal \FIFO_D30_wire\ : std_logic;
signal \DATA0_wire\ : std_logic;
signal \clock_inst.pll_config_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    FIFO_BE1 <= \FIFO_BE1_wire\;
    VALID <= \VALID_wire\;
    FIFO_D14 <= \FIFO_D14_wire\;
    FIFO_CLK <= \FIFO_CLK_wire\;
    DATA30 <= \DATA30_wire\;
    DEBUG_9 <= \DEBUG_9_wire\;
    FIFO_D8 <= \FIFO_D8_wire\;
    DATA7 <= \DATA7_wire\;
    DEBUG_1 <= \DEBUG_1_wire\;
    DATA4 <= \DATA4_wire\;
    FIFO_D26 <= \FIFO_D26_wire\;
    DATA24 <= \DATA24_wire\;
    DTR <= \DTR_wire\;
    DATA29 <= \DATA29_wire\;
    FIFO_D16 <= \FIFO_D16_wire\;
    FT_SIWU <= \FT_SIWU_wire\;
    DEBUG_6 <= \DEBUG_6_wire\;
    DATA17 <= \DATA17_wire\;
    DATA21 <= \DATA21_wire\;
    SYNC <= \SYNC_wire\;
    SCK <= \SCK_wire\;
    UPDATE <= \UPDATE_wire\;
    DATA3 <= \DATA3_wire\;
    DATA18 <= \DATA18_wire\;
    DATA25 <= \DATA25_wire\;
    DEBUG_5 <= \DEBUG_5_wire\;
    RESET <= \RESET_wire\;
    DATA22 <= \DATA22_wire\;
    DSR <= \DSR_wire\;
    FT_WR <= \FT_WR_wire\;
    FIFO_D0 <= \FIFO_D0_wire\;
    DATA12 <= \DATA12_wire\;
    FIFO_D31 <= \FIFO_D31_wire\;
    DATA11 <= \DATA11_wire\;
    DATA26 <= \DATA26_wire\;
    FT_RD <= \FT_RD_wire\;
    DATA1 <= \DATA1_wire\;
    DATA31 <= \DATA31_wire\;
    FIFO_D10 <= \FIFO_D10_wire\;
    DATA5 <= \DATA5_wire\;
    INVERT <= \INVERT_wire\;
    FIFO_D13 <= \FIFO_D13_wire\;
    ICE_CREST <= \ICE_CREST_wire\;
    DEBUG_3 <= \DEBUG_3_wire\;
    FIFO_D17 <= \FIFO_D17_wire\;
    DATA8 <= \DATA8_wire\;
    FIFO_D27 <= \FIFO_D27_wire\;
    FIFO_D1 <= \FIFO_D1_wire\;
    DATA15 <= \DATA15_wire\;
    DATA20 <= \DATA20_wire\;
    \SOUT_wire\ <= SOUT;
    DATA16 <= \DATA16_wire\;
    DATA28 <= \DATA28_wire\;
    FIFO_D23 <= \FIFO_D23_wire\;
    ICE_CLK <= \ICE_CLK_wire\;
    CTS <= \CTS_wire\;
    SLM_CLK <= \SLM_CLK_wire\;
    FIFO_D20 <= \FIFO_D20_wire\;
    FT_OE <= \FT_OE_wire\;
    FT_TXE <= \FT_TXE_wire\;
    FIFO_BE3 <= \FIFO_BE3_wire\;
    FIFO_D19 <= \FIFO_D19_wire\;
    FIFO_D7 <= \FIFO_D7_wire\;
    \UART_RX_wire\ <= UART_RX;
    FIFO_D6 <= \FIFO_D6_wire\;
    SDAT <= \SDAT_wire\;
    FIFO_BE0 <= \FIFO_BE0_wire\;
    DATA19 <= \DATA19_wire\;
    FIFO_D28 <= \FIFO_D28_wire\;
    DATA14 <= \DATA14_wire\;
    DATA10 <= \DATA10_wire\;
    DATA6 <= \DATA6_wire\;
    FIFO_BE2 <= \FIFO_BE2_wire\;
    FIFO_D11 <= \FIFO_D11_wire\;
    FIFO_D3 <= \FIFO_D3_wire\;
    RST <= \RST_wire\;
    FIFO_D25 <= \FIFO_D25_wire\;
    ICE_CDONE <= \ICE_CDONE_wire\;
    SEN <= \SEN_wire\;
    DCD <= \DCD_wire\;
    FIFO_D9 <= \FIFO_D9_wire\;
    DATA9 <= \DATA9_wire\;
    FIFO_D12 <= \FIFO_D12_wire\;
    DATA27 <= \DATA27_wire\;
    DEBUG_0 <= \DEBUG_0_wire\;
    DATA2 <= \DATA2_wire\;
    FIFO_D24 <= \FIFO_D24_wire\;
    FIFO_D2 <= \FIFO_D2_wire\;
    FIFO_D22 <= \FIFO_D22_wire\;
    UART_TX <= \UART_TX_wire\;
    FIFO_D29 <= \FIFO_D29_wire\;
    FIFO_D21 <= \FIFO_D21_wire\;
    FR_RXF <= \FR_RXF_wire\;
    DEBUG_8 <= \DEBUG_8_wire\;
    FIFO_D15 <= \FIFO_D15_wire\;
    DEBUG_2 <= \DEBUG_2_wire\;
    DATA13 <= \DATA13_wire\;
    FIFO_D5 <= \FIFO_D5_wire\;
    FIFO_D4 <= \FIFO_D4_wire\;
    FIFO_D18 <= \FIFO_D18_wire\;
    DATA23 <= \DATA23_wire\;
    \ICE_SYSCLK_wire\ <= ICE_SYSCLK;
    FIFO_D30 <= \FIFO_D30_wire\;
    DATA0 <= \DATA0_wire\;
    \clock_inst.pll_config_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';

    \clock_inst.pll_config\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0001",
            DIVQ => "100",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__5166\,
            RESETB => \N__11869\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \clock_inst.pll_config_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => pll_clk_unbuf
        );

    \FIFO_BE1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13369\,
            DIN => \N__13368\,
            DOUT => \N__13367\,
            PACKAGEPIN => \FIFO_BE1_wire\
        );

    \FIFO_BE1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13369\,
            PADOUT => \N__13368\,
            PADIN => \N__13367\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VALID_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13360\,
            DIN => \N__13359\,
            DOUT => \N__13358\,
            PACKAGEPIN => \VALID_wire\
        );

    \VALID_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13360\,
            PADOUT => \N__13359\,
            PADIN => \N__13358\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D14_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13351\,
            DIN => \N__13350\,
            DOUT => \N__13349\,
            PACKAGEPIN => \FIFO_D14_wire\
        );

    \FIFO_D14_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13351\,
            PADOUT => \N__13350\,
            PADIN => \N__13349\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13342\,
            DIN => \N__13341\,
            DOUT => \N__13340\,
            PACKAGEPIN => \FIFO_CLK_wire\
        );

    \FIFO_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13342\,
            PADOUT => \N__13341\,
            PADIN => \N__13340\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA30_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13333\,
            DIN => \N__13332\,
            DOUT => \N__13331\,
            PACKAGEPIN => \DATA30_wire\
        );

    \DATA30_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13333\,
            PADOUT => \N__13332\,
            PADIN => \N__13331\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11928\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_9_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13324\,
            DIN => \N__13323\,
            DOUT => \N__13322\,
            PACKAGEPIN => \DEBUG_9_wire\
        );

    \DEBUG_9_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13324\,
            PADOUT => \N__13323\,
            PADIN => \N__13322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10589\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13315\,
            DIN => \N__13314\,
            DOUT => \N__13313\,
            PACKAGEPIN => \FIFO_D8_wire\
        );

    \FIFO_D8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13315\,
            PADOUT => \N__13314\,
            PADIN => \N__13313\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13306\,
            DIN => \N__13305\,
            DOUT => \N__13304\,
            PACKAGEPIN => \DATA7_wire\
        );

    \DATA7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13306\,
            PADOUT => \N__13305\,
            PADIN => \N__13304\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11981\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13297\,
            DIN => \N__13296\,
            DOUT => \N__13295\,
            PACKAGEPIN => \DEBUG_1_wire\
        );

    \DEBUG_1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13297\,
            PADOUT => \N__13296\,
            PADIN => \N__13295\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11577\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA4_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13288\,
            DIN => \N__13287\,
            DOUT => \N__13286\,
            PACKAGEPIN => \DATA4_wire\
        );

    \DATA4_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13288\,
            PADOUT => \N__13287\,
            PADIN => \N__13286\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11964\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D26_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13279\,
            DIN => \N__13278\,
            DOUT => \N__13277\,
            PACKAGEPIN => \FIFO_D26_wire\
        );

    \FIFO_D26_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13279\,
            PADOUT => \N__13278\,
            PADIN => \N__13277\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA24_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13270\,
            DIN => \N__13269\,
            DOUT => \N__13268\,
            PACKAGEPIN => \DATA24_wire\
        );

    \DATA24_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13270\,
            PADOUT => \N__13269\,
            PADIN => \N__13268\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11930\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DTR_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13261\,
            DIN => \N__13260\,
            DOUT => \N__13259\,
            PACKAGEPIN => \DTR_wire\
        );

    \DTR_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13261\,
            PADOUT => \N__13260\,
            PADIN => \N__13259\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA29_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13252\,
            DIN => \N__13251\,
            DOUT => \N__13250\,
            PACKAGEPIN => \DATA29_wire\
        );

    \DATA29_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13252\,
            PADOUT => \N__13251\,
            PADIN => \N__13250\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11925\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D16_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13243\,
            DIN => \N__13242\,
            DOUT => \N__13241\,
            PACKAGEPIN => \FIFO_D16_wire\
        );

    \FIFO_D16_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13243\,
            PADOUT => \N__13242\,
            PADIN => \N__13241\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_SIWU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13234\,
            DIN => \N__13233\,
            DOUT => \N__13232\,
            PACKAGEPIN => \FT_SIWU_wire\
        );

    \FT_SIWU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13234\,
            PADOUT => \N__13233\,
            PADIN => \N__13232\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_6_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13225\,
            DIN => \N__13224\,
            DOUT => \N__13223\,
            PACKAGEPIN => \DEBUG_6_wire\
        );

    \DEBUG_6_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13225\,
            PADOUT => \N__13224\,
            PADIN => \N__13223\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10532\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA17_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13216\,
            DIN => \N__13215\,
            DOUT => \N__13214\,
            PACKAGEPIN => \DATA17_wire\
        );

    \DATA17_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13216\,
            PADOUT => \N__13215\,
            PADIN => \N__13214\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11985\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA21_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13207\,
            DIN => \N__13206\,
            DOUT => \N__13205\,
            PACKAGEPIN => \DATA21_wire\
        );

    \DATA21_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13207\,
            PADOUT => \N__13206\,
            PADIN => \N__13205\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11966\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13198\,
            DIN => \N__13197\,
            DOUT => \N__13196\,
            PACKAGEPIN => \SYNC_wire\
        );

    \SYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13198\,
            PADOUT => \N__13197\,
            PADIN => \N__13196\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13189\,
            DIN => \N__13188\,
            DOUT => \N__13187\,
            PACKAGEPIN => \SCK_wire\
        );

    \SCK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13189\,
            PADOUT => \N__13188\,
            PADIN => \N__13187\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10542\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UPDATE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13180\,
            DIN => \N__13179\,
            DOUT => \N__13178\,
            PACKAGEPIN => \UPDATE_wire\
        );

    \UPDATE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13180\,
            PADOUT => \N__13179\,
            PADIN => \N__13178\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13171\,
            DIN => \N__13170\,
            DOUT => \N__13169\,
            PACKAGEPIN => \DATA3_wire\
        );

    \DATA3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13171\,
            PADOUT => \N__13170\,
            PADIN => \N__13169\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11863\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA18_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13162\,
            DIN => \N__13161\,
            DOUT => \N__13160\,
            PACKAGEPIN => \DATA18_wire\
        );

    \DATA18_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13162\,
            PADOUT => \N__13161\,
            PADIN => \N__13160\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11984\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA25_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13153\,
            DIN => \N__13152\,
            DOUT => \N__13151\,
            PACKAGEPIN => \DATA25_wire\
        );

    \DATA25_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13153\,
            PADOUT => \N__13152\,
            PADIN => \N__13151\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11862\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_5_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13144\,
            DIN => \N__13143\,
            DOUT => \N__13142\,
            PACKAGEPIN => \DEBUG_5_wire\
        );

    \DEBUG_5_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13144\,
            PADOUT => \N__13143\,
            PADIN => \N__13142\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10233\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESET_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13135\,
            DIN => \N__13134\,
            DOUT => \N__13133\,
            PACKAGEPIN => \RESET_wire\
        );

    \RESET_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13135\,
            PADOUT => \N__13134\,
            PADIN => \N__13133\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5241\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA22_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13126\,
            DIN => \N__13125\,
            DOUT => \N__13124\,
            PACKAGEPIN => \DATA22_wire\
        );

    \DATA22_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13126\,
            PADOUT => \N__13125\,
            PADIN => \N__13124\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11965\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DSR_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13117\,
            DIN => \N__13116\,
            DOUT => \N__13115\,
            PACKAGEPIN => \DSR_wire\
        );

    \DSR_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13117\,
            PADOUT => \N__13116\,
            PADIN => \N__13115\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_WR_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13108\,
            DIN => \N__13107\,
            DOUT => \N__13106\,
            PACKAGEPIN => \FT_WR_wire\
        );

    \FT_WR_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13108\,
            PADOUT => \N__13107\,
            PADIN => \N__13106\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D0_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13099\,
            DIN => \N__13098\,
            DOUT => \N__13097\,
            PACKAGEPIN => \FIFO_D0_wire\
        );

    \FIFO_D0_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13099\,
            PADOUT => \N__13098\,
            PADIN => \N__13097\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA12_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13090\,
            DIN => \N__13089\,
            DOUT => \N__13088\,
            PACKAGEPIN => \DATA12_wire\
        );

    \DATA12_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13090\,
            PADOUT => \N__13089\,
            PADIN => \N__13088\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11832\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D31_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13081\,
            DIN => \N__13080\,
            DOUT => \N__13079\,
            PACKAGEPIN => \FIFO_D31_wire\
        );

    \FIFO_D31_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13081\,
            PADOUT => \N__13080\,
            PADIN => \N__13079\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA11_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13072\,
            DIN => \N__13071\,
            DOUT => \N__13070\,
            PACKAGEPIN => \DATA11_wire\
        );

    \DATA11_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13072\,
            PADOUT => \N__13071\,
            PADIN => \N__13070\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11831\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA26_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13063\,
            DIN => \N__13062\,
            DOUT => \N__13061\,
            PACKAGEPIN => \DATA26_wire\
        );

    \DATA26_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13063\,
            PADOUT => \N__13062\,
            PADIN => \N__13061\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11861\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_RD_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13054\,
            DIN => \N__13053\,
            DOUT => \N__13052\,
            PACKAGEPIN => \FT_RD_wire\
        );

    \FT_RD_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13054\,
            PADOUT => \N__13053\,
            PADIN => \N__13052\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13045\,
            DIN => \N__13044\,
            DOUT => \N__13043\,
            PACKAGEPIN => \DATA1_wire\
        );

    \DATA1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13045\,
            PADOUT => \N__13044\,
            PADIN => \N__13043\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11926\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA31_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13036\,
            DIN => \N__13035\,
            DOUT => \N__13034\,
            PACKAGEPIN => \DATA31_wire\
        );

    \DATA31_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13036\,
            PADOUT => \N__13035\,
            PADIN => \N__13034\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11927\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D10_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13027\,
            DIN => \N__13026\,
            DOUT => \N__13025\,
            PACKAGEPIN => \FIFO_D10_wire\
        );

    \FIFO_D10_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13027\,
            PADOUT => \N__13026\,
            PADIN => \N__13025\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA5_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13018\,
            DIN => \N__13017\,
            DOUT => \N__13016\,
            PACKAGEPIN => \DATA5_wire\
        );

    \DATA5_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13018\,
            PADOUT => \N__13017\,
            PADIN => \N__13016\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11833\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \INVERT_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13009\,
            DIN => \N__13008\,
            DOUT => \N__13007\,
            PACKAGEPIN => \INVERT_wire\
        );

    \INVERT_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13009\,
            PADOUT => \N__13008\,
            PADIN => \N__13007\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D13_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13000\,
            DIN => \N__12999\,
            DOUT => \N__12998\,
            PACKAGEPIN => \FIFO_D13_wire\
        );

    \FIFO_D13_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13000\,
            PADOUT => \N__12999\,
            PADIN => \N__12998\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ICE_CREST_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12991\,
            DIN => \N__12990\,
            DOUT => \N__12989\,
            PACKAGEPIN => \ICE_CREST_wire\
        );

    \ICE_CREST_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12991\,
            PADOUT => \N__12990\,
            PADIN => \N__12989\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12982\,
            DIN => \N__12981\,
            DOUT => \N__12980\,
            PACKAGEPIN => \DEBUG_3_wire\
        );

    \DEBUG_3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12982\,
            PADOUT => \N__12981\,
            PADIN => \N__12980\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D17_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12973\,
            DIN => \N__12972\,
            DOUT => \N__12971\,
            PACKAGEPIN => \FIFO_D17_wire\
        );

    \FIFO_D17_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12973\,
            PADOUT => \N__12972\,
            PADIN => \N__12971\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12964\,
            DIN => \N__12963\,
            DOUT => \N__12962\,
            PACKAGEPIN => \DATA8_wire\
        );

    \DATA8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12964\,
            PADOUT => \N__12963\,
            PADIN => \N__12962\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11801\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D27_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12955\,
            DIN => \N__12954\,
            DOUT => \N__12953\,
            PACKAGEPIN => \FIFO_D27_wire\
        );

    \FIFO_D27_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12955\,
            PADOUT => \N__12954\,
            PADIN => \N__12953\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12946\,
            DIN => \N__12945\,
            DOUT => \N__12944\,
            PACKAGEPIN => \FIFO_D1_wire\
        );

    \FIFO_D1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12946\,
            PADOUT => \N__12945\,
            PADIN => \N__12944\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA15_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12937\,
            DIN => \N__12936\,
            DOUT => \N__12935\,
            PACKAGEPIN => \DATA15_wire\
        );

    \DATA15_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12937\,
            PADOUT => \N__12936\,
            PADIN => \N__12935\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11979\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA20_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12928\,
            DIN => \N__12927\,
            DOUT => \N__12926\,
            PACKAGEPIN => \DATA20_wire\
        );

    \DATA20_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12928\,
            PADOUT => \N__12927\,
            PADIN => \N__12926\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11834\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_5_c_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12919\,
            DIN => \N__12918\,
            DOUT => \N__12917\,
            PACKAGEPIN => \SOUT_wire\
        );

    \DEBUG_5_c_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12919\,
            PADOUT => \N__12918\,
            PADIN => \N__12917\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_5_c_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA16_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12910\,
            DIN => \N__12909\,
            DOUT => \N__12908\,
            PACKAGEPIN => \DATA16_wire\
        );

    \DATA16_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12910\,
            PADOUT => \N__12909\,
            PADIN => \N__12908\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11980\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA28_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12901\,
            DIN => \N__12900\,
            DOUT => \N__12899\,
            PACKAGEPIN => \DATA28_wire\
        );

    \DATA28_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12901\,
            PADOUT => \N__12900\,
            PADIN => \N__12899\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11881\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D23_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12892\,
            DIN => \N__12891\,
            DOUT => \N__12890\,
            PACKAGEPIN => \FIFO_D23_wire\
        );

    \FIFO_D23_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12892\,
            PADOUT => \N__12891\,
            PADIN => \N__12890\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ICE_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12883\,
            DIN => \N__12882\,
            DOUT => \N__12881\,
            PACKAGEPIN => \ICE_CLK_wire\
        );

    \ICE_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12883\,
            PADOUT => \N__12882\,
            PADIN => \N__12881\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CTS_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12874\,
            DIN => \N__12873\,
            DOUT => \N__12872\,
            PACKAGEPIN => \CTS_wire\
        );

    \CTS_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12874\,
            PADOUT => \N__12873\,
            PADIN => \N__12872\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SLM_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12865\,
            DIN => \N__12864\,
            DOUT => \N__12863\,
            PACKAGEPIN => \SLM_CLK_wire\
        );

    \SLM_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12865\,
            PADOUT => \N__12864\,
            PADIN => \N__12863\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12153\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D20_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12856\,
            DIN => \N__12855\,
            DOUT => \N__12854\,
            PACKAGEPIN => \FIFO_D20_wire\
        );

    \FIFO_D20_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12856\,
            PADOUT => \N__12855\,
            PADIN => \N__12854\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_OE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12847\,
            DIN => \N__12846\,
            DOUT => \N__12845\,
            PACKAGEPIN => \FT_OE_wire\
        );

    \FT_OE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12847\,
            PADOUT => \N__12846\,
            PADIN => \N__12845\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_TXE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12838\,
            DIN => \N__12837\,
            DOUT => \N__12836\,
            PACKAGEPIN => \FT_TXE_wire\
        );

    \FT_TXE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12838\,
            PADOUT => \N__12837\,
            PADIN => \N__12836\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_BE3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12829\,
            DIN => \N__12828\,
            DOUT => \N__12827\,
            PACKAGEPIN => \FIFO_BE3_wire\
        );

    \FIFO_BE3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12829\,
            PADOUT => \N__12828\,
            PADIN => \N__12827\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D19_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12820\,
            DIN => \N__12819\,
            DOUT => \N__12818\,
            PACKAGEPIN => \FIFO_D19_wire\
        );

    \FIFO_D19_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12820\,
            PADOUT => \N__12819\,
            PADIN => \N__12818\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12811\,
            DIN => \N__12810\,
            DOUT => \N__12809\,
            PACKAGEPIN => \FIFO_D7_wire\
        );

    \FIFO_D7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12811\,
            PADOUT => \N__12810\,
            PADIN => \N__12809\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UART_RX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12802\,
            DIN => \N__12801\,
            DOUT => \N__12800\,
            PACKAGEPIN => \UART_RX_wire\
        );

    \UART_RX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12802\,
            PADOUT => \N__12801\,
            PADIN => \N__12800\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \UART_RX_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D6_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12793\,
            DIN => \N__12792\,
            DOUT => \N__12791\,
            PACKAGEPIN => \FIFO_D6_wire\
        );

    \FIFO_D6_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12793\,
            PADOUT => \N__12792\,
            PADIN => \N__12791\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SDAT_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12784\,
            DIN => \N__12783\,
            DOUT => \N__12782\,
            PACKAGEPIN => \SDAT_wire\
        );

    \SDAT_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12784\,
            PADOUT => \N__12783\,
            PADIN => \N__12782\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7674\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_BE0_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12775\,
            DIN => \N__12774\,
            DOUT => \N__12773\,
            PACKAGEPIN => \FIFO_BE0_wire\
        );

    \FIFO_BE0_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12775\,
            PADOUT => \N__12774\,
            PADIN => \N__12773\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA19_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12766\,
            DIN => \N__12765\,
            DOUT => \N__12764\,
            PACKAGEPIN => \DATA19_wire\
        );

    \DATA19_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12766\,
            PADOUT => \N__12765\,
            PADIN => \N__12764\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11982\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D28_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12757\,
            DIN => \N__12756\,
            DOUT => \N__12755\,
            PACKAGEPIN => \FIFO_D28_wire\
        );

    \FIFO_D28_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12757\,
            PADOUT => \N__12756\,
            PADIN => \N__12755\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA14_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12748\,
            DIN => \N__12747\,
            DOUT => \N__12746\,
            PACKAGEPIN => \DATA14_wire\
        );

    \DATA14_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12748\,
            PADOUT => \N__12747\,
            PADIN => \N__12746\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11953\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA10_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12739\,
            DIN => \N__12738\,
            DOUT => \N__12737\,
            PACKAGEPIN => \DATA10_wire\
        );

    \DATA10_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12739\,
            PADOUT => \N__12738\,
            PADIN => \N__12737\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11870\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA6_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12730\,
            DIN => \N__12729\,
            DOUT => \N__12728\,
            PACKAGEPIN => \DATA6_wire\
        );

    \DATA6_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12730\,
            PADOUT => \N__12729\,
            PADIN => \N__12728\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11983\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_BE2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12721\,
            DIN => \N__12720\,
            DOUT => \N__12719\,
            PACKAGEPIN => \FIFO_BE2_wire\
        );

    \FIFO_BE2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12721\,
            PADOUT => \N__12720\,
            PADIN => \N__12719\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D11_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12712\,
            DIN => \N__12711\,
            DOUT => \N__12710\,
            PACKAGEPIN => \FIFO_D11_wire\
        );

    \FIFO_D11_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12712\,
            PADOUT => \N__12711\,
            PADIN => \N__12710\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12703\,
            DIN => \N__12702\,
            DOUT => \N__12701\,
            PACKAGEPIN => \FIFO_D3_wire\
        );

    \FIFO_D3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12703\,
            PADOUT => \N__12702\,
            PADIN => \N__12701\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12694\,
            DIN => \N__12693\,
            DOUT => \N__12692\,
            PACKAGEPIN => \RST_wire\
        );

    \RST_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12694\,
            PADOUT => \N__12693\,
            PADIN => \N__12692\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D25_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12685\,
            DIN => \N__12684\,
            DOUT => \N__12683\,
            PACKAGEPIN => \FIFO_D25_wire\
        );

    \FIFO_D25_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12685\,
            PADOUT => \N__12684\,
            PADIN => \N__12683\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ICE_CDONE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12676\,
            DIN => \N__12675\,
            DOUT => \N__12674\,
            PACKAGEPIN => \ICE_CDONE_wire\
        );

    \ICE_CDONE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12676\,
            PADOUT => \N__12675\,
            PADIN => \N__12674\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SEN_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12667\,
            DIN => \N__12666\,
            DOUT => \N__12665\,
            PACKAGEPIN => \SEN_wire\
        );

    \SEN_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12667\,
            PADOUT => \N__12666\,
            PADIN => \N__12665\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DCD_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12658\,
            DIN => \N__12657\,
            DOUT => \N__12656\,
            PACKAGEPIN => \DCD_wire\
        );

    \DCD_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12658\,
            PADOUT => \N__12657\,
            PADIN => \N__12656\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D9_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12649\,
            DIN => \N__12648\,
            DOUT => \N__12647\,
            PACKAGEPIN => \FIFO_D9_wire\
        );

    \FIFO_D9_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12649\,
            PADOUT => \N__12648\,
            PADIN => \N__12647\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA9_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12640\,
            DIN => \N__12639\,
            DOUT => \N__12638\,
            PACKAGEPIN => \DATA9_wire\
        );

    \DATA9_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12640\,
            PADOUT => \N__12639\,
            PADIN => \N__12638\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11911\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D12_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12631\,
            DIN => \N__12630\,
            DOUT => \N__12629\,
            PACKAGEPIN => \FIFO_D12_wire\
        );

    \FIFO_D12_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12631\,
            PADOUT => \N__12630\,
            PADIN => \N__12629\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA27_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12622\,
            DIN => \N__12621\,
            DOUT => \N__12620\,
            PACKAGEPIN => \DATA27_wire\
        );

    \DATA27_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12622\,
            PADOUT => \N__12621\,
            PADIN => \N__12620\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11846\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_0_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12613\,
            DIN => \N__12612\,
            DOUT => \N__12611\,
            PACKAGEPIN => \DEBUG_0_wire\
        );

    \DEBUG_0_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12613\,
            PADOUT => \N__12612\,
            PADIN => \N__12611\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12366\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12604\,
            DIN => \N__12603\,
            DOUT => \N__12602\,
            PACKAGEPIN => \DATA2_wire\
        );

    \DATA2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12604\,
            PADOUT => \N__12603\,
            PADIN => \N__12602\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11734\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D24_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12595\,
            DIN => \N__12594\,
            DOUT => \N__12593\,
            PACKAGEPIN => \FIFO_D24_wire\
        );

    \FIFO_D24_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12595\,
            PADOUT => \N__12594\,
            PADIN => \N__12593\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12586\,
            DIN => \N__12585\,
            DOUT => \N__12584\,
            PACKAGEPIN => \FIFO_D2_wire\
        );

    \FIFO_D2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12586\,
            PADOUT => \N__12585\,
            PADIN => \N__12584\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D22_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12577\,
            DIN => \N__12576\,
            DOUT => \N__12575\,
            PACKAGEPIN => \FIFO_D22_wire\
        );

    \FIFO_D22_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12577\,
            PADOUT => \N__12576\,
            PADIN => \N__12575\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UART_TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12568\,
            DIN => \N__12567\,
            DOUT => \N__12566\,
            PACKAGEPIN => \UART_TX_wire\
        );

    \UART_TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12568\,
            PADOUT => \N__12567\,
            PADIN => \N__12566\,
            CLOCKENABLE => \N__10716\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7062\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__12338\
        );

    \FIFO_D29_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12559\,
            DIN => \N__12558\,
            DOUT => \N__12557\,
            PACKAGEPIN => \FIFO_D29_wire\
        );

    \FIFO_D29_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12559\,
            PADOUT => \N__12558\,
            PADIN => \N__12557\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D21_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12550\,
            DIN => \N__12549\,
            DOUT => \N__12548\,
            PACKAGEPIN => \FIFO_D21_wire\
        );

    \FIFO_D21_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12550\,
            PADOUT => \N__12549\,
            PADIN => \N__12548\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FR_RXF_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12541\,
            DIN => \N__12540\,
            DOUT => \N__12539\,
            PACKAGEPIN => \FR_RXF_wire\
        );

    \FR_RXF_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12541\,
            PADOUT => \N__12540\,
            PADIN => \N__12539\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12532\,
            DIN => \N__12531\,
            DOUT => \N__12530\,
            PACKAGEPIN => \DEBUG_8_wire\
        );

    \DEBUG_8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12532\,
            PADOUT => \N__12531\,
            PADIN => \N__12530\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7670\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D15_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12523\,
            DIN => \N__12522\,
            DOUT => \N__12521\,
            PACKAGEPIN => \FIFO_D15_wire\
        );

    \FIFO_D15_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12523\,
            PADOUT => \N__12522\,
            PADIN => \N__12521\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12514\,
            DIN => \N__12513\,
            DOUT => \N__12512\,
            PACKAGEPIN => \DEBUG_2_wire\
        );

    \DEBUG_2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12514\,
            PADOUT => \N__12513\,
            PADIN => \N__12512\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11535\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA13_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12505\,
            DIN => \N__12504\,
            DOUT => \N__12503\,
            PACKAGEPIN => \DATA13_wire\
        );

    \DATA13_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12505\,
            PADOUT => \N__12504\,
            PADIN => \N__12503\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11952\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D5_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12496\,
            DIN => \N__12495\,
            DOUT => \N__12494\,
            PACKAGEPIN => \FIFO_D5_wire\
        );

    \FIFO_D5_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12496\,
            PADOUT => \N__12495\,
            PADIN => \N__12494\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D4_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12487\,
            DIN => \N__12486\,
            DOUT => \N__12485\,
            PACKAGEPIN => \FIFO_D4_wire\
        );

    \FIFO_D4_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12487\,
            PADOUT => \N__12486\,
            PADIN => \N__12485\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D18_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12478\,
            DIN => \N__12477\,
            DOUT => \N__12476\,
            PACKAGEPIN => \FIFO_D18_wire\
        );

    \FIFO_D18_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12478\,
            PADOUT => \N__12477\,
            PADIN => \N__12476\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA23_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12469\,
            DIN => \N__12468\,
            DOUT => \N__12467\,
            PACKAGEPIN => \DATA23_wire\
        );

    \DATA23_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12469\,
            PADOUT => \N__12468\,
            PADIN => \N__12467\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11963\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ICE_SYSCLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12460\,
            DIN => \N__12459\,
            DOUT => \N__12458\,
            PACKAGEPIN => \ICE_SYSCLK_wire\
        );

    \ICE_SYSCLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12460\,
            PADOUT => \N__12459\,
            PADIN => \N__12458\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ICE_SYSCLK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D30_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12451\,
            DIN => \N__12450\,
            DOUT => \N__12449\,
            PACKAGEPIN => \FIFO_D30_wire\
        );

    \FIFO_D30_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12451\,
            PADOUT => \N__12450\,
            PADIN => \N__12449\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA0_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12442\,
            DIN => \N__12441\,
            DOUT => \N__12440\,
            PACKAGEPIN => \DATA0_wire\
        );

    \DATA0_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12442\,
            PADOUT => \N__12441\,
            PADIN => \N__12440\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11929\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2869\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12420\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__12420\,
            I => n7
        );

    \I__2867\ : InMux
    port map (
            O => \N__12417\,
            I => n3095
        );

    \I__2866\ : InMux
    port map (
            O => \N__12414\,
            I => \N__12411\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__12411\,
            I => n6_adj_491
        );

    \I__2864\ : InMux
    port map (
            O => \N__12408\,
            I => n3096
        );

    \I__2863\ : InMux
    port map (
            O => \N__12405\,
            I => \N__12402\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__12402\,
            I => n5
        );

    \I__2861\ : InMux
    port map (
            O => \N__12399\,
            I => n3097
        );

    \I__2860\ : InMux
    port map (
            O => \N__12396\,
            I => \N__12393\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__12393\,
            I => n4_adj_492
        );

    \I__2858\ : InMux
    port map (
            O => \N__12390\,
            I => n3098
        );

    \I__2857\ : InMux
    port map (
            O => \N__12387\,
            I => \N__12384\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__12384\,
            I => n3
        );

    \I__2855\ : InMux
    port map (
            O => \N__12381\,
            I => n3099
        );

    \I__2854\ : InMux
    port map (
            O => \N__12378\,
            I => \N__12375\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__12375\,
            I => n2
        );

    \I__2852\ : InMux
    port map (
            O => \N__12372\,
            I => n3100
        );

    \I__2851\ : InMux
    port map (
            O => \N__12369\,
            I => \bfn_24_11_0_\
        );

    \I__2850\ : IoInMux
    port map (
            O => \N__12366\,
            I => \N__12363\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__12363\,
            I => \N__12360\
        );

    \I__2848\ : Span4Mux_s3_h
    port map (
            O => \N__12360\,
            I => \N__12357\
        );

    \I__2847\ : Span4Mux_v
    port map (
            O => \N__12357\,
            I => \N__12354\
        );

    \I__2846\ : Span4Mux_v
    port map (
            O => \N__12354\,
            I => \N__12350\
        );

    \I__2845\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12347\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__12350\,
            I => \DEBUG_0_c_24\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__12347\,
            I => \DEBUG_0_c_24\
        );

    \I__2842\ : InMux
    port map (
            O => \N__12342\,
            I => \N__12339\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__12339\,
            I => \N__12328\
        );

    \I__2840\ : ClkMux
    port map (
            O => \N__12338\,
            I => \N__12159\
        );

    \I__2839\ : ClkMux
    port map (
            O => \N__12337\,
            I => \N__12159\
        );

    \I__2838\ : ClkMux
    port map (
            O => \N__12336\,
            I => \N__12159\
        );

    \I__2837\ : ClkMux
    port map (
            O => \N__12335\,
            I => \N__12159\
        );

    \I__2836\ : ClkMux
    port map (
            O => \N__12334\,
            I => \N__12159\
        );

    \I__2835\ : ClkMux
    port map (
            O => \N__12333\,
            I => \N__12159\
        );

    \I__2834\ : ClkMux
    port map (
            O => \N__12332\,
            I => \N__12159\
        );

    \I__2833\ : ClkMux
    port map (
            O => \N__12331\,
            I => \N__12159\
        );

    \I__2832\ : Glb2LocalMux
    port map (
            O => \N__12328\,
            I => \N__12159\
        );

    \I__2831\ : ClkMux
    port map (
            O => \N__12327\,
            I => \N__12159\
        );

    \I__2830\ : ClkMux
    port map (
            O => \N__12326\,
            I => \N__12159\
        );

    \I__2829\ : ClkMux
    port map (
            O => \N__12325\,
            I => \N__12159\
        );

    \I__2828\ : ClkMux
    port map (
            O => \N__12324\,
            I => \N__12159\
        );

    \I__2827\ : ClkMux
    port map (
            O => \N__12323\,
            I => \N__12159\
        );

    \I__2826\ : ClkMux
    port map (
            O => \N__12322\,
            I => \N__12159\
        );

    \I__2825\ : ClkMux
    port map (
            O => \N__12321\,
            I => \N__12159\
        );

    \I__2824\ : ClkMux
    port map (
            O => \N__12320\,
            I => \N__12159\
        );

    \I__2823\ : ClkMux
    port map (
            O => \N__12319\,
            I => \N__12159\
        );

    \I__2822\ : ClkMux
    port map (
            O => \N__12318\,
            I => \N__12159\
        );

    \I__2821\ : ClkMux
    port map (
            O => \N__12317\,
            I => \N__12159\
        );

    \I__2820\ : ClkMux
    port map (
            O => \N__12316\,
            I => \N__12159\
        );

    \I__2819\ : ClkMux
    port map (
            O => \N__12315\,
            I => \N__12159\
        );

    \I__2818\ : ClkMux
    port map (
            O => \N__12314\,
            I => \N__12159\
        );

    \I__2817\ : ClkMux
    port map (
            O => \N__12313\,
            I => \N__12159\
        );

    \I__2816\ : ClkMux
    port map (
            O => \N__12312\,
            I => \N__12159\
        );

    \I__2815\ : ClkMux
    port map (
            O => \N__12311\,
            I => \N__12159\
        );

    \I__2814\ : ClkMux
    port map (
            O => \N__12310\,
            I => \N__12159\
        );

    \I__2813\ : ClkMux
    port map (
            O => \N__12309\,
            I => \N__12159\
        );

    \I__2812\ : ClkMux
    port map (
            O => \N__12308\,
            I => \N__12159\
        );

    \I__2811\ : ClkMux
    port map (
            O => \N__12307\,
            I => \N__12159\
        );

    \I__2810\ : ClkMux
    port map (
            O => \N__12306\,
            I => \N__12159\
        );

    \I__2809\ : ClkMux
    port map (
            O => \N__12305\,
            I => \N__12159\
        );

    \I__2808\ : ClkMux
    port map (
            O => \N__12304\,
            I => \N__12159\
        );

    \I__2807\ : ClkMux
    port map (
            O => \N__12303\,
            I => \N__12159\
        );

    \I__2806\ : ClkMux
    port map (
            O => \N__12302\,
            I => \N__12159\
        );

    \I__2805\ : ClkMux
    port map (
            O => \N__12301\,
            I => \N__12159\
        );

    \I__2804\ : ClkMux
    port map (
            O => \N__12300\,
            I => \N__12159\
        );

    \I__2803\ : ClkMux
    port map (
            O => \N__12299\,
            I => \N__12159\
        );

    \I__2802\ : ClkMux
    port map (
            O => \N__12298\,
            I => \N__12159\
        );

    \I__2801\ : ClkMux
    port map (
            O => \N__12297\,
            I => \N__12159\
        );

    \I__2800\ : ClkMux
    port map (
            O => \N__12296\,
            I => \N__12159\
        );

    \I__2799\ : ClkMux
    port map (
            O => \N__12295\,
            I => \N__12159\
        );

    \I__2798\ : ClkMux
    port map (
            O => \N__12294\,
            I => \N__12159\
        );

    \I__2797\ : ClkMux
    port map (
            O => \N__12293\,
            I => \N__12159\
        );

    \I__2796\ : ClkMux
    port map (
            O => \N__12292\,
            I => \N__12159\
        );

    \I__2795\ : ClkMux
    port map (
            O => \N__12291\,
            I => \N__12159\
        );

    \I__2794\ : ClkMux
    port map (
            O => \N__12290\,
            I => \N__12159\
        );

    \I__2793\ : ClkMux
    port map (
            O => \N__12289\,
            I => \N__12159\
        );

    \I__2792\ : ClkMux
    port map (
            O => \N__12288\,
            I => \N__12159\
        );

    \I__2791\ : ClkMux
    port map (
            O => \N__12287\,
            I => \N__12159\
        );

    \I__2790\ : ClkMux
    port map (
            O => \N__12286\,
            I => \N__12159\
        );

    \I__2789\ : ClkMux
    port map (
            O => \N__12285\,
            I => \N__12159\
        );

    \I__2788\ : ClkMux
    port map (
            O => \N__12284\,
            I => \N__12159\
        );

    \I__2787\ : ClkMux
    port map (
            O => \N__12283\,
            I => \N__12159\
        );

    \I__2786\ : ClkMux
    port map (
            O => \N__12282\,
            I => \N__12159\
        );

    \I__2785\ : ClkMux
    port map (
            O => \N__12281\,
            I => \N__12159\
        );

    \I__2784\ : ClkMux
    port map (
            O => \N__12280\,
            I => \N__12159\
        );

    \I__2783\ : ClkMux
    port map (
            O => \N__12279\,
            I => \N__12159\
        );

    \I__2782\ : ClkMux
    port map (
            O => \N__12278\,
            I => \N__12159\
        );

    \I__2781\ : GlobalMux
    port map (
            O => \N__12159\,
            I => \N__12156\
        );

    \I__2780\ : gio2CtrlBuf
    port map (
            O => \N__12156\,
            I => \SLM_CLK_c\
        );

    \I__2779\ : IoInMux
    port map (
            O => \N__12153\,
            I => \N__12150\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__12150\,
            I => \N__12147\
        );

    \I__2777\ : IoSpan4Mux
    port map (
            O => \N__12147\,
            I => \N__12144\
        );

    \I__2776\ : Span4Mux_s3_h
    port map (
            O => \N__12144\,
            I => \N__12141\
        );

    \I__2775\ : Odrv4
    port map (
            O => \N__12141\,
            I => \GB_BUFFER_SLM_CLK_c_THRU_CO\
        );

    \I__2774\ : InMux
    port map (
            O => \N__12138\,
            I => \N__12135\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__12135\,
            I => n16
        );

    \I__2772\ : InMux
    port map (
            O => \N__12132\,
            I => n3086
        );

    \I__2771\ : InMux
    port map (
            O => \N__12129\,
            I => \N__12126\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__12126\,
            I => n15
        );

    \I__2769\ : InMux
    port map (
            O => \N__12123\,
            I => n3087
        );

    \I__2768\ : InMux
    port map (
            O => \N__12120\,
            I => \N__12117\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__12117\,
            I => n14
        );

    \I__2766\ : InMux
    port map (
            O => \N__12114\,
            I => n3088
        );

    \I__2765\ : InMux
    port map (
            O => \N__12111\,
            I => \N__12108\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__12108\,
            I => n13
        );

    \I__2763\ : InMux
    port map (
            O => \N__12105\,
            I => n3089
        );

    \I__2762\ : InMux
    port map (
            O => \N__12102\,
            I => \N__12099\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__12099\,
            I => n12
        );

    \I__2760\ : InMux
    port map (
            O => \N__12096\,
            I => n3090
        );

    \I__2759\ : InMux
    port map (
            O => \N__12093\,
            I => \N__12090\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__12090\,
            I => n11
        );

    \I__2757\ : InMux
    port map (
            O => \N__12087\,
            I => n3091
        );

    \I__2756\ : InMux
    port map (
            O => \N__12084\,
            I => \N__12081\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__12081\,
            I => n10
        );

    \I__2754\ : InMux
    port map (
            O => \N__12078\,
            I => n3092
        );

    \I__2753\ : InMux
    port map (
            O => \N__12075\,
            I => \N__12072\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__12072\,
            I => n9
        );

    \I__2751\ : InMux
    port map (
            O => \N__12069\,
            I => \bfn_24_10_0_\
        );

    \I__2750\ : InMux
    port map (
            O => \N__12066\,
            I => \N__12063\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__12063\,
            I => n8_adj_490
        );

    \I__2748\ : InMux
    port map (
            O => \N__12060\,
            I => n3094
        );

    \I__2747\ : InMux
    port map (
            O => \N__12057\,
            I => \N__12054\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__12054\,
            I => n24
        );

    \I__2745\ : InMux
    port map (
            O => \N__12051\,
            I => n3078
        );

    \I__2744\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12045\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__12045\,
            I => n23
        );

    \I__2742\ : InMux
    port map (
            O => \N__12042\,
            I => n3079
        );

    \I__2741\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12036\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__12036\,
            I => n22
        );

    \I__2739\ : InMux
    port map (
            O => \N__12033\,
            I => n3080
        );

    \I__2738\ : InMux
    port map (
            O => \N__12030\,
            I => \N__12027\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__12027\,
            I => n21
        );

    \I__2736\ : InMux
    port map (
            O => \N__12024\,
            I => n3081
        );

    \I__2735\ : InMux
    port map (
            O => \N__12021\,
            I => \N__12018\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__12018\,
            I => n20
        );

    \I__2733\ : InMux
    port map (
            O => \N__12015\,
            I => n3082
        );

    \I__2732\ : InMux
    port map (
            O => \N__12012\,
            I => \N__12009\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__12009\,
            I => n19
        );

    \I__2730\ : InMux
    port map (
            O => \N__12006\,
            I => n3083
        );

    \I__2729\ : InMux
    port map (
            O => \N__12003\,
            I => \N__12000\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__12000\,
            I => n18
        );

    \I__2727\ : InMux
    port map (
            O => \N__11997\,
            I => n3084
        );

    \I__2726\ : InMux
    port map (
            O => \N__11994\,
            I => \N__11991\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__11991\,
            I => n17
        );

    \I__2724\ : InMux
    port map (
            O => \N__11988\,
            I => \bfn_24_9_0_\
        );

    \I__2723\ : IoInMux
    port map (
            O => \N__11985\,
            I => \N__11976\
        );

    \I__2722\ : IoInMux
    port map (
            O => \N__11984\,
            I => \N__11973\
        );

    \I__2721\ : IoInMux
    port map (
            O => \N__11983\,
            I => \N__11970\
        );

    \I__2720\ : IoInMux
    port map (
            O => \N__11982\,
            I => \N__11967\
        );

    \I__2719\ : IoInMux
    port map (
            O => \N__11981\,
            I => \N__11960\
        );

    \I__2718\ : IoInMux
    port map (
            O => \N__11980\,
            I => \N__11957\
        );

    \I__2717\ : IoInMux
    port map (
            O => \N__11979\,
            I => \N__11954\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__11976\,
            I => \N__11943\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__11973\,
            I => \N__11943\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__11970\,
            I => \N__11943\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__11967\,
            I => \N__11943\
        );

    \I__2712\ : IoInMux
    port map (
            O => \N__11966\,
            I => \N__11940\
        );

    \I__2711\ : IoInMux
    port map (
            O => \N__11965\,
            I => \N__11937\
        );

    \I__2710\ : IoInMux
    port map (
            O => \N__11964\,
            I => \N__11934\
        );

    \I__2709\ : IoInMux
    port map (
            O => \N__11963\,
            I => \N__11931\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__11960\,
            I => \N__11918\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11957\,
            I => \N__11918\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__11954\,
            I => \N__11918\
        );

    \I__2705\ : IoInMux
    port map (
            O => \N__11953\,
            I => \N__11915\
        );

    \I__2704\ : IoInMux
    port map (
            O => \N__11952\,
            I => \N__11912\
        );

    \I__2703\ : IoSpan4Mux
    port map (
            O => \N__11943\,
            I => \N__11900\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__11940\,
            I => \N__11900\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__11937\,
            I => \N__11900\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__11934\,
            I => \N__11900\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__11931\,
            I => \N__11900\
        );

    \I__2698\ : IoInMux
    port map (
            O => \N__11930\,
            I => \N__11897\
        );

    \I__2697\ : IoInMux
    port map (
            O => \N__11929\,
            I => \N__11894\
        );

    \I__2696\ : IoInMux
    port map (
            O => \N__11928\,
            I => \N__11891\
        );

    \I__2695\ : IoInMux
    port map (
            O => \N__11927\,
            I => \N__11888\
        );

    \I__2694\ : IoInMux
    port map (
            O => \N__11926\,
            I => \N__11885\
        );

    \I__2693\ : IoInMux
    port map (
            O => \N__11925\,
            I => \N__11882\
        );

    \I__2692\ : IoSpan4Mux
    port map (
            O => \N__11918\,
            I => \N__11874\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__11915\,
            I => \N__11874\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__11912\,
            I => \N__11874\
        );

    \I__2689\ : IoInMux
    port map (
            O => \N__11911\,
            I => \N__11871\
        );

    \I__2688\ : IoSpan4Mux
    port map (
            O => \N__11900\,
            I => \N__11864\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__11897\,
            I => \N__11864\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__11894\,
            I => \N__11850\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__11891\,
            I => \N__11850\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__11888\,
            I => \N__11850\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11885\,
            I => \N__11850\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__11882\,
            I => \N__11850\
        );

    \I__2681\ : IoInMux
    port map (
            O => \N__11881\,
            I => \N__11847\
        );

    \I__2680\ : IoSpan4Mux
    port map (
            O => \N__11874\,
            I => \N__11841\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__11871\,
            I => \N__11841\
        );

    \I__2678\ : IoInMux
    port map (
            O => \N__11870\,
            I => \N__11838\
        );

    \I__2677\ : IoInMux
    port map (
            O => \N__11869\,
            I => \N__11835\
        );

    \I__2676\ : IoSpan4Mux
    port map (
            O => \N__11864\,
            I => \N__11828\
        );

    \I__2675\ : IoInMux
    port map (
            O => \N__11863\,
            I => \N__11825\
        );

    \I__2674\ : IoInMux
    port map (
            O => \N__11862\,
            I => \N__11822\
        );

    \I__2673\ : IoInMux
    port map (
            O => \N__11861\,
            I => \N__11819\
        );

    \I__2672\ : IoSpan4Mux
    port map (
            O => \N__11850\,
            I => \N__11814\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__11847\,
            I => \N__11814\
        );

    \I__2670\ : IoInMux
    port map (
            O => \N__11846\,
            I => \N__11811\
        );

    \I__2669\ : IoSpan4Mux
    port map (
            O => \N__11841\,
            I => \N__11806\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__11838\,
            I => \N__11806\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__11835\,
            I => \N__11798\
        );

    \I__2666\ : IoInMux
    port map (
            O => \N__11834\,
            I => \N__11795\
        );

    \I__2665\ : IoInMux
    port map (
            O => \N__11833\,
            I => \N__11792\
        );

    \I__2664\ : IoInMux
    port map (
            O => \N__11832\,
            I => \N__11789\
        );

    \I__2663\ : IoInMux
    port map (
            O => \N__11831\,
            I => \N__11786\
        );

    \I__2662\ : IoSpan4Mux
    port map (
            O => \N__11828\,
            I => \N__11777\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__11825\,
            I => \N__11777\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__11822\,
            I => \N__11777\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__11819\,
            I => \N__11777\
        );

    \I__2658\ : IoSpan4Mux
    port map (
            O => \N__11814\,
            I => \N__11772\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__11811\,
            I => \N__11772\
        );

    \I__2656\ : Span4Mux_s3_h
    port map (
            O => \N__11806\,
            I => \N__11769\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__11805\,
            I => \N__11766\
        );

    \I__2654\ : CascadeMux
    port map (
            O => \N__11804\,
            I => \N__11763\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__11803\,
            I => \N__11759\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__11802\,
            I => \N__11756\
        );

    \I__2651\ : IoInMux
    port map (
            O => \N__11801\,
            I => \N__11753\
        );

    \I__2650\ : IoSpan4Mux
    port map (
            O => \N__11798\,
            I => \N__11750\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__11795\,
            I => \N__11745\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__11792\,
            I => \N__11745\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__11789\,
            I => \N__11740\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__11786\,
            I => \N__11740\
        );

    \I__2645\ : IoSpan4Mux
    port map (
            O => \N__11777\,
            I => \N__11735\
        );

    \I__2644\ : IoSpan4Mux
    port map (
            O => \N__11772\,
            I => \N__11735\
        );

    \I__2643\ : Span4Mux_h
    port map (
            O => \N__11769\,
            I => \N__11731\
        );

    \I__2642\ : InMux
    port map (
            O => \N__11766\,
            I => \N__11726\
        );

    \I__2641\ : InMux
    port map (
            O => \N__11763\,
            I => \N__11726\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11762\,
            I => \N__11719\
        );

    \I__2639\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11719\
        );

    \I__2638\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11719\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__11753\,
            I => \N__11716\
        );

    \I__2636\ : Span4Mux_s2_v
    port map (
            O => \N__11750\,
            I => \N__11713\
        );

    \I__2635\ : Span12Mux_s11_v
    port map (
            O => \N__11745\,
            I => \N__11708\
        );

    \I__2634\ : Span12Mux_s3_h
    port map (
            O => \N__11740\,
            I => \N__11708\
        );

    \I__2633\ : Span4Mux_s3_v
    port map (
            O => \N__11735\,
            I => \N__11705\
        );

    \I__2632\ : IoInMux
    port map (
            O => \N__11734\,
            I => \N__11702\
        );

    \I__2631\ : Span4Mux_v
    port map (
            O => \N__11731\,
            I => \N__11695\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__11726\,
            I => \N__11695\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__11719\,
            I => \N__11695\
        );

    \I__2628\ : Span12Mux_s3_h
    port map (
            O => \N__11716\,
            I => \N__11692\
        );

    \I__2627\ : Span4Mux_v
    port map (
            O => \N__11713\,
            I => \N__11689\
        );

    \I__2626\ : Span12Mux_h
    port map (
            O => \N__11708\,
            I => \N__11682\
        );

    \I__2625\ : Sp12to4
    port map (
            O => \N__11705\,
            I => \N__11682\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__11702\,
            I => \N__11682\
        );

    \I__2623\ : Span4Mux_h
    port map (
            O => \N__11695\,
            I => \N__11679\
        );

    \I__2622\ : Span12Mux_v
    port map (
            O => \N__11692\,
            I => \N__11676\
        );

    \I__2621\ : Sp12to4
    port map (
            O => \N__11689\,
            I => \N__11671\
        );

    \I__2620\ : Span12Mux_s11_v
    port map (
            O => \N__11682\,
            I => \N__11671\
        );

    \I__2619\ : Span4Mux_h
    port map (
            O => \N__11679\,
            I => \N__11668\
        );

    \I__2618\ : Odrv12
    port map (
            O => \N__11676\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2617\ : Odrv12
    port map (
            O => \N__11671\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__11668\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2615\ : InMux
    port map (
            O => \N__11661\,
            I => \spi0.n3059\
        );

    \I__2614\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11654\
        );

    \I__2613\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11651\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__11654\,
            I => \spi0.spi_clk_counter_5\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__11651\,
            I => \spi0.spi_clk_counter_5\
        );

    \I__2610\ : SRMux
    port map (
            O => \N__11646\,
            I => \N__11643\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__11643\,
            I => \N__11640\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__11640\,
            I => \N__11637\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__11637\,
            I => \spi0.n1931\
        );

    \I__2606\ : InMux
    port map (
            O => \N__11634\,
            I => \N__11631\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__11631\,
            I => start_transfer_prev
        );

    \I__2604\ : InMux
    port map (
            O => \N__11628\,
            I => \N__11625\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__11625\,
            I => \N__11621\
        );

    \I__2602\ : InMux
    port map (
            O => \N__11624\,
            I => \N__11618\
        );

    \I__2601\ : Odrv12
    port map (
            O => \N__11621\,
            I => n5_adj_496
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__11618\,
            I => n5_adj_496
        );

    \I__2599\ : InMux
    port map (
            O => \N__11613\,
            I => \N__11610\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__11610\,
            I => \N__11606\
        );

    \I__2597\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11603\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__11606\,
            I => start_transfer_edge
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__11603\,
            I => start_transfer_edge
        );

    \I__2594\ : InMux
    port map (
            O => \N__11598\,
            I => \N__11595\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__11595\,
            I => \N__11592\
        );

    \I__2592\ : Span12Mux_v
    port map (
            O => \N__11592\,
            I => \N__11589\
        );

    \I__2591\ : Odrv12
    port map (
            O => \N__11589\,
            I => \UART_RX_c\
        );

    \I__2590\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11583\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__11583\,
            I => \N__11580\
        );

    \I__2588\ : Odrv12
    port map (
            O => \N__11580\,
            I => \pc_rx.r_Rx_Data_R\
        );

    \I__2587\ : IoInMux
    port map (
            O => \N__11577\,
            I => \N__11574\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__11574\,
            I => \N__11571\
        );

    \I__2585\ : Span4Mux_s2_h
    port map (
            O => \N__11571\,
            I => \N__11566\
        );

    \I__2584\ : InMux
    port map (
            O => \N__11570\,
            I => \N__11561\
        );

    \I__2583\ : InMux
    port map (
            O => \N__11569\,
            I => \N__11561\
        );

    \I__2582\ : Span4Mux_v
    port map (
            O => \N__11566\,
            I => \N__11558\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__11561\,
            I => \N__11555\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__11558\,
            I => \N__11549\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__11555\,
            I => \N__11549\
        );

    \I__2578\ : InMux
    port map (
            O => \N__11554\,
            I => \N__11546\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__11549\,
            I => \DEBUG_1_c\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__11546\,
            I => \DEBUG_1_c\
        );

    \I__2575\ : InMux
    port map (
            O => \N__11541\,
            I => \N__11538\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__11538\,
            I => uart_rx_complete_prev
        );

    \I__2573\ : IoInMux
    port map (
            O => \N__11535\,
            I => \N__11532\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__11532\,
            I => \N__11529\
        );

    \I__2571\ : IoSpan4Mux
    port map (
            O => \N__11529\,
            I => \N__11525\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__11528\,
            I => \N__11521\
        );

    \I__2569\ : Span4Mux_s2_h
    port map (
            O => \N__11525\,
            I => \N__11518\
        );

    \I__2568\ : InMux
    port map (
            O => \N__11524\,
            I => \N__11513\
        );

    \I__2567\ : InMux
    port map (
            O => \N__11521\,
            I => \N__11513\
        );

    \I__2566\ : Span4Mux_h
    port map (
            O => \N__11518\,
            I => \N__11510\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__11513\,
            I => \N__11507\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__11510\,
            I => \DEBUG_2_c\
        );

    \I__2563\ : Odrv4
    port map (
            O => \N__11507\,
            I => \DEBUG_2_c\
        );

    \I__2562\ : InMux
    port map (
            O => \N__11502\,
            I => \N__11493\
        );

    \I__2561\ : InMux
    port map (
            O => \N__11501\,
            I => \N__11490\
        );

    \I__2560\ : InMux
    port map (
            O => \N__11500\,
            I => \N__11487\
        );

    \I__2559\ : InMux
    port map (
            O => \N__11499\,
            I => \N__11484\
        );

    \I__2558\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11479\
        );

    \I__2557\ : InMux
    port map (
            O => \N__11497\,
            I => \N__11479\
        );

    \I__2556\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11476\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__11493\,
            I => \N__11471\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__11490\,
            I => \N__11462\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__11487\,
            I => \N__11462\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__11484\,
            I => \N__11462\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__11479\,
            I => \N__11462\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__11476\,
            I => \N__11451\
        );

    \I__2549\ : InMux
    port map (
            O => \N__11475\,
            I => \N__11448\
        );

    \I__2548\ : InMux
    port map (
            O => \N__11474\,
            I => \N__11444\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__11471\,
            I => \N__11439\
        );

    \I__2546\ : Span4Mux_v
    port map (
            O => \N__11462\,
            I => \N__11439\
        );

    \I__2545\ : InMux
    port map (
            O => \N__11461\,
            I => \N__11434\
        );

    \I__2544\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11434\
        );

    \I__2543\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11431\
        );

    \I__2542\ : InMux
    port map (
            O => \N__11458\,
            I => \N__11426\
        );

    \I__2541\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11426\
        );

    \I__2540\ : InMux
    port map (
            O => \N__11456\,
            I => \N__11423\
        );

    \I__2539\ : InMux
    port map (
            O => \N__11455\,
            I => \N__11420\
        );

    \I__2538\ : InMux
    port map (
            O => \N__11454\,
            I => \N__11417\
        );

    \I__2537\ : Span4Mux_h
    port map (
            O => \N__11451\,
            I => \N__11412\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__11448\,
            I => \N__11412\
        );

    \I__2535\ : InMux
    port map (
            O => \N__11447\,
            I => \N__11409\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__11444\,
            I => \N__11394\
        );

    \I__2533\ : Sp12to4
    port map (
            O => \N__11439\,
            I => \N__11394\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__11434\,
            I => \N__11394\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__11431\,
            I => \N__11394\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__11426\,
            I => \N__11394\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__11423\,
            I => \N__11394\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__11420\,
            I => \N__11394\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__11417\,
            I => \N__11391\
        );

    \I__2526\ : Span4Mux_h
    port map (
            O => \N__11412\,
            I => \N__11386\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__11409\,
            I => \N__11386\
        );

    \I__2524\ : Odrv12
    port map (
            O => \N__11394\,
            I => uart_rx_complete_rising_edge
        );

    \I__2523\ : Odrv12
    port map (
            O => \N__11391\,
            I => uart_rx_complete_rising_edge
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__11386\,
            I => uart_rx_complete_rising_edge
        );

    \I__2521\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11375\
        );

    \I__2520\ : InMux
    port map (
            O => \N__11378\,
            I => \N__11372\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__11375\,
            I => even_byte_flag
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__11372\,
            I => even_byte_flag
        );

    \I__2517\ : InMux
    port map (
            O => \N__11367\,
            I => \N__11364\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__11364\,
            I => n25
        );

    \I__2515\ : InMux
    port map (
            O => \N__11361\,
            I => \bfn_24_8_0_\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__11358\,
            I => \spi0.n10_cascade_\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__11355\,
            I => \spi0.n1931_cascade_\
        );

    \I__2512\ : ClkMux
    port map (
            O => \N__11352\,
            I => \N__11345\
        );

    \I__2511\ : ClkMux
    port map (
            O => \N__11351\,
            I => \N__11342\
        );

    \I__2510\ : ClkMux
    port map (
            O => \N__11350\,
            I => \N__11339\
        );

    \I__2509\ : ClkMux
    port map (
            O => \N__11349\,
            I => \N__11334\
        );

    \I__2508\ : ClkMux
    port map (
            O => \N__11348\,
            I => \N__11329\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__11345\,
            I => \N__11324\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__11342\,
            I => \N__11324\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__11339\,
            I => \N__11321\
        );

    \I__2504\ : ClkMux
    port map (
            O => \N__11338\,
            I => \N__11318\
        );

    \I__2503\ : ClkMux
    port map (
            O => \N__11337\,
            I => \N__11311\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__11334\,
            I => \N__11308\
        );

    \I__2501\ : ClkMux
    port map (
            O => \N__11333\,
            I => \N__11305\
        );

    \I__2500\ : ClkMux
    port map (
            O => \N__11332\,
            I => \N__11302\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__11329\,
            I => \N__11296\
        );

    \I__2498\ : Span4Mux_v
    port map (
            O => \N__11324\,
            I => \N__11296\
        );

    \I__2497\ : Span4Mux_h
    port map (
            O => \N__11321\,
            I => \N__11293\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__11318\,
            I => \N__11290\
        );

    \I__2495\ : ClkMux
    port map (
            O => \N__11317\,
            I => \N__11287\
        );

    \I__2494\ : ClkMux
    port map (
            O => \N__11316\,
            I => \N__11284\
        );

    \I__2493\ : InMux
    port map (
            O => \N__11315\,
            I => \N__11281\
        );

    \I__2492\ : ClkMux
    port map (
            O => \N__11314\,
            I => \N__11278\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__11311\,
            I => \N__11275\
        );

    \I__2490\ : Span4Mux_v
    port map (
            O => \N__11308\,
            I => \N__11268\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__11305\,
            I => \N__11268\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__11302\,
            I => \N__11268\
        );

    \I__2487\ : ClkMux
    port map (
            O => \N__11301\,
            I => \N__11265\
        );

    \I__2486\ : Span4Mux_h
    port map (
            O => \N__11296\,
            I => \N__11261\
        );

    \I__2485\ : Span4Mux_v
    port map (
            O => \N__11293\,
            I => \N__11258\
        );

    \I__2484\ : Span4Mux_v
    port map (
            O => \N__11290\,
            I => \N__11253\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__11287\,
            I => \N__11253\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__11284\,
            I => \N__11246\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__11281\,
            I => \N__11246\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__11278\,
            I => \N__11246\
        );

    \I__2479\ : Span4Mux_v
    port map (
            O => \N__11275\,
            I => \N__11239\
        );

    \I__2478\ : Span4Mux_h
    port map (
            O => \N__11268\,
            I => \N__11239\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__11265\,
            I => \N__11239\
        );

    \I__2476\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11236\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__11261\,
            I => \spi0.spi_clk\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__11258\,
            I => \spi0.spi_clk\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__11253\,
            I => \spi0.spi_clk\
        );

    \I__2472\ : Odrv4
    port map (
            O => \N__11246\,
            I => \spi0.spi_clk\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__11239\,
            I => \spi0.spi_clk\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__11236\,
            I => \spi0.spi_clk\
        );

    \I__2469\ : InMux
    port map (
            O => \N__11223\,
            I => \N__11219\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__11222\,
            I => \N__11215\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__11219\,
            I => \N__11208\
        );

    \I__2466\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11205\
        );

    \I__2465\ : InMux
    port map (
            O => \N__11215\,
            I => \N__11200\
        );

    \I__2464\ : InMux
    port map (
            O => \N__11214\,
            I => \N__11200\
        );

    \I__2463\ : InMux
    port map (
            O => \N__11213\,
            I => \N__11197\
        );

    \I__2462\ : InMux
    port map (
            O => \N__11212\,
            I => \N__11194\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__11211\,
            I => \N__11182\
        );

    \I__2460\ : Span4Mux_h
    port map (
            O => \N__11208\,
            I => \N__11177\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__11205\,
            I => \N__11177\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__11200\,
            I => \N__11174\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__11197\,
            I => \N__11169\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__11194\,
            I => \N__11169\
        );

    \I__2455\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11160\
        );

    \I__2454\ : InMux
    port map (
            O => \N__11192\,
            I => \N__11160\
        );

    \I__2453\ : InMux
    port map (
            O => \N__11191\,
            I => \N__11160\
        );

    \I__2452\ : InMux
    port map (
            O => \N__11190\,
            I => \N__11160\
        );

    \I__2451\ : InMux
    port map (
            O => \N__11189\,
            I => \N__11151\
        );

    \I__2450\ : InMux
    port map (
            O => \N__11188\,
            I => \N__11151\
        );

    \I__2449\ : InMux
    port map (
            O => \N__11187\,
            I => \N__11151\
        );

    \I__2448\ : InMux
    port map (
            O => \N__11186\,
            I => \N__11151\
        );

    \I__2447\ : InMux
    port map (
            O => \N__11185\,
            I => \N__11146\
        );

    \I__2446\ : InMux
    port map (
            O => \N__11182\,
            I => \N__11146\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__11177\,
            I => state_reg_2
        );

    \I__2444\ : Odrv4
    port map (
            O => \N__11174\,
            I => state_reg_2
        );

    \I__2443\ : Odrv4
    port map (
            O => \N__11169\,
            I => state_reg_2
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__11160\,
            I => state_reg_2
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__11151\,
            I => state_reg_2
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__11146\,
            I => state_reg_2
        );

    \I__2439\ : InMux
    port map (
            O => \N__11133\,
            I => \N__11128\
        );

    \I__2438\ : InMux
    port map (
            O => \N__11132\,
            I => \N__11120\
        );

    \I__2437\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11120\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__11128\,
            I => \N__11116\
        );

    \I__2435\ : InMux
    port map (
            O => \N__11127\,
            I => \N__11113\
        );

    \I__2434\ : InMux
    port map (
            O => \N__11126\,
            I => \N__11108\
        );

    \I__2433\ : InMux
    port map (
            O => \N__11125\,
            I => \N__11108\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__11120\,
            I => \N__11099\
        );

    \I__2431\ : InMux
    port map (
            O => \N__11119\,
            I => \N__11096\
        );

    \I__2430\ : Span4Mux_h
    port map (
            O => \N__11116\,
            I => \N__11089\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__11113\,
            I => \N__11089\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__11108\,
            I => \N__11089\
        );

    \I__2427\ : InMux
    port map (
            O => \N__11107\,
            I => \N__11082\
        );

    \I__2426\ : InMux
    port map (
            O => \N__11106\,
            I => \N__11082\
        );

    \I__2425\ : InMux
    port map (
            O => \N__11105\,
            I => \N__11082\
        );

    \I__2424\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11079\
        );

    \I__2423\ : InMux
    port map (
            O => \N__11103\,
            I => \N__11074\
        );

    \I__2422\ : InMux
    port map (
            O => \N__11102\,
            I => \N__11074\
        );

    \I__2421\ : Odrv4
    port map (
            O => \N__11099\,
            I => state_reg_0
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__11096\,
            I => state_reg_0
        );

    \I__2419\ : Odrv4
    port map (
            O => \N__11089\,
            I => state_reg_0
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__11082\,
            I => state_reg_0
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__11079\,
            I => state_reg_0
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__11074\,
            I => state_reg_0
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__11061\,
            I => \N__11049\
        );

    \I__2414\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11046\
        );

    \I__2413\ : SRMux
    port map (
            O => \N__11059\,
            I => \N__11043\
        );

    \I__2412\ : InMux
    port map (
            O => \N__11058\,
            I => \N__11031\
        );

    \I__2411\ : InMux
    port map (
            O => \N__11057\,
            I => \N__11031\
        );

    \I__2410\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11028\
        );

    \I__2409\ : InMux
    port map (
            O => \N__11055\,
            I => \N__11005\
        );

    \I__2408\ : InMux
    port map (
            O => \N__11054\,
            I => \N__11005\
        );

    \I__2407\ : InMux
    port map (
            O => \N__11053\,
            I => \N__11005\
        );

    \I__2406\ : InMux
    port map (
            O => \N__11052\,
            I => \N__11005\
        );

    \I__2405\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11002\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__11046\,
            I => \N__10997\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__11043\,
            I => \N__10997\
        );

    \I__2402\ : InMux
    port map (
            O => \N__11042\,
            I => \N__10982\
        );

    \I__2401\ : InMux
    port map (
            O => \N__11041\,
            I => \N__10982\
        );

    \I__2400\ : InMux
    port map (
            O => \N__11040\,
            I => \N__10982\
        );

    \I__2399\ : InMux
    port map (
            O => \N__11039\,
            I => \N__10982\
        );

    \I__2398\ : InMux
    port map (
            O => \N__11038\,
            I => \N__10982\
        );

    \I__2397\ : InMux
    port map (
            O => \N__11037\,
            I => \N__10982\
        );

    \I__2396\ : InMux
    port map (
            O => \N__11036\,
            I => \N__10982\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__11031\,
            I => \N__10977\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__11028\,
            I => \N__10977\
        );

    \I__2393\ : InMux
    port map (
            O => \N__11027\,
            I => \N__10972\
        );

    \I__2392\ : InMux
    port map (
            O => \N__11026\,
            I => \N__10972\
        );

    \I__2391\ : InMux
    port map (
            O => \N__11025\,
            I => \N__10969\
        );

    \I__2390\ : InMux
    port map (
            O => \N__11024\,
            I => \N__10960\
        );

    \I__2389\ : InMux
    port map (
            O => \N__11023\,
            I => \N__10960\
        );

    \I__2388\ : InMux
    port map (
            O => \N__11022\,
            I => \N__10960\
        );

    \I__2387\ : InMux
    port map (
            O => \N__11021\,
            I => \N__10960\
        );

    \I__2386\ : InMux
    port map (
            O => \N__11020\,
            I => \N__10949\
        );

    \I__2385\ : InMux
    port map (
            O => \N__11019\,
            I => \N__10949\
        );

    \I__2384\ : InMux
    port map (
            O => \N__11018\,
            I => \N__10949\
        );

    \I__2383\ : InMux
    port map (
            O => \N__11017\,
            I => \N__10949\
        );

    \I__2382\ : InMux
    port map (
            O => \N__11016\,
            I => \N__10949\
        );

    \I__2381\ : InMux
    port map (
            O => \N__11015\,
            I => \N__10944\
        );

    \I__2380\ : InMux
    port map (
            O => \N__11014\,
            I => \N__10944\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__11005\,
            I => state_reg_1
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__11002\,
            I => state_reg_1
        );

    \I__2377\ : Odrv12
    port map (
            O => \N__10997\,
            I => state_reg_1
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__10982\,
            I => state_reg_1
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__10977\,
            I => state_reg_1
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__10972\,
            I => state_reg_1
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__10969\,
            I => state_reg_1
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10960\,
            I => state_reg_1
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10949\,
            I => state_reg_1
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__10944\,
            I => state_reg_1
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__10923\,
            I => \N__10920\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10920\,
            I => \N__10916\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10913\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__10916\,
            I => \spi0.spi_clk_counter_0\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__10913\,
            I => \spi0.spi_clk_counter_0\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10908\,
            I => \bfn_19_10_0_\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10905\,
            I => \N__10901\
        );

    \I__2362\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10898\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__10901\,
            I => \spi0.spi_clk_counter_1\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__10898\,
            I => \spi0.spi_clk_counter_1\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10893\,
            I => \spi0.n3055\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10890\,
            I => \N__10886\
        );

    \I__2357\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10883\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10886\,
            I => \spi0.spi_clk_counter_2\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__10883\,
            I => \spi0.spi_clk_counter_2\
        );

    \I__2354\ : InMux
    port map (
            O => \N__10878\,
            I => \spi0.n3056\
        );

    \I__2353\ : InMux
    port map (
            O => \N__10875\,
            I => \N__10871\
        );

    \I__2352\ : InMux
    port map (
            O => \N__10874\,
            I => \N__10868\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__10871\,
            I => \spi0.spi_clk_counter_3\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10868\,
            I => \spi0.spi_clk_counter_3\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10863\,
            I => \spi0.n3057\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10860\,
            I => \N__10856\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10853\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10856\,
            I => \spi0.spi_clk_counter_4\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10853\,
            I => \spi0.spi_clk_counter_4\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10848\,
            I => \spi0.n3058\
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__10845\,
            I => \N__10842\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10842\,
            I => \N__10838\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10841\,
            I => \N__10835\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__10838\,
            I => \pc_tx.r_Clock_Count_2\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10835\,
            I => \pc_tx.r_Clock_Count_2\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10830\,
            I => \pc_tx.n3070\
        );

    \I__2337\ : InMux
    port map (
            O => \N__10827\,
            I => \N__10823\
        );

    \I__2336\ : InMux
    port map (
            O => \N__10826\,
            I => \N__10820\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__10823\,
            I => \pc_tx.r_Clock_Count_3\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__10820\,
            I => \pc_tx.r_Clock_Count_3\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10815\,
            I => \pc_tx.n3071\
        );

    \I__2332\ : InMux
    port map (
            O => \N__10812\,
            I => \N__10808\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10811\,
            I => \N__10805\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__10808\,
            I => \pc_tx.r_Clock_Count_4\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10805\,
            I => \pc_tx.r_Clock_Count_4\
        );

    \I__2328\ : InMux
    port map (
            O => \N__10800\,
            I => \pc_tx.n3072\
        );

    \I__2327\ : InMux
    port map (
            O => \N__10797\,
            I => \N__10793\
        );

    \I__2326\ : InMux
    port map (
            O => \N__10796\,
            I => \N__10790\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10793\,
            I => \pc_tx.r_Clock_Count_5\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__10790\,
            I => \pc_tx.r_Clock_Count_5\
        );

    \I__2323\ : InMux
    port map (
            O => \N__10785\,
            I => \pc_tx.n3073\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10782\,
            I => \N__10778\
        );

    \I__2321\ : InMux
    port map (
            O => \N__10781\,
            I => \N__10775\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__10778\,
            I => \pc_tx.r_Clock_Count_6\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__10775\,
            I => \pc_tx.r_Clock_Count_6\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10770\,
            I => \pc_tx.n3074\
        );

    \I__2317\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10763\
        );

    \I__2316\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10760\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__10763\,
            I => \pc_tx.r_Clock_Count_7\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__10760\,
            I => \pc_tx.r_Clock_Count_7\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10755\,
            I => \pc_tx.n3075\
        );

    \I__2312\ : InMux
    port map (
            O => \N__10752\,
            I => \N__10749\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__10749\,
            I => \N__10745\
        );

    \I__2310\ : InMux
    port map (
            O => \N__10748\,
            I => \N__10742\
        );

    \I__2309\ : Odrv4
    port map (
            O => \N__10745\,
            I => \pc_tx.r_Clock_Count_8\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__10742\,
            I => \pc_tx.r_Clock_Count_8\
        );

    \I__2307\ : InMux
    port map (
            O => \N__10737\,
            I => \bfn_19_8_0_\
        );

    \I__2306\ : InMux
    port map (
            O => \N__10734\,
            I => \pc_tx.n3077\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10731\,
            I => \N__10728\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__10728\,
            I => \N__10724\
        );

    \I__2303\ : InMux
    port map (
            O => \N__10727\,
            I => \N__10721\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__10724\,
            I => \pc_tx.r_Clock_Count_9\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10721\,
            I => \pc_tx.r_Clock_Count_9\
        );

    \I__2300\ : CEMux
    port map (
            O => \N__10716\,
            I => \N__10713\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__10713\,
            I => \N__10710\
        );

    \I__2298\ : Span4Mux_s3_h
    port map (
            O => \N__10710\,
            I => \N__10705\
        );

    \I__2297\ : CEMux
    port map (
            O => \N__10709\,
            I => \N__10702\
        );

    \I__2296\ : CEMux
    port map (
            O => \N__10708\,
            I => \N__10699\
        );

    \I__2295\ : Sp12to4
    port map (
            O => \N__10705\,
            I => \N__10696\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__10702\,
            I => \N__10693\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__10699\,
            I => \N__10690\
        );

    \I__2292\ : Span12Mux_s11_v
    port map (
            O => \N__10696\,
            I => \N__10687\
        );

    \I__2291\ : Span4Mux_v
    port map (
            O => \N__10693\,
            I => \N__10684\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__10690\,
            I => \N__10681\
        );

    \I__2289\ : Odrv12
    port map (
            O => \N__10687\,
            I => \pc_tx.n1\
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__10684\,
            I => \pc_tx.n1\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__10681\,
            I => \pc_tx.n1\
        );

    \I__2286\ : SRMux
    port map (
            O => \N__10674\,
            I => \N__10670\
        );

    \I__2285\ : SRMux
    port map (
            O => \N__10673\,
            I => \N__10667\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__10670\,
            I => \N__10664\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__10667\,
            I => \N__10661\
        );

    \I__2282\ : Span4Mux_h
    port map (
            O => \N__10664\,
            I => \N__10658\
        );

    \I__2281\ : Span4Mux_h
    port map (
            O => \N__10661\,
            I => \N__10655\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__10658\,
            I => \pc_tx.n1930\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__10655\,
            I => \pc_tx.n1930\
        );

    \I__2278\ : InMux
    port map (
            O => \N__10650\,
            I => \N__10647\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__10647\,
            I => \N__10644\
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__10644\,
            I => \spi0.CS_w\
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__10641\,
            I => \N__10638\
        );

    \I__2274\ : InMux
    port map (
            O => \N__10638\,
            I => \N__10635\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__10635\,
            I => \N__10631\
        );

    \I__2272\ : InMux
    port map (
            O => \N__10634\,
            I => \N__10628\
        );

    \I__2271\ : Span4Mux_h
    port map (
            O => \N__10631\,
            I => \N__10624\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__10628\,
            I => \N__10621\
        );

    \I__2269\ : InMux
    port map (
            O => \N__10627\,
            I => \N__10618\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__10624\,
            I => tx_data_byte_1
        );

    \I__2267\ : Odrv12
    port map (
            O => \N__10621\,
            I => tx_data_byte_1
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__10618\,
            I => tx_data_byte_1
        );

    \I__2265\ : InMux
    port map (
            O => \N__10611\,
            I => \N__10608\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__10608\,
            I => \N__10605\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__10605\,
            I => \N__10601\
        );

    \I__2262\ : InMux
    port map (
            O => \N__10604\,
            I => \N__10598\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__10601\,
            I => tx_addr_byte_1
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__10598\,
            I => tx_addr_byte_1
        );

    \I__2259\ : IoInMux
    port map (
            O => \N__10593\,
            I => \N__10590\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__10590\,
            I => \N__10586\
        );

    \I__2257\ : IoInMux
    port map (
            O => \N__10589\,
            I => \N__10583\
        );

    \I__2256\ : Span4Mux_s0_v
    port map (
            O => \N__10586\,
            I => \N__10580\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__10583\,
            I => \N__10577\
        );

    \I__2254\ : Span4Mux_h
    port map (
            O => \N__10580\,
            I => \N__10574\
        );

    \I__2253\ : Span4Mux_s3_v
    port map (
            O => \N__10577\,
            I => \N__10571\
        );

    \I__2252\ : Sp12to4
    port map (
            O => \N__10574\,
            I => \N__10568\
        );

    \I__2251\ : Span4Mux_v
    port map (
            O => \N__10571\,
            I => \N__10565\
        );

    \I__2250\ : Span12Mux_h
    port map (
            O => \N__10568\,
            I => \N__10562\
        );

    \I__2249\ : Span4Mux_v
    port map (
            O => \N__10565\,
            I => \N__10559\
        );

    \I__2248\ : Span12Mux_v
    port map (
            O => \N__10562\,
            I => \N__10555\
        );

    \I__2247\ : Span4Mux_h
    port map (
            O => \N__10559\,
            I => \N__10552\
        );

    \I__2246\ : InMux
    port map (
            O => \N__10558\,
            I => \N__10549\
        );

    \I__2245\ : Odrv12
    port map (
            O => \N__10555\,
            I => \DEBUG_9_c\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__10552\,
            I => \DEBUG_9_c\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__10549\,
            I => \DEBUG_9_c\
        );

    \I__2242\ : IoInMux
    port map (
            O => \N__10542\,
            I => \N__10539\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__10539\,
            I => \N__10536\
        );

    \I__2240\ : Span4Mux_s1_v
    port map (
            O => \N__10536\,
            I => \N__10533\
        );

    \I__2239\ : Span4Mux_v
    port map (
            O => \N__10533\,
            I => \N__10529\
        );

    \I__2238\ : IoInMux
    port map (
            O => \N__10532\,
            I => \N__10526\
        );

    \I__2237\ : Sp12to4
    port map (
            O => \N__10529\,
            I => \N__10523\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__10526\,
            I => \N__10520\
        );

    \I__2235\ : Span12Mux_s10_h
    port map (
            O => \N__10523\,
            I => \N__10517\
        );

    \I__2234\ : IoSpan4Mux
    port map (
            O => \N__10520\,
            I => \N__10514\
        );

    \I__2233\ : Span12Mux_v
    port map (
            O => \N__10517\,
            I => \N__10511\
        );

    \I__2232\ : Sp12to4
    port map (
            O => \N__10514\,
            I => \N__10508\
        );

    \I__2231\ : Span12Mux_h
    port map (
            O => \N__10511\,
            I => \N__10503\
        );

    \I__2230\ : Span12Mux_s9_h
    port map (
            O => \N__10508\,
            I => \N__10503\
        );

    \I__2229\ : Odrv12
    port map (
            O => \N__10503\,
            I => \DEBUG_6_c\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__10500\,
            I => \pc_tx.n3125_cascade_\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__10497\,
            I => \pc_tx.n29_cascade_\
        );

    \I__2226\ : InMux
    port map (
            O => \N__10494\,
            I => \N__10486\
        );

    \I__2225\ : InMux
    port map (
            O => \N__10493\,
            I => \N__10483\
        );

    \I__2224\ : InMux
    port map (
            O => \N__10492\,
            I => \N__10478\
        );

    \I__2223\ : InMux
    port map (
            O => \N__10491\,
            I => \N__10478\
        );

    \I__2222\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10473\
        );

    \I__2221\ : InMux
    port map (
            O => \N__10489\,
            I => \N__10473\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__10486\,
            I => \N__10465\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__10483\,
            I => \N__10465\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__10478\,
            I => \N__10465\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__10473\,
            I => \N__10462\
        );

    \I__2216\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10459\
        );

    \I__2215\ : Span4Mux_h
    port map (
            O => \N__10465\,
            I => \N__10456\
        );

    \I__2214\ : Span4Mux_h
    port map (
            O => \N__10462\,
            I => \N__10453\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__10459\,
            I => \N__10450\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__10456\,
            I => \r_SM_Main_2_N_180_1\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__10453\,
            I => \r_SM_Main_2_N_180_1\
        );

    \I__2210\ : Odrv12
    port map (
            O => \N__10450\,
            I => \r_SM_Main_2_N_180_1\
        );

    \I__2209\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10439\
        );

    \I__2208\ : InMux
    port map (
            O => \N__10442\,
            I => \N__10436\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__10439\,
            I => \pc_tx.r_Clock_Count_0\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__10436\,
            I => \pc_tx.r_Clock_Count_0\
        );

    \I__2205\ : InMux
    port map (
            O => \N__10431\,
            I => \bfn_19_7_0_\
        );

    \I__2204\ : InMux
    port map (
            O => \N__10428\,
            I => \N__10424\
        );

    \I__2203\ : InMux
    port map (
            O => \N__10427\,
            I => \N__10421\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__10424\,
            I => \pc_tx.r_Clock_Count_1\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__10421\,
            I => \pc_tx.r_Clock_Count_1\
        );

    \I__2200\ : InMux
    port map (
            O => \N__10416\,
            I => \pc_tx.n3069\
        );

    \I__2199\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10407\
        );

    \I__2198\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10407\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__10407\,
            I => \N__10402\
        );

    \I__2196\ : InMux
    port map (
            O => \N__10406\,
            I => \N__10397\
        );

    \I__2195\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10397\
        );

    \I__2194\ : Span4Mux_v
    port map (
            O => \N__10402\,
            I => \N__10394\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__10397\,
            I => \N__10391\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__10394\,
            I => \N__10387\
        );

    \I__2191\ : Span4Mux_v
    port map (
            O => \N__10391\,
            I => \N__10384\
        );

    \I__2190\ : InMux
    port map (
            O => \N__10390\,
            I => \N__10381\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__10387\,
            I => rx_buf_byte_3
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__10384\,
            I => rx_buf_byte_3
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__10381\,
            I => rx_buf_byte_3
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__10374\,
            I => \N__10371\
        );

    \I__2185\ : InMux
    port map (
            O => \N__10371\,
            I => \N__10367\
        );

    \I__2184\ : InMux
    port map (
            O => \N__10370\,
            I => \N__10363\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__10367\,
            I => \N__10360\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__10366\,
            I => \N__10356\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__10363\,
            I => \N__10353\
        );

    \I__2180\ : Span4Mux_v
    port map (
            O => \N__10360\,
            I => \N__10350\
        );

    \I__2179\ : InMux
    port map (
            O => \N__10359\,
            I => \N__10347\
        );

    \I__2178\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10344\
        );

    \I__2177\ : Span4Mux_v
    port map (
            O => \N__10353\,
            I => \N__10340\
        );

    \I__2176\ : Sp12to4
    port map (
            O => \N__10350\,
            I => \N__10333\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__10347\,
            I => \N__10333\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__10344\,
            I => \N__10333\
        );

    \I__2173\ : InMux
    port map (
            O => \N__10343\,
            I => \N__10330\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__10340\,
            I => rx_buf_byte_1
        );

    \I__2171\ : Odrv12
    port map (
            O => \N__10333\,
            I => rx_buf_byte_1
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__10330\,
            I => rx_buf_byte_1
        );

    \I__2169\ : InMux
    port map (
            O => \N__10323\,
            I => \N__10308\
        );

    \I__2168\ : InMux
    port map (
            O => \N__10322\,
            I => \N__10308\
        );

    \I__2167\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10308\
        );

    \I__2166\ : InMux
    port map (
            O => \N__10320\,
            I => \N__10308\
        );

    \I__2165\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10301\
        );

    \I__2164\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10301\
        );

    \I__2163\ : InMux
    port map (
            O => \N__10317\,
            I => \N__10301\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__10308\,
            I => \rx_shift_reg_15__N_315\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__10301\,
            I => \rx_shift_reg_15__N_315\
        );

    \I__2160\ : InMux
    port map (
            O => \N__10296\,
            I => \N__10291\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__10295\,
            I => \N__10288\
        );

    \I__2158\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10284\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__10291\,
            I => \N__10281\
        );

    \I__2156\ : InMux
    port map (
            O => \N__10288\,
            I => \N__10276\
        );

    \I__2155\ : InMux
    port map (
            O => \N__10287\,
            I => \N__10276\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__10284\,
            I => \N__10273\
        );

    \I__2153\ : Span4Mux_v
    port map (
            O => \N__10281\,
            I => \N__10268\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__10276\,
            I => \N__10268\
        );

    \I__2151\ : Span4Mux_h
    port map (
            O => \N__10273\,
            I => \N__10262\
        );

    \I__2150\ : Span4Mux_h
    port map (
            O => \N__10268\,
            I => \N__10262\
        );

    \I__2149\ : InMux
    port map (
            O => \N__10267\,
            I => \N__10259\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__10262\,
            I => rx_buf_byte_0
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__10259\,
            I => rx_buf_byte_0
        );

    \I__2146\ : InMux
    port map (
            O => \N__10254\,
            I => \N__10248\
        );

    \I__2145\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10248\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__10248\,
            I => rx_shift_reg_4
        );

    \I__2143\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10241\
        );

    \I__2142\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10238\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__10241\,
            I => rx_shift_reg_5
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__10238\,
            I => rx_shift_reg_5
        );

    \I__2139\ : IoInMux
    port map (
            O => \N__10233\,
            I => \N__10229\
        );

    \I__2138\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10226\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__10229\,
            I => \N__10223\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__10226\,
            I => \N__10220\
        );

    \I__2135\ : Span12Mux_s2_h
    port map (
            O => \N__10223\,
            I => \N__10217\
        );

    \I__2134\ : Span4Mux_v
    port map (
            O => \N__10220\,
            I => \N__10214\
        );

    \I__2133\ : Span12Mux_h
    port map (
            O => \N__10217\,
            I => \N__10211\
        );

    \I__2132\ : Span4Mux_h
    port map (
            O => \N__10214\,
            I => \N__10208\
        );

    \I__2131\ : Span12Mux_h
    port map (
            O => \N__10211\,
            I => \N__10205\
        );

    \I__2130\ : Sp12to4
    port map (
            O => \N__10208\,
            I => \N__10202\
        );

    \I__2129\ : Span12Mux_v
    port map (
            O => \N__10205\,
            I => \N__10197\
        );

    \I__2128\ : Span12Mux_h
    port map (
            O => \N__10202\,
            I => \N__10197\
        );

    \I__2127\ : Span12Mux_v
    port map (
            O => \N__10197\,
            I => \N__10194\
        );

    \I__2126\ : Odrv12
    port map (
            O => \N__10194\,
            I => \DEBUG_5_c_c\
        );

    \I__2125\ : InMux
    port map (
            O => \N__10191\,
            I => \N__10188\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__10188\,
            I => rx_shift_reg_0
        );

    \I__2123\ : InMux
    port map (
            O => \N__10185\,
            I => \N__10181\
        );

    \I__2122\ : InMux
    port map (
            O => \N__10184\,
            I => \N__10178\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__10181\,
            I => rx_shift_reg_3
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__10178\,
            I => rx_shift_reg_3
        );

    \I__2119\ : InMux
    port map (
            O => \N__10173\,
            I => \N__10169\
        );

    \I__2118\ : InMux
    port map (
            O => \N__10172\,
            I => \N__10166\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__10169\,
            I => rx_shift_reg_1
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__10166\,
            I => rx_shift_reg_1
        );

    \I__2115\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10148\
        );

    \I__2114\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10148\
        );

    \I__2113\ : InMux
    port map (
            O => \N__10159\,
            I => \N__10148\
        );

    \I__2112\ : InMux
    port map (
            O => \N__10158\,
            I => \N__10141\
        );

    \I__2111\ : InMux
    port map (
            O => \N__10157\,
            I => \N__10141\
        );

    \I__2110\ : InMux
    port map (
            O => \N__10156\,
            I => \N__10136\
        );

    \I__2109\ : InMux
    port map (
            O => \N__10155\,
            I => \N__10136\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__10148\,
            I => \N__10133\
        );

    \I__2107\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10114\
        );

    \I__2106\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10114\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__10141\,
            I => \N__10109\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__10136\,
            I => \N__10109\
        );

    \I__2103\ : Span4Mux_h
    port map (
            O => \N__10133\,
            I => \N__10106\
        );

    \I__2102\ : InMux
    port map (
            O => \N__10132\,
            I => \N__10101\
        );

    \I__2101\ : InMux
    port map (
            O => \N__10131\,
            I => \N__10101\
        );

    \I__2100\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10088\
        );

    \I__2099\ : InMux
    port map (
            O => \N__10129\,
            I => \N__10088\
        );

    \I__2098\ : InMux
    port map (
            O => \N__10128\,
            I => \N__10088\
        );

    \I__2097\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10088\
        );

    \I__2096\ : InMux
    port map (
            O => \N__10126\,
            I => \N__10088\
        );

    \I__2095\ : InMux
    port map (
            O => \N__10125\,
            I => \N__10088\
        );

    \I__2094\ : InMux
    port map (
            O => \N__10124\,
            I => \N__10077\
        );

    \I__2093\ : InMux
    port map (
            O => \N__10123\,
            I => \N__10077\
        );

    \I__2092\ : InMux
    port map (
            O => \N__10122\,
            I => \N__10077\
        );

    \I__2091\ : InMux
    port map (
            O => \N__10121\,
            I => \N__10077\
        );

    \I__2090\ : InMux
    port map (
            O => \N__10120\,
            I => \N__10077\
        );

    \I__2089\ : InMux
    port map (
            O => \N__10119\,
            I => \N__10074\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__10114\,
            I => n3418
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__10109\,
            I => n3418
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__10106\,
            I => n3418
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__10101\,
            I => n3418
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__10088\,
            I => n3418
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__10077\,
            I => n3418
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__10074\,
            I => n3418
        );

    \I__2081\ : InMux
    port map (
            O => \N__10059\,
            I => \N__10055\
        );

    \I__2080\ : InMux
    port map (
            O => \N__10058\,
            I => \N__10052\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__10055\,
            I => rx_shift_reg_2
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__10052\,
            I => rx_shift_reg_2
        );

    \I__2077\ : InMux
    port map (
            O => \N__10047\,
            I => \N__10044\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__10044\,
            I => \pc_rx.n1798\
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__10041\,
            I => \N__10029\
        );

    \I__2074\ : InMux
    port map (
            O => \N__10040\,
            I => \N__10022\
        );

    \I__2073\ : InMux
    port map (
            O => \N__10039\,
            I => \N__10022\
        );

    \I__2072\ : InMux
    port map (
            O => \N__10038\,
            I => \N__10017\
        );

    \I__2071\ : InMux
    port map (
            O => \N__10037\,
            I => \N__10017\
        );

    \I__2070\ : InMux
    port map (
            O => \N__10036\,
            I => \N__10012\
        );

    \I__2069\ : InMux
    port map (
            O => \N__10035\,
            I => \N__10012\
        );

    \I__2068\ : InMux
    port map (
            O => \N__10034\,
            I => \N__10005\
        );

    \I__2067\ : InMux
    port map (
            O => \N__10033\,
            I => \N__10005\
        );

    \I__2066\ : InMux
    port map (
            O => \N__10032\,
            I => \N__10005\
        );

    \I__2065\ : InMux
    port map (
            O => \N__10029\,
            I => \N__10002\
        );

    \I__2064\ : InMux
    port map (
            O => \N__10028\,
            I => \N__9997\
        );

    \I__2063\ : InMux
    port map (
            O => \N__10027\,
            I => \N__9997\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__10022\,
            I => \pc_rx.r_SM_Main_1\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__10017\,
            I => \pc_rx.r_SM_Main_1\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__10012\,
            I => \pc_rx.r_SM_Main_1\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__10005\,
            I => \pc_rx.r_SM_Main_1\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__10002\,
            I => \pc_rx.r_SM_Main_1\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__9997\,
            I => \pc_rx.r_SM_Main_1\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9984\,
            I => \N__9977\
        );

    \I__2055\ : InMux
    port map (
            O => \N__9983\,
            I => \N__9968\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9982\,
            I => \N__9968\
        );

    \I__2053\ : InMux
    port map (
            O => \N__9981\,
            I => \N__9968\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9968\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__9977\,
            I => \N__9962\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9968\,
            I => \N__9962\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9959\
        );

    \I__2048\ : Span4Mux_v
    port map (
            O => \N__9962\,
            I => \N__9951\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9959\,
            I => \N__9951\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9958\,
            I => \N__9948\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9957\,
            I => \N__9942\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9956\,
            I => \N__9942\
        );

    \I__2043\ : Span4Mux_h
    port map (
            O => \N__9951\,
            I => \N__9937\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9948\,
            I => \N__9937\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9947\,
            I => \N__9934\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9942\,
            I => \pc_rx.r_SM_Main_2_N_104_2\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__9937\,
            I => \pc_rx.r_SM_Main_2_N_104_2\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9934\,
            I => \pc_rx.r_SM_Main_2_N_104_2\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__9927\,
            I => \N__9922\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__9926\,
            I => \N__9916\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__9925\,
            I => \N__9913\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9922\,
            I => \N__9906\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9921\,
            I => \N__9903\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9920\,
            I => \N__9898\
        );

    \I__2031\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9898\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9916\,
            I => \N__9891\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9913\,
            I => \N__9891\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9912\,
            I => \N__9891\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9886\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9910\,
            I => \N__9886\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9909\,
            I => \N__9883\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9906\,
            I => \pc_rx.r_SM_Main_0\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9903\,
            I => \pc_rx.r_SM_Main_0\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__9898\,
            I => \pc_rx.r_SM_Main_0\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9891\,
            I => \pc_rx.r_SM_Main_0\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__9886\,
            I => \pc_rx.r_SM_Main_0\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__9883\,
            I => \pc_rx.r_SM_Main_0\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9870\,
            I => \N__9863\
        );

    \I__2017\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9863\
        );

    \I__2016\ : SRMux
    port map (
            O => \N__9868\,
            I => \N__9860\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9863\,
            I => \N__9853\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__9860\,
            I => \N__9853\
        );

    \I__2013\ : InMux
    port map (
            O => \N__9859\,
            I => \N__9850\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__9858\,
            I => \N__9843\
        );

    \I__2011\ : Span4Mux_h
    port map (
            O => \N__9853\,
            I => \N__9840\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__9850\,
            I => \N__9837\
        );

    \I__2009\ : InMux
    port map (
            O => \N__9849\,
            I => \N__9832\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9848\,
            I => \N__9832\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9829\
        );

    \I__2006\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9826\
        );

    \I__2005\ : InMux
    port map (
            O => \N__9843\,
            I => \N__9823\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__9840\,
            I => \pc_rx.r_SM_Main_2\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__9837\,
            I => \pc_rx.r_SM_Main_2\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9832\,
            I => \pc_rx.r_SM_Main_2\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9829\,
            I => \pc_rx.r_SM_Main_2\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9826\,
            I => \pc_rx.r_SM_Main_2\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__9823\,
            I => \pc_rx.r_SM_Main_2\
        );

    \I__1998\ : InMux
    port map (
            O => \N__9810\,
            I => \N__9806\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9809\,
            I => \N__9801\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__9806\,
            I => \N__9798\
        );

    \I__1995\ : InMux
    port map (
            O => \N__9805\,
            I => \N__9793\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9804\,
            I => \N__9793\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9801\,
            I => \N__9790\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__9798\,
            I => \N__9787\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__9793\,
            I => \N__9784\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__9790\,
            I => n1787
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__9787\,
            I => n1787
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__9784\,
            I => n1787
        );

    \I__1987\ : InMux
    port map (
            O => \N__9777\,
            I => \N__9763\
        );

    \I__1986\ : InMux
    port map (
            O => \N__9776\,
            I => \N__9763\
        );

    \I__1985\ : InMux
    port map (
            O => \N__9775\,
            I => \N__9763\
        );

    \I__1984\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9755\
        );

    \I__1983\ : InMux
    port map (
            O => \N__9773\,
            I => \N__9755\
        );

    \I__1982\ : InMux
    port map (
            O => \N__9772\,
            I => \N__9755\
        );

    \I__1981\ : InMux
    port map (
            O => \N__9771\,
            I => \N__9750\
        );

    \I__1980\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9750\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__9763\,
            I => \N__9747\
        );

    \I__1978\ : InMux
    port map (
            O => \N__9762\,
            I => \N__9744\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__9755\,
            I => \N__9741\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__9750\,
            I => \N__9738\
        );

    \I__1975\ : Span4Mux_v
    port map (
            O => \N__9747\,
            I => \N__9732\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__9744\,
            I => \N__9729\
        );

    \I__1973\ : Span4Mux_v
    port map (
            O => \N__9741\,
            I => \N__9724\
        );

    \I__1972\ : Span4Mux_v
    port map (
            O => \N__9738\,
            I => \N__9724\
        );

    \I__1971\ : InMux
    port map (
            O => \N__9737\,
            I => \N__9721\
        );

    \I__1970\ : InMux
    port map (
            O => \N__9736\,
            I => \N__9716\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9735\,
            I => \N__9716\
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__9732\,
            I => \r_Rx_Data\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__9729\,
            I => \r_Rx_Data\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__9724\,
            I => \r_Rx_Data\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__9721\,
            I => \r_Rx_Data\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__9716\,
            I => \r_Rx_Data\
        );

    \I__1963\ : InMux
    port map (
            O => \N__9705\,
            I => \N__9701\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9698\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__9701\,
            I => \N__9695\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__9698\,
            I => n4
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__9695\,
            I => n4
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__9690\,
            I => \N__9686\
        );

    \I__1957\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9683\
        );

    \I__1956\ : InMux
    port map (
            O => \N__9686\,
            I => \N__9680\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__9683\,
            I => pc_data_rx_1
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__9680\,
            I => pc_data_rx_1
        );

    \I__1953\ : SRMux
    port map (
            O => \N__9675\,
            I => \N__9666\
        );

    \I__1952\ : InMux
    port map (
            O => \N__9674\,
            I => \N__9653\
        );

    \I__1951\ : InMux
    port map (
            O => \N__9673\,
            I => \N__9653\
        );

    \I__1950\ : SRMux
    port map (
            O => \N__9672\,
            I => \N__9653\
        );

    \I__1949\ : SRMux
    port map (
            O => \N__9671\,
            I => \N__9650\
        );

    \I__1948\ : SRMux
    port map (
            O => \N__9670\,
            I => \N__9647\
        );

    \I__1947\ : SRMux
    port map (
            O => \N__9669\,
            I => \N__9644\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__9666\,
            I => \N__9637\
        );

    \I__1945\ : InMux
    port map (
            O => \N__9665\,
            I => \N__9628\
        );

    \I__1944\ : InMux
    port map (
            O => \N__9664\,
            I => \N__9628\
        );

    \I__1943\ : InMux
    port map (
            O => \N__9663\,
            I => \N__9625\
        );

    \I__1942\ : InMux
    port map (
            O => \N__9662\,
            I => \N__9618\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9618\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9618\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__9653\,
            I => \N__9614\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__9650\,
            I => \N__9609\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__9647\,
            I => \N__9609\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__9644\,
            I => \N__9606\
        );

    \I__1935\ : SRMux
    port map (
            O => \N__9643\,
            I => \N__9603\
        );

    \I__1934\ : InMux
    port map (
            O => \N__9642\,
            I => \N__9596\
        );

    \I__1933\ : InMux
    port map (
            O => \N__9641\,
            I => \N__9596\
        );

    \I__1932\ : InMux
    port map (
            O => \N__9640\,
            I => \N__9596\
        );

    \I__1931\ : Span4Mux_v
    port map (
            O => \N__9637\,
            I => \N__9593\
        );

    \I__1930\ : InMux
    port map (
            O => \N__9636\,
            I => \N__9588\
        );

    \I__1929\ : InMux
    port map (
            O => \N__9635\,
            I => \N__9588\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9583\
        );

    \I__1927\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9583\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__9628\,
            I => \N__9576\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__9625\,
            I => \N__9576\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9618\,
            I => \N__9576\
        );

    \I__1923\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9573\
        );

    \I__1922\ : Span4Mux_v
    port map (
            O => \N__9614\,
            I => \N__9562\
        );

    \I__1921\ : Span4Mux_v
    port map (
            O => \N__9609\,
            I => \N__9562\
        );

    \I__1920\ : Span4Mux_h
    port map (
            O => \N__9606\,
            I => \N__9562\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__9603\,
            I => \N__9562\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__9596\,
            I => \N__9559\
        );

    \I__1917\ : Span4Mux_h
    port map (
            O => \N__9593\,
            I => \N__9555\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__9588\,
            I => \N__9552\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__9583\,
            I => \N__9549\
        );

    \I__1914\ : Span4Mux_v
    port map (
            O => \N__9576\,
            I => \N__9546\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__9573\,
            I => \N__9543\
        );

    \I__1912\ : InMux
    port map (
            O => \N__9572\,
            I => \N__9538\
        );

    \I__1911\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9538\
        );

    \I__1910\ : Span4Mux_h
    port map (
            O => \N__9562\,
            I => \N__9533\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__9559\,
            I => \N__9533\
        );

    \I__1908\ : InMux
    port map (
            O => \N__9558\,
            I => \N__9530\
        );

    \I__1907\ : Span4Mux_h
    port map (
            O => \N__9555\,
            I => \N__9523\
        );

    \I__1906\ : Span4Mux_v
    port map (
            O => \N__9552\,
            I => \N__9523\
        );

    \I__1905\ : Span4Mux_v
    port map (
            O => \N__9549\,
            I => \N__9523\
        );

    \I__1904\ : Span4Mux_h
    port map (
            O => \N__9546\,
            I => \N__9518\
        );

    \I__1903\ : Span4Mux_v
    port map (
            O => \N__9543\,
            I => \N__9518\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__9538\,
            I => \N__9515\
        );

    \I__1901\ : Span4Mux_h
    port map (
            O => \N__9533\,
            I => \N__9510\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__9530\,
            I => \N__9510\
        );

    \I__1899\ : Odrv4
    port map (
            O => \N__9523\,
            I => reset_all_w
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__9518\,
            I => reset_all_w
        );

    \I__1897\ : Odrv12
    port map (
            O => \N__9515\,
            I => reset_all_w
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__9510\,
            I => reset_all_w
        );

    \I__1895\ : InMux
    port map (
            O => \N__9501\,
            I => \N__9495\
        );

    \I__1894\ : InMux
    port map (
            O => \N__9500\,
            I => \N__9495\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__9495\,
            I => rx_shift_reg_6
        );

    \I__1892\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9489\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__9489\,
            I => \N__9483\
        );

    \I__1890\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9478\
        );

    \I__1889\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9478\
        );

    \I__1888\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9475\
        );

    \I__1887\ : Span4Mux_v
    port map (
            O => \N__9483\,
            I => \N__9472\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__9478\,
            I => \N__9467\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__9475\,
            I => \N__9467\
        );

    \I__1884\ : Span4Mux_h
    port map (
            O => \N__9472\,
            I => \N__9463\
        );

    \I__1883\ : Span12Mux_h
    port map (
            O => \N__9467\,
            I => \N__9460\
        );

    \I__1882\ : InMux
    port map (
            O => \N__9466\,
            I => \N__9457\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__9463\,
            I => rx_buf_byte_2
        );

    \I__1880\ : Odrv12
    port map (
            O => \N__9460\,
            I => rx_buf_byte_2
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__9457\,
            I => rx_buf_byte_2
        );

    \I__1878\ : InMux
    port map (
            O => \N__9450\,
            I => \N__9443\
        );

    \I__1877\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9440\
        );

    \I__1876\ : InMux
    port map (
            O => \N__9448\,
            I => \N__9435\
        );

    \I__1875\ : InMux
    port map (
            O => \N__9447\,
            I => \N__9435\
        );

    \I__1874\ : InMux
    port map (
            O => \N__9446\,
            I => \N__9432\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__9443\,
            I => n888
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__9440\,
            I => n888
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__9435\,
            I => n888
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__9432\,
            I => n888
        );

    \I__1869\ : InMux
    port map (
            O => \N__9423\,
            I => \N__9417\
        );

    \I__1868\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9410\
        );

    \I__1867\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9410\
        );

    \I__1866\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9410\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__9417\,
            I => \spi0.n1458\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__9410\,
            I => \spi0.n1458\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__9405\,
            I => \spi0.n13_cascade_\
        );

    \I__1862\ : InMux
    port map (
            O => \N__9402\,
            I => \N__9399\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__9399\,
            I => \spi0.state_next_0\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__9396\,
            I => \N__9393\
        );

    \I__1859\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9390\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__9390\,
            I => \spi0.n499\
        );

    \I__1857\ : InMux
    port map (
            O => \N__9387\,
            I => \N__9384\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__9384\,
            I => \spi0.n498\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__9381\,
            I => \N__9378\
        );

    \I__1854\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9375\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__9375\,
            I => \spi0.n502\
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__9372\,
            I => \N__9367\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__9371\,
            I => \N__9364\
        );

    \I__1850\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9358\
        );

    \I__1849\ : InMux
    port map (
            O => \N__9367\,
            I => \N__9358\
        );

    \I__1848\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9355\
        );

    \I__1847\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9352\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__9358\,
            I => \N__9347\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__9355\,
            I => \N__9347\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__9352\,
            I => \state_next_2__N_308\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__9347\,
            I => \state_next_2__N_308\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__9342\,
            I => \N__9338\
        );

    \I__1841\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9335\
        );

    \I__1840\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9332\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__9335\,
            I => \spi0.n911\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__9332\,
            I => \spi0.n911\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__9327\,
            I => \N__9324\
        );

    \I__1836\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9321\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__9321\,
            I => \spi0.n503\
        );

    \I__1834\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9313\
        );

    \I__1833\ : InMux
    port map (
            O => \N__9317\,
            I => \N__9310\
        );

    \I__1832\ : InMux
    port map (
            O => \N__9316\,
            I => \N__9307\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__9313\,
            I => \spi0.state_next_2__N_306\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__9310\,
            I => \spi0.state_next_2__N_306\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__9307\,
            I => \spi0.state_next_2__N_306\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__9300\,
            I => \N__9292\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__9299\,
            I => \N__9285\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__9298\,
            I => \N__9281\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__9297\,
            I => \N__9277\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__9296\,
            I => \N__9274\
        );

    \I__1823\ : CascadeMux
    port map (
            O => \N__9295\,
            I => \N__9271\
        );

    \I__1822\ : InMux
    port map (
            O => \N__9292\,
            I => \N__9263\
        );

    \I__1821\ : InMux
    port map (
            O => \N__9291\,
            I => \N__9263\
        );

    \I__1820\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9252\
        );

    \I__1819\ : InMux
    port map (
            O => \N__9289\,
            I => \N__9252\
        );

    \I__1818\ : InMux
    port map (
            O => \N__9288\,
            I => \N__9252\
        );

    \I__1817\ : InMux
    port map (
            O => \N__9285\,
            I => \N__9252\
        );

    \I__1816\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9252\
        );

    \I__1815\ : InMux
    port map (
            O => \N__9281\,
            I => \N__9247\
        );

    \I__1814\ : InMux
    port map (
            O => \N__9280\,
            I => \N__9247\
        );

    \I__1813\ : InMux
    port map (
            O => \N__9277\,
            I => \N__9234\
        );

    \I__1812\ : InMux
    port map (
            O => \N__9274\,
            I => \N__9234\
        );

    \I__1811\ : InMux
    port map (
            O => \N__9271\,
            I => \N__9234\
        );

    \I__1810\ : InMux
    port map (
            O => \N__9270\,
            I => \N__9234\
        );

    \I__1809\ : InMux
    port map (
            O => \N__9269\,
            I => \N__9234\
        );

    \I__1808\ : InMux
    port map (
            O => \N__9268\,
            I => \N__9234\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__9263\,
            I => \N__9231\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__9252\,
            I => \N__9226\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__9247\,
            I => \N__9226\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__9234\,
            I => \spi0.state_next_1\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__9231\,
            I => \spi0.state_next_1\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__9226\,
            I => \spi0.state_next_1\
        );

    \I__1801\ : InMux
    port map (
            O => \N__9219\,
            I => \N__9194\
        );

    \I__1800\ : InMux
    port map (
            O => \N__9218\,
            I => \N__9194\
        );

    \I__1799\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9194\
        );

    \I__1798\ : InMux
    port map (
            O => \N__9216\,
            I => \N__9194\
        );

    \I__1797\ : InMux
    port map (
            O => \N__9215\,
            I => \N__9194\
        );

    \I__1796\ : InMux
    port map (
            O => \N__9214\,
            I => \N__9189\
        );

    \I__1795\ : InMux
    port map (
            O => \N__9213\,
            I => \N__9189\
        );

    \I__1794\ : InMux
    port map (
            O => \N__9212\,
            I => \N__9174\
        );

    \I__1793\ : InMux
    port map (
            O => \N__9211\,
            I => \N__9174\
        );

    \I__1792\ : InMux
    port map (
            O => \N__9210\,
            I => \N__9174\
        );

    \I__1791\ : InMux
    port map (
            O => \N__9209\,
            I => \N__9174\
        );

    \I__1790\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9174\
        );

    \I__1789\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9174\
        );

    \I__1788\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9174\
        );

    \I__1787\ : InMux
    port map (
            O => \N__9205\,
            I => \N__9171\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__9194\,
            I => \spi0.n4\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__9189\,
            I => \spi0.n4\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__9174\,
            I => \spi0.n4\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__9171\,
            I => \spi0.n4\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__9162\,
            I => \N__9159\
        );

    \I__1781\ : InMux
    port map (
            O => \N__9159\,
            I => \N__9156\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__9156\,
            I => \spi0.n504\
        );

    \I__1779\ : InMux
    port map (
            O => \N__9153\,
            I => \N__9150\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__9150\,
            I => \pc_rx.n1\
        );

    \I__1777\ : InMux
    port map (
            O => \N__9147\,
            I => \N__9143\
        );

    \I__1776\ : InMux
    port map (
            O => \N__9146\,
            I => \N__9140\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__9143\,
            I => \N__9133\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__9140\,
            I => \N__9133\
        );

    \I__1773\ : InMux
    port map (
            O => \N__9139\,
            I => \N__9128\
        );

    \I__1772\ : InMux
    port map (
            O => \N__9138\,
            I => \N__9128\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__9133\,
            I => \pc_rx.r_SM_Main_2_N_110_0\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__9128\,
            I => \pc_rx.r_SM_Main_2_N_110_0\
        );

    \I__1769\ : CascadeMux
    port map (
            O => \N__9123\,
            I => \N__9120\
        );

    \I__1768\ : InMux
    port map (
            O => \N__9120\,
            I => \N__9117\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__9117\,
            I => \pc_rx.n4\
        );

    \I__1766\ : InMux
    port map (
            O => \N__9114\,
            I => \N__9110\
        );

    \I__1765\ : InMux
    port map (
            O => \N__9113\,
            I => \N__9107\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__9110\,
            I => \N__9101\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__9107\,
            I => \N__9098\
        );

    \I__1762\ : InMux
    port map (
            O => \N__9106\,
            I => \N__9095\
        );

    \I__1761\ : InMux
    port map (
            O => \N__9105\,
            I => \N__9092\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__9104\,
            I => \N__9088\
        );

    \I__1759\ : Span4Mux_h
    port map (
            O => \N__9101\,
            I => \N__9082\
        );

    \I__1758\ : Span4Mux_v
    port map (
            O => \N__9098\,
            I => \N__9082\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__9095\,
            I => \N__9077\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__9092\,
            I => \N__9077\
        );

    \I__1755\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9074\
        );

    \I__1754\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9069\
        );

    \I__1753\ : InMux
    port map (
            O => \N__9087\,
            I => \N__9069\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__9082\,
            I => fifo_read_cmd
        );

    \I__1751\ : Odrv4
    port map (
            O => \N__9077\,
            I => fifo_read_cmd
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__9074\,
            I => fifo_read_cmd
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__9069\,
            I => fifo_read_cmd
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__9060\,
            I => \N__9056\
        );

    \I__1747\ : InMux
    port map (
            O => \N__9059\,
            I => \N__9053\
        );

    \I__1746\ : InMux
    port map (
            O => \N__9056\,
            I => \N__9050\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__9053\,
            I => \N__9046\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__9050\,
            I => \N__9043\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__9049\,
            I => \N__9039\
        );

    \I__1742\ : Span4Mux_h
    port map (
            O => \N__9046\,
            I => \N__9032\
        );

    \I__1741\ : Span4Mux_h
    port map (
            O => \N__9043\,
            I => \N__9029\
        );

    \I__1740\ : InMux
    port map (
            O => \N__9042\,
            I => \N__9024\
        );

    \I__1739\ : InMux
    port map (
            O => \N__9039\,
            I => \N__9024\
        );

    \I__1738\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9019\
        );

    \I__1737\ : InMux
    port map (
            O => \N__9037\,
            I => \N__9019\
        );

    \I__1736\ : InMux
    port map (
            O => \N__9036\,
            I => \N__9014\
        );

    \I__1735\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9014\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__9032\,
            I => is_fifo_empty_flag
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__9029\,
            I => is_fifo_empty_flag
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__9024\,
            I => is_fifo_empty_flag
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__9019\,
            I => is_fifo_empty_flag
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__9014\,
            I => is_fifo_empty_flag
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__9003\,
            I => \N__8997\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__9002\,
            I => \N__8994\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__9001\,
            I => \N__8987\
        );

    \I__1726\ : InMux
    port map (
            O => \N__9000\,
            I => \N__8981\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8981\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8978\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8974\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__8992\,
            I => \N__8971\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8967\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8964\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8987\,
            I => \N__8961\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8958\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8981\,
            I => \N__8955\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__8978\,
            I => \N__8952\
        );

    \I__1715\ : CascadeMux
    port map (
            O => \N__8977\,
            I => \N__8948\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8974\,
            I => \N__8944\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8939\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8939\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8967\,
            I => \N__8929\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8964\,
            I => \N__8929\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__8961\,
            I => \N__8929\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__8958\,
            I => \N__8929\
        );

    \I__1707\ : Span4Mux_h
    port map (
            O => \N__8955\,
            I => \N__8924\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__8952\,
            I => \N__8924\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8917\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8948\,
            I => \N__8917\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8917\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__8944\,
            I => \N__8914\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8939\,
            I => \N__8911\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__8938\,
            I => \N__8908\
        );

    \I__1699\ : Span12Mux_h
    port map (
            O => \N__8929\,
            I => \N__8905\
        );

    \I__1698\ : Sp12to4
    port map (
            O => \N__8924\,
            I => \N__8900\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8917\,
            I => \N__8900\
        );

    \I__1696\ : Span4Mux_h
    port map (
            O => \N__8914\,
            I => \N__8895\
        );

    \I__1695\ : Span4Mux_v
    port map (
            O => \N__8911\,
            I => \N__8895\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8892\
        );

    \I__1693\ : Odrv12
    port map (
            O => \N__8905\,
            I => rd_addr_r_0
        );

    \I__1692\ : Odrv12
    port map (
            O => \N__8900\,
            I => rd_addr_r_0
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__8895\,
            I => rd_addr_r_0
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__8892\,
            I => rd_addr_r_0
        );

    \I__1689\ : SRMux
    port map (
            O => \N__8883\,
            I => \N__8880\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8880\,
            I => \N__8877\
        );

    \I__1687\ : Span4Mux_h
    port map (
            O => \N__8877\,
            I => \N__8874\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__8874\,
            I => \spi0.n895\
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__8871\,
            I => \n888_cascade_\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__8868\,
            I => \N__8865\
        );

    \I__1683\ : InMux
    port map (
            O => \N__8865\,
            I => \N__8862\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__8862\,
            I => \spi0.n507\
        );

    \I__1681\ : InMux
    port map (
            O => \N__8859\,
            I => \N__8853\
        );

    \I__1680\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8853\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8853\,
            I => \spi0.state_next_2__N_307\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__8850\,
            I => \spi0.n3476_cascade_\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8844\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__8844\,
            I => \spi0.n25\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8838\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8838\,
            I => \spi0.n13\
        );

    \I__1673\ : CascadeMux
    port map (
            O => \N__8835\,
            I => \rx_shift_reg_15__N_315_cascade_\
        );

    \I__1672\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8828\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__8831\,
            I => \N__8825\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8828\,
            I => \N__8821\
        );

    \I__1669\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8818\
        );

    \I__1668\ : InMux
    port map (
            O => \N__8824\,
            I => \N__8815\
        );

    \I__1667\ : Span4Mux_v
    port map (
            O => \N__8821\,
            I => \N__8809\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__8818\,
            I => \N__8809\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8815\,
            I => \N__8806\
        );

    \I__1664\ : InMux
    port map (
            O => \N__8814\,
            I => \N__8803\
        );

    \I__1663\ : Span4Mux_h
    port map (
            O => \N__8809\,
            I => \N__8797\
        );

    \I__1662\ : Span4Mux_v
    port map (
            O => \N__8806\,
            I => \N__8797\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__8803\,
            I => \N__8794\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8802\,
            I => \N__8791\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__8797\,
            I => rx_buf_byte_7
        );

    \I__1658\ : Odrv12
    port map (
            O => \N__8794\,
            I => rx_buf_byte_7
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__8791\,
            I => rx_buf_byte_7
        );

    \I__1656\ : InMux
    port map (
            O => \N__8784\,
            I => \N__8781\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__8781\,
            I => rx_shift_reg_8
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__8778\,
            I => \N__8774\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__8777\,
            I => \N__8770\
        );

    \I__1652\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8760\
        );

    \I__1651\ : InMux
    port map (
            O => \N__8773\,
            I => \N__8760\
        );

    \I__1650\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8760\
        );

    \I__1649\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8760\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__8760\,
            I => \N__8756\
        );

    \I__1647\ : InMux
    port map (
            O => \N__8759\,
            I => \N__8753\
        );

    \I__1646\ : Odrv12
    port map (
            O => \N__8756\,
            I => rx_buf_byte_5
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__8753\,
            I => rx_buf_byte_5
        );

    \I__1644\ : InMux
    port map (
            O => \N__8748\,
            I => \N__8742\
        );

    \I__1643\ : InMux
    port map (
            O => \N__8747\,
            I => \N__8742\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__8742\,
            I => rx_shift_reg_7
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__8739\,
            I => \N__8733\
        );

    \I__1640\ : InMux
    port map (
            O => \N__8738\,
            I => \N__8726\
        );

    \I__1639\ : InMux
    port map (
            O => \N__8737\,
            I => \N__8726\
        );

    \I__1638\ : InMux
    port map (
            O => \N__8736\,
            I => \N__8726\
        );

    \I__1637\ : InMux
    port map (
            O => \N__8733\,
            I => \N__8723\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__8726\,
            I => \N__8720\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__8723\,
            I => \N__8717\
        );

    \I__1634\ : Span4Mux_h
    port map (
            O => \N__8720\,
            I => \N__8713\
        );

    \I__1633\ : Span4Mux_v
    port map (
            O => \N__8717\,
            I => \N__8710\
        );

    \I__1632\ : InMux
    port map (
            O => \N__8716\,
            I => \N__8707\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__8713\,
            I => rx_buf_byte_6
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__8710\,
            I => rx_buf_byte_6
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__8707\,
            I => rx_buf_byte_6
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__8700\,
            I => \N__8697\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8689\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8696\,
            I => \N__8689\
        );

    \I__1625\ : InMux
    port map (
            O => \N__8695\,
            I => \N__8686\
        );

    \I__1624\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8683\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8689\,
            I => \N__8677\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__8686\,
            I => \N__8677\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__8683\,
            I => \N__8674\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8682\,
            I => \N__8671\
        );

    \I__1619\ : Odrv12
    port map (
            O => \N__8677\,
            I => rx_buf_byte_4
        );

    \I__1618\ : Odrv4
    port map (
            O => \N__8674\,
            I => rx_buf_byte_4
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__8671\,
            I => rx_buf_byte_4
        );

    \I__1616\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8658\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8658\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__8658\,
            I => \N__8655\
        );

    \I__1613\ : Odrv4
    port map (
            O => \N__8655\,
            I => spi_busy
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__8652\,
            I => \N__8649\
        );

    \I__1611\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8646\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__8646\,
            I => \N__8638\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8631\
        );

    \I__1608\ : InMux
    port map (
            O => \N__8644\,
            I => \N__8631\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8643\,
            I => \N__8631\
        );

    \I__1606\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8626\
        );

    \I__1605\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8626\
        );

    \I__1604\ : Odrv12
    port map (
            O => \N__8638\,
            I => is_tx_fifo_full_flag
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__8631\,
            I => is_tx_fifo_full_flag
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__8626\,
            I => is_tx_fifo_full_flag
        );

    \I__1601\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8615\
        );

    \I__1600\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8612\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__8615\,
            I => \N__8609\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__8612\,
            I => \N__8606\
        );

    \I__1597\ : Span4Mux_h
    port map (
            O => \N__8609\,
            I => \N__8598\
        );

    \I__1596\ : Span4Mux_h
    port map (
            O => \N__8606\,
            I => \N__8598\
        );

    \I__1595\ : InMux
    port map (
            O => \N__8605\,
            I => \N__8595\
        );

    \I__1594\ : InMux
    port map (
            O => \N__8604\,
            I => \N__8590\
        );

    \I__1593\ : InMux
    port map (
            O => \N__8603\,
            I => \N__8590\
        );

    \I__1592\ : Odrv4
    port map (
            O => \N__8598\,
            I => fifo_write_cmd
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__8595\,
            I => fifo_write_cmd
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__8590\,
            I => fifo_write_cmd
        );

    \I__1589\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8577\
        );

    \I__1588\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8577\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__8577\,
            I => \N__8572\
        );

    \I__1586\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8569\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__8575\,
            I => \N__8566\
        );

    \I__1584\ : Span4Mux_h
    port map (
            O => \N__8572\,
            I => \N__8557\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__8569\,
            I => \N__8557\
        );

    \I__1582\ : InMux
    port map (
            O => \N__8566\,
            I => \N__8550\
        );

    \I__1581\ : InMux
    port map (
            O => \N__8565\,
            I => \N__8550\
        );

    \I__1580\ : InMux
    port map (
            O => \N__8564\,
            I => \N__8550\
        );

    \I__1579\ : InMux
    port map (
            O => \N__8563\,
            I => \N__8545\
        );

    \I__1578\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8545\
        );

    \I__1577\ : Sp12to4
    port map (
            O => \N__8557\,
            I => \N__8537\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__8550\,
            I => \N__8537\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__8545\,
            I => \N__8537\
        );

    \I__1574\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8534\
        );

    \I__1573\ : Odrv12
    port map (
            O => \N__8537\,
            I => wr_addr_r_0
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__8534\,
            I => wr_addr_r_0
        );

    \I__1571\ : InMux
    port map (
            O => \N__8529\,
            I => \N__8519\
        );

    \I__1570\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8519\
        );

    \I__1569\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8516\
        );

    \I__1568\ : InMux
    port map (
            O => \N__8526\,
            I => \N__8513\
        );

    \I__1567\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8508\
        );

    \I__1566\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8508\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__8519\,
            I => \r_Bit_Index_0\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__8516\,
            I => \r_Bit_Index_0\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__8513\,
            I => \r_Bit_Index_0\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__8508\,
            I => \r_Bit_Index_0\
        );

    \I__1561\ : CEMux
    port map (
            O => \N__8499\,
            I => \N__8496\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__8496\,
            I => \pc_rx.n3432\
        );

    \I__1559\ : SRMux
    port map (
            O => \N__8493\,
            I => \N__8490\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__8490\,
            I => \N__8487\
        );

    \I__1557\ : Span4Mux_v
    port map (
            O => \N__8487\,
            I => \N__8483\
        );

    \I__1556\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8480\
        );

    \I__1555\ : Odrv4
    port map (
            O => \N__8483\,
            I => n3191
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__8480\,
            I => n3191
        );

    \I__1553\ : SRMux
    port map (
            O => \N__8475\,
            I => \N__8469\
        );

    \I__1552\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8464\
        );

    \I__1551\ : InMux
    port map (
            O => \N__8473\,
            I => \N__8464\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__8472\,
            I => \N__8459\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__8469\,
            I => \N__8455\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__8464\,
            I => \N__8452\
        );

    \I__1547\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8449\
        );

    \I__1546\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8442\
        );

    \I__1545\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8442\
        );

    \I__1544\ : InMux
    port map (
            O => \N__8458\,
            I => \N__8442\
        );

    \I__1543\ : Odrv4
    port map (
            O => \N__8455\,
            I => \r_SM_Main_2\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__8452\,
            I => \r_SM_Main_2\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__8449\,
            I => \r_SM_Main_2\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__8442\,
            I => \r_SM_Main_2\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__8433\,
            I => \N__8426\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__8432\,
            I => \N__8423\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__8431\,
            I => \N__8420\
        );

    \I__1536\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8410\
        );

    \I__1535\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8410\
        );

    \I__1534\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8407\
        );

    \I__1533\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8402\
        );

    \I__1532\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8402\
        );

    \I__1531\ : InMux
    port map (
            O => \N__8419\,
            I => \N__8393\
        );

    \I__1530\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8393\
        );

    \I__1529\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8393\
        );

    \I__1528\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8393\
        );

    \I__1527\ : InMux
    port map (
            O => \N__8415\,
            I => \N__8390\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__8410\,
            I => \r_SM_Main_1\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__8407\,
            I => \r_SM_Main_1\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__8402\,
            I => \r_SM_Main_1\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__8393\,
            I => \r_SM_Main_1\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__8390\,
            I => \r_SM_Main_1\
        );

    \I__1521\ : CascadeMux
    port map (
            O => \N__8379\,
            I => \N__8371\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__8378\,
            I => \N__8368\
        );

    \I__1519\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8363\
        );

    \I__1518\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8356\
        );

    \I__1517\ : InMux
    port map (
            O => \N__8375\,
            I => \N__8356\
        );

    \I__1516\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8356\
        );

    \I__1515\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8351\
        );

    \I__1514\ : InMux
    port map (
            O => \N__8368\,
            I => \N__8351\
        );

    \I__1513\ : InMux
    port map (
            O => \N__8367\,
            I => \N__8346\
        );

    \I__1512\ : InMux
    port map (
            O => \N__8366\,
            I => \N__8346\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__8363\,
            I => \r_SM_Main_0\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__8356\,
            I => \r_SM_Main_0\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__8351\,
            I => \r_SM_Main_0\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__8346\,
            I => \r_SM_Main_0\
        );

    \I__1507\ : InMux
    port map (
            O => \N__8337\,
            I => \N__8331\
        );

    \I__1506\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8331\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__8331\,
            I => n4_adj_495
        );

    \I__1504\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8325\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__8325\,
            I => \N__8321\
        );

    \I__1502\ : InMux
    port map (
            O => \N__8324\,
            I => \N__8318\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__8321\,
            I => n4_adj_494
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__8318\,
            I => n4_adj_494
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__8313\,
            I => \N__8310\
        );

    \I__1498\ : InMux
    port map (
            O => \N__8310\,
            I => \N__8307\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__8307\,
            I => \N__8304\
        );

    \I__1496\ : Span4Mux_h
    port map (
            O => \N__8304\,
            I => \N__8301\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__8301\,
            I => n2527
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__8298\,
            I => \n2527_cascade_\
        );

    \I__1493\ : InMux
    port map (
            O => \N__8295\,
            I => \N__8286\
        );

    \I__1492\ : InMux
    port map (
            O => \N__8294\,
            I => \N__8277\
        );

    \I__1491\ : InMux
    port map (
            O => \N__8293\,
            I => \N__8277\
        );

    \I__1490\ : InMux
    port map (
            O => \N__8292\,
            I => \N__8277\
        );

    \I__1489\ : InMux
    port map (
            O => \N__8291\,
            I => \N__8277\
        );

    \I__1488\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8272\
        );

    \I__1487\ : InMux
    port map (
            O => \N__8289\,
            I => \N__8272\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__8286\,
            I => \pc_rx.r_Bit_Index_1\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__8277\,
            I => \pc_rx.r_Bit_Index_1\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__8272\,
            I => \pc_rx.r_Bit_Index_1\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__8265\,
            I => \N__8262\
        );

    \I__1482\ : InMux
    port map (
            O => \N__8262\,
            I => \N__8259\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__8259\,
            I => \N__8251\
        );

    \I__1480\ : InMux
    port map (
            O => \N__8258\,
            I => \N__8242\
        );

    \I__1479\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8242\
        );

    \I__1478\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8242\
        );

    \I__1477\ : InMux
    port map (
            O => \N__8255\,
            I => \N__8242\
        );

    \I__1476\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8239\
        );

    \I__1475\ : Odrv12
    port map (
            O => \N__8251\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__8242\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__8239\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__1472\ : InMux
    port map (
            O => \N__8232\,
            I => \N__8226\
        );

    \I__1471\ : InMux
    port map (
            O => \N__8231\,
            I => \N__8226\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__8226\,
            I => pc_data_rx_7
        );

    \I__1469\ : InMux
    port map (
            O => \N__8223\,
            I => \N__8220\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__8220\,
            I => \N__8216\
        );

    \I__1467\ : InMux
    port map (
            O => \N__8219\,
            I => \N__8213\
        );

    \I__1466\ : Span4Mux_h
    port map (
            O => \N__8216\,
            I => \N__8207\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__8213\,
            I => \N__8207\
        );

    \I__1464\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8204\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__8207\,
            I => tx_data_byte_7
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__8204\,
            I => tx_data_byte_7
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__8199\,
            I => \pc_rx.r_SM_Main_2_N_107_0_cascade_\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__8196\,
            I => \n1801_cascade_\
        );

    \I__1459\ : CascadeMux
    port map (
            O => \N__8193\,
            I => \N__8189\
        );

    \I__1458\ : InMux
    port map (
            O => \N__8192\,
            I => \N__8186\
        );

    \I__1457\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8183\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__8186\,
            I => n6
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__8183\,
            I => n6
        );

    \I__1454\ : InMux
    port map (
            O => \N__8178\,
            I => \N__8175\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__8175\,
            I => \pc_rx.r_SM_Main_2_N_107_0\
        );

    \I__1452\ : InMux
    port map (
            O => \N__8172\,
            I => \N__8169\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__8169\,
            I => \pc_rx.n2615\
        );

    \I__1450\ : InMux
    port map (
            O => \N__8166\,
            I => \N__8163\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__8163\,
            I => \spi0.n500\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__8160\,
            I => \spi0.n4_cascade_\
        );

    \I__1447\ : InMux
    port map (
            O => \N__8157\,
            I => \N__8154\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__8154\,
            I => \spi0.n492\
        );

    \I__1445\ : CascadeMux
    port map (
            O => \N__8151\,
            I => \spi0.state_next_1_cascade_\
        );

    \I__1444\ : InMux
    port map (
            O => \N__8148\,
            I => \N__8145\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__8145\,
            I => \spi0.n493\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__8142\,
            I => \N__8139\
        );

    \I__1441\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8136\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__8136\,
            I => \spi0.n494\
        );

    \I__1439\ : InMux
    port map (
            O => \N__8133\,
            I => \N__8130\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__8130\,
            I => \spi0.n495\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__8127\,
            I => \N__8124\
        );

    \I__1436\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8121\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__8121\,
            I => \spi0.n496\
        );

    \I__1434\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8115\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__8115\,
            I => \spi0.n497\
        );

    \I__1432\ : InMux
    port map (
            O => \N__8112\,
            I => \N__8109\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__8109\,
            I => \N__8105\
        );

    \I__1430\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8102\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__8105\,
            I => tx_addr_byte_2
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__8102\,
            I => tx_addr_byte_2
        );

    \I__1427\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8094\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__8094\,
            I => tx_shift_reg_9
        );

    \I__1425\ : CascadeMux
    port map (
            O => \N__8091\,
            I => \n3418_cascade_\
        );

    \I__1424\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8085\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__8085\,
            I => tx_shift_reg_10
        );

    \I__1422\ : InMux
    port map (
            O => \N__8082\,
            I => \N__8075\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__8081\,
            I => \N__8067\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__8080\,
            I => \N__8064\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__8079\,
            I => \N__8061\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__8078\,
            I => \N__8058\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__8075\,
            I => \N__8051\
        );

    \I__1416\ : InMux
    port map (
            O => \N__8074\,
            I => \N__8040\
        );

    \I__1415\ : InMux
    port map (
            O => \N__8073\,
            I => \N__8040\
        );

    \I__1414\ : InMux
    port map (
            O => \N__8072\,
            I => \N__8040\
        );

    \I__1413\ : InMux
    port map (
            O => \N__8071\,
            I => \N__8040\
        );

    \I__1412\ : InMux
    port map (
            O => \N__8070\,
            I => \N__8040\
        );

    \I__1411\ : InMux
    port map (
            O => \N__8067\,
            I => \N__8025\
        );

    \I__1410\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8025\
        );

    \I__1409\ : InMux
    port map (
            O => \N__8061\,
            I => \N__8025\
        );

    \I__1408\ : InMux
    port map (
            O => \N__8058\,
            I => \N__8025\
        );

    \I__1407\ : InMux
    port map (
            O => \N__8057\,
            I => \N__8025\
        );

    \I__1406\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8025\
        );

    \I__1405\ : InMux
    port map (
            O => \N__8055\,
            I => \N__8025\
        );

    \I__1404\ : InMux
    port map (
            O => \N__8054\,
            I => \N__8022\
        );

    \I__1403\ : Span4Mux_h
    port map (
            O => \N__8051\,
            I => \N__8019\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__8040\,
            I => n1763
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__8025\,
            I => n1763
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__8022\,
            I => n1763
        );

    \I__1399\ : Odrv4
    port map (
            O => \N__8019\,
            I => n1763
        );

    \I__1398\ : InMux
    port map (
            O => \N__8010\,
            I => \N__8007\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__8007\,
            I => tx_shift_reg_7
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__8004\,
            I => \N__8001\
        );

    \I__1395\ : InMux
    port map (
            O => \N__8001\,
            I => \N__7997\
        );

    \I__1394\ : InMux
    port map (
            O => \N__8000\,
            I => \N__7994\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7997\,
            I => tx_addr_byte_0
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7994\,
            I => tx_addr_byte_0
        );

    \I__1391\ : CascadeMux
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7983\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7983\,
            I => tx_shift_reg_8
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__7980\,
            I => \N__7977\
        );

    \I__1387\ : InMux
    port map (
            O => \N__7977\,
            I => \N__7974\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7974\,
            I => \spi0.n3467\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__7971\,
            I => \spi0.n3467_cascade_\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__7968\,
            I => \spi0.state_next_2_cascade_\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__7965\,
            I => \N__7961\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7958\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7955\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7958\,
            I => pc_data_rx_2
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__7955\,
            I => pc_data_rx_2
        );

    \I__1378\ : InMux
    port map (
            O => \N__7950\,
            I => \N__7947\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7947\,
            I => \N__7943\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7940\
        );

    \I__1375\ : Span4Mux_v
    port map (
            O => \N__7943\,
            I => \N__7934\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7940\,
            I => \N__7934\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7931\
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__7934\,
            I => tx_data_byte_2
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7931\,
            I => tx_data_byte_2
        );

    \I__1370\ : InMux
    port map (
            O => \N__7926\,
            I => \N__7922\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__7925\,
            I => \N__7919\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7922\,
            I => \N__7916\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7913\
        );

    \I__1366\ : Odrv4
    port map (
            O => \N__7916\,
            I => pc_data_rx_5
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__7913\,
            I => pc_data_rx_5
        );

    \I__1364\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7903\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7907\,
            I => \N__7900\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7906\,
            I => \N__7897\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7903\,
            I => tx_data_byte_0
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__7900\,
            I => tx_data_byte_0
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7897\,
            I => tx_data_byte_0
        );

    \I__1358\ : InMux
    port map (
            O => \N__7890\,
            I => \N__7887\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7887\,
            I => \N__7884\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__7884\,
            I => tx_shift_reg_6
        );

    \I__1355\ : CascadeMux
    port map (
            O => \N__7881\,
            I => \n1763_cascade_\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7875\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__7875\,
            I => \N__7872\
        );

    \I__1352\ : Odrv4
    port map (
            O => \N__7872\,
            I => tx_shift_reg_0
        );

    \I__1351\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7866\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__7866\,
            I => tx_shift_reg_1
        );

    \I__1349\ : CascadeMux
    port map (
            O => \N__7863\,
            I => \N__7860\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7860\,
            I => \N__7857\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__7857\,
            I => \N__7853\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7856\,
            I => \N__7850\
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__7853\,
            I => tx_addr_byte_3
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7850\,
            I => tx_addr_byte_3
        );

    \I__1343\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7842\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7842\,
            I => tx_shift_reg_11
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__7839\,
            I => \pc_rx.n6_adj_487_cascade_\
        );

    \I__1340\ : CEMux
    port map (
            O => \N__7836\,
            I => \N__7833\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__7833\,
            I => \N__7829\
        );

    \I__1338\ : CEMux
    port map (
            O => \N__7832\,
            I => \N__7826\
        );

    \I__1337\ : Span4Mux_v
    port map (
            O => \N__7829\,
            I => \N__7823\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7826\,
            I => \N__7820\
        );

    \I__1335\ : Span4Mux_h
    port map (
            O => \N__7823\,
            I => \N__7817\
        );

    \I__1334\ : Sp12to4
    port map (
            O => \N__7820\,
            I => \N__7814\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__7817\,
            I => \pc_rx.n1849\
        );

    \I__1332\ : Odrv12
    port map (
            O => \N__7814\,
            I => \pc_rx.n1849\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__7809\,
            I => \n6_cascade_\
        );

    \I__1330\ : InMux
    port map (
            O => \N__7806\,
            I => \N__7803\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__7803\,
            I => \pc_tx.n1518\
        );

    \I__1328\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7790\
        );

    \I__1327\ : InMux
    port map (
            O => \N__7799\,
            I => \N__7790\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7790\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7797\,
            I => \N__7787\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__7790\,
            I => \N__7784\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__7787\,
            I => \N__7781\
        );

    \I__1322\ : Odrv4
    port map (
            O => \N__7784\,
            I => n1782
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__7781\,
            I => n1782
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__7776\,
            I => \N__7773\
        );

    \I__1319\ : InMux
    port map (
            O => \N__7773\,
            I => \N__7770\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__7770\,
            I => \N__7767\
        );

    \I__1317\ : Sp12to4
    port map (
            O => \N__7767\,
            I => \N__7762\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7766\,
            I => \N__7757\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7765\,
            I => \N__7757\
        );

    \I__1314\ : Odrv12
    port map (
            O => \N__7762\,
            I => tx_data_byte_3
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__7757\,
            I => tx_data_byte_3
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__7752\,
            I => \N__7748\
        );

    \I__1311\ : CascadeMux
    port map (
            O => \N__7751\,
            I => \N__7745\
        );

    \I__1310\ : InMux
    port map (
            O => \N__7748\,
            I => \N__7740\
        );

    \I__1309\ : InMux
    port map (
            O => \N__7745\,
            I => \N__7740\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__7740\,
            I => pc_data_rx_3
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__7737\,
            I => \N__7734\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7734\,
            I => \N__7730\
        );

    \I__1305\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7727\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__7730\,
            I => \N__7721\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__7727\,
            I => \N__7721\
        );

    \I__1302\ : InMux
    port map (
            O => \N__7726\,
            I => \N__7718\
        );

    \I__1301\ : Odrv4
    port map (
            O => \N__7721\,
            I => tx_data_byte_5
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7718\,
            I => tx_data_byte_5
        );

    \I__1299\ : InMux
    port map (
            O => \N__7713\,
            I => \N__7710\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__7710\,
            I => tx_shift_reg_5
        );

    \I__1297\ : InMux
    port map (
            O => \N__7707\,
            I => \N__7704\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__7704\,
            I => tx_shift_reg_3
        );

    \I__1295\ : InMux
    port map (
            O => \N__7701\,
            I => \N__7698\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__7698\,
            I => tx_shift_reg_4
        );

    \I__1293\ : InMux
    port map (
            O => \N__7695\,
            I => \N__7692\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__7692\,
            I => tx_shift_reg_14
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__7689\,
            I => \N__7686\
        );

    \I__1290\ : InMux
    port map (
            O => \N__7686\,
            I => \N__7682\
        );

    \I__1289\ : InMux
    port map (
            O => \N__7685\,
            I => \N__7679\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__7682\,
            I => tx_addr_byte_7
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__7679\,
            I => tx_addr_byte_7
        );

    \I__1286\ : IoInMux
    port map (
            O => \N__7674\,
            I => \N__7671\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__7671\,
            I => \N__7667\
        );

    \I__1284\ : IoInMux
    port map (
            O => \N__7670\,
            I => \N__7664\
        );

    \I__1283\ : Span4Mux_s1_v
    port map (
            O => \N__7667\,
            I => \N__7661\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__7664\,
            I => \N__7658\
        );

    \I__1281\ : Span4Mux_v
    port map (
            O => \N__7661\,
            I => \N__7655\
        );

    \I__1280\ : IoSpan4Mux
    port map (
            O => \N__7658\,
            I => \N__7652\
        );

    \I__1279\ : Sp12to4
    port map (
            O => \N__7655\,
            I => \N__7649\
        );

    \I__1278\ : Span4Mux_s0_v
    port map (
            O => \N__7652\,
            I => \N__7646\
        );

    \I__1277\ : Span12Mux_h
    port map (
            O => \N__7649\,
            I => \N__7643\
        );

    \I__1276\ : Sp12to4
    port map (
            O => \N__7646\,
            I => \N__7640\
        );

    \I__1275\ : Span12Mux_v
    port map (
            O => \N__7643\,
            I => \N__7635\
        );

    \I__1274\ : Span12Mux_v
    port map (
            O => \N__7640\,
            I => \N__7635\
        );

    \I__1273\ : Odrv12
    port map (
            O => \N__7635\,
            I => \DEBUG_8_c\
        );

    \I__1272\ : InMux
    port map (
            O => \N__7632\,
            I => \N__7629\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__7629\,
            I => \N__7625\
        );

    \I__1270\ : InMux
    port map (
            O => \N__7628\,
            I => \N__7622\
        );

    \I__1269\ : Span4Mux_v
    port map (
            O => \N__7625\,
            I => \N__7617\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__7622\,
            I => \N__7617\
        );

    \I__1267\ : Span4Mux_v
    port map (
            O => \N__7617\,
            I => \N__7613\
        );

    \I__1266\ : InMux
    port map (
            O => \N__7616\,
            I => \N__7610\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__7613\,
            I => tx_data_byte_4
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__7610\,
            I => tx_data_byte_4
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__7605\,
            I => \N__7602\
        );

    \I__1262\ : InMux
    port map (
            O => \N__7602\,
            I => \N__7599\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__7599\,
            I => \N__7595\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7598\,
            I => \N__7592\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__7595\,
            I => tx_addr_byte_4
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__7592\,
            I => tx_addr_byte_4
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__7587\,
            I => \pc_rx.n3412_cascade_\
        );

    \I__1256\ : SRMux
    port map (
            O => \N__7584\,
            I => \N__7580\
        );

    \I__1255\ : SRMux
    port map (
            O => \N__7583\,
            I => \N__7577\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__7580\,
            I => \N__7574\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__7577\,
            I => \N__7571\
        );

    \I__1252\ : Span4Mux_v
    port map (
            O => \N__7574\,
            I => \N__7568\
        );

    \I__1251\ : Span4Mux_h
    port map (
            O => \N__7571\,
            I => \N__7565\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__7568\,
            I => \pc_rx.n1946\
        );

    \I__1249\ : Odrv4
    port map (
            O => \N__7565\,
            I => \pc_rx.n1946\
        );

    \I__1248\ : InMux
    port map (
            O => \N__7560\,
            I => \N__7557\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__7557\,
            I => \N__7554\
        );

    \I__1246\ : Span4Mux_v
    port map (
            O => \N__7554\,
            I => \N__7549\
        );

    \I__1245\ : InMux
    port map (
            O => \N__7553\,
            I => \N__7546\
        );

    \I__1244\ : InMux
    port map (
            O => \N__7552\,
            I => \N__7543\
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__7549\,
            I => tx_uart_active_flag
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__7546\,
            I => tx_uart_active_flag
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__7543\,
            I => tx_uart_active_flag
        );

    \I__1240\ : InMux
    port map (
            O => \N__7536\,
            I => \N__7533\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__7533\,
            I => \N__7527\
        );

    \I__1238\ : InMux
    port map (
            O => \N__7532\,
            I => \N__7522\
        );

    \I__1237\ : InMux
    port map (
            O => \N__7531\,
            I => \N__7522\
        );

    \I__1236\ : InMux
    port map (
            O => \N__7530\,
            I => \N__7519\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__7527\,
            I => \r_SM_Main_2_N_183_0\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__7522\,
            I => \r_SM_Main_2_N_183_0\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__7519\,
            I => \r_SM_Main_2_N_183_0\
        );

    \I__1232\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7509\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__7509\,
            I => spi_busy_prev
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__7506\,
            I => \N__7503\
        );

    \I__1229\ : InMux
    port map (
            O => \N__7503\,
            I => \N__7500\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__7500\,
            I => \N__7497\
        );

    \I__1227\ : Span4Mux_v
    port map (
            O => \N__7497\,
            I => \N__7493\
        );

    \I__1226\ : InMux
    port map (
            O => \N__7496\,
            I => \N__7490\
        );

    \I__1225\ : Span4Mux_h
    port map (
            O => \N__7493\,
            I => \N__7484\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__7490\,
            I => \N__7484\
        );

    \I__1223\ : InMux
    port map (
            O => \N__7489\,
            I => \N__7481\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__7484\,
            I => tx_data_byte_6
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__7481\,
            I => tx_data_byte_6
        );

    \I__1220\ : InMux
    port map (
            O => \N__7476\,
            I => \N__7472\
        );

    \I__1219\ : InMux
    port map (
            O => \N__7475\,
            I => \N__7469\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__7472\,
            I => tx_addr_byte_5
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__7469\,
            I => tx_addr_byte_5
        );

    \I__1216\ : InMux
    port map (
            O => \N__7464\,
            I => \N__7461\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__7461\,
            I => tx_shift_reg_12
        );

    \I__1214\ : InMux
    port map (
            O => \N__7458\,
            I => \N__7455\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__7455\,
            I => \N__7452\
        );

    \I__1212\ : Span12Mux_h
    port map (
            O => \N__7452\,
            I => \N__7448\
        );

    \I__1211\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7445\
        );

    \I__1210\ : Odrv12
    port map (
            O => \N__7448\,
            I => tx_addr_byte_6
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__7445\,
            I => tx_addr_byte_6
        );

    \I__1208\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7437\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__7437\,
            I => tx_shift_reg_13
        );

    \I__1206\ : InMux
    port map (
            O => \N__7434\,
            I => \N__7431\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__7431\,
            I => tx_shift_reg_2
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__7428\,
            I => \N__7424\
        );

    \I__1203\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7421\
        );

    \I__1202\ : InMux
    port map (
            O => \N__7424\,
            I => \N__7418\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__7421\,
            I => pc_data_rx_4
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__7418\,
            I => pc_data_rx_4
        );

    \I__1199\ : InMux
    port map (
            O => \N__7413\,
            I => \N__7409\
        );

    \I__1198\ : InMux
    port map (
            O => \N__7412\,
            I => \N__7404\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__7409\,
            I => \N__7401\
        );

    \I__1196\ : InMux
    port map (
            O => \N__7408\,
            I => \N__7396\
        );

    \I__1195\ : InMux
    port map (
            O => \N__7407\,
            I => \N__7396\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__7404\,
            I => \N__7393\
        );

    \I__1193\ : Span4Mux_v
    port map (
            O => \N__7401\,
            I => \N__7386\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__7396\,
            I => \N__7386\
        );

    \I__1191\ : Span4Mux_v
    port map (
            O => \N__7393\,
            I => \N__7382\
        );

    \I__1190\ : InMux
    port map (
            O => \N__7392\,
            I => \N__7379\
        );

    \I__1189\ : InMux
    port map (
            O => \N__7391\,
            I => \N__7376\
        );

    \I__1188\ : Span4Mux_h
    port map (
            O => \N__7386\,
            I => \N__7373\
        );

    \I__1187\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7370\
        );

    \I__1186\ : Span4Mux_h
    port map (
            O => \N__7382\,
            I => \N__7366\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__7379\,
            I => \N__7361\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__7376\,
            I => \N__7361\
        );

    \I__1183\ : Span4Mux_v
    port map (
            O => \N__7373\,
            I => \N__7356\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__7370\,
            I => \N__7356\
        );

    \I__1181\ : InMux
    port map (
            O => \N__7369\,
            I => \N__7353\
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__7366\,
            I => n1697
        );

    \I__1179\ : Odrv12
    port map (
            O => \N__7361\,
            I => n1697
        );

    \I__1178\ : Odrv4
    port map (
            O => \N__7356\,
            I => n1697
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__7353\,
            I => n1697
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__7344\,
            I => \n3381_cascade_\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__7341\,
            I => \N__7337\
        );

    \I__1174\ : InMux
    port map (
            O => \N__7340\,
            I => \N__7334\
        );

    \I__1173\ : InMux
    port map (
            O => \N__7337\,
            I => \N__7331\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__7334\,
            I => pc_data_rx_0
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__7331\,
            I => pc_data_rx_0
        );

    \I__1170\ : InMux
    port map (
            O => \N__7326\,
            I => \N__7323\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__7323\,
            I => \N__7319\
        );

    \I__1168\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7316\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__7319\,
            I => pc_data_rx_6
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__7316\,
            I => pc_data_rx_6
        );

    \I__1165\ : InMux
    port map (
            O => \N__7311\,
            I => \N__7308\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__7308\,
            I => spi_busy_falling_edge
        );

    \I__1163\ : InMux
    port map (
            O => \N__7305\,
            I => \N__7300\
        );

    \I__1162\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7297\
        );

    \I__1161\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7294\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__7300\,
            I => \pc_rx.r_Clock_Count_0\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__7297\,
            I => \pc_rx.r_Clock_Count_0\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__7294\,
            I => \pc_rx.r_Clock_Count_0\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__7287\,
            I => \N__7284\
        );

    \I__1156\ : InMux
    port map (
            O => \N__7284\,
            I => \N__7277\
        );

    \I__1155\ : InMux
    port map (
            O => \N__7283\,
            I => \N__7277\
        );

    \I__1154\ : InMux
    port map (
            O => \N__7282\,
            I => \N__7274\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__7277\,
            I => \pc_rx.r_Clock_Count_3\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__7274\,
            I => \pc_rx.r_Clock_Count_3\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__7269\,
            I => \N__7265\
        );

    \I__1150\ : InMux
    port map (
            O => \N__7268\,
            I => \N__7259\
        );

    \I__1149\ : InMux
    port map (
            O => \N__7265\,
            I => \N__7259\
        );

    \I__1148\ : InMux
    port map (
            O => \N__7264\,
            I => \N__7256\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__7259\,
            I => \pc_rx.r_Clock_Count_2\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__7256\,
            I => \pc_rx.r_Clock_Count_2\
        );

    \I__1145\ : InMux
    port map (
            O => \N__7251\,
            I => \N__7246\
        );

    \I__1144\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7243\
        );

    \I__1143\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7240\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__7246\,
            I => \pc_rx.r_Clock_Count_1\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__7243\,
            I => \pc_rx.r_Clock_Count_1\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__7240\,
            I => \pc_rx.r_Clock_Count_1\
        );

    \I__1139\ : InMux
    port map (
            O => \N__7233\,
            I => \N__7226\
        );

    \I__1138\ : InMux
    port map (
            O => \N__7232\,
            I => \N__7226\
        );

    \I__1137\ : InMux
    port map (
            O => \N__7231\,
            I => \N__7223\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__7226\,
            I => \pc_rx.r_Clock_Count_5\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__7223\,
            I => \pc_rx.r_Clock_Count_5\
        );

    \I__1134\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7211\
        );

    \I__1133\ : InMux
    port map (
            O => \N__7217\,
            I => \N__7211\
        );

    \I__1132\ : InMux
    port map (
            O => \N__7216\,
            I => \N__7208\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__7211\,
            I => \pc_rx.r_Clock_Count_6\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__7208\,
            I => \pc_rx.r_Clock_Count_6\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__7203\,
            I => \pc_rx.n3400_cascade_\
        );

    \I__1128\ : InMux
    port map (
            O => \N__7200\,
            I => \N__7193\
        );

    \I__1127\ : InMux
    port map (
            O => \N__7199\,
            I => \N__7193\
        );

    \I__1126\ : InMux
    port map (
            O => \N__7198\,
            I => \N__7190\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__7193\,
            I => \pc_rx.r_Clock_Count_4\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__7190\,
            I => \pc_rx.r_Clock_Count_4\
        );

    \I__1123\ : InMux
    port map (
            O => \N__7185\,
            I => \N__7178\
        );

    \I__1122\ : InMux
    port map (
            O => \N__7184\,
            I => \N__7178\
        );

    \I__1121\ : InMux
    port map (
            O => \N__7183\,
            I => \N__7175\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__7178\,
            I => \pc_rx.r_Clock_Count_8\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__7175\,
            I => \pc_rx.r_Clock_Count_8\
        );

    \I__1118\ : InMux
    port map (
            O => \N__7170\,
            I => \N__7163\
        );

    \I__1117\ : InMux
    port map (
            O => \N__7169\,
            I => \N__7163\
        );

    \I__1116\ : InMux
    port map (
            O => \N__7168\,
            I => \N__7160\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__7163\,
            I => \pc_rx.r_Clock_Count_9\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__7160\,
            I => \pc_rx.r_Clock_Count_9\
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__7155\,
            I => \pc_rx.n2605_cascade_\
        );

    \I__1112\ : InMux
    port map (
            O => \N__7152\,
            I => \N__7145\
        );

    \I__1111\ : InMux
    port map (
            O => \N__7151\,
            I => \N__7145\
        );

    \I__1110\ : InMux
    port map (
            O => \N__7150\,
            I => \N__7142\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__7145\,
            I => \pc_rx.r_Clock_Count_7\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__7142\,
            I => \pc_rx.r_Clock_Count_7\
        );

    \I__1107\ : InMux
    port map (
            O => \N__7137\,
            I => \N__7132\
        );

    \I__1106\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7127\
        );

    \I__1105\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7124\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__7132\,
            I => \N__7121\
        );

    \I__1103\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7116\
        );

    \I__1102\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7116\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__7127\,
            I => \N__7111\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__7124\,
            I => \N__7108\
        );

    \I__1099\ : Span4Mux_h
    port map (
            O => \N__7121\,
            I => \N__7103\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__7116\,
            I => \N__7103\
        );

    \I__1097\ : InMux
    port map (
            O => \N__7115\,
            I => \N__7098\
        );

    \I__1096\ : InMux
    port map (
            O => \N__7114\,
            I => \N__7098\
        );

    \I__1095\ : Span12Mux_v
    port map (
            O => \N__7111\,
            I => \N__7094\
        );

    \I__1094\ : Span4Mux_h
    port map (
            O => \N__7108\,
            I => \N__7091\
        );

    \I__1093\ : Span4Mux_v
    port map (
            O => \N__7103\,
            I => \N__7086\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__7098\,
            I => \N__7086\
        );

    \I__1091\ : InMux
    port map (
            O => \N__7097\,
            I => \N__7083\
        );

    \I__1090\ : Odrv12
    port map (
            O => \N__7094\,
            I => \r_Bit_Index_0_adj_489\
        );

    \I__1089\ : Odrv4
    port map (
            O => \N__7091\,
            I => \r_Bit_Index_0_adj_489\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__7086\,
            I => \r_Bit_Index_0_adj_489\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__7083\,
            I => \r_Bit_Index_0_adj_489\
        );

    \I__1086\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7071\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__7071\,
            I => \N__7068\
        );

    \I__1084\ : Span4Mux_v
    port map (
            O => \N__7068\,
            I => \N__7065\
        );

    \I__1083\ : Odrv4
    port map (
            O => \N__7065\,
            I => \pc_tx.o_Tx_Serial_N_212\
        );

    \I__1082\ : IoInMux
    port map (
            O => \N__7062\,
            I => \N__7059\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__7059\,
            I => \N__7056\
        );

    \I__1080\ : IoSpan4Mux
    port map (
            O => \N__7056\,
            I => \N__7053\
        );

    \I__1079\ : IoSpan4Mux
    port map (
            O => \N__7053\,
            I => \N__7050\
        );

    \I__1078\ : Sp12to4
    port map (
            O => \N__7050\,
            I => \N__7047\
        );

    \I__1077\ : Span12Mux_s7_h
    port map (
            O => \N__7047\,
            I => \N__7044\
        );

    \I__1076\ : Odrv12
    port map (
            O => \N__7044\,
            I => \pc_tx.n3\
        );

    \I__1075\ : CEMux
    port map (
            O => \N__7041\,
            I => \N__7038\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__7038\,
            I => \N__7035\
        );

    \I__1073\ : Sp12to4
    port map (
            O => \N__7035\,
            I => \N__7031\
        );

    \I__1072\ : InMux
    port map (
            O => \N__7034\,
            I => \N__7028\
        );

    \I__1071\ : Odrv12
    port map (
            O => \N__7031\,
            I => n1851
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__7028\,
            I => n1851
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__7023\,
            I => \N__7019\
        );

    \I__1068\ : InMux
    port map (
            O => \N__7022\,
            I => \N__7014\
        );

    \I__1067\ : InMux
    port map (
            O => \N__7019\,
            I => \N__7014\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__7014\,
            I => \N__7011\
        );

    \I__1065\ : Span4Mux_v
    port map (
            O => \N__7011\,
            I => \N__7008\
        );

    \I__1064\ : Odrv4
    port map (
            O => \N__7008\,
            I => \pc_tx.n2597\
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__7005\,
            I => \n1851_cascade_\
        );

    \I__1062\ : SRMux
    port map (
            O => \N__7002\,
            I => \N__6999\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__6999\,
            I => \N__6996\
        );

    \I__1060\ : Sp12to4
    port map (
            O => \N__6996\,
            I => \N__6992\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6989\
        );

    \I__1058\ : Odrv12
    port map (
            O => \N__6992\,
            I => n1934
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6989\,
            I => n1934
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__6984\,
            I => \tx_fifo.lscc_fifo_inst.n4_cascade_\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__6981\,
            I => \N__6978\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6978\,
            I => \N__6974\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6971\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6974\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6971\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__6966\,
            I => \N__6963\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6963\,
            I => \N__6959\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__6962\,
            I => \N__6956\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6959\,
            I => \N__6953\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6956\,
            I => \N__6950\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__6953\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__6950\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__6945\,
            I => \N__6940\
        );

    \I__1042\ : CascadeMux
    port map (
            O => \N__6944\,
            I => \N__6937\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__6943\,
            I => \N__6934\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6930\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6926\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6923\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__6933\,
            I => \N__6920\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6930\,
            I => \N__6916\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6929\,
            I => \N__6913\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6926\,
            I => \N__6908\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6923\,
            I => \N__6908\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6920\,
            I => \N__6905\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__6919\,
            I => \N__6900\
        );

    \I__1030\ : Span4Mux_h
    port map (
            O => \N__6916\,
            I => \N__6888\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6913\,
            I => \N__6888\
        );

    \I__1028\ : Span4Mux_v
    port map (
            O => \N__6908\,
            I => \N__6883\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__6905\,
            I => \N__6883\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6904\,
            I => \N__6876\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6903\,
            I => \N__6876\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6876\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6899\,
            I => \N__6867\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6898\,
            I => \N__6867\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6897\,
            I => \N__6867\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6896\,
            I => \N__6867\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6895\,
            I => \N__6862\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6894\,
            I => \N__6862\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6859\
        );

    \I__1016\ : Odrv4
    port map (
            O => \N__6888\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__1015\ : Odrv4
    port map (
            O => \N__6883\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__6876\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__6867\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6862\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__6859\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__6846\,
            I => \N__6842\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6845\,
            I => \N__6839\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6836\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6839\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6836\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6831\,
            I => \N__6822\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6830\,
            I => \N__6813\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6829\,
            I => \N__6813\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6828\,
            I => \N__6813\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6827\,
            I => \N__6813\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__6826\,
            I => \N__6808\
        );

    \I__999\ : InMux
    port map (
            O => \N__6825\,
            I => \N__6796\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__6822\,
            I => \N__6791\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__6813\,
            I => \N__6791\
        );

    \I__996\ : InMux
    port map (
            O => \N__6812\,
            I => \N__6784\
        );

    \I__995\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6784\
        );

    \I__994\ : InMux
    port map (
            O => \N__6808\,
            I => \N__6784\
        );

    \I__993\ : InMux
    port map (
            O => \N__6807\,
            I => \N__6759\
        );

    \I__992\ : InMux
    port map (
            O => \N__6806\,
            I => \N__6759\
        );

    \I__991\ : InMux
    port map (
            O => \N__6805\,
            I => \N__6752\
        );

    \I__990\ : InMux
    port map (
            O => \N__6804\,
            I => \N__6752\
        );

    \I__989\ : InMux
    port map (
            O => \N__6803\,
            I => \N__6752\
        );

    \I__988\ : InMux
    port map (
            O => \N__6802\,
            I => \N__6743\
        );

    \I__987\ : InMux
    port map (
            O => \N__6801\,
            I => \N__6743\
        );

    \I__986\ : InMux
    port map (
            O => \N__6800\,
            I => \N__6743\
        );

    \I__985\ : InMux
    port map (
            O => \N__6799\,
            I => \N__6743\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__6796\,
            I => \N__6740\
        );

    \I__983\ : Span4Mux_v
    port map (
            O => \N__6791\,
            I => \N__6735\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__6784\,
            I => \N__6735\
        );

    \I__981\ : InMux
    port map (
            O => \N__6783\,
            I => \N__6720\
        );

    \I__980\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6720\
        );

    \I__979\ : InMux
    port map (
            O => \N__6781\,
            I => \N__6720\
        );

    \I__978\ : InMux
    port map (
            O => \N__6780\,
            I => \N__6720\
        );

    \I__977\ : InMux
    port map (
            O => \N__6779\,
            I => \N__6720\
        );

    \I__976\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6720\
        );

    \I__975\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6720\
        );

    \I__974\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6709\
        );

    \I__973\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6709\
        );

    \I__972\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6709\
        );

    \I__971\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6709\
        );

    \I__970\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6709\
        );

    \I__969\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6702\
        );

    \I__968\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6702\
        );

    \I__967\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6702\
        );

    \I__966\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6697\
        );

    \I__965\ : InMux
    port map (
            O => \N__6767\,
            I => \N__6697\
        );

    \I__964\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6690\
        );

    \I__963\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6690\
        );

    \I__962\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6690\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__6759\,
            I => wr_addr_r_1
        );

    \I__960\ : LocalMux
    port map (
            O => \N__6752\,
            I => wr_addr_r_1
        );

    \I__959\ : LocalMux
    port map (
            O => \N__6743\,
            I => wr_addr_r_1
        );

    \I__958\ : Odrv4
    port map (
            O => \N__6740\,
            I => wr_addr_r_1
        );

    \I__957\ : Odrv4
    port map (
            O => \N__6735\,
            I => wr_addr_r_1
        );

    \I__956\ : LocalMux
    port map (
            O => \N__6720\,
            I => wr_addr_r_1
        );

    \I__955\ : LocalMux
    port map (
            O => \N__6709\,
            I => wr_addr_r_1
        );

    \I__954\ : LocalMux
    port map (
            O => \N__6702\,
            I => wr_addr_r_1
        );

    \I__953\ : LocalMux
    port map (
            O => \N__6697\,
            I => wr_addr_r_1
        );

    \I__952\ : LocalMux
    port map (
            O => \N__6690\,
            I => wr_addr_r_1
        );

    \I__951\ : InMux
    port map (
            O => \N__6669\,
            I => \N__6656\
        );

    \I__950\ : InMux
    port map (
            O => \N__6668\,
            I => \N__6656\
        );

    \I__949\ : InMux
    port map (
            O => \N__6667\,
            I => \N__6656\
        );

    \I__948\ : InMux
    port map (
            O => \N__6666\,
            I => \N__6653\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__6665\,
            I => \N__6643\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__6664\,
            I => \N__6640\
        );

    \I__945\ : CascadeMux
    port map (
            O => \N__6663\,
            I => \N__6637\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__6656\,
            I => \N__6634\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__6653\,
            I => \N__6631\
        );

    \I__942\ : InMux
    port map (
            O => \N__6652\,
            I => \N__6628\
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__6651\,
            I => \N__6625\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__6650\,
            I => \N__6622\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__6649\,
            I => \N__6619\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__6648\,
            I => \N__6616\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__6647\,
            I => \N__6613\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__6646\,
            I => \N__6610\
        );

    \I__935\ : InMux
    port map (
            O => \N__6643\,
            I => \N__6603\
        );

    \I__934\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6603\
        );

    \I__933\ : InMux
    port map (
            O => \N__6637\,
            I => \N__6603\
        );

    \I__932\ : Span4Mux_v
    port map (
            O => \N__6634\,
            I => \N__6599\
        );

    \I__931\ : Span4Mux_v
    port map (
            O => \N__6631\,
            I => \N__6596\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__6628\,
            I => \N__6593\
        );

    \I__929\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6586\
        );

    \I__928\ : InMux
    port map (
            O => \N__6622\,
            I => \N__6586\
        );

    \I__927\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6586\
        );

    \I__926\ : InMux
    port map (
            O => \N__6616\,
            I => \N__6581\
        );

    \I__925\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6581\
        );

    \I__924\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6578\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__6603\,
            I => \N__6575\
        );

    \I__922\ : InMux
    port map (
            O => \N__6602\,
            I => \N__6572\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__6599\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__920\ : Odrv4
    port map (
            O => \N__6596\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__919\ : Odrv12
    port map (
            O => \N__6593\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__6586\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__6581\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__6578\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__915\ : Odrv4
    port map (
            O => \N__6575\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__6572\,
            I => \tx_fifo.lscc_fifo_inst.n3\
        );

    \I__913\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6551\
        );

    \I__912\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6548\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__6551\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_3\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__6548\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_3\
        );

    \I__909\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6540\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__6540\,
            I => \pc_rx.n6\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__6537\,
            I => \pc_rx.n3399_cascade_\
        );

    \I__906\ : InMux
    port map (
            O => \N__6534\,
            I => \N__6531\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__6531\,
            I => \pc_rx.n3430\
        );

    \I__904\ : InMux
    port map (
            O => \N__6528\,
            I => \N__6525\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__6525\,
            I => \N__6522\
        );

    \I__902\ : Odrv12
    port map (
            O => \N__6522\,
            I => \tx_fifo.lscc_fifo_inst.n3552\
        );

    \I__901\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6516\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__6516\,
            I => \N__6512\
        );

    \I__899\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6509\
        );

    \I__898\ : Odrv4
    port map (
            O => \N__6512\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_4\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__6509\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_4\
        );

    \I__896\ : InMux
    port map (
            O => \N__6504\,
            I => \N__6498\
        );

    \I__895\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6498\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__6498\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__6495\,
            I => \N__6492\
        );

    \I__892\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6489\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__6489\,
            I => \N__6485\
        );

    \I__890\ : InMux
    port map (
            O => \N__6488\,
            I => \N__6482\
        );

    \I__889\ : Odrv4
    port map (
            O => \N__6485\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_0\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__6482\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_0\
        );

    \I__887\ : InMux
    port map (
            O => \N__6477\,
            I => \N__6471\
        );

    \I__886\ : InMux
    port map (
            O => \N__6476\,
            I => \N__6471\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__6471\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_7\
        );

    \I__884\ : CascadeMux
    port map (
            O => \N__6468\,
            I => \tx_fifo.lscc_fifo_inst.n3_cascade_\
        );

    \I__883\ : InMux
    port map (
            O => \N__6465\,
            I => \N__6462\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__6462\,
            I => \N__6459\
        );

    \I__881\ : Span4Mux_v
    port map (
            O => \N__6459\,
            I => \N__6455\
        );

    \I__880\ : InMux
    port map (
            O => \N__6458\,
            I => \N__6452\
        );

    \I__879\ : Odrv4
    port map (
            O => \N__6455\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_2\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__6452\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_2\
        );

    \I__877\ : InMux
    port map (
            O => \N__6447\,
            I => \N__6443\
        );

    \I__876\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6440\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__6443\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_6\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__6440\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_6\
        );

    \I__873\ : InMux
    port map (
            O => \N__6435\,
            I => \pc_rx.n3065\
        );

    \I__872\ : InMux
    port map (
            O => \N__6432\,
            I => \pc_rx.n3066\
        );

    \I__871\ : InMux
    port map (
            O => \N__6429\,
            I => \bfn_14_4_0_\
        );

    \I__870\ : InMux
    port map (
            O => \N__6426\,
            I => \pc_rx.n3068\
        );

    \I__869\ : InMux
    port map (
            O => \N__6423\,
            I => \N__6420\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__6420\,
            I => \N__6416\
        );

    \I__867\ : InMux
    port map (
            O => \N__6419\,
            I => \N__6413\
        );

    \I__866\ : Odrv4
    port map (
            O => \N__6416\,
            I => fifo_temp_output_0
        );

    \I__865\ : LocalMux
    port map (
            O => \N__6413\,
            I => fifo_temp_output_0
        );

    \I__864\ : InMux
    port map (
            O => \N__6408\,
            I => \N__6404\
        );

    \I__863\ : InMux
    port map (
            O => \N__6407\,
            I => \N__6401\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__6404\,
            I => \r_Tx_Data_0\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__6401\,
            I => \r_Tx_Data_0\
        );

    \I__860\ : InMux
    port map (
            O => \N__6396\,
            I => \N__6392\
        );

    \I__859\ : InMux
    port map (
            O => \N__6395\,
            I => \N__6389\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__6392\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_0\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__6389\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_0\
        );

    \I__856\ : InMux
    port map (
            O => \N__6384\,
            I => \N__6381\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__6381\,
            I => \N__6378\
        );

    \I__854\ : Odrv4
    port map (
            O => \N__6378\,
            I => \tx_fifo.lscc_fifo_inst.n3564\
        );

    \I__853\ : CascadeMux
    port map (
            O => \N__6375\,
            I => \N__6368\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__6374\,
            I => \N__6362\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__6373\,
            I => \N__6358\
        );

    \I__850\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6353\
        );

    \I__849\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6353\
        );

    \I__848\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6348\
        );

    \I__847\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6348\
        );

    \I__846\ : InMux
    port map (
            O => \N__6366\,
            I => \N__6345\
        );

    \I__845\ : InMux
    port map (
            O => \N__6365\,
            I => \N__6340\
        );

    \I__844\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6340\
        );

    \I__843\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6336\
        );

    \I__842\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6333\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__6353\,
            I => \N__6330\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__6348\,
            I => \N__6327\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__6345\,
            I => \N__6324\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__6340\,
            I => \N__6321\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__6339\,
            I => \N__6315\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__6336\,
            I => \N__6302\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__6333\,
            I => \N__6302\
        );

    \I__834\ : Span4Mux_v
    port map (
            O => \N__6330\,
            I => \N__6294\
        );

    \I__833\ : Span4Mux_v
    port map (
            O => \N__6327\,
            I => \N__6294\
        );

    \I__832\ : Span4Mux_v
    port map (
            O => \N__6324\,
            I => \N__6294\
        );

    \I__831\ : Span4Mux_h
    port map (
            O => \N__6321\,
            I => \N__6291\
        );

    \I__830\ : InMux
    port map (
            O => \N__6320\,
            I => \N__6288\
        );

    \I__829\ : InMux
    port map (
            O => \N__6319\,
            I => \N__6285\
        );

    \I__828\ : InMux
    port map (
            O => \N__6318\,
            I => \N__6276\
        );

    \I__827\ : InMux
    port map (
            O => \N__6315\,
            I => \N__6276\
        );

    \I__826\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6276\
        );

    \I__825\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6276\
        );

    \I__824\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6273\
        );

    \I__823\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6268\
        );

    \I__822\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6268\
        );

    \I__821\ : InMux
    port map (
            O => \N__6309\,
            I => \N__6261\
        );

    \I__820\ : InMux
    port map (
            O => \N__6308\,
            I => \N__6261\
        );

    \I__819\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6261\
        );

    \I__818\ : Span4Mux_h
    port map (
            O => \N__6302\,
            I => \N__6258\
        );

    \I__817\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6255\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__6294\,
            I => rd_addr_r_1
        );

    \I__815\ : Odrv4
    port map (
            O => \N__6291\,
            I => rd_addr_r_1
        );

    \I__814\ : LocalMux
    port map (
            O => \N__6288\,
            I => rd_addr_r_1
        );

    \I__813\ : LocalMux
    port map (
            O => \N__6285\,
            I => rd_addr_r_1
        );

    \I__812\ : LocalMux
    port map (
            O => \N__6276\,
            I => rd_addr_r_1
        );

    \I__811\ : LocalMux
    port map (
            O => \N__6273\,
            I => rd_addr_r_1
        );

    \I__810\ : LocalMux
    port map (
            O => \N__6268\,
            I => rd_addr_r_1
        );

    \I__809\ : LocalMux
    port map (
            O => \N__6261\,
            I => rd_addr_r_1
        );

    \I__808\ : Odrv4
    port map (
            O => \N__6258\,
            I => rd_addr_r_1
        );

    \I__807\ : LocalMux
    port map (
            O => \N__6255\,
            I => rd_addr_r_1
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__6234\,
            I => \N__6231\
        );

    \I__805\ : InMux
    port map (
            O => \N__6231\,
            I => \N__6228\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__6228\,
            I => \N__6225\
        );

    \I__803\ : Odrv4
    port map (
            O => \N__6225\,
            I => \mem_LUT_data_raw_r_6\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__6222\,
            I => \N__6218\
        );

    \I__801\ : InMux
    port map (
            O => \N__6221\,
            I => \N__6215\
        );

    \I__800\ : InMux
    port map (
            O => \N__6218\,
            I => \N__6212\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__6215\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__6212\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3\
        );

    \I__797\ : InMux
    port map (
            O => \N__6207\,
            I => \N__6204\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__6204\,
            I => \tx_fifo.lscc_fifo_inst.n3540\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__6201\,
            I => \N__6198\
        );

    \I__794\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6194\
        );

    \I__793\ : InMux
    port map (
            O => \N__6197\,
            I => \N__6191\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__6194\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_3\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__6191\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_3\
        );

    \I__790\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6183\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__6183\,
            I => \N__6180\
        );

    \I__788\ : Odrv4
    port map (
            O => \N__6180\,
            I => \mem_LUT_data_raw_r_3\
        );

    \I__787\ : CEMux
    port map (
            O => \N__6177\,
            I => \N__6174\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6170\
        );

    \I__785\ : CEMux
    port map (
            O => \N__6173\,
            I => \N__6167\
        );

    \I__784\ : Span4Mux_v
    port map (
            O => \N__6170\,
            I => \N__6162\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__6167\,
            I => \N__6162\
        );

    \I__782\ : Span4Mux_h
    port map (
            O => \N__6162\,
            I => \N__6156\
        );

    \I__781\ : CEMux
    port map (
            O => \N__6161\,
            I => \N__6153\
        );

    \I__780\ : InMux
    port map (
            O => \N__6160\,
            I => \N__6150\
        );

    \I__779\ : CEMux
    port map (
            O => \N__6159\,
            I => \N__6147\
        );

    \I__778\ : Odrv4
    port map (
            O => \N__6156\,
            I => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__6153\,
            I => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__6150\,
            I => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__6147\,
            I => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w\
        );

    \I__774\ : InMux
    port map (
            O => \N__6138\,
            I => \bfn_14_3_0_\
        );

    \I__773\ : InMux
    port map (
            O => \N__6135\,
            I => \pc_rx.n3060\
        );

    \I__772\ : InMux
    port map (
            O => \N__6132\,
            I => \pc_rx.n3061\
        );

    \I__771\ : InMux
    port map (
            O => \N__6129\,
            I => \pc_rx.n3062\
        );

    \I__770\ : InMux
    port map (
            O => \N__6126\,
            I => \pc_rx.n3063\
        );

    \I__769\ : InMux
    port map (
            O => \N__6123\,
            I => \pc_rx.n3064\
        );

    \I__768\ : InMux
    port map (
            O => \N__6120\,
            I => \N__6117\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__6117\,
            I => n3414
        );

    \I__766\ : InMux
    port map (
            O => \N__6114\,
            I => \N__6111\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__6111\,
            I => n15_adj_498
        );

    \I__764\ : InMux
    port map (
            O => \N__6108\,
            I => \N__6099\
        );

    \I__763\ : InMux
    port map (
            O => \N__6107\,
            I => \N__6099\
        );

    \I__762\ : InMux
    port map (
            O => \N__6106\,
            I => \N__6099\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__6099\,
            I => wr_fifo_en_w
        );

    \I__760\ : InMux
    port map (
            O => \N__6096\,
            I => \N__6090\
        );

    \I__759\ : InMux
    port map (
            O => \N__6095\,
            I => \N__6090\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__6090\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6\
        );

    \I__757\ : InMux
    port map (
            O => \N__6087\,
            I => \N__6084\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__6084\,
            I => \tx_fifo.lscc_fifo_inst.n3546\
        );

    \I__755\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6077\
        );

    \I__754\ : InMux
    port map (
            O => \N__6080\,
            I => \N__6074\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__6077\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_6\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__6074\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_6\
        );

    \I__751\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6065\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__6068\,
            I => \N__6062\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__6065\,
            I => \N__6059\
        );

    \I__748\ : InMux
    port map (
            O => \N__6062\,
            I => \N__6056\
        );

    \I__747\ : Odrv4
    port map (
            O => \N__6059\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__6056\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6\
        );

    \I__745\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6047\
        );

    \I__744\ : InMux
    port map (
            O => \N__6050\,
            I => \N__6044\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__6047\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__6044\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5\
        );

    \I__741\ : InMux
    port map (
            O => \N__6039\,
            I => \N__6033\
        );

    \I__740\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6033\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__6033\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_5\
        );

    \I__738\ : InMux
    port map (
            O => \N__6030\,
            I => \N__6024\
        );

    \I__737\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6024\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__6024\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5\
        );

    \I__735\ : InMux
    port map (
            O => \N__6021\,
            I => \N__6018\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__6018\,
            I => \tx_fifo.lscc_fifo_inst.n3558\
        );

    \I__733\ : InMux
    port map (
            O => \N__6015\,
            I => \N__6010\
        );

    \I__732\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6005\
        );

    \I__731\ : InMux
    port map (
            O => \N__6013\,
            I => \N__6005\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__6010\,
            I => \tx_fifo.lscc_fifo_inst.rd_addr_r_2\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__6005\,
            I => \tx_fifo.lscc_fifo_inst.rd_addr_r_2\
        );

    \I__728\ : InMux
    port map (
            O => \N__6000\,
            I => \N__5997\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__5997\,
            I => n1
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__5994\,
            I => \n3110_cascade_\
        );

    \I__725\ : InMux
    port map (
            O => \N__5991\,
            I => \N__5988\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5988\,
            I => wr_addr_p1_w_2
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__5985\,
            I => \wr_addr_p1_w_2_cascade_\
        );

    \I__722\ : InMux
    port map (
            O => \N__5982\,
            I => \N__5977\
        );

    \I__721\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5974\
        );

    \I__720\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5971\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__5977\,
            I => wr_addr_r_2
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5974\,
            I => wr_addr_r_2
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5971\,
            I => wr_addr_r_2
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__5964\,
            I => \N__5961\
        );

    \I__715\ : InMux
    port map (
            O => \N__5961\,
            I => \N__5958\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__5958\,
            I => \tx_fifo.lscc_fifo_inst.n2\
        );

    \I__713\ : CascadeMux
    port map (
            O => \N__5955\,
            I => \N__5951\
        );

    \I__712\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5948\
        );

    \I__711\ : InMux
    port map (
            O => \N__5951\,
            I => \N__5945\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5948\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__5945\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0\
        );

    \I__708\ : InMux
    port map (
            O => \N__5940\,
            I => \N__5930\
        );

    \I__707\ : InMux
    port map (
            O => \N__5939\,
            I => \N__5930\
        );

    \I__706\ : InMux
    port map (
            O => \N__5938\,
            I => \N__5930\
        );

    \I__705\ : InMux
    port map (
            O => \N__5937\,
            I => \N__5927\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5930\,
            I => \pc_tx.r_Bit_Index_2\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5927\,
            I => \pc_tx.r_Bit_Index_2\
        );

    \I__702\ : InMux
    port map (
            O => \N__5922\,
            I => \N__5919\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5919\,
            I => \N__5916\
        );

    \I__700\ : Span12Mux_h
    port map (
            O => \N__5916\,
            I => \N__5913\
        );

    \I__699\ : Odrv12
    port map (
            O => \N__5913\,
            I => \pc_tx.n3456\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__5910\,
            I => \N__5907\
        );

    \I__697\ : InMux
    port map (
            O => \N__5907\,
            I => \N__5904\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5904\,
            I => \N__5901\
        );

    \I__695\ : Span4Mux_h
    port map (
            O => \N__5901\,
            I => \N__5898\
        );

    \I__694\ : Odrv4
    port map (
            O => \N__5898\,
            I => \pc_tx.n3455\
        );

    \I__693\ : InMux
    port map (
            O => \N__5895\,
            I => \N__5889\
        );

    \I__692\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5889\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__5889\,
            I => \N__5884\
        );

    \I__690\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5879\
        );

    \I__689\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5879\
        );

    \I__688\ : Odrv4
    port map (
            O => \N__5884\,
            I => \pc_tx.r_Bit_Index_1\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__5879\,
            I => \pc_tx.r_Bit_Index_1\
        );

    \I__686\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5871\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__5871\,
            I => \N__5868\
        );

    \I__684\ : Odrv4
    port map (
            O => \N__5868\,
            I => \pc_tx.n3522\
        );

    \I__683\ : InMux
    port map (
            O => \N__5865\,
            I => \N__5861\
        );

    \I__682\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5858\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5861\,
            I => \N__5855\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5858\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1\
        );

    \I__679\ : Odrv4
    port map (
            O => \N__5855\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__5850\,
            I => \N__5846\
        );

    \I__677\ : InMux
    port map (
            O => \N__5849\,
            I => \N__5843\
        );

    \I__676\ : InMux
    port map (
            O => \N__5846\,
            I => \N__5840\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5843\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__5840\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__5835\,
            I => \N__5832\
        );

    \I__672\ : InMux
    port map (
            O => \N__5832\,
            I => \N__5828\
        );

    \I__671\ : InMux
    port map (
            O => \N__5831\,
            I => \N__5825\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__5828\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_5\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5825\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_5\
        );

    \I__668\ : InMux
    port map (
            O => \N__5820\,
            I => \N__5816\
        );

    \I__667\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5813\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__5816\,
            I => rd_addr_p1_w_1
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5813\,
            I => rd_addr_p1_w_1
        );

    \I__664\ : InMux
    port map (
            O => \N__5808\,
            I => \N__5804\
        );

    \I__663\ : InMux
    port map (
            O => \N__5807\,
            I => \N__5801\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__5804\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5801\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2\
        );

    \I__660\ : InMux
    port map (
            O => \N__5796\,
            I => \N__5790\
        );

    \I__659\ : InMux
    port map (
            O => \N__5795\,
            I => \N__5790\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__5790\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_1\
        );

    \I__657\ : InMux
    port map (
            O => \N__5787\,
            I => \N__5784\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__5784\,
            I => \N__5781\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__5781\,
            I => \tx_fifo.lscc_fifo_inst.n3528\
        );

    \I__654\ : InMux
    port map (
            O => \N__5778\,
            I => \N__5774\
        );

    \I__653\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5771\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__5774\,
            I => \r_Tx_Data_1\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__5771\,
            I => \r_Tx_Data_1\
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__5766\,
            I => \pc_tx.n3461_cascade_\
        );

    \I__649\ : InMux
    port map (
            O => \N__5763\,
            I => \N__5760\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__5760\,
            I => \N__5757\
        );

    \I__647\ : Odrv4
    port map (
            O => \N__5757\,
            I => \pc_tx.n3462\
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__5754\,
            I => \N__5750\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__5753\,
            I => \N__5747\
        );

    \I__644\ : InMux
    port map (
            O => \N__5750\,
            I => \N__5744\
        );

    \I__643\ : InMux
    port map (
            O => \N__5747\,
            I => \N__5741\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__5744\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_1\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__5741\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_1\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__5736\,
            I => \N__5733\
        );

    \I__639\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5730\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__5730\,
            I => \mem_LUT_data_raw_r_1\
        );

    \I__637\ : InMux
    port map (
            O => \N__5727\,
            I => \N__5724\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__5724\,
            I => \tx_fifo.lscc_fifo_inst.n3570\
        );

    \I__635\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5718\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__5718\,
            I => \N__5715\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__5715\,
            I => \N__5712\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__5712\,
            I => \mem_LUT_data_raw_r_4\
        );

    \I__631\ : CascadeMux
    port map (
            O => \N__5709\,
            I => \N__5706\
        );

    \I__630\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5703\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__5703\,
            I => \N__5700\
        );

    \I__628\ : Span4Mux_h
    port map (
            O => \N__5700\,
            I => \N__5697\
        );

    \I__627\ : Odrv4
    port map (
            O => \N__5697\,
            I => \mem_LUT_data_raw_r_5\
        );

    \I__626\ : CascadeMux
    port map (
            O => \N__5694\,
            I => \rd_addr_p1_w_2_cascade_\
        );

    \I__625\ : InMux
    port map (
            O => \N__5691\,
            I => \N__5688\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__5688\,
            I => n3428
        );

    \I__623\ : InMux
    port map (
            O => \N__5685\,
            I => \N__5682\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__5682\,
            I => rd_addr_p1_w_2
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__5679\,
            I => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w_cascade_\
        );

    \I__620\ : CascadeMux
    port map (
            O => \N__5676\,
            I => \n1_cascade_\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__5673\,
            I => \n32_cascade_\
        );

    \I__618\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5667\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__5667\,
            I => n4_adj_500
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__5664\,
            I => \n24_adj_499_cascade_\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__5661\,
            I => \N__5657\
        );

    \I__614\ : InMux
    port map (
            O => \N__5660\,
            I => \N__5654\
        );

    \I__613\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5651\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__5654\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_2\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__5651\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_2\
        );

    \I__610\ : CascadeMux
    port map (
            O => \N__5646\,
            I => \N__5643\
        );

    \I__609\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5639\
        );

    \I__608\ : InMux
    port map (
            O => \N__5642\,
            I => \N__5636\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__5639\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__5636\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2\
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__5631\,
            I => \tx_fifo.lscc_fifo_inst.n3534_cascade_\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__5628\,
            I => \N__5625\
        );

    \I__603\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5622\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5622\,
            I => \mem_LUT_data_raw_r_2\
        );

    \I__601\ : InMux
    port map (
            O => \N__5619\,
            I => \N__5611\
        );

    \I__600\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5611\
        );

    \I__599\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5608\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__5616\,
            I => \N__5604\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__5611\,
            I => \N__5600\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__5608\,
            I => \N__5597\
        );

    \I__595\ : InMux
    port map (
            O => \N__5607\,
            I => \N__5592\
        );

    \I__594\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5592\
        );

    \I__593\ : CascadeMux
    port map (
            O => \N__5603\,
            I => \N__5588\
        );

    \I__592\ : Span4Mux_v
    port map (
            O => \N__5600\,
            I => \N__5582\
        );

    \I__591\ : Span4Mux_v
    port map (
            O => \N__5597\,
            I => \N__5582\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__5592\,
            I => \N__5579\
        );

    \I__589\ : InMux
    port map (
            O => \N__5591\,
            I => \N__5574\
        );

    \I__588\ : InMux
    port map (
            O => \N__5588\,
            I => \N__5574\
        );

    \I__587\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5571\
        );

    \I__586\ : Odrv4
    port map (
            O => \N__5582\,
            I => n1827
        );

    \I__585\ : Odrv4
    port map (
            O => \N__5579\,
            I => n1827
        );

    \I__584\ : LocalMux
    port map (
            O => \N__5574\,
            I => n1827
        );

    \I__583\ : LocalMux
    port map (
            O => \N__5571\,
            I => n1827
        );

    \I__582\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5558\
        );

    \I__581\ : InMux
    port map (
            O => \N__5561\,
            I => \N__5555\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__5558\,
            I => fifo_temp_output_1
        );

    \I__579\ : LocalMux
    port map (
            O => \N__5555\,
            I => fifo_temp_output_1
        );

    \I__578\ : CascadeMux
    port map (
            O => \N__5550\,
            I => \N__5547\
        );

    \I__577\ : InMux
    port map (
            O => \N__5547\,
            I => \N__5544\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__5544\,
            I => \N__5541\
        );

    \I__575\ : Odrv4
    port map (
            O => \N__5541\,
            I => \mem_LUT_data_raw_r_0\
        );

    \I__574\ : CascadeMux
    port map (
            O => \N__5538\,
            I => \N__5535\
        );

    \I__573\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5531\
        );

    \I__572\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5528\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__5531\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_7\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__5528\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_7\
        );

    \I__569\ : CascadeMux
    port map (
            O => \N__5523\,
            I => \N__5520\
        );

    \I__568\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5514\
        );

    \I__567\ : InMux
    port map (
            O => \N__5519\,
            I => \N__5514\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__5514\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4\
        );

    \I__565\ : InMux
    port map (
            O => \N__5511\,
            I => \N__5505\
        );

    \I__564\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5505\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__5505\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_4\
        );

    \I__562\ : InMux
    port map (
            O => \N__5502\,
            I => \N__5499\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__5499\,
            I => \N__5495\
        );

    \I__560\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5492\
        );

    \I__559\ : Odrv12
    port map (
            O => \N__5495\,
            I => fifo_temp_output_2
        );

    \I__558\ : LocalMux
    port map (
            O => \N__5492\,
            I => fifo_temp_output_2
        );

    \I__557\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5483\
        );

    \I__556\ : InMux
    port map (
            O => \N__5486\,
            I => \N__5480\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__5483\,
            I => fifo_temp_output_4
        );

    \I__554\ : LocalMux
    port map (
            O => \N__5480\,
            I => fifo_temp_output_4
        );

    \I__553\ : InMux
    port map (
            O => \N__5475\,
            I => \N__5471\
        );

    \I__552\ : InMux
    port map (
            O => \N__5474\,
            I => \N__5468\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__5471\,
            I => \r_Tx_Data_4\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__5468\,
            I => \r_Tx_Data_4\
        );

    \I__549\ : InMux
    port map (
            O => \N__5463\,
            I => \N__5460\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__5460\,
            I => \N__5456\
        );

    \I__547\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5453\
        );

    \I__546\ : Odrv12
    port map (
            O => \N__5456\,
            I => fifo_temp_output_3
        );

    \I__545\ : LocalMux
    port map (
            O => \N__5453\,
            I => fifo_temp_output_3
        );

    \I__544\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5444\
        );

    \I__543\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5441\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__5444\,
            I => fifo_temp_output_7
        );

    \I__541\ : LocalMux
    port map (
            O => \N__5441\,
            I => fifo_temp_output_7
        );

    \I__540\ : InMux
    port map (
            O => \N__5436\,
            I => \N__5432\
        );

    \I__539\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5429\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__5432\,
            I => fifo_temp_output_6
        );

    \I__537\ : LocalMux
    port map (
            O => \N__5429\,
            I => fifo_temp_output_6
        );

    \I__536\ : InMux
    port map (
            O => \N__5424\,
            I => \N__5420\
        );

    \I__535\ : InMux
    port map (
            O => \N__5423\,
            I => \N__5417\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__5420\,
            I => \r_Tx_Data_7\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__5417\,
            I => \r_Tx_Data_7\
        );

    \I__532\ : InMux
    port map (
            O => \N__5412\,
            I => \N__5406\
        );

    \I__531\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5406\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__5406\,
            I => \r_Tx_Data_6\
        );

    \I__529\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5399\
        );

    \I__528\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5396\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__5399\,
            I => \r_Tx_Data_3\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__5396\,
            I => \r_Tx_Data_3\
        );

    \I__525\ : InMux
    port map (
            O => \N__5391\,
            I => \N__5385\
        );

    \I__524\ : InMux
    port map (
            O => \N__5390\,
            I => \N__5385\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__5385\,
            I => \r_Tx_Data_2\
        );

    \I__522\ : InMux
    port map (
            O => \N__5382\,
            I => \N__5378\
        );

    \I__521\ : InMux
    port map (
            O => \N__5381\,
            I => \N__5375\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__5378\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__5375\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7\
        );

    \I__518\ : InMux
    port map (
            O => \N__5370\,
            I => \N__5362\
        );

    \I__517\ : InMux
    port map (
            O => \N__5369\,
            I => \N__5351\
        );

    \I__516\ : InMux
    port map (
            O => \N__5368\,
            I => \N__5351\
        );

    \I__515\ : InMux
    port map (
            O => \N__5367\,
            I => \N__5351\
        );

    \I__514\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5351\
        );

    \I__513\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5351\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__5362\,
            I => reset_clk_counter_0
        );

    \I__511\ : LocalMux
    port map (
            O => \N__5351\,
            I => reset_clk_counter_0
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__5346\,
            I => \N__5341\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__5345\,
            I => \N__5336\
        );

    \I__508\ : InMux
    port map (
            O => \N__5344\,
            I => \N__5333\
        );

    \I__507\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5328\
        );

    \I__506\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5328\
        );

    \I__505\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5323\
        );

    \I__504\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5323\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__5333\,
            I => reset_clk_counter_1
        );

    \I__502\ : LocalMux
    port map (
            O => \N__5328\,
            I => reset_clk_counter_1
        );

    \I__501\ : LocalMux
    port map (
            O => \N__5323\,
            I => reset_clk_counter_1
        );

    \I__500\ : InMux
    port map (
            O => \N__5316\,
            I => \N__5307\
        );

    \I__499\ : InMux
    port map (
            O => \N__5315\,
            I => \N__5307\
        );

    \I__498\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5307\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__5307\,
            I => \reset_all_w_N_61\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__5304\,
            I => \N__5301\
        );

    \I__495\ : InMux
    port map (
            O => \N__5301\,
            I => \N__5295\
        );

    \I__494\ : InMux
    port map (
            O => \N__5300\,
            I => \N__5288\
        );

    \I__493\ : InMux
    port map (
            O => \N__5299\,
            I => \N__5288\
        );

    \I__492\ : InMux
    port map (
            O => \N__5298\,
            I => \N__5288\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__5295\,
            I => reset_clk_counter_2
        );

    \I__490\ : LocalMux
    port map (
            O => \N__5288\,
            I => reset_clk_counter_2
        );

    \I__489\ : InMux
    port map (
            O => \N__5283\,
            I => \N__5277\
        );

    \I__488\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5277\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__5277\,
            I => fifo_temp_output_5
        );

    \I__486\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5271\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__5271\,
            I => \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r\
        );

    \I__484\ : CascadeMux
    port map (
            O => \N__5268\,
            I => \N__5265\
        );

    \I__483\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5262\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__5262\,
            I => \N__5259\
        );

    \I__481\ : Odrv12
    port map (
            O => \N__5259\,
            I => \mem_LUT_data_raw_r_7\
        );

    \I__480\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5253\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__5253\,
            I => \N__5249\
        );

    \I__478\ : InMux
    port map (
            O => \N__5252\,
            I => \N__5246\
        );

    \I__477\ : Odrv4
    port map (
            O => \N__5249\,
            I => \r_Tx_Data_5\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__5246\,
            I => \r_Tx_Data_5\
        );

    \I__475\ : IoInMux
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__5238\,
            I => \N__5235\
        );

    \I__473\ : IoSpan4Mux
    port map (
            O => \N__5235\,
            I => \N__5232\
        );

    \I__472\ : Span4Mux_s2_v
    port map (
            O => \N__5232\,
            I => \N__5229\
        );

    \I__471\ : Span4Mux_v
    port map (
            O => \N__5229\,
            I => \N__5226\
        );

    \I__470\ : Sp12to4
    port map (
            O => \N__5226\,
            I => \N__5223\
        );

    \I__469\ : Odrv12
    port map (
            O => \N__5223\,
            I => \RESET_c\
        );

    \I__468\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5217\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__5217\,
            I => \N__5214\
        );

    \I__466\ : Glb2LocalMux
    port map (
            O => \N__5214\,
            I => \N__5211\
        );

    \I__465\ : GlobalMux
    port map (
            O => \N__5211\,
            I => pll_clk_unbuf
        );

    \I__464\ : IoInMux
    port map (
            O => \N__5208\,
            I => \N__5205\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__5205\,
            I => \N__5202\
        );

    \I__462\ : IoSpan4Mux
    port map (
            O => \N__5202\,
            I => \N__5199\
        );

    \I__461\ : Span4Mux_s3_h
    port map (
            O => \N__5199\,
            I => \N__5196\
        );

    \I__460\ : Span4Mux_h
    port map (
            O => \N__5196\,
            I => \N__5193\
        );

    \I__459\ : Span4Mux_v
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__458\ : Odrv4
    port map (
            O => \N__5190\,
            I => \GB_BUFFER_pll_clk_unbuf_THRU_CO\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__5187\,
            I => \reset_all_w_N_61_cascade_\
        );

    \I__456\ : CascadeMux
    port map (
            O => \N__5184\,
            I => \n2_adj_493_cascade_\
        );

    \I__455\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5176\
        );

    \I__454\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5171\
        );

    \I__453\ : InMux
    port map (
            O => \N__5179\,
            I => \N__5171\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__5176\,
            I => reset_clk_counter_3
        );

    \I__451\ : LocalMux
    port map (
            O => \N__5171\,
            I => reset_clk_counter_3
        );

    \I__450\ : IoInMux
    port map (
            O => \N__5166\,
            I => \N__5163\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__5163\,
            I => \N__5160\
        );

    \I__448\ : Span4Mux_s3_v
    port map (
            O => \N__5160\,
            I => \N__5157\
        );

    \I__447\ : Sp12to4
    port map (
            O => \N__5157\,
            I => \N__5154\
        );

    \I__446\ : Span12Mux_h
    port map (
            O => \N__5154\,
            I => \N__5151\
        );

    \I__445\ : Span12Mux_v
    port map (
            O => \N__5151\,
            I => \N__5148\
        );

    \I__444\ : Odrv12
    port map (
            O => \N__5148\,
            I => \ICE_SYSCLK_c\
        );

    \INVspi0.tx_shift_reg_i7C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i7C_net\,
            I => \N__11351\
        );

    \INVspi0.tx_shift_reg_i0C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i0C_net\,
            I => \N__11338\
        );

    \INVspi0.tx_shift_reg_i15C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i15C_net\,
            I => \N__11333\
        );

    \INVspi0.tx_shift_reg_i6C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i6C_net\,
            I => \N__11352\
        );

    \IN_MUX_bfv_19_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_10_0_\
        );

    \IN_MUX_bfv_19_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_7_0_\
        );

    \IN_MUX_bfv_19_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pc_tx.n3076\,
            carryinitout => \bfn_19_8_0_\
        );

    \IN_MUX_bfv_14_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_3_0_\
        );

    \IN_MUX_bfv_14_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pc_rx.n3067\,
            carryinitout => \bfn_14_4_0_\
        );

    \IN_MUX_bfv_24_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_8_0_\
        );

    \IN_MUX_bfv_24_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n3085,
            carryinitout => \bfn_24_9_0_\
        );

    \IN_MUX_bfv_24_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n3093,
            carryinitout => \bfn_24_10_0_\
        );

    \IN_MUX_bfv_24_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n3101,
            carryinitout => \bfn_24_11_0_\
        );

    \clk_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5208\,
            GLOBALBUFFEROUTPUT => \SLM_CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i1759_1_lut_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9617\,
            lcout => \RESET_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_pll_clk_unbuf_THRU_LUT4_0_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5220\,
            lcout => \GB_BUFFER_pll_clk_unbuf_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_all_r_207_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5181\,
            in1 => \N__5344\,
            in2 => \N__5304\,
            in3 => \N__5370\,
            lcout => reset_all_w,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_clk_counter_i3_584__i1_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__5340\,
            in1 => \N__5368\,
            in2 => \_gnd_net_\,
            in3 => \N__5315\,
            lcout => reset_clk_counter_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5366\,
            in1 => \N__5179\,
            in2 => \N__5345\,
            in3 => \N__5298\,
            lcout => \reset_all_w_N_61\,
            ltout => \reset_all_w_N_61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2690_2_lut_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5187\,
            in3 => \N__5365\,
            lcout => OPEN,
            ltout => \n2_adj_493_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_clk_counter_i3_584__i3_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001001"
        )
    port map (
            in0 => \N__5339\,
            in1 => \N__5180\,
            in2 => \N__5184\,
            in3 => \N__5300\,
            lcout => reset_clk_counter_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_clk_counter_i3_584__i0_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5367\,
            in2 => \_gnd_net_\,
            in3 => \N__5314\,
            lcout => reset_clk_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_clk_counter_i3_584__i2_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100110101010"
        )
    port map (
            in0 => \N__5299\,
            in1 => \N__5369\,
            in2 => \N__5346\,
            in3 => \N__5316\,
            lcout => reset_clk_counter_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i5_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__5617\,
            in1 => \N__9558\,
            in2 => \N__5709\,
            in3 => \N__5283\,
            lcout => fifo_temp_output_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12281\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i5_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5282\,
            in1 => \N__5252\,
            in2 => \_gnd_net_\,
            in3 => \N__7413\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12281\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i3_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5463\,
            in1 => \N__5402\,
            in2 => \_gnd_net_\,
            in3 => \N__7392\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i8_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__6319\,
            in1 => \N__6528\,
            in2 => \N__5538\,
            in3 => \N__5382\,
            lcout => \mem_LUT_data_raw_r_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12286\,
            ce => \N__6173\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r_86_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__9634\,
            in1 => \N__9106\,
            in2 => \_gnd_net_\,
            in3 => \N__9042\,
            lcout => \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12284\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i1_2_lut_3_lut_4_lut_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101110"
        )
    port map (
            in0 => \N__5274\,
            in1 => \N__9633\,
            in2 => \N__9049\,
            in3 => \N__9105\,
            lcout => n1827,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i4_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__5486\,
            in1 => \N__9571\,
            in2 => \N__5603\,
            in3 => \N__5721\,
            lcout => fifo_temp_output_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12283\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i7_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__9572\,
            in1 => \N__5591\,
            in2 => \N__5268\,
            in3 => \N__5447\,
            lcout => fifo_temp_output_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12283\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i3068_3_lut_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7137\,
            in1 => \N__5256\,
            in2 => \_gnd_net_\,
            in3 => \N__5475\,
            lcout => \pc_tx.n3455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i4_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5487\,
            in1 => \N__5474\,
            in2 => \_gnd_net_\,
            in3 => \N__7407\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i6_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__9636\,
            in1 => \N__5607\,
            in2 => \N__6234\,
            in3 => \N__5435\,
            lcout => fifo_temp_output_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i3_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__6186\,
            in1 => \N__9635\,
            in2 => \N__5616\,
            in3 => \N__5459\,
            lcout => fifo_temp_output_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i7_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5423\,
            in1 => \N__7408\,
            in2 => \_gnd_net_\,
            in3 => \N__5448\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i6_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5412\,
            in1 => \N__7412\,
            in2 => \_gnd_net_\,
            in3 => \N__5436\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i3069_3_lut_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5424\,
            in1 => \N__5411\,
            in2 => \_gnd_net_\,
            in3 => \N__7136\,
            lcout => \pc_tx.n3456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i3075_3_lut_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7135\,
            in1 => \N__5403\,
            in2 => \_gnd_net_\,
            in3 => \N__5390\,
            lcout => \pc_tx.n3462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i2_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7391\,
            in1 => \N__5391\,
            in2 => \_gnd_net_\,
            in3 => \N__5502\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i59_60_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__8832\,
            in1 => \N__6831\,
            in2 => \N__6944\,
            in3 => \N__5381\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i155_156_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__6668\,
            in1 => \N__6828\,
            in2 => \N__8831\,
            in3 => \N__5534\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i242_243_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__5519\,
            in1 => \N__6829\,
            in2 => \N__6943\,
            in3 => \N__8696\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i137_138_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__6827\,
            in1 => \N__10359\,
            in2 => \N__5753\,
            in3 => \N__6667\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__5511\,
            in1 => \N__6312\,
            in2 => \N__5523\,
            in3 => \N__8993\,
            lcout => \tx_fifo.lscc_fifo_inst.n3570\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i338_339_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__6830\,
            in1 => \N__6669\,
            in2 => \N__8700\,
            in3 => \N__5510\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i332_333_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__9488\,
            in1 => \N__6652\,
            in2 => \N__5661\,
            in3 => \N__6812\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i2_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__5498\,
            in1 => \N__9661\,
            in2 => \N__5628\,
            in3 => \N__5587\,
            lcout => fifo_temp_output_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__9035\,
            in1 => \N__8582\,
            in2 => \N__9003\,
            in3 => \N__9091\,
            lcout => n4_adj_500,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r__i1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__5820\,
            in1 => \N__6160\,
            in2 => \N__6373\,
            in3 => \N__9662\,
            lcout => rd_addr_r_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i236_237_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__9487\,
            in1 => \N__6811\,
            in2 => \N__6933\,
            in3 => \N__5642\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__8583\,
            in1 => \N__9000\,
            in2 => \N__6826\,
            in3 => \N__6301\,
            lcout => OPEN,
            ltout => \n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__9036\,
            in1 => \_gnd_net_\,
            in2 => \N__5673\,
            in3 => \N__8618\,
            lcout => OPEN,
            ltout => \n24_adj_499_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.empty_r_85_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__5670\,
            in1 => \N__9660\,
            in2 => \N__5664\,
            in3 => \N__5691\,
            lcout => is_fifo_empty_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3151_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__6311\,
            in1 => \N__5660\,
            in2 => \N__5646\,
            in3 => \N__8991\,
            lcout => OPEN,
            ltout => \tx_fifo.lscc_fifo_inst.n3534_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i3_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__5808\,
            in1 => \N__6465\,
            in2 => \N__5631\,
            in3 => \N__6310\,
            lcout => \mem_LUT_data_raw_r_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12285\,
            ce => \N__6161\,
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i1_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5561\,
            in1 => \N__7385\,
            in2 => \_gnd_net_\,
            in3 => \N__5777\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i0_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__6419\,
            in1 => \N__9664\,
            in2 => \N__5550\,
            in3 => \N__5618\,
            lcout => fifo_temp_output_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i1_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__5562\,
            in1 => \N__9665\,
            in2 => \N__5736\,
            in3 => \N__5619\,
            lcout => fifo_temp_output_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i1_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__6384\,
            in1 => \N__5954\,
            in2 => \N__6495\,
            in3 => \N__6313\,
            lcout => \mem_LUT_data_raw_r_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12295\,
            ce => \N__6159\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i2_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__6314\,
            in1 => \N__5787\,
            in2 => \N__5754\,
            in3 => \N__5864\,
            lcout => \mem_LUT_data_raw_r_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12295\,
            ce => \N__6159\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i5_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110110101000"
        )
    port map (
            in0 => \N__5727\,
            in1 => \N__6519\,
            in2 => \N__6339\,
            in3 => \N__5849\,
            lcout => \mem_LUT_data_raw_r_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12295\,
            ce => \N__6159\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i6_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__6318\,
            in1 => \N__6021\,
            in2 => \N__5835\,
            in3 => \N__6051\,
            lcout => \mem_LUT_data_raw_r_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12295\,
            ce => \N__6159\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i781_3_lut_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__6013\,
            in1 => \_gnd_net_\,
            in2 => \N__8977\,
            in3 => \N__6309\,
            lcout => rd_addr_p1_w_2,
            ltout => \rd_addr_p1_w_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3041_4_lut_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__5982\,
            in1 => \N__6768\,
            in2 => \N__5694\,
            in3 => \N__5819\,
            lcout => n3428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_en_i_I_0_2_lut_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9104\,
            in3 => \N__9038\,
            lcout => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w\,
            ltout => \tx_fifo.lscc_fifo_inst.rd_fifo_en_w_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r__i2_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__5685\,
            in1 => \N__6014\,
            in2 => \N__5679\,
            in3 => \N__9663\,
            lcout => \tx_fifo.lscc_fifo_inst.rd_addr_r_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_r_1__I_0_i1_2_lut_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__8951\,
            in1 => \N__8576\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n1,
            ltout => \n1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3028_4_lut_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__6307\,
            in1 => \N__6767\,
            in2 => \N__5676\,
            in3 => \N__9087\,
            lcout => n3414,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_read_cmd_212_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9037\,
            in2 => \_gnd_net_\,
            in3 => \N__7560\,
            lcout => fifo_read_cmd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i774_2_lut_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__6308\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8947\,
            lcout => rd_addr_p1_w_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i329_330_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__6806\,
            in1 => \N__6666\,
            in2 => \N__10374\,
            in3 => \N__5795\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12288\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i44_45_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__5807\,
            in1 => \N__6807\,
            in2 => \N__6945\,
            in3 => \N__9492\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12288\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3146_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__5796\,
            in1 => \N__6320\,
            in2 => \N__6966\,
            in3 => \N__8990\,
            lcout => \tx_fifo.lscc_fifo_inst.n3528\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Bit_Index_i1_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__7114\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5887\,
            lcout => \pc_tx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12304\,
            ce => \N__7041\,
            sr => \N__7002\
        );

    \pc_tx.r_Bit_Index_i2_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__5888\,
            in1 => \N__7115\,
            in2 => \_gnd_net_\,
            in3 => \N__5937\,
            lcout => \pc_tx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12304\,
            ce => \N__7041\,
            sr => \N__7002\
        );

    \pc_tx.i3074_3_lut_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7131\,
            in1 => \N__5778\,
            in2 => \_gnd_net_\,
            in3 => \N__6408\,
            lcout => OPEN,
            ltout => \pc_tx.n3461_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.n3522_bdd_4_lut_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010011000"
        )
    port map (
            in0 => \N__5874\,
            in1 => \N__5939\,
            in2 => \N__5766\,
            in3 => \N__5763\,
            lcout => \pc_tx.o_Tx_Serial_N_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i6_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7326\,
            in1 => \N__11474\,
            in2 => \_gnd_net_\,
            in3 => \N__7489\,
            lcout => tx_data_byte_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2_2_lut_3_lut_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5894\,
            in1 => \N__7130\,
            in2 => \_gnd_net_\,
            in3 => \N__5938\,
            lcout => \pc_tx.n2597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i38_39_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__6825\,
            in1 => \N__6929\,
            in2 => \N__5955\,
            in3 => \N__10296\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Bit_Index_1__bdd_4_lut_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__5940\,
            in1 => \N__5922\,
            in2 => \N__5910\,
            in3 => \N__5895\,
            lcout => \pc_tx.n3522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i41_42_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__6897\,
            in1 => \N__6781\,
            in2 => \N__10366\,
            in3 => \N__5865\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i245_246_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__6778\,
            in1 => \N__6896\,
            in2 => \N__8777\,
            in3 => \N__6029\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i341_342_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__6038\,
            in1 => \N__6780\,
            in2 => \N__6651\,
            in3 => \N__8773\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i50_51_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__6782\,
            in1 => \N__6898\,
            in2 => \N__5850\,
            in3 => \N__8695\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i149_150_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__5831\,
            in1 => \N__6777\,
            in2 => \N__6649\,
            in3 => \N__8769\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i53_54_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__6783\,
            in1 => \N__6899\,
            in2 => \N__8778\,
            in3 => \N__6050\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i326_327_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__10294\,
            in1 => \N__6779\,
            in2 => \N__6650\,
            in3 => \N__6395\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3171_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101011010000"
        )
    port map (
            in0 => \N__6366\,
            in1 => \N__6039\,
            in2 => \N__9002\,
            in3 => \N__6030\,
            lcout => \tx_fifo.lscc_fifo_inst.n3558\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i1_4_lut_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000000"
        )
    port map (
            in0 => \N__5991\,
            in1 => \N__6015\,
            in2 => \N__5964\,
            in3 => \N__6000\,
            lcout => OPEN,
            ltout => \n3110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.full_r_84_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100000"
        )
    port map (
            in0 => \N__6106\,
            in1 => \N__9640\,
            in2 => \N__5994\,
            in3 => \N__6114\,
            lcout => is_tx_fifo_full_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i759_3_lut_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__6764\,
            in1 => \N__5980\,
            in2 => \_gnd_net_\,
            in3 => \N__8564\,
            lcout => wr_addr_p1_w_2,
            ltout => \wr_addr_p1_w_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_r__i2_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__6108\,
            in1 => \N__9642\,
            in2 => \N__5985\,
            in3 => \N__5981\,
            lcout => wr_addr_r_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_p1_w_1__I_0_i2_2_lut_3_lut_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__6765\,
            in1 => \N__8565\,
            in2 => \_gnd_net_\,
            in3 => \N__6361\,
            lcout => \tx_fifo.lscc_fifo_inst.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_en_i_I_0_2_lut_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8642\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8605\,
            lcout => wr_fifo_en_w,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__6120\,
            in1 => \N__8641\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n15_adj_498,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_r__i1_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__6107\,
            in1 => \N__9641\,
            in2 => \N__8575\,
            in3 => \N__6766\,
            lcout => wr_addr_r_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3161_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010110000"
        )
    port map (
            in0 => \N__6447\,
            in1 => \N__6365\,
            in2 => \N__9001\,
            in3 => \N__6096\,
            lcout => \tx_fifo.lscc_fifo_inst.n3546\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3156_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__8986\,
            in1 => \N__6555\,
            in2 => \N__6374\,
            in3 => \N__6845\,
            lcout => \tx_fifo.lscc_fifo_inst.n3540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i248_249_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__8737\,
            in1 => \N__6774\,
            in2 => \N__6919\,
            in3 => \N__6095\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i56_57_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__6776\,
            in1 => \N__6904\,
            in2 => \N__6068\,
            in3 => \N__8738\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i143_144_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__10412\,
            in1 => \N__6772\,
            in2 => \N__6647\,
            in3 => \N__6197\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i47_48_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__6775\,
            in1 => \N__6903\,
            in2 => \N__6222\,
            in3 => \N__10413\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i152_153_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__8736\,
            in1 => \N__6773\,
            in2 => \N__6648\,
            in3 => \N__6080\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i7_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110110101000"
        )
    port map (
            in0 => \N__6087\,
            in1 => \N__6081\,
            in2 => \N__6375\,
            in3 => \N__6069\,
            lcout => \mem_LUT_data_raw_r_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12289\,
            ce => \N__6177\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i4_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__6221\,
            in1 => \N__6207\,
            in2 => \N__6201\,
            in3 => \N__6367\,
            lcout => \mem_LUT_data_raw_r_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12289\,
            ce => \N__6177\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Clock_Count_586__i0_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7303\,
            in2 => \_gnd_net_\,
            in3 => \N__6138\,
            lcout => \pc_rx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_14_3_0_\,
            carryout => \pc_rx.n3060\,
            clk => \N__12316\,
            ce => \N__7832\,
            sr => \N__7583\
        );

    \pc_rx.r_Clock_Count_586__i1_LC_14_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7249\,
            in2 => \_gnd_net_\,
            in3 => \N__6135\,
            lcout => \pc_rx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \pc_rx.n3060\,
            carryout => \pc_rx.n3061\,
            clk => \N__12316\,
            ce => \N__7832\,
            sr => \N__7583\
        );

    \pc_rx.r_Clock_Count_586__i2_LC_14_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7264\,
            in2 => \_gnd_net_\,
            in3 => \N__6132\,
            lcout => \pc_rx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \pc_rx.n3061\,
            carryout => \pc_rx.n3062\,
            clk => \N__12316\,
            ce => \N__7832\,
            sr => \N__7583\
        );

    \pc_rx.r_Clock_Count_586__i3_LC_14_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7282\,
            in2 => \_gnd_net_\,
            in3 => \N__6129\,
            lcout => \pc_rx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \pc_rx.n3062\,
            carryout => \pc_rx.n3063\,
            clk => \N__12316\,
            ce => \N__7832\,
            sr => \N__7583\
        );

    \pc_rx.r_Clock_Count_586__i4_LC_14_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7198\,
            in2 => \_gnd_net_\,
            in3 => \N__6126\,
            lcout => \pc_rx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \pc_rx.n3063\,
            carryout => \pc_rx.n3064\,
            clk => \N__12316\,
            ce => \N__7832\,
            sr => \N__7583\
        );

    \pc_rx.r_Clock_Count_586__i5_LC_14_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7231\,
            in2 => \_gnd_net_\,
            in3 => \N__6123\,
            lcout => \pc_rx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \pc_rx.n3064\,
            carryout => \pc_rx.n3065\,
            clk => \N__12316\,
            ce => \N__7832\,
            sr => \N__7583\
        );

    \pc_rx.r_Clock_Count_586__i6_LC_14_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7216\,
            in2 => \_gnd_net_\,
            in3 => \N__6435\,
            lcout => \pc_rx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \pc_rx.n3065\,
            carryout => \pc_rx.n3066\,
            clk => \N__12316\,
            ce => \N__7832\,
            sr => \N__7583\
        );

    \pc_rx.r_Clock_Count_586__i7_LC_14_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7150\,
            in2 => \_gnd_net_\,
            in3 => \N__6432\,
            lcout => \pc_rx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \pc_rx.n3066\,
            carryout => \pc_rx.n3067\,
            clk => \N__12316\,
            ce => \N__7832\,
            sr => \N__7583\
        );

    \pc_rx.r_Clock_Count_586__i8_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7183\,
            in2 => \_gnd_net_\,
            in3 => \N__6429\,
            lcout => \pc_rx.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \bfn_14_4_0_\,
            carryout => \pc_rx.n3068\,
            clk => \N__12312\,
            ce => \N__7836\,
            sr => \N__7584\
        );

    \pc_rx.r_Clock_Count_586__i9_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__7168\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6426\,
            lcout => \pc_rx.r_Clock_Count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12312\,
            ce => \N__7836\,
            sr => \N__7584\
        );

    \tx_data_byte_r_i0_i4_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7427\,
            in1 => \N__11496\,
            in2 => \_gnd_net_\,
            in3 => \N__7616\,
            lcout => tx_data_byte_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i6_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7451\,
            in1 => \N__11460\,
            in2 => \_gnd_net_\,
            in3 => \N__7496\,
            lcout => tx_addr_byte_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i0_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7369\,
            in1 => \N__6407\,
            in2 => \_gnd_net_\,
            in3 => \N__6423\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i5_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11461\,
            in1 => \N__7726\,
            in2 => \_gnd_net_\,
            in3 => \N__7926\,
            lcout => tx_data_byte_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3176_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011110000"
        )
    port map (
            in0 => \N__6396\,
            in1 => \N__6504\,
            in2 => \N__8992\,
            in3 => \N__6372\,
            lcout => \tx_fifo.lscc_fifo_inst.n3564\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3166_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__8970\,
            in1 => \N__6477\,
            in2 => \N__6981\,
            in3 => \N__6371\,
            lcout => \tx_fifo.lscc_fifo_inst.n3552\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i146_147_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__8694\,
            in1 => \N__6800\,
            in2 => \N__6664\,
            in3 => \N__6515\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i230_231_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__6801\,
            in1 => \N__6893\,
            in2 => \N__10295\,
            in3 => \N__6503\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i134_135_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__6488\,
            in1 => \N__6799\,
            in2 => \N__6663\,
            in3 => \N__10287\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i347_348_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__6476\,
            in1 => \N__6802\,
            in2 => \N__6665\,
            in3 => \N__8814\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i3_2_lut_3_lut_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8603\,
            in1 => \N__8644\,
            in2 => \_gnd_net_\,
            in3 => \N__8562\,
            lcout => \tx_fifo.lscc_fifo_inst.n3\,
            ltout => \tx_fifo.lscc_fifo_inst.n3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i140_141_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__6458\,
            in1 => \N__6769\,
            in2 => \N__6468\,
            in3 => \N__9486\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i344_345_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__6771\,
            in1 => \N__6602\,
            in2 => \N__8739\,
            in3 => \N__6446\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_write_cmd_211_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__8643\,
            in1 => \N__7311\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => fifo_write_cmd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i4_2_lut_3_lut_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__8604\,
            in1 => \N__8645\,
            in2 => \_gnd_net_\,
            in3 => \N__8563\,
            lcout => \tx_fifo.lscc_fifo_inst.n4\,
            ltout => \tx_fifo.lscc_fifo_inst.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i251_252_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__6977\,
            in1 => \N__6770\,
            in2 => \N__6984\,
            in3 => \N__8824\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i233_234_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__6894\,
            in1 => \N__6803\,
            in2 => \N__6962\,
            in3 => \N__10370\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i239_240_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__6804\,
            in1 => \N__6895\,
            in2 => \N__6846\,
            in3 => \N__10405\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i7_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11501\,
            in1 => \N__8223\,
            in2 => \_gnd_net_\,
            in3 => \N__7685\,
            lcout => tx_addr_byte_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i335_336_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__10406\,
            in1 => \N__6805\,
            in2 => \N__6646\,
            in3 => \N__6554\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_adj_16_LC_15_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7184\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7232\,
            lcout => \pc_rx.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_3_lut_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7305\,
            in1 => \N__7251\,
            in2 => \_gnd_net_\,
            in3 => \N__7268\,
            lcout => OPEN,
            ltout => \pc_rx.n3399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i4_4_lut_LC_15_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__6543\,
            in1 => \N__7170\,
            in2 => \N__6537\,
            in3 => \N__6534\,
            lcout => \pc_rx.r_SM_Main_2_N_110_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i3043_4_lut_LC_15_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7152\,
            in1 => \N__7218\,
            in2 => \N__7287\,
            in3 => \N__7200\,
            lcout => \pc_rx.n3430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_4_lut_adj_17_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7304\,
            in1 => \N__7283\,
            in2 => \N__7269\,
            in3 => \N__7250\,
            lcout => OPEN,
            ltout => \pc_rx.n3400_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2252_4_lut_LC_15_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__7233\,
            in1 => \N__7217\,
            in2 => \N__7203\,
            in3 => \N__7199\,
            lcout => OPEN,
            ltout => \pc_rx.n2605_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2256_4_lut_LC_15_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__7185\,
            in1 => \N__7169\,
            in2 => \N__7155\,
            in3 => \N__7151\,
            lcout => \pc_rx.r_SM_Main_2_N_104_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Bit_Index_i0_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6995\,
            in1 => \N__7097\,
            in2 => \_gnd_net_\,
            in3 => \N__7034\,
            lcout => \r_Bit_Index_0_adj_489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_SM_Main_2__I_0_55_i3_3_lut_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100101"
        )
    port map (
            in0 => \N__8419\,
            in1 => \_gnd_net_\,
            in2 => \N__8379\,
            in3 => \N__7074\,
            lcout => \pc_tx.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i1163_4_lut_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__7536\,
            in1 => \N__10493\,
            in2 => \N__7023\,
            in3 => \N__8416\,
            lcout => \pc_tx.n1518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i1_3_lut_4_lut_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__8418\,
            in1 => \N__10494\,
            in2 => \N__8378\,
            in3 => \N__8463\,
            lcout => n1851,
            ltout => \n1851_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i1579_3_lut_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__7022\,
            in1 => \_gnd_net_\,
            in2 => \N__7005\,
            in3 => \N__8417\,
            lcout => n1934,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_SM_Main_i2_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__10490\,
            in1 => \N__8429\,
            in2 => \N__8472\,
            in3 => \N__8376\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i4_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__7799\,
            in1 => \N__9776\,
            in2 => \N__7428\,
            in3 => \N__8328\,
            lcout => pc_data_rx_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2_3_lut_4_lut_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8458\,
            in1 => \N__7531\,
            in2 => \N__8431\,
            in3 => \N__8374\,
            lcout => n1697,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i0_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__7798\,
            in1 => \N__9775\,
            in2 => \N__7341\,
            in3 => \N__9705\,
            lcout => pc_data_rx_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i3103_4_lut_4_lut_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000001100"
        )
    port map (
            in0 => \N__10489\,
            in1 => \N__7532\,
            in2 => \N__8432\,
            in3 => \N__8375\,
            lcout => OPEN,
            ltout => \n3381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Active_46_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011100"
        )
    port map (
            in0 => \N__8430\,
            in1 => \N__7552\,
            in2 => \N__7344\,
            in3 => \N__8462\,
            lcout => tx_uart_active_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i0_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7340\,
            in1 => \N__11459\,
            in2 => \_gnd_net_\,
            in3 => \N__7906\,
            lcout => tx_data_byte_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i6_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__7800\,
            in1 => \N__9777\,
            in2 => \N__8313\,
            in3 => \N__7322\,
            lcout => pc_data_rx_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_busy_falling_edge_209_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8663\,
            in2 => \_gnd_net_\,
            in3 => \N__7512\,
            lcout => spi_busy_falling_edge,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i0_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8000\,
            in1 => \N__11497\,
            in2 => \_gnd_net_\,
            in3 => \N__7907\,
            lcout => tx_addr_byte_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \start_tx_213_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__7530\,
            in1 => \N__7553\,
            in2 => \N__9060\,
            in3 => \N__9113\,
            lcout => \r_SM_Main_2_N_183_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i5_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11498\,
            in1 => \N__7733\,
            in2 => \_gnd_net_\,
            in3 => \N__7475\,
            lcout => tx_addr_byte_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_busy_prev_210_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8664\,
            lcout => spi_busy_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i6_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__8082\,
            in1 => \N__10128\,
            in2 => \N__7506\,
            in3 => \N__7713\,
            lcout => tx_shift_reg_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i13_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__10125\,
            in1 => \N__7476\,
            in2 => \N__8078\,
            in3 => \N__7464\,
            lcout => tx_shift_reg_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i12_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__7845\,
            in1 => \N__8055\,
            in2 => \N__7605\,
            in3 => \N__10129\,
            lcout => tx_shift_reg_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i14_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__10126\,
            in1 => \N__7458\,
            in2 => \N__8079\,
            in3 => \N__7440\,
            lcout => tx_shift_reg_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i3_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__7434\,
            in1 => \N__8056\,
            in2 => \N__7776\,
            in3 => \N__10130\,
            lcout => tx_shift_reg_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i2_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__7946\,
            in1 => \N__10131\,
            in2 => \N__8080\,
            in3 => \N__7869\,
            lcout => tx_shift_reg_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i5_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__10132\,
            in1 => \N__8057\,
            in2 => \N__7737\,
            in3 => \N__7701\,
            lcout => tx_shift_reg_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i4_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__10127\,
            in1 => \N__7628\,
            in2 => \N__8081\,
            in3 => \N__7707\,
            lcout => tx_shift_reg_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i15_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__7695\,
            in1 => \N__8054\,
            in2 => \N__7689\,
            in3 => \N__10119\,
            lcout => \DEBUG_8_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i15C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i4_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11500\,
            in1 => \N__7632\,
            in2 => \_gnd_net_\,
            in3 => \N__7598\,
            lcout => tx_addr_byte_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i2_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7950\,
            in1 => \N__11499\,
            in2 => \_gnd_net_\,
            in3 => \N__8108\,
            lcout => tx_addr_byte_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i3026_2_lut_3_lut_LC_16_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__9139\,
            in1 => \N__9771\,
            in2 => \_gnd_net_\,
            in3 => \N__9919\,
            lcout => OPEN,
            ltout => \pc_rx.n3412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_4_lut_LC_16_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000101"
        )
    port map (
            in0 => \N__9869\,
            in1 => \N__9947\,
            in2 => \N__7587\,
            in3 => \N__10035\,
            lcout => \pc_rx.n1946\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2_2_lut_adj_12_LC_16_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__9770\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9138\,
            lcout => OPEN,
            ltout => \pc_rx.n6_adj_487_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i3119_4_lut_LC_16_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__10036\,
            in1 => \N__9870\,
            in2 => \N__7839\,
            in3 => \N__9920\,
            lcout => \pc_rx.n1849\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2_2_lut_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9921\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9859\,
            lcout => n6,
            ltout => \n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_4_lut_adj_11_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__10037\,
            in1 => \N__8526\,
            in2 => \N__7809\,
            in3 => \N__9956\,
            lcout => n1787,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_4_lut_adj_13_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__9957\,
            in1 => \N__8527\,
            in2 => \N__8193\,
            in3 => \N__10038\,
            lcout => n1782,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_SM_Main_i1_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__10492\,
            in1 => \N__8415\,
            in2 => \_gnd_net_\,
            in3 => \N__8367\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12317\,
            ce => 'H',
            sr => \N__8475\
        );

    \pc_tx.r_SM_Main_i0_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__8366\,
            in1 => \N__10491\,
            in2 => \_gnd_net_\,
            in3 => \N__7806\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12317\,
            ce => 'H',
            sr => \N__8475\
        );

    \pc_rx.r_Rx_Byte_i2_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__8336\,
            in1 => \N__9772\,
            in2 => \N__7965\,
            in3 => \N__7797\,
            lcout => pc_data_rx_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i3_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__7766\,
            in1 => \_gnd_net_\,
            in2 => \N__7752\,
            in3 => \N__11458\,
            lcout => tx_data_byte_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i3_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7856\,
            in1 => \N__11456\,
            in2 => \_gnd_net_\,
            in3 => \N__7765\,
            lcout => tx_addr_byte_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i3_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__9773\,
            in1 => \N__8337\,
            in2 => \N__7751\,
            in3 => \N__9804\,
            lcout => pc_data_rx_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i2_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7964\,
            in1 => \N__11457\,
            in2 => \_gnd_net_\,
            in3 => \N__7939\,
            lcout => tx_data_byte_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i5_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__9805\,
            in1 => \N__9774\,
            in2 => \N__7925\,
            in3 => \N__8324\,
            lcout => pc_data_rx_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i0_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7908\,
            in1 => \N__11212\,
            in2 => \_gnd_net_\,
            in3 => \N__11056\,
            lcout => tx_shift_reg_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i0C_net\,
            ce => 'H',
            sr => \N__8883\
        );

    \spi0.i1_2_lut_3_lut_adj_18_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__11014\,
            in1 => \_gnd_net_\,
            in2 => \N__11211\,
            in3 => \N__11103\,
            lcout => n1763,
            ltout => \n1763_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i7_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__8219\,
            in1 => \N__7890\,
            in2 => \N__7881\,
            in3 => \N__10123\,
            lcout => tx_shift_reg_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i7C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i1_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__10120\,
            in1 => \N__7878\,
            in2 => \N__10641\,
            in3 => \N__8073\,
            lcout => tx_shift_reg_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i7C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i11_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__8070\,
            in1 => \N__8088\,
            in2 => \N__7863\,
            in3 => \N__10122\,
            lcout => tx_shift_reg_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i7C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i9_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__10121\,
            in1 => \N__10611\,
            in2 => \N__7989\,
            in3 => \N__8074\,
            lcout => tx_shift_reg_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i7C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i19_3_lut_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110011"
        )
    port map (
            in0 => \N__11102\,
            in1 => \N__11185\,
            in2 => \_gnd_net_\,
            in3 => \N__11015\,
            lcout => n3418,
            ltout => \n3418_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i10_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__8112\,
            in1 => \N__8097\,
            in2 => \N__8091\,
            in3 => \N__8072\,
            lcout => tx_shift_reg_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i7C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i8_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__8071\,
            in1 => \N__8010\,
            in2 => \N__8004\,
            in3 => \N__10124\,
            lcout => tx_shift_reg_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i7C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.state_reg_i2_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__11193\,
            in1 => \N__9422\,
            in2 => \N__7980\,
            in3 => \N__9450\,
            lcout => state_reg_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11317\,
            ce => 'H',
            sr => \N__9643\
        );

    \spi0.i1104_2_lut_4_lut_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001001100"
        )
    port map (
            in0 => \N__11105\,
            in1 => \N__11190\,
            in2 => \N__9372\,
            in3 => \N__11021\,
            lcout => \spi0.n1458\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i7_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__11023\,
            in1 => \N__9370\,
            in2 => \N__9300\,
            in3 => \N__9205\,
            lcout => \spi0.n500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11317\,
            ce => 'H',
            sr => \N__9643\
        );

    \spi0.state_reg_i0_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__9421\,
            in1 => \N__8841\,
            in2 => \_gnd_net_\,
            in3 => \N__9448\,
            lcout => state_reg_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11317\,
            ce => 'H',
            sr => \N__9643\
        );

    \spi0.i3099_2_lut_3_lut_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__11022\,
            in1 => \N__11106\,
            in2 => \_gnd_net_\,
            in3 => \N__9317\,
            lcout => \spi0.n3467\,
            ltout => \spi0.n3467_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.mux_514_i3_4_lut_4_lut_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__9420\,
            in1 => \N__11191\,
            in2 => \N__7971\,
            in3 => \N__9447\,
            lcout => OPEN,
            ltout => \spi0.state_next_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i1_4_lut_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__11192\,
            in1 => \N__11107\,
            in2 => \N__7968\,
            in3 => \N__9402\,
            lcout => \spi0.n4\,
            ltout => \spi0.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i8_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000010"
        )
    port map (
            in0 => \N__8166\,
            in1 => \N__9291\,
            in2 => \N__8160\,
            in3 => \N__11024\,
            lcout => \spi0.n499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11317\,
            ce => 'H',
            sr => \N__9643\
        );

    \spi0.t_FSM_i15_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__11040\,
            in1 => \N__8148\,
            in2 => \N__9297\,
            in3 => \N__9212\,
            lcout => \spi0.n492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11348\,
            ce => 'H',
            sr => \N__9670\
        );

    \spi0.mux_514_i2_4_lut_4_lut_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__9449\,
            in1 => \N__11213\,
            in2 => \N__9342\,
            in3 => \N__11036\,
            lcout => \spi0.state_next_1\,
            ltout => \spi0.state_next_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i0_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111011110"
        )
    port map (
            in0 => \N__11037\,
            in1 => \N__8157\,
            in2 => \N__8151\,
            in3 => \N__9206\,
            lcout => \spi0.n507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11348\,
            ce => 'H',
            sr => \N__9670\
        );

    \spi0.t_FSM_i14_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000010000"
        )
    port map (
            in0 => \N__9211\,
            in1 => \N__9270\,
            in2 => \N__8142\,
            in3 => \N__11042\,
            lcout => \spi0.n493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11348\,
            ce => 'H',
            sr => \N__9670\
        );

    \spi0.t_FSM_i13_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__11039\,
            in1 => \N__8133\,
            in2 => \N__9296\,
            in3 => \N__9210\,
            lcout => \spi0.n494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11348\,
            ce => 'H',
            sr => \N__9670\
        );

    \spi0.t_FSM_i12_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000010000"
        )
    port map (
            in0 => \N__9209\,
            in1 => \N__9269\,
            in2 => \N__8127\,
            in3 => \N__11041\,
            lcout => \spi0.n495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11348\,
            ce => 'H',
            sr => \N__9670\
        );

    \spi0.t_FSM_i11_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__11038\,
            in1 => \N__8118\,
            in2 => \N__9295\,
            in3 => \N__9208\,
            lcout => \spi0.n496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11348\,
            ce => 'H',
            sr => \N__9670\
        );

    \spi0.t_FSM_i10_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100000000"
        )
    port map (
            in0 => \N__9207\,
            in1 => \N__9268\,
            in2 => \N__11061\,
            in3 => \N__9387\,
            lcout => \spi0.n497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11348\,
            ce => 'H',
            sr => \N__9670\
        );

    \pc_rx.r_SM_Main_i0_LC_17_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__10027\,
            in1 => \N__8172\,
            in2 => \_gnd_net_\,
            in3 => \N__9153\,
            lcout => \pc_rx.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12331\,
            ce => 'H',
            sr => \N__9868\
        );

    \pc_rx.r_SM_Main_i1_LC_17_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100001010"
        )
    port map (
            in0 => \N__9909\,
            in1 => \N__9958\,
            in2 => \N__9123\,
            in3 => \N__10028\,
            lcout => \pc_rx.r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12331\,
            ce => 'H',
            sr => \N__9868\
        );

    \pc_rx.i1_3_lut_4_lut_LC_17_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8295\,
            in1 => \N__8524\,
            in2 => \N__8265\,
            in3 => \N__9981\,
            lcout => \pc_rx.r_SM_Main_2_N_107_0\,
            ltout => \pc_rx.r_SM_Main_2_N_107_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_3_lut_4_lut_adj_15_LC_17_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__9912\,
            in1 => \N__9848\,
            in2 => \N__8199\,
            in3 => \N__10033\,
            lcout => n3191,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i3133_3_lut_4_lut_LC_17_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__9982\,
            in1 => \N__9849\,
            in2 => \N__9925\,
            in3 => \N__10034\,
            lcout => \pc_rx.n3432\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_adj_10_LC_17_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9980\,
            lcout => OPEN,
            ltout => \n1801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Bit_Index_i0_LC_17_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010010"
        )
    port map (
            in0 => \N__8525\,
            in1 => \N__8486\,
            in2 => \N__8196\,
            in3 => \N__8192\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_LC_17_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110100011"
        )
    port map (
            in0 => \N__9983\,
            in1 => \N__8178\,
            in2 => \N__9926\,
            in3 => \_gnd_net_\,
            lcout => \pc_rx.n2615\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Bit_Index_i2_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8290\,
            in1 => \N__8529\,
            in2 => \_gnd_net_\,
            in3 => \N__8254\,
            lcout => \pc_rx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12321\,
            ce => \N__8499\,
            sr => \N__8493\
        );

    \pc_rx.r_Bit_Index_i1_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8289\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8528\,
            lcout => \pc_rx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12321\,
            ce => \N__8499\,
            sr => \N__8493\
        );

    \pc_tx.i1_1_lut_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8473\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pc_tx.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i3129_4_lut_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100011"
        )
    port map (
            in0 => \N__10472\,
            in1 => \N__8474\,
            in2 => \N__8433\,
            in3 => \N__8377\,
            lcout => \pc_tx.n1930\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.equal_260_i4_2_lut_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__8292\,
            in1 => \N__8256\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n4_adj_495,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.equal_259_i4_2_lut_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__8255\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8291\,
            lcout => n4_adj_494,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2175_2_lut_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__8294\,
            in1 => \N__8258\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n2527,
            ltout => \n2527_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i7_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__8231\,
            in1 => \N__9762\,
            in2 => \N__8298\,
            in3 => \N__9809\,
            lcout => pc_data_rx_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.equal_263_i4_2_lut_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__8293\,
            in1 => \N__8257\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i7_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8232\,
            in1 => \N__11455\,
            in2 => \_gnd_net_\,
            in3 => \N__8212\,
            lcout => tx_data_byte_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.state_reg_2__I_0_108_i5_3_lut_3_lut_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__11131\,
            in1 => \N__11214\,
            in2 => \_gnd_net_\,
            in3 => \N__11057\,
            lcout => \rx_shift_reg_15__N_315\,
            ltout => \rx_shift_reg_15__N_315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i7_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8784\,
            in2 => \N__8835\,
            in3 => \N__8802\,
            lcout => rx_buf_byte_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i8_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9500\,
            in2 => \_gnd_net_\,
            in3 => \N__10147\,
            lcout => rx_shift_reg_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i9_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__10146\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8747\,
            lcout => rx_shift_reg_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i5_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8759\,
            in1 => \N__9501\,
            in2 => \_gnd_net_\,
            in3 => \N__10318\,
            lcout => rx_buf_byte_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i6_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10319\,
            in1 => \N__8716\,
            in2 => \_gnd_net_\,
            in3 => \N__8748\,
            lcout => rx_buf_byte_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i4_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8682\,
            in1 => \N__10245\,
            in2 => \_gnd_net_\,
            in3 => \N__10317\,
            lcout => rx_buf_byte_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.busy_86_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__11058\,
            in1 => \_gnd_net_\,
            in2 => \N__11222\,
            in3 => \N__11132\,
            lcout => spi_busy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_r__i0_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110001101100110"
        )
    port map (
            in0 => \N__9674\,
            in1 => \N__8544\,
            in2 => \N__8652\,
            in3 => \N__8619\,
            lcout => wr_addr_r_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12310\,
            ce => 'H',
            sr => \N__9672\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r__i0_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000011110"
        )
    port map (
            in0 => \N__9114\,
            in1 => \N__9673\,
            in2 => \N__8938\,
            in3 => \N__9059\,
            lcout => rd_addr_r_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12310\,
            ce => 'H',
            sr => \N__9672\
        );

    \spi0.i1_1_lut_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11104\,
            lcout => \spi0.n895\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i531_4_lut_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__11186\,
            in1 => \N__11126\,
            in2 => \N__9371\,
            in3 => \N__11025\,
            lcout => n888,
            ltout => \n888_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.state_reg_i1_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__11018\,
            in1 => \N__11189\,
            in2 => \N__8871\,
            in3 => \N__9341\,
            lcout => state_reg_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11332\,
            ce => 'H',
            sr => \N__9669\
        );

    \spi0.t_FSM_i2_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100000000"
        )
    port map (
            in0 => \N__9214\,
            in1 => \N__11020\,
            in2 => \N__9298\,
            in3 => \N__8859\,
            lcout => \spi0.state_next_2__N_306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11332\,
            ce => 'H',
            sr => \N__9669\
        );

    \spi0.t_FSM_i1_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__11019\,
            in1 => \N__9280\,
            in2 => \N__8868\,
            in3 => \N__9213\,
            lcout => \spi0.state_next_2__N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11332\,
            ce => 'H',
            sr => \N__9669\
        );

    \spi0.i29_3_lut_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11613\,
            in1 => \N__11016\,
            in2 => \_gnd_net_\,
            in3 => \N__8858\,
            lcout => \spi0.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i3100_3_lut_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__11017\,
            in1 => \N__11187\,
            in2 => \_gnd_net_\,
            in3 => \N__9316\,
            lcout => OPEN,
            ltout => \spi0.n3476_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i28_4_lut_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110011"
        )
    port map (
            in0 => \N__11188\,
            in1 => \N__11125\,
            in2 => \N__8850\,
            in3 => \N__8847\,
            lcout => \spi0.n13\,
            ltout => \spi0.n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.mux_514_i1_3_lut_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__9446\,
            in1 => \N__9423\,
            in2 => \N__9405\,
            in3 => \_gnd_net_\,
            lcout => \spi0.state_next_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i9_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000010000"
        )
    port map (
            in0 => \N__9219\,
            in1 => \N__11055\,
            in2 => \N__9396\,
            in3 => \N__9290\,
            lcout => \spi0.n498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11350\,
            ce => 'H',
            sr => \N__9671\
        );

    \spi0.t_FSM_i5_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__9284\,
            in1 => \N__11027\,
            in2 => \N__9327\,
            in3 => \N__9217\,
            lcout => \spi0.n502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11350\,
            ce => 'H',
            sr => \N__9671\
        );

    \spi0.t_FSM_i6_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000010000"
        )
    port map (
            in0 => \N__9218\,
            in1 => \N__11054\,
            in2 => \N__9381\,
            in3 => \N__9289\,
            lcout => \state_next_2__N_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11350\,
            ce => 'H',
            sr => \N__9671\
        );

    \spi0.i1_2_lut_3_lut_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__9363\,
            in1 => \N__11119\,
            in2 => \_gnd_net_\,
            in3 => \N__11026\,
            lcout => \spi0.n911\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i4_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000010000"
        )
    port map (
            in0 => \N__9216\,
            in1 => \N__11053\,
            in2 => \N__9162\,
            in3 => \N__9288\,
            lcout => \spi0.n503\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11350\,
            ce => 'H',
            sr => \N__9671\
        );

    \spi0.t_FSM_i3_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__11052\,
            in1 => \N__9318\,
            in2 => \N__9299\,
            in3 => \N__9215\,
            lcout => \spi0.n504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11350\,
            ce => 'H',
            sr => \N__9671\
        );

    \pc_rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_18_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__9736\,
            in1 => \N__9147\,
            in2 => \_gnd_net_\,
            in3 => \N__9911\,
            lcout => \pc_rx.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_LC_18_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9735\,
            in2 => \_gnd_net_\,
            in3 => \N__9146\,
            lcout => \pc_rx.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i13_3_lut_4_lut_LC_18_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000001111"
        )
    port map (
            in0 => \N__9967\,
            in1 => \N__9847\,
            in2 => \N__10041\,
            in3 => \N__9910\,
            lcout => \pc_rx.n1798\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Data_50_LC_18_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11586\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_DV_52_LC_18_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__10039\,
            in1 => \N__11554\,
            in2 => \N__9858\,
            in3 => \N__10047\,
            lcout => \DEBUG_1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_SM_Main_i2_LC_18_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__10040\,
            in1 => \N__9984\,
            in2 => \N__9927\,
            in3 => \N__9846\,
            lcout => \pc_rx.r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i1_LC_18_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11475\,
            in1 => \N__10627\,
            in2 => \_gnd_net_\,
            in3 => \N__9689\,
            lcout => tx_data_byte_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i1_LC_18_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__9810\,
            in1 => \N__9737\,
            in2 => \N__9690\,
            in3 => \N__9704\,
            lcout => pc_data_rx_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.CS_81_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10650\,
            lcout => \DEBUG_9_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11316\,
            ce => 'H',
            sr => \N__9675\
        );

    \spi0.rx__5_i7_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__10161\,
            in1 => \N__10244\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rx_shift_reg_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i2_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10322\,
            in1 => \N__9466\,
            in2 => \_gnd_net_\,
            in3 => \N__10185\,
            lcout => rx_buf_byte_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i5_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__10160\,
            in1 => \N__10184\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rx_shift_reg_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i3_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10323\,
            in1 => \N__10390\,
            in2 => \_gnd_net_\,
            in3 => \N__10254\,
            lcout => rx_buf_byte_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i1_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10343\,
            in1 => \N__10059\,
            in2 => \_gnd_net_\,
            in3 => \N__10321\,
            lcout => rx_buf_byte_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i0_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10267\,
            in1 => \N__10173\,
            in2 => \_gnd_net_\,
            in3 => \N__10320\,
            lcout => rx_buf_byte_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i6_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10159\,
            in2 => \_gnd_net_\,
            in3 => \N__10253\,
            lcout => rx_shift_reg_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i2_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10155\,
            in2 => \_gnd_net_\,
            in3 => \N__10191\,
            lcout => rx_shift_reg_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i1_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__10232\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10157\,
            lcout => rx_shift_reg_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i4_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10156\,
            in2 => \_gnd_net_\,
            in3 => \N__10058\,
            lcout => rx_shift_reg_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i3_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10172\,
            in2 => \_gnd_net_\,
            in3 => \N__10158\,
            lcout => rx_shift_reg_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.CS_w_79_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11127\,
            in2 => \_gnd_net_\,
            in3 => \N__11218\,
            lcout => \spi0.CS_w\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11301\,
            ce => 'H',
            sr => \N__11059\
        );

    \tx_addr_byte_r_i0_i1_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10634\,
            in1 => \N__11502\,
            in2 => \_gnd_net_\,
            in3 => \N__10604\,
            lcout => tx_addr_byte_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i2_3_lut_LC_19_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11315\,
            in1 => \N__10558\,
            in2 => \_gnd_net_\,
            in3 => \N__11628\,
            lcout => \DEBUG_6_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i3_4_lut_LC_19_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10827\,
            in1 => \N__10428\,
            in2 => \N__10845\,
            in3 => \N__10443\,
            lcout => OPEN,
            ltout => \pc_tx.n3125_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i1_4_lut_LC_19_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__10782\,
            in1 => \N__10797\,
            in2 => \N__10500\,
            in3 => \N__10812\,
            lcout => OPEN,
            ltout => \pc_tx.n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2231_4_lut_LC_19_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__10767\,
            in1 => \N__10731\,
            in2 => \N__10497\,
            in3 => \N__10752\,
            lcout => \r_SM_Main_2_N_180_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Clock_Count_588__i0_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10442\,
            in2 => \_gnd_net_\,
            in3 => \N__10431\,
            lcout => \pc_tx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_19_7_0_\,
            carryout => \pc_tx.n3069\,
            clk => \N__12322\,
            ce => \N__10708\,
            sr => \N__10673\
        );

    \pc_tx.r_Clock_Count_588__i1_LC_19_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10427\,
            in2 => \_gnd_net_\,
            in3 => \N__10416\,
            lcout => \pc_tx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \pc_tx.n3069\,
            carryout => \pc_tx.n3070\,
            clk => \N__12322\,
            ce => \N__10708\,
            sr => \N__10673\
        );

    \pc_tx.r_Clock_Count_588__i2_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10841\,
            in2 => \_gnd_net_\,
            in3 => \N__10830\,
            lcout => \pc_tx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \pc_tx.n3070\,
            carryout => \pc_tx.n3071\,
            clk => \N__12322\,
            ce => \N__10708\,
            sr => \N__10673\
        );

    \pc_tx.r_Clock_Count_588__i3_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10826\,
            in2 => \_gnd_net_\,
            in3 => \N__10815\,
            lcout => \pc_tx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \pc_tx.n3071\,
            carryout => \pc_tx.n3072\,
            clk => \N__12322\,
            ce => \N__10708\,
            sr => \N__10673\
        );

    \pc_tx.r_Clock_Count_588__i4_LC_19_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10811\,
            in2 => \_gnd_net_\,
            in3 => \N__10800\,
            lcout => \pc_tx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \pc_tx.n3072\,
            carryout => \pc_tx.n3073\,
            clk => \N__12322\,
            ce => \N__10708\,
            sr => \N__10673\
        );

    \pc_tx.r_Clock_Count_588__i5_LC_19_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10796\,
            in2 => \_gnd_net_\,
            in3 => \N__10785\,
            lcout => \pc_tx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \pc_tx.n3073\,
            carryout => \pc_tx.n3074\,
            clk => \N__12322\,
            ce => \N__10708\,
            sr => \N__10673\
        );

    \pc_tx.r_Clock_Count_588__i6_LC_19_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10781\,
            in2 => \_gnd_net_\,
            in3 => \N__10770\,
            lcout => \pc_tx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \pc_tx.n3074\,
            carryout => \pc_tx.n3075\,
            clk => \N__12322\,
            ce => \N__10708\,
            sr => \N__10673\
        );

    \pc_tx.r_Clock_Count_588__i7_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10766\,
            in2 => \_gnd_net_\,
            in3 => \N__10755\,
            lcout => \pc_tx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \pc_tx.n3075\,
            carryout => \pc_tx.n3076\,
            clk => \N__12322\,
            ce => \N__10708\,
            sr => \N__10673\
        );

    \pc_tx.r_Clock_Count_588__i8_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10748\,
            in2 => \_gnd_net_\,
            in3 => \N__10737\,
            lcout => \pc_tx.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \bfn_19_8_0_\,
            carryout => \pc_tx.n3077\,
            clk => \N__12319\,
            ce => \N__10709\,
            sr => \N__10674\
        );

    \pc_tx.r_Clock_Count_588__i9_LC_19_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__10727\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10734\,
            lcout => \pc_tx.r_Clock_Count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12319\,
            ce => \N__10709\,
            sr => \N__10674\
        );

    \spi0.i4_4_lut_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__11658\,
            in1 => \N__10905\,
            in2 => \N__10923\,
            in3 => \N__10890\,
            lcout => OPEN,
            ltout => \spi0.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i3125_3_lut_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__10875\,
            in1 => \_gnd_net_\,
            in2 => \N__11358\,
            in3 => \N__10860\,
            lcout => \spi0.n1931\,
            ltout => \spi0.n1931_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.spi_clk_76_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__11264\,
            in1 => \_gnd_net_\,
            in2 => \N__11355\,
            in3 => \_gnd_net_\,
            lcout => \spi0.spi_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.state_reg_2__I_0_101_i5_2_lut_3_lut_LC_19_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__11223\,
            in1 => \N__11133\,
            in2 => \_gnd_net_\,
            in3 => \N__11060\,
            lcout => n5_adj_496,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.spi_clk_counter_589__i0_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10919\,
            in2 => \_gnd_net_\,
            in3 => \N__10908\,
            lcout => \spi0.spi_clk_counter_0\,
            ltout => OPEN,
            carryin => \bfn_19_10_0_\,
            carryout => \spi0.n3055\,
            clk => \N__12311\,
            ce => 'H',
            sr => \N__11646\
        );

    \spi0.spi_clk_counter_589__i1_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10904\,
            in2 => \N__11802\,
            in3 => \N__10893\,
            lcout => \spi0.spi_clk_counter_1\,
            ltout => OPEN,
            carryin => \spi0.n3055\,
            carryout => \spi0.n3056\,
            clk => \N__12311\,
            ce => 'H',
            sr => \N__11646\
        );

    \spi0.spi_clk_counter_589__i2_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10889\,
            in2 => \N__11804\,
            in3 => \N__10878\,
            lcout => \spi0.spi_clk_counter_2\,
            ltout => OPEN,
            carryin => \spi0.n3056\,
            carryout => \spi0.n3057\,
            clk => \N__12311\,
            ce => 'H',
            sr => \N__11646\
        );

    \spi0.spi_clk_counter_589__i3_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10874\,
            in2 => \N__11803\,
            in3 => \N__10863\,
            lcout => \spi0.spi_clk_counter_3\,
            ltout => OPEN,
            carryin => \spi0.n3057\,
            carryout => \spi0.n3058\,
            clk => \N__12311\,
            ce => 'H',
            sr => \N__11646\
        );

    \spi0.spi_clk_counter_589__i4_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10859\,
            in2 => \N__11805\,
            in3 => \N__10848\,
            lcout => \spi0.spi_clk_counter_4\,
            ltout => OPEN,
            carryin => \spi0.n3058\,
            carryout => \spi0.n3059\,
            clk => \N__12311\,
            ce => 'H',
            sr => \N__11646\
        );

    \spi0.spi_clk_counter_589__i5_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11762\,
            in1 => \N__11657\,
            in2 => \_gnd_net_\,
            in3 => \N__11661\,
            lcout => \spi0.spi_clk_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12311\,
            ce => 'H',
            sr => \N__11646\
        );

    \spi0.start_transfer_prev_74_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => start_transfer_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.start_transfer_edge_73_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__11634\,
            in1 => \N__11609\,
            in2 => \N__11528\,
            in3 => \N__11624\,
            lcout => start_transfer_edge,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Data_R_49_LC_22_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11598\,
            lcout => \pc_rx.r_Rx_Data_R\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_complete_rising_edge_214_LC_22_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__11541\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11570\,
            lcout => uart_rx_complete_rising_edge,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_complete_prev_215_LC_22_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11569\,
            lcout => uart_rx_complete_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debug_check_218_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11379\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11447\,
            lcout => \DEBUG_2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \even_byte_flag_221_LC_22_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11454\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11378\,
            lcout => even_byte_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12323\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i0_LC_24_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11367\,
            in2 => \_gnd_net_\,
            in3 => \N__11361\,
            lcout => n25,
            ltout => OPEN,
            carryin => \bfn_24_8_0_\,
            carryout => n3078,
            clk => \N__12336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i1_LC_24_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12057\,
            in2 => \_gnd_net_\,
            in3 => \N__12051\,
            lcout => n24,
            ltout => OPEN,
            carryin => n3078,
            carryout => n3079,
            clk => \N__12336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i2_LC_24_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12048\,
            in2 => \_gnd_net_\,
            in3 => \N__12042\,
            lcout => n23,
            ltout => OPEN,
            carryin => n3079,
            carryout => n3080,
            clk => \N__12336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i3_LC_24_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12039\,
            in2 => \_gnd_net_\,
            in3 => \N__12033\,
            lcout => n22,
            ltout => OPEN,
            carryin => n3080,
            carryout => n3081,
            clk => \N__12336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i4_LC_24_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12030\,
            in2 => \_gnd_net_\,
            in3 => \N__12024\,
            lcout => n21,
            ltout => OPEN,
            carryin => n3081,
            carryout => n3082,
            clk => \N__12336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i5_LC_24_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12021\,
            in2 => \_gnd_net_\,
            in3 => \N__12015\,
            lcout => n20,
            ltout => OPEN,
            carryin => n3082,
            carryout => n3083,
            clk => \N__12336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i6_LC_24_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12012\,
            in2 => \_gnd_net_\,
            in3 => \N__12006\,
            lcout => n19,
            ltout => OPEN,
            carryin => n3083,
            carryout => n3084,
            clk => \N__12336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i7_LC_24_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12003\,
            in2 => \_gnd_net_\,
            in3 => \N__11997\,
            lcout => n18,
            ltout => OPEN,
            carryin => n3084,
            carryout => n3085,
            clk => \N__12336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i8_LC_24_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11994\,
            in2 => \_gnd_net_\,
            in3 => \N__11988\,
            lcout => n17,
            ltout => OPEN,
            carryin => \bfn_24_9_0_\,
            carryout => n3086,
            clk => \N__12334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i9_LC_24_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12138\,
            in2 => \_gnd_net_\,
            in3 => \N__12132\,
            lcout => n16,
            ltout => OPEN,
            carryin => n3086,
            carryout => n3087,
            clk => \N__12334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i10_LC_24_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12129\,
            in2 => \_gnd_net_\,
            in3 => \N__12123\,
            lcout => n15,
            ltout => OPEN,
            carryin => n3087,
            carryout => n3088,
            clk => \N__12334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i11_LC_24_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12120\,
            in2 => \_gnd_net_\,
            in3 => \N__12114\,
            lcout => n14,
            ltout => OPEN,
            carryin => n3088,
            carryout => n3089,
            clk => \N__12334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i12_LC_24_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12111\,
            in2 => \_gnd_net_\,
            in3 => \N__12105\,
            lcout => n13,
            ltout => OPEN,
            carryin => n3089,
            carryout => n3090,
            clk => \N__12334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i13_LC_24_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12102\,
            in2 => \_gnd_net_\,
            in3 => \N__12096\,
            lcout => n12,
            ltout => OPEN,
            carryin => n3090,
            carryout => n3091,
            clk => \N__12334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i14_LC_24_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12093\,
            in2 => \_gnd_net_\,
            in3 => \N__12087\,
            lcout => n11,
            ltout => OPEN,
            carryin => n3091,
            carryout => n3092,
            clk => \N__12334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i15_LC_24_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12084\,
            in2 => \_gnd_net_\,
            in3 => \N__12078\,
            lcout => n10,
            ltout => OPEN,
            carryin => n3092,
            carryout => n3093,
            clk => \N__12334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i16_LC_24_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12075\,
            in2 => \_gnd_net_\,
            in3 => \N__12069\,
            lcout => n9,
            ltout => OPEN,
            carryin => \bfn_24_10_0_\,
            carryout => n3094,
            clk => \N__12333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i17_LC_24_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12066\,
            in2 => \_gnd_net_\,
            in3 => \N__12060\,
            lcout => n8_adj_490,
            ltout => OPEN,
            carryin => n3094,
            carryout => n3095,
            clk => \N__12333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i18_LC_24_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12423\,
            in2 => \_gnd_net_\,
            in3 => \N__12417\,
            lcout => n7,
            ltout => OPEN,
            carryin => n3095,
            carryout => n3096,
            clk => \N__12333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i19_LC_24_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12414\,
            in2 => \_gnd_net_\,
            in3 => \N__12408\,
            lcout => n6_adj_491,
            ltout => OPEN,
            carryin => n3096,
            carryout => n3097,
            clk => \N__12333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i20_LC_24_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12405\,
            in2 => \_gnd_net_\,
            in3 => \N__12399\,
            lcout => n5,
            ltout => OPEN,
            carryin => n3097,
            carryout => n3098,
            clk => \N__12333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i21_LC_24_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12396\,
            in2 => \_gnd_net_\,
            in3 => \N__12390\,
            lcout => n4_adj_492,
            ltout => OPEN,
            carryin => n3098,
            carryout => n3099,
            clk => \N__12333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i22_LC_24_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12387\,
            in2 => \_gnd_net_\,
            in3 => \N__12381\,
            lcout => n3,
            ltout => OPEN,
            carryin => n3099,
            carryout => n3100,
            clk => \N__12333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i23_LC_24_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12378\,
            in2 => \_gnd_net_\,
            in3 => \N__12372\,
            lcout => n2,
            ltout => OPEN,
            carryin => n3100,
            carryout => n3101,
            clk => \N__12333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_583_790__i24_LC_24_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12353\,
            in2 => \_gnd_net_\,
            in3 => \N__12369\,
            lcout => \DEBUG_0_c_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_SLM_CLK_c_THRU_LUT4_0_LC_24_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12342\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_SLM_CLK_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

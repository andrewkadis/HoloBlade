// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Jun 03 01:59:42 2020
//
// Verilog Description of module top
//

module top (ICE_SYSCLK, DCD, DSR, DTR, CTS, RST, UART_RX, UART_TX, 
            SEN, SCK, SOUT, SDAT, UPDATE, RESET, SLM_CLK, INVERT, 
            SYNC, VALID, DATA31, DATA0, DATA30, DATA29, DATA1, 
            DATA28, DATA27, DATA2, DATA26, DATA25, DATA3, DATA24, 
            DATA23, DATA4, DATA22, DATA21, DATA5, DATA20, DATA19, 
            DATA6, DATA18, DATA17, DATA7, DATA16, DATA15, DATA8, 
            DATA14, DATA13, DATA12, DATA11, DATA9, DATA10, FT_OE, 
            FT_RD, FT_WR, FT_SIWU, FR_RXF, FT_TXE, FIFO_BE3, FIFO_BE2, 
            FIFO_BE1, FIFO_BE0, FIFO_D31, FIFO_D30, FIFO_D29, FIFO_D28, 
            FIFO_D27, FIFO_CLK, FIFO_D26, FIFO_D25, FIFO_D24, FIFO_D23, 
            FIFO_D22, FIFO_D21, FIFO_D20, FIFO_D19, FIFO_D18, FIFO_D17, 
            FIFO_D16, FIFO_D15, FIFO_D14, FIFO_D13, FIFO_D12, FIFO_D11, 
            FIFO_D10, FIFO_D9, FIFO_D8, FIFO_D7, FIFO_D6, FIFO_D5, 
            FIFO_D4, FIFO_D3, FIFO_D2, FIFO_D1, FIFO_D0, DEBUG_0, 
            DEBUG_1, DEBUG_2, DEBUG_3, DEBUG_5, DEBUG_6, DEBUG_8, 
            DEBUG_9, ICE_CLK, ICE_CDONE, ICE_CREST) /* synthesis syn_module_defined=1 */ ;   // src/top.v(5[8:11])
    input ICE_SYSCLK;   // src/top.v(8[11:21])
    output DCD;   // src/top.v(11[12:15])
    output DSR;   // src/top.v(12[12:15])
    output DTR;   // src/top.v(13[12:15])
    output CTS;   // src/top.v(14[12:15])
    output RST;   // src/top.v(15[12:15])
    input UART_RX;   // src/top.v(16[12:19])
    output UART_TX;   // src/top.v(17[12:19])
    output SEN;   // src/top.v(20[12:15])
    output SCK;   // src/top.v(21[12:15])
    input SOUT;   // src/top.v(22[12:16])
    output SDAT;   // src/top.v(23[12:16])
    output UPDATE;   // src/top.v(27[12:18])
    output RESET;   // src/top.v(28[12:17])
    output SLM_CLK;   // src/top.v(29[12:19])
    output INVERT;   // src/top.v(30[12:18])
    output SYNC;   // src/top.v(31[12:16])
    output VALID;   // src/top.v(32[12:17])
    output DATA31;   // src/top.v(34[12:18])
    output DATA0;   // src/top.v(35[12:17])
    output DATA30;   // src/top.v(36[12:18])
    output DATA29;   // src/top.v(37[12:18])
    output DATA1;   // src/top.v(38[12:17])
    output DATA28;   // src/top.v(39[12:18])
    output DATA27;   // src/top.v(40[12:18])
    output DATA2;   // src/top.v(41[12:17])
    output DATA26;   // src/top.v(42[12:18])
    output DATA25;   // src/top.v(43[12:18])
    output DATA3;   // src/top.v(44[12:17])
    output DATA24;   // src/top.v(45[12:18])
    output DATA23;   // src/top.v(46[12:18])
    output DATA4;   // src/top.v(47[12:17])
    output DATA22;   // src/top.v(48[12:18])
    output DATA21;   // src/top.v(49[12:18])
    output DATA5;   // src/top.v(50[12:17])
    output DATA20;   // src/top.v(51[12:18])
    output DATA19;   // src/top.v(52[12:18])
    output DATA6;   // src/top.v(53[12:17])
    output DATA18;   // src/top.v(54[12:18])
    output DATA17;   // src/top.v(55[12:18])
    output DATA7;   // src/top.v(56[12:17])
    output DATA16;   // src/top.v(57[12:18])
    output DATA15;   // src/top.v(58[12:18])
    output DATA8;   // src/top.v(59[12:17])
    output DATA14;   // src/top.v(60[12:18])
    output DATA13;   // src/top.v(61[12:18])
    output DATA12;   // src/top.v(62[12:18])
    output DATA11;   // src/top.v(63[12:18])
    output DATA9;   // src/top.v(64[12:17])
    output DATA10;   // src/top.v(65[12:18])
    output FT_OE;   // src/top.v(69[12:17])
    output FT_RD;   // src/top.v(70[12:17])
    output FT_WR;   // src/top.v(71[12:17])
    output FT_SIWU;   // src/top.v(72[12:19])
    input FR_RXF;   // src/top.v(73[12:18])
    input FT_TXE;   // src/top.v(74[12:18])
    input FIFO_BE3;   // src/top.v(75[12:20])
    input FIFO_BE2;   // src/top.v(76[12:20])
    input FIFO_BE1;   // src/top.v(77[12:20])
    input FIFO_BE0;   // src/top.v(78[12:20])
    input FIFO_D31;   // src/top.v(79[12:20])
    input FIFO_D30;   // src/top.v(80[12:20])
    input FIFO_D29;   // src/top.v(81[12:20])
    input FIFO_D28;   // src/top.v(82[12:20])
    input FIFO_D27;   // src/top.v(83[12:20])
    input FIFO_CLK;   // src/top.v(84[12:20])
    input FIFO_D26;   // src/top.v(85[12:20])
    input FIFO_D25;   // src/top.v(86[12:20])
    input FIFO_D24;   // src/top.v(87[12:20])
    input FIFO_D23;   // src/top.v(88[12:20])
    input FIFO_D22;   // src/top.v(89[12:20])
    input FIFO_D21;   // src/top.v(90[12:20])
    input FIFO_D20;   // src/top.v(91[12:20])
    input FIFO_D19;   // src/top.v(92[12:20])
    input FIFO_D18;   // src/top.v(93[12:20])
    input FIFO_D17;   // src/top.v(94[12:20])
    input FIFO_D16;   // src/top.v(95[12:20])
    input FIFO_D15;   // src/top.v(97[11:19])
    input FIFO_D14;   // src/top.v(98[11:19])
    input FIFO_D13;   // src/top.v(99[11:19])
    input FIFO_D12;   // src/top.v(100[11:19])
    input FIFO_D11;   // src/top.v(101[11:19])
    input FIFO_D10;   // src/top.v(102[11:19])
    input FIFO_D9;   // src/top.v(103[11:18])
    input FIFO_D8;   // src/top.v(104[11:18])
    input FIFO_D7;   // src/top.v(105[11:18])
    input FIFO_D6;   // src/top.v(106[11:18])
    input FIFO_D5;   // src/top.v(107[11:18])
    input FIFO_D4;   // src/top.v(108[11:18])
    input FIFO_D3;   // src/top.v(109[11:18])
    input FIFO_D2;   // src/top.v(110[11:18])
    input FIFO_D1;   // src/top.v(111[11:18])
    input FIFO_D0;   // src/top.v(112[11:18])
    output DEBUG_0;   // src/top.v(115[12:19])
    output DEBUG_1;   // src/top.v(116[12:19])
    output DEBUG_2;   // src/top.v(117[12:19])
    output DEBUG_3;   // src/top.v(118[12:19])
    output DEBUG_5;   // src/top.v(119[12:19])
    output DEBUG_6;   // src/top.v(120[12:19])
    output DEBUG_8;   // src/top.v(121[12:19])
    output DEBUG_9;   // src/top.v(122[12:19])
    output ICE_CLK;   // src/top.v(125[12:19])
    output ICE_CDONE;   // src/top.v(126[12:21])
    output ICE_CREST;   // src/top.v(127[12:21])
    
    wire DEBUG_6_c /* synthesis SET_AS_NETWORK=DEBUG_6_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    
    wire GND_net, VCC_net, ICE_SYSCLK_c, UART_RX_c, UART_TX_c, SEN_c_1, 
        SCK_c_0, SOUT_c, SDAT_c_15, UPDATE_c_2, RESET_c, INVERT_c_3, 
        DEBUG_3_c, DEBUG_9_c, DATA15_c, DEBUG_5_c, DATA14_c, DATA13_c, 
        DATA17_c, DATA12_c, DATA11_c, DATA18_c, DATA10_c, DATA9_c, 
        DATA19_c, DATA8_c, DATA7_c, DATA20_c, DATA6_c, DATA5_c, 
        FT_OE_c, FT_RD_c, FR_RXF_c, FIFO_D15_c_15, FIFO_D14_c_14, 
        FIFO_D13_c_13, FIFO_D12_c_12, FIFO_D11_c_11, FIFO_D10_c_10, 
        FIFO_D9_c_9, FIFO_D8_c_8, FIFO_D7_c_7, FIFO_D6_c_6, FIFO_D5_c_5, 
        FIFO_D4_c_4, FIFO_D3_c_3, FIFO_D2_c_2, FIFO_D1_c_1, FIFO_D0_c_0, 
        DEBUG_0_c_24, DEBUG_1_c, DEBUG_2_c, debug_led3, n6602, reset_all_w;
    wire [3:0]reset_clk_counter;   // src/top.v(242[10:27])
    
    wire write_to_dc32_fifo;
    wire [3:0]state;   // src/timing_controller.v(44[11:16])
    
    wire dc32_fifo_is_full, \REG.mem_8_12 , \REG.mem_8_11 , \REG.mem_8_10 , 
        \REG.mem_8_9 , \REG.mem_8_8 , \REG.mem_8_7 , \REG.mem_8_6 , 
        \REG.mem_8_5 , \REG.mem_8_4 , \REG.mem_8_3 , \REG.mem_8_2 , 
        \REG.mem_8_1 , \REG.mem_8_0 ;
    wire [31:0]fifo_data_out;   // src/top.v(473[12:25])
    wire [6:0]num_words_in_buffer;   // src/top.v(474[12:31])
    
    wire reset_all, buffer_switch_done;
    wire [7:0]pc_data_rx;   // src/top.v(643[11:21])
    
    wire \REG.mem_10_10 , tx_uart_active_flag, spi_start_transfer_r, multi_byte_spi_trans_flag_r;
    wire [7:0]tx_addr_byte;   // src/top.v(765[11:23])
    wire [7:0]tx_data_byte;   // src/top.v(767[11:23])
    wire [7:0]rx_buf_byte;   // src/top.v(774[11:22])
    
    wire is_tx_fifo_full_flag, fifo_write_cmd, spi_rx_byte_ready, fifo_read_cmd, 
        is_fifo_empty_flag;
    wire [31:0]fifo_temp_output;   // src/top.v(864[12:28])
    
    wire even_byte_flag, uart_rx_complete_rising_edge, uart_rx_complete_prev, 
        reset_all_w_N_61, start_tx_N_64, pll_clk_unbuf, \REG.mem_15_15 , 
        multi_byte_spi_trans_flag_r_N_72, \REG.mem_7_15 , \REG.mem_7_14 , 
        \REG.mem_7_13 , \REG.mem_15_14 , \REG.mem_15_13 , \REG.mem_15_12 , 
        \REG.mem_15_11 , \REG.mem_15_10 , \REG.mem_15_9 , \REG.mem_15_8 , 
        \REG.mem_15_7 , \REG.mem_15_6 , \REG.mem_15_5 , \REG.mem_15_4 , 
        \REG.mem_15_3 , \REG.mem_15_2 , \REG.mem_15_1 , \REG.mem_15_0 , 
        \REG.mem_14_15 , \REG.mem_14_14 , \REG.mem_14_13 , \REG.mem_14_12 , 
        \REG.mem_14_11 , \REG.mem_14_10 , \REG.mem_14_9 , \REG.mem_14_8 , 
        \REG.mem_14_7 , \REG.mem_14_6 , \REG.mem_14_5 , \REG.mem_14_4 , 
        \REG.mem_14_3 , \REG.mem_14_2 , \REG.mem_14_1 , \REG.mem_14_0 , 
        \REG.mem_13_15 , \REG.mem_13_14 , \REG.mem_13_13 , \REG.mem_13_12 , 
        \REG.mem_13_11 , \REG.mem_13_10 , \REG.mem_13_9 , \REG.mem_13_8 , 
        \REG.mem_13_7 , \REG.mem_13_6 , \REG.mem_13_5 , \REG.mem_13_4 , 
        \REG.mem_13_3 , \REG.mem_13_2 , \REG.mem_13_1 , \REG.mem_13_0 , 
        \REG.mem_12_15 , \REG.mem_12_14 , \REG.mem_12_13 , \REG.mem_12_12 , 
        \REG.mem_12_11 , \REG.mem_12_10 , \REG.mem_12_9 , \REG.mem_12_8 , 
        \REG.mem_12_7 , \REG.mem_12_6 , \REG.mem_12_5 , \REG.mem_12_4 , 
        \REG.mem_12_3 , \REG.mem_12_2 , \REG.mem_12_1 , \REG.mem_12_0 , 
        \REG.mem_11_15 , \REG.mem_11_14 , \REG.mem_11_13 , \REG.mem_11_12 , 
        \REG.mem_11_11 , \REG.mem_11_10 , \REG.mem_11_9 , \REG.mem_11_8 , 
        \REG.mem_11_7 , \REG.mem_11_6 , \REG.mem_11_5 , \REG.mem_11_4 , 
        \REG.mem_11_3 , \REG.mem_11_2 , \REG.mem_11_1 , \REG.mem_11_0 , 
        n2414, n1586, \REG.mem_7_12 , \REG.mem_7_11 , \REG.mem_7_10 , 
        \REG.mem_7_9 , \REG.mem_7_8 , \REG.mem_7_7 , \REG.mem_7_6 , 
        \REG.mem_7_5 , \REG.mem_7_4 , \REG.mem_7_3 , \REG.mem_7_2 , 
        \REG.mem_7_1 , \REG.mem_7_0 , \REG.mem_6_15 , \REG.mem_6_14 , 
        \REG.mem_6_13 , \REG.mem_9_12 , \REG.mem_9_11 , \REG.mem_9_10 , 
        \REG.mem_9_9 , \REG.mem_9_8 , \REG.mem_9_7 , \REG.mem_9_6 , 
        \REG.mem_9_5 , \REG.mem_9_4 , n4, \REG.mem_9_3 , \REG.mem_9_2 , 
        \REG.mem_9_1 , \REG.mem_9_0 , n4169, n4168, n4167, n4166, 
        n4165, n4164, \REG.mem_6_12 , \REG.mem_6_11 , \REG.mem_6_10 , 
        \REG.mem_6_9 , \REG.mem_6_8 , \REG.mem_6_7 , \REG.mem_6_6 , 
        \REG.mem_6_5 , r_Rx_Data;
    wire [2:0]r_Bit_Index;   // src/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // src/uart_rx.v(36[17:26])
    
    wire n1431, \REG.mem_10_9 , n4163, n4162, n4161, n6572, \REG.mem_10_8 , 
        n4160, n4159, n4158, n4157, n4156, n4155;
    wire [2:0]r_SM_Main_adj_1138;   // src/uart_tx.v(31[16:25])
    wire [7:0]r_Tx_Data;   // src/uart_tx.v(34[16:25])
    wire [2:0]r_SM_Main_2__N_728;
    wire [2:0]r_SM_Main_2__N_725;
    
    wire \REG.mem_10_7 , \REG.mem_10_6 , n4154, \REG.mem_10_15 ;
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    wire [15:0]rx_shift_reg;   // src/spi.v(72[12:24])
    
    wire \REG.mem_10_5 , \REG.mem_10_14 , \REG.mem_10_4 , n4145, \REG.mem_10_13 , 
        \REG.mem_10_12 , \REG.mem_10_11 , n4_adj_1098, n131, \REG.mem_8_15 , 
        n3533, \REG.mem_10_3 , n4144, n4143, n4137, n4135, \REG.mem_6_4 , 
        \REG.mem_6_3 , \REG.mem_6_2 , \REG.mem_6_1 , \REG.mem_6_0 , 
        \REG.mem_8_14 , \REG.mem_10_2 , \REG.mem_8_13 , n3151, n4_adj_1099, 
        \REG.mem_5_15 , \REG.mem_5_14 , \REG.mem_5_13 , \REG.mem_5_12 , 
        \REG.mem_5_11 , \REG.mem_5_10 , \REG.mem_5_9 , \REG.mem_5_8 , 
        \REG.mem_5_7 , \REG.mem_5_6 , \REG.mem_5_5 , \REG.mem_5_4 , 
        \REG.mem_5_3 , \REG.mem_5_2 , \REG.mem_5_1 , \REG.mem_5_0 ;
    wire [6:0]wr_addr_r;   // src/fifo_dc_32_lut_gen.v(194[29:38])
    wire [6:0]wr_addr_nxt_c;   // src/fifo_dc_32_lut_gen.v(196[29:42])
    wire [6:0]rp_sync1_r;   // src/fifo_dc_32_lut_gen.v(199[37:47])
    wire [6:0]wr_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(202[37:51])
    wire [6:0]rd_addr_r;   // src/fifo_dc_32_lut_gen.v(215[29:38])
    
    wire \REG.mem_9_13 , \REG.mem_9_14 , \REG.mem_9_15 ;
    wire [6:0]wp_sync1_r;   // src/fifo_dc_32_lut_gen.v(220[37:47])
    wire [6:0]rd_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(223[37:51])
    
    wire t_rd_fifo_en_w;
    wire [31:0]\REG.out_raw ;   // src/fifo_dc_32_lut_gen.v(877[47:54])
    
    wire \REG.mem_2_2 , \REG.mem_2_1 , \REG.mem_2_0 , n4130;
    wire [6:0]rd_addr_nxt_c_6__N_176;
    
    wire n8, n4129, n8_adj_1100, n4123, rd_fifo_en_w, rd_fifo_en_prev_r;
    wire [2:0]wr_addr_r_adj_1162;   // src/fifo_quad_word_mod.v(65[31:40])
    wire [2:0]wr_addr_p1_w_adj_1164;   // src/fifo_quad_word_mod.v(67[32:44])
    wire [2:0]rd_addr_r_adj_1165;   // src/fifo_quad_word_mod.v(69[31:40])
    wire [2:0]rd_addr_p1_w_adj_1167;   // src/fifo_quad_word_mod.v(71[32:44])
    
    wire full_nxt_r, n32, n24;
    wire [31:0]\mem_LUT.data_raw_r ;   // src/fifo_quad_word_mod.v(449[42:52])
    
    wire n4115, n15, n8987, n5353, n2326, \REG.mem_2_15 , \REG.mem_2_14 , 
        \REG.mem_2_13 , \REG.mem_2_12 , \REG.mem_2_11 , \REG.mem_2_10 , 
        \REG.mem_2_9 , \REG.mem_2_8 , \REG.mem_2_7 , \REG.mem_2_6 , 
        \REG.mem_2_5 , \REG.mem_2_4 , \REG.mem_2_3 , n2410, n4111, 
        n5349, n5348, n5347, n5345, n5344, n5339, n5338, n5337, 
        n3785, n1638, n4108, \REG.mem_10_1 , \REG.mem_10_0 , n4107, 
        n1326, \REG.mem_18_0 , \REG.mem_18_1 , \REG.mem_18_2 , \REG.mem_18_3 , 
        \REG.mem_18_4 , \REG.mem_18_5 , \REG.mem_18_6 , \REG.mem_18_7 , 
        \REG.mem_18_8 , \REG.mem_18_9 , \REG.mem_18_10 , \REG.mem_18_11 , 
        \REG.mem_18_12 , \REG.mem_18_13 , \REG.mem_18_14 , \REG.mem_18_15 , 
        \REG.mem_19_0 , \REG.mem_19_1 , \REG.mem_19_2 , \REG.mem_19_3 , 
        \REG.mem_19_4 , \REG.mem_19_5 , \REG.mem_19_6 , \REG.mem_19_7 , 
        \REG.mem_19_8 , \REG.mem_19_9 , \REG.mem_19_10 , \REG.mem_19_11 , 
        \REG.mem_19_12 , \REG.mem_19_13 , \REG.mem_19_14 , \REG.mem_19_15 , 
        n4103, n3525, n5330, \REG.mem_21_0 , \REG.mem_21_1 , \REG.mem_21_2 , 
        \REG.mem_21_3 , \REG.mem_21_4 , \REG.mem_21_5 , \REG.mem_21_6 , 
        \REG.mem_21_7 , \REG.mem_21_8 , \REG.mem_21_9 , \REG.mem_21_10 , 
        \REG.mem_21_11 , \REG.mem_21_12 , \REG.mem_21_13 , \REG.mem_21_14 , 
        \REG.mem_21_15 , \REG.mem_22_0 , \REG.mem_22_1 , \REG.mem_22_2 , 
        \REG.mem_22_3 , \REG.mem_22_4 , \REG.mem_22_5 , \REG.mem_22_6 , 
        \REG.mem_22_7 , \REG.mem_22_8 , \REG.mem_22_9 , \REG.mem_22_10 , 
        \REG.mem_22_11 , \REG.mem_22_12 , \REG.mem_22_13 , \REG.mem_22_14 , 
        \REG.mem_22_15 , \REG.mem_23_0 , \REG.mem_23_1 , \REG.mem_23_2 , 
        \REG.mem_23_3 , \REG.mem_23_4 , \REG.mem_23_5 , \REG.mem_23_6 , 
        \REG.mem_23_7 , \REG.mem_23_8 , \REG.mem_23_9 , \REG.mem_23_10 , 
        \REG.mem_23_11 , \REG.mem_23_12 , \REG.mem_23_13 , \REG.mem_23_14 , 
        \REG.mem_23_15 , \REG.mem_24_0 , \REG.mem_24_1 , \REG.mem_24_2 , 
        \REG.mem_24_3 , \REG.mem_24_4 , \REG.mem_24_5 , \REG.mem_24_6 , 
        \REG.mem_24_7 , \REG.mem_24_8 , \REG.mem_24_9 , \REG.mem_24_10 , 
        \REG.mem_24_11 , \REG.mem_24_12 , \REG.mem_24_13 , \REG.mem_24_14 , 
        \REG.mem_24_15 , \REG.mem_25_0 , \REG.mem_25_1 , \REG.mem_25_2 , 
        \REG.mem_25_3 , \REG.mem_25_4 , \REG.mem_25_5 , \REG.mem_25_6 , 
        \REG.mem_25_7 , \REG.mem_25_8 , \REG.mem_25_9 , \REG.mem_25_10 , 
        \REG.mem_25_11 , \REG.mem_25_12 , \REG.mem_25_13 , \REG.mem_25_14 , 
        \REG.mem_25_15 , \REG.mem_26_0 , \REG.mem_26_1 , \REG.mem_26_2 , 
        \REG.mem_26_3 , \REG.mem_26_4 , \REG.mem_26_5 , \REG.mem_26_6 , 
        \REG.mem_26_7 , \REG.mem_26_8 , \REG.mem_26_9 , \REG.mem_26_10 , 
        \REG.mem_26_11 , \REG.mem_26_12 , \REG.mem_26_13 , \REG.mem_26_14 , 
        \REG.mem_26_15 , \REG.mem_28_0 , \REG.mem_28_1 , \REG.mem_28_2 , 
        \REG.mem_28_3 , \REG.mem_28_4 , \REG.mem_28_5 , \REG.mem_28_6 , 
        \REG.mem_28_7 , \REG.mem_28_8 , \REG.mem_28_9 , \REG.mem_28_10 , 
        \REG.mem_28_11 , \REG.mem_28_12 , \REG.mem_28_13 , \REG.mem_28_14 , 
        \REG.mem_28_15 , \REG.mem_29_0 , \REG.mem_29_1 , \REG.mem_29_2 , 
        \REG.mem_29_3 , \REG.mem_29_4 , \REG.mem_29_5 , \REG.mem_29_6 , 
        \REG.mem_29_7 , \REG.mem_29_8 , \REG.mem_29_9 , \REG.mem_29_10 , 
        \REG.mem_29_11 , \REG.mem_29_12 , \REG.mem_29_13 , \REG.mem_29_14 , 
        \REG.mem_29_15 , \REG.mem_30_0 , \REG.mem_30_1 , \REG.mem_30_2 , 
        \REG.mem_30_3 , \REG.mem_30_4 , \REG.mem_30_5 , \REG.mem_30_6 , 
        \REG.mem_30_7 , \REG.mem_30_8 , \REG.mem_30_9 , \REG.mem_30_10 , 
        \REG.mem_30_11 , \REG.mem_30_12 , \REG.mem_30_13 , \REG.mem_30_14 , 
        \REG.mem_30_15 , n5327, \REG.mem_34_0 , \REG.mem_34_1 , \REG.mem_34_2 , 
        \REG.mem_34_3 , \REG.mem_34_4 , \REG.mem_34_5 , \REG.mem_34_6 , 
        \REG.mem_34_7 , \REG.mem_34_8 , \REG.mem_34_9 , \REG.mem_34_10 , 
        \REG.mem_34_11 , \REG.mem_34_12 , \REG.mem_34_13 , \REG.mem_34_14 , 
        \REG.mem_34_15 , n10552, \REG.mem_37_0 , \REG.mem_37_1 , \REG.mem_37_2 , 
        \REG.mem_37_3 , \REG.mem_37_4 , \REG.mem_37_5 , \REG.mem_37_6 , 
        \REG.mem_37_7 , \REG.mem_37_8 , \REG.mem_37_9 , \REG.mem_37_10 , 
        \REG.mem_37_11 , \REG.mem_37_12 , \REG.mem_37_13 , \REG.mem_37_14 , 
        \REG.mem_37_15 , \REG.mem_38_0 , \REG.mem_38_1 , \REG.mem_38_2 , 
        \REG.mem_38_3 , \REG.mem_38_4 , \REG.mem_38_5 , \REG.mem_38_6 , 
        \REG.mem_38_7 , \REG.mem_38_8 , \REG.mem_38_9 , \REG.mem_38_10 , 
        \REG.mem_38_11 , \REG.mem_38_12 , \REG.mem_38_13 , \REG.mem_38_14 , 
        \REG.mem_38_15 , \REG.mem_39_0 , \REG.mem_39_1 , \REG.mem_39_2 , 
        \REG.mem_39_3 , \REG.mem_39_4 , \REG.mem_39_5 , \REG.mem_39_6 , 
        \REG.mem_39_7 , \REG.mem_39_8 , \REG.mem_39_9 , \REG.mem_39_10 , 
        \REG.mem_39_11 , \REG.mem_39_12 , \REG.mem_39_13 , \REG.mem_39_14 , 
        \REG.mem_39_15 , \REG.mem_40_0 , \REG.mem_40_1 , \REG.mem_40_2 , 
        \REG.mem_40_3 , \REG.mem_40_4 , \REG.mem_40_5 , \REG.mem_40_6 , 
        \REG.mem_40_7 , \REG.mem_40_8 , \REG.mem_40_9 , \REG.mem_40_10 , 
        \REG.mem_40_11 , \REG.mem_40_12 , \REG.mem_40_13 , \REG.mem_40_14 , 
        \REG.mem_40_15 , n3734, \REG.mem_41_0 , \REG.mem_41_1 , \REG.mem_41_2 , 
        \REG.mem_41_3 , \REG.mem_41_4 , \REG.mem_41_5 , \REG.mem_41_6 , 
        \REG.mem_41_7 , \REG.mem_41_8 , \REG.mem_41_9 , \REG.mem_41_10 , 
        \REG.mem_41_11 , \REG.mem_41_12 , \REG.mem_41_13 , \REG.mem_41_14 , 
        \REG.mem_41_15 , n9299, \REG.mem_42_0 , \REG.mem_42_1 , \REG.mem_42_2 , 
        \REG.mem_42_3 , \REG.mem_42_4 , \REG.mem_42_5 , \REG.mem_42_6 , 
        \REG.mem_42_7 , \REG.mem_42_8 , \REG.mem_42_9 , \REG.mem_42_10 , 
        \REG.mem_42_11 , \REG.mem_42_12 , \REG.mem_42_13 , \REG.mem_42_14 , 
        \REG.mem_42_15 , \REG.mem_43_0 , \REG.mem_43_1 , \REG.mem_43_2 , 
        \REG.mem_43_3 , \REG.mem_43_4 , \REG.mem_43_5 , \REG.mem_43_6 , 
        \REG.mem_43_7 , \REG.mem_43_8 , \REG.mem_43_9 , \REG.mem_43_10 , 
        \REG.mem_43_11 , \REG.mem_43_12 , \REG.mem_43_13 , \REG.mem_43_14 , 
        \REG.mem_43_15 , n8963, \REG.mem_44_0 , \REG.mem_44_1 , \REG.mem_44_2 , 
        \REG.mem_44_3 , \REG.mem_44_4 , \REG.mem_44_5 , \REG.mem_44_6 , 
        \REG.mem_44_7 , \REG.mem_44_8 , \REG.mem_44_9 , \REG.mem_44_10 , 
        \REG.mem_44_11 , \REG.mem_44_12 , \REG.mem_44_13 , \REG.mem_44_14 , 
        \REG.mem_44_15 , n9355, \REG.mem_45_0 , \REG.mem_45_1 , \REG.mem_45_2 , 
        \REG.mem_45_3 , \REG.mem_45_4 , \REG.mem_45_5 , \REG.mem_45_6 , 
        \REG.mem_45_7 , \REG.mem_45_8 , \REG.mem_45_9 , \REG.mem_45_10 , 
        \REG.mem_45_11 , \REG.mem_45_12 , \REG.mem_45_13 , \REG.mem_45_14 , 
        \REG.mem_45_15 , n2851, n9345, n4101, \REG.mem_46_0 , \REG.mem_46_1 , 
        \REG.mem_46_2 , \REG.mem_46_3 , \REG.mem_46_4 , \REG.mem_46_5 , 
        \REG.mem_46_6 , \REG.mem_46_7 , \REG.mem_46_8 , \REG.mem_46_9 , 
        \REG.mem_46_10 , \REG.mem_46_11 , \REG.mem_46_12 , \REG.mem_46_13 , 
        \REG.mem_46_14 , \REG.mem_46_15 , \REG.mem_47_0 , \REG.mem_47_1 , 
        \REG.mem_47_2 , \REG.mem_47_3 , \REG.mem_47_4 , \REG.mem_47_5 , 
        \REG.mem_47_6 , \REG.mem_47_7 , \REG.mem_47_8 , \REG.mem_47_9 , 
        \REG.mem_47_10 , \REG.mem_47_11 , \REG.mem_47_12 , \REG.mem_47_13 , 
        \REG.mem_47_14 , \REG.mem_47_15 , n5317, \REG.mem_50_0 , \REG.mem_50_1 , 
        \REG.mem_50_2 , \REG.mem_50_3 , \REG.mem_50_4 , \REG.mem_50_5 , 
        \REG.mem_50_6 , \REG.mem_50_7 , \REG.mem_50_8 , \REG.mem_50_9 , 
        \REG.mem_50_10 , \REG.mem_50_11 , \REG.mem_50_12 , \REG.mem_50_13 , 
        \REG.mem_50_14 , \REG.mem_50_15 , \REG.mem_51_0 , \REG.mem_51_1 , 
        \REG.mem_51_2 , \REG.mem_51_3 , \REG.mem_51_4 , \REG.mem_51_5 , 
        \REG.mem_51_6 , \REG.mem_51_7 , \REG.mem_51_8 , \REG.mem_51_9 , 
        \REG.mem_51_10 , \REG.mem_51_11 , \REG.mem_51_12 , \REG.mem_51_13 , 
        \REG.mem_51_14 , \REG.mem_51_15 , n5314, \REG.mem_53_0 , \REG.mem_53_1 , 
        \REG.mem_53_2 , \REG.mem_53_3 , \REG.mem_53_4 , \REG.mem_53_5 , 
        \REG.mem_53_6 , \REG.mem_53_7 , \REG.mem_53_8 , \REG.mem_53_9 , 
        \REG.mem_53_10 , \REG.mem_53_11 , \REG.mem_53_12 , \REG.mem_53_13 , 
        \REG.mem_53_14 , \REG.mem_53_15 , \REG.mem_54_0 , \REG.mem_54_1 , 
        \REG.mem_54_2 , \REG.mem_54_3 , \REG.mem_54_4 , \REG.mem_54_5 , 
        \REG.mem_54_6 , \REG.mem_54_7 , \REG.mem_54_8 , \REG.mem_54_9 , 
        \REG.mem_54_10 , \REG.mem_54_11 , \REG.mem_54_12 , \REG.mem_54_13 , 
        \REG.mem_54_14 , \REG.mem_54_15 , \REG.mem_55_0 , \REG.mem_55_1 , 
        \REG.mem_55_2 , \REG.mem_55_3 , \REG.mem_55_4 , \REG.mem_55_5 , 
        \REG.mem_55_6 , \REG.mem_55_7 , \REG.mem_55_8 , \REG.mem_55_9 , 
        \REG.mem_55_10 , \REG.mem_55_11 , \REG.mem_55_12 , \REG.mem_55_13 , 
        \REG.mem_55_14 , \REG.mem_55_15 , \REG.mem_56_0 , \REG.mem_56_1 , 
        \REG.mem_56_2 , \REG.mem_56_3 , \REG.mem_56_4 , \REG.mem_56_5 , 
        \REG.mem_56_6 , \REG.mem_56_7 , \REG.mem_56_8 , \REG.mem_56_9 , 
        \REG.mem_56_10 , \REG.mem_56_11 , \REG.mem_56_12 , \REG.mem_56_13 , 
        \REG.mem_56_14 , \REG.mem_56_15 , \REG.mem_57_0 , \REG.mem_57_1 , 
        \REG.mem_57_2 , \REG.mem_57_3 , \REG.mem_57_4 , \REG.mem_57_5 , 
        \REG.mem_57_6 , \REG.mem_57_7 , \REG.mem_57_8 , \REG.mem_57_9 , 
        \REG.mem_57_10 , \REG.mem_57_11 , \REG.mem_57_12 , \REG.mem_57_13 , 
        \REG.mem_57_14 , \REG.mem_57_15 , \REG.mem_58_0 , \REG.mem_58_1 , 
        \REG.mem_58_2 , \REG.mem_58_3 , \REG.mem_58_4 , \REG.mem_58_5 , 
        \REG.mem_58_6 , \REG.mem_58_7 , \REG.mem_58_8 , \REG.mem_58_9 , 
        \REG.mem_58_10 , \REG.mem_58_11 , \REG.mem_58_12 , \REG.mem_58_13 , 
        \REG.mem_58_14 , \REG.mem_58_15 , \REG.mem_60_0 , \REG.mem_60_1 , 
        \REG.mem_60_2 , \REG.mem_60_3 , \REG.mem_60_4 , \REG.mem_60_5 , 
        \REG.mem_60_6 , \REG.mem_60_7 , \REG.mem_60_8 , \REG.mem_60_9 , 
        \REG.mem_60_10 , \REG.mem_60_11 , \REG.mem_60_12 , \REG.mem_60_13 , 
        \REG.mem_60_14 , \REG.mem_60_15 , \REG.mem_61_0 , \REG.mem_61_1 , 
        \REG.mem_61_2 , \REG.mem_61_3 , \REG.mem_61_4 , \REG.mem_61_5 , 
        \REG.mem_61_6 , \REG.mem_61_7 , \REG.mem_61_8 , \REG.mem_61_9 , 
        \REG.mem_61_10 , \REG.mem_61_11 , \REG.mem_61_12 , \REG.mem_61_13 , 
        \REG.mem_61_14 , \REG.mem_61_15 , \REG.mem_62_0 , \REG.mem_62_1 , 
        \REG.mem_62_2 , \REG.mem_62_3 , \REG.mem_62_4 , \REG.mem_62_5 , 
        \REG.mem_62_6 , \REG.mem_62_7 , \REG.mem_62_8 , \REG.mem_62_9 , 
        \REG.mem_62_10 , \REG.mem_62_11 , \REG.mem_62_12 , \REG.mem_62_13 , 
        \REG.mem_62_14 , \REG.mem_62_15 , n3, n4_adj_1101, n5, n7, 
        n8_adj_1102, n9, n10, n11, n12, n14, n15_adj_1103, n18, 
        n19, n20, n21, n22, n23, n24_adj_1104, n25, n26, n27, 
        n28, n31, n35, n36, n37, n39, n40, n41, n42, n43, 
        n44, n46, n47, n50, n51, n52, n53, n54, n55, n56, 
        n57, n58, n59, n60, n63, n5311, n5308, n5305, n5302, 
        n5299, n5296, n63_adj_1105, n5293, n5290, n5287, n5286, 
        n5285, n5276, n5275, n5274, n5265, n5255, n5252, n5249, 
        n5236, n5233, n5230, n5212, n5208, n5207, n5206, n5205, 
        n5204, n5203, n5202, n5201, n5200, n5199, n5198, n5197, 
        n5196, n5195, n5194, n5193, n5192, n5191, n5190, n5189, 
        n5188, n5187, n5186, n5185, n5184, n5183, n5182, n5181, 
        n5180, n5179, n5178, n5177, n5176, n5175, n5174, n5173, 
        n5172, n5171, n5170, n5169, n5168, n5167, n5166, n5165, 
        n5164, n5163, n5162, n5161, n5144, n5143, n5142, n5141, 
        n5140, n5139, n5138, n5137, n5136, n5135, n5134, n5133, 
        n5132, n5131, n5130, n5129, n5128, n5127, n5126, n5125, 
        n5124, n5123, n5122, n5121, n5120, n5119, n5118, n5117, 
        n5116, n5115, n5114, n5113, n5110, n5109, n5108, n5107, 
        n5106, n5105, n5104, n5103, n5102, n5101, n5100, n5099, 
        n5098, n5097, n5096, n5095, n5094, n5091, n5090, n5089, 
        n5088, n5087, n5086, n5085, n5084, n5083, n5082, n5081, 
        n5080, n5079, n5078, n5077, n5076, n5075, n5074, n5073, 
        n5072, n5071, n5070, n5069, n5068, n5067, n5066, n5065, 
        n5064, n5063, n5062, n5061, n5060, n5057, n5056, n5055, 
        n5054, n5053, n5052, n5051, n5050, n5049, n5048, n5047, 
        n5046, n5045, n5044, n5043, n5042, n5041, n5024, n5023, 
        n5022, n5021, n5020, n5019, n5018, n5017, n5016, n5015, 
        n5014, n5013, n5012, n5011, n5010, n5008, n5007, n5006, 
        n5005, n5004, n5003, n5002, n5001, n5000, n4999, n4998, 
        n4997, n4996, n4995, n4994, n4993, n4992, n4974, n4973, 
        n4972, n4971, n4970, n9482, n4969, n4967, n4946, n4945, 
        n4944, n4943, n4942, n4941, n4940, n4939, n4938, n4937, 
        n4936, n4935, n4934, n4933, n4932, n4929, n4928, n4927, 
        n4926, n4925, n4924, n4923, n4922, n8776, n4921, n4920, 
        n4919, n4918, n4917, n4916, n4915, n4914, n4913, n4912, 
        n4911, n4910, n4909, n4908, n4907, n4906, n4905, n4904, 
        n4903, n4902, n4901, n4900, n4899, n4898, n4897, n4896, 
        n4895, n4894, n4893, n4892, n4891, n4890, n8775, n4889, 
        n4888, n4887, n4886, n4885, n4884, n4883, n4882, n4880, 
        n4879, n4878, n4877, n4876, n4875, n4874, n8774, n8773, 
        n8772, n8771, n8770, n4873, n4872, n4871, n4870, n4869, 
        n4868, n4867, n4866, n4865, n4864, n4863, n4862, n4861, 
        n4860, n4859, n4858, n8769, n8768, n8767, n4857, n4856, 
        n4855, n4854, n4853, n4852, n4851, n4850, n4849, n4848, 
        n4847, n4846, n4845, n4844, n4843, n4842, n8766, n8765, 
        n4841, n4840, n4839, n4838, n4837, n4836, n4835, n4834, 
        n4833, n4832, n4831, n4830, n4829, n4828, n4827, n4826, 
        n4825, n4824, n4823, n4822, n4821, n4820, n4819, n4818, 
        n4817, n4814, n4813, n4812, n4811, n4810, n4809, n4808, 
        n4807, n4806, n4805, n4804, n4803, n4802, n4801, n4800, 
        n4799, n4798, n4797, n4796, n4795, n4794, n4793, n4792, 
        n4791, n4790, n4789, n4788, n4787, n4786, n4785, n4784, 
        n4783, n4782, n4781, n4780, n4779, n4778, n4777, n4776, 
        n4775, n4774, n4773, n4772, n4771, n4770, n4769, n4768, 
        n4767, n4766, n4733, n4732, n4731, n4730, n4729, n4728, 
        n4727, n4726, n4725, n4724, n4723, n4722, n4721, n4720, 
        n4719, n4718, n8764, n4701, n4699, n12410, n4683, n4682, 
        n4681, n4680, n4679, n4678, n4677, n4676, n4675, n4674, 
        n4673, n4672, n4655, n4654, n4653, n4652, n4651, n4650, 
        n4649, n4648, n4647, n4646, n4645, n4644, n4643, n4642, 
        n4641, n4640, n4639, n4638, n4637, n4636, n4635, n4634, 
        n4633, n4631, n4629, n4627, n4626, n4625, n4624, n4623, 
        n4622, n4621, n4620, n4619, n4618, n4617, n4616, n8763, 
        n4615, n8762, n8824, n4614, n4613, n4612, n4611, n4610, 
        n4609, n4608, n4607, n4606, n4605, n4604, n4603, n4602, 
        n4601, n4600, n4599, n130, n129, n128, n127, n126, n125, 
        n124, n123, n122, n121, n120, n119, n118, n4598, n4597, 
        n4596, n117, n116, n115, n114, n113, n112, n111, n110, 
        n109, n108, n107, n106, n4579, n4578, n4577, n4576, 
        n4575, n4574, n4573, n4572, n4571, n4570, n4569, n4568, 
        n4567, n8761, n4566, n4565, n4564, n4563, n4562, n4561, 
        n4560, n4559, n4558, n4557, n4556, n4555, n4554, n4553, 
        n4552, n4551, n8760, n8759, n8661, n4550, n4549, n4548, 
        n4547, n4546, n4545, n4544, n4543, n4542, n4541, n4540, 
        n4539, n4538, n4537, n4536, n4535, n8758, n4534, n4533, 
        n4532, n4531, n4530, n4529, n4528, n4527, n4526, n4525, 
        n4524, n4523, n4522, n4521, n4520, n4519, n8757, n4518, 
        n4517, n4516, n4515, n4514, n4513, n4512, n4511, n4510, 
        n4509, n4508, n4507, n4506, n4505, n4504, n4503, n8756, 
        n25_adj_1106, n24_adj_1107, n23_adj_1108, n22_adj_1109, n21_adj_1110, 
        n20_adj_1111, n19_adj_1112, n4502, n4501, n4500, n4499, 
        n4498, n4497, n4496, n4495, n4494, n4493, n4492, n4491, 
        n4490, n4489, n4488, n4487, n18_adj_1113, n17, n16, n15_adj_1114, 
        n14_adj_1115, n13, n12_adj_1116, n11_adj_1117, n10_adj_1118, 
        n9_adj_1119, n8_adj_1120, n7_adj_1121, n6, n5_adj_1122, n4_adj_1123, 
        n3_adj_1124, n4486, n4485, n4484, n4483, n4482, n4481, 
        n4480, n4479, n4478, n4477, n4476, n4475, n4474, n4473, 
        n4472, n2, n25_adj_1125, n4455, n8755, n8754, n4454, n4453, 
        n4452, n4451, n4450, n4449, n4448, n4447, n4446, n4445, 
        n4444, n4443, n4442, n4441, n4440, n4439, n4438, n4437, 
        n4436, n4435, n4434, n4433, n4432, n4431, n4430, n4429, 
        n4099, n4098, n4096, n4093, n4091, n4428, n4427, n4426, 
        n4425, n4424, n8753, n4391, n4390, n4389, n4388, n4387, 
        n4386, n4385, n4384, n4383, n4382, n4381, n4380, n4379, 
        n4378, n4377, n4376, n4375, n4374, n4373, n4372, n4371, 
        n4370, n4369, n4368, n4367, n4366, n4365, n4364, n4363, 
        n4362, n4361, n4360, n4359, n4358, n4357, n4356, n4355, 
        n4090, n4089, n4086, n4082, n4081, n4354, n4353, n4352, 
        n4351, n4350, n4349, n4348, n4347, n4346, n4345, n4344, 
        n4343, n4342, n4341, n4340, n4339, n4338, n4337, n4336, 
        n4335, n4334, n4333, n4332, n4331, n4330, n4329, n4328, 
        n4327, n4326, n4325, n4324, n4323, n9440, n4322, n4321, 
        n4320, n4319, n4318, n4317, n4316, n4315, n4314, n4313, 
        n4312, n4311, n4310, n4309, n4308, n4307, n4306, n4305, 
        n4304, n4303, n4302, n4301, n4300, n4299, n4298, n4297, 
        n4296, n4295, n4294, n4293, n4292, n4291, n4290, n4289, 
        n4288, n4287, n4286, n4285, n4284, n4283, n4282, n4281, 
        n4080, n4079, n4073, n4280, n4279, n4278, n4277, n4276, 
        n4275, n4274, n4273, n4272, n4270, n4268, n4265, n4264, 
        n4263, n4262, n4261, n4260, n4259, n4258, n4257, n4256, 
        n4255, n4254, n4253, n4252, n4251, n4250, n4249, n4_adj_1126, 
        n9073, n4248, n4247, n4246, n4245, n4244, n4243, n4242, 
        n4241, n4240, n4239, n4238, n4237, n9398, n4236, n4235, 
        n4234, n4233, n4232, n4231, n4230, n4229, n4228, n4227, 
        n4226, n4225, n4224, n4223, n9406, n4222, n4221, n4220, 
        n4219, n4218, n4217, n4216, n4215, n4214, n4213, n4212, 
        n4211, n4210, n4209, n4208, n4207, n4206, n4205, n3642, 
        n6392, n4204, n4203, n4202, n3629, n3626, n3935, n4_adj_1127, 
        n9057, n8863, n8861, n8859, n1, n3474;
    
    VCC i2 (.Y(VCC_net));
    timing_controller timing_controller_inst (.state({state}), .DEBUG_6_c(DEBUG_6_c), 
            .\num_words_in_buffer[4] (num_words_in_buffer[4]), .\num_words_in_buffer[6] (num_words_in_buffer[6]), 
            .\num_words_in_buffer[5] (num_words_in_buffer[5]), .\num_words_in_buffer[3] (num_words_in_buffer[3]), 
            .DEBUG_2_c(DEBUG_2_c), .n9057(n9057), .buffer_switch_done(buffer_switch_done), 
            .n63(n63_adj_1105), .GND_net(GND_net), .n9355(n9355), .VCC_net(VCC_net), 
            .n1326(n1326), .n1431(n1431), .n6392(n6392), .n6602(n6602), 
            .n6572(n6572), .n3474(n3474), .INVERT_c_3(INVERT_c_3), .reset_all(reset_all), 
            .UPDATE_c_2(UPDATE_c_2)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(507[19] 518[2])
    SB_LUT4 i3705_3_lut (.I0(\REG.mem_38_12 ), .I1(FIFO_D12_c_12), .I2(n27), 
            .I3(GND_net), .O(n4794));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3706_3_lut (.I0(\REG.mem_38_13 ), .I1(FIFO_D13_c_13), .I2(n27), 
            .I3(GND_net), .O(n4795));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3707_3_lut (.I0(\REG.mem_38_14 ), .I1(FIFO_D14_c_14), .I2(n27), 
            .I3(GND_net), .O(n4796));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3560_3_lut (.I0(\REG.mem_30_15 ), .I1(FIFO_D15_c_15), .I2(n35), 
            .I3(GND_net), .O(n4649));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3561_2_lut (.I0(reset_all), .I1(rp_sync1_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n4650));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3561_2_lut.LUT_INIT = 16'h4444;
    bluejay_data bluejay_data_inst (.DEBUG_6_c(DEBUG_6_c), .GND_net(GND_net), 
            .DEBUG_9_c(DEBUG_9_c), .DEBUG_3_c(DEBUG_3_c), .buffer_switch_done(buffer_switch_done), 
            .DEBUG_2_c(DEBUG_2_c), .DEBUG_5_c(DEBUG_5_c), .VCC_net(VCC_net), 
            .DATA15_c(DATA15_c), .DATA14_c(DATA14_c), .DATA13_c(DATA13_c), 
            .DATA12_c(DATA12_c), .DATA11_c(DATA11_c), .DATA10_c(DATA10_c), 
            .DATA9_c(DATA9_c), .DATA8_c(DATA8_c), .DATA7_c(DATA7_c), .DATA6_c(DATA6_c), 
            .DATA5_c(DATA5_c), .DATA20_c(DATA20_c), .DATA19_c(DATA19_c), 
            .DATA18_c(DATA18_c), .\fifo_data_out[1] (fifo_data_out[1]), 
            .\fifo_data_out[2] (fifo_data_out[2]), .\fifo_data_out[0] (fifo_data_out[0]), 
            .\fifo_data_out[5] (fifo_data_out[5]), .\fifo_data_out[6] (fifo_data_out[6]), 
            .\fifo_data_out[7] (fifo_data_out[7]), .\fifo_data_out[8] (fifo_data_out[8]), 
            .\fifo_data_out[9] (fifo_data_out[9]), .\fifo_data_out[10] (fifo_data_out[10]), 
            .\fifo_data_out[11] (fifo_data_out[11]), .\fifo_data_out[12] (fifo_data_out[12]), 
            .\fifo_data_out[13] (fifo_data_out[13]), .\fifo_data_out[14] (fifo_data_out[14]), 
            .\fifo_data_out[15] (fifo_data_out[15]), .\fifo_data_out[3] (fifo_data_out[3]), 
            .\fifo_data_out[4] (fifo_data_out[4]), .DATA17_c(DATA17_c)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(584[14] 597[2])
    SB_DFF uart_rx_complete_prev_81 (.Q(uart_rx_complete_prev), .C(DEBUG_6_c), 
           .D(debug_led3));   // src/top.v(1023[8] 1029[4])
    SB_GB clk_gb (.GLOBAL_BUFFER_OUTPUT(DEBUG_6_c), .USER_SIGNAL_TO_GLOBAL_BUFFER(pll_clk_unbuf)) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/clock.v(82[7:96])
    SB_LUT4 i3708_3_lut (.I0(\REG.mem_38_15 ), .I1(FIFO_D15_c_15), .I2(n27), 
            .I3(GND_net), .O(n4797));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3709_3_lut (.I0(\REG.mem_39_0 ), .I1(FIFO_D0_c_0), .I2(n26), 
            .I3(GND_net), .O(n4798));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3709_3_lut.LUT_INIT = 16'hcaca;
    SB_IO UART_TX_pad (.PACKAGE_PIN(UART_TX), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UART_TX_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_TX_pad.PIN_TYPE = 6'b011001;
    defparam UART_TX_pad.PULLUP = 1'b0;
    defparam UART_TX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_TX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i3710_3_lut (.I0(\REG.mem_39_1 ), .I1(FIFO_D1_c_1), .I2(n26), 
            .I3(GND_net), .O(n4799));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3711_3_lut (.I0(\REG.mem_39_2 ), .I1(FIFO_D2_c_2), .I2(n26), 
            .I3(GND_net), .O(n4800));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3712_3_lut (.I0(\REG.mem_39_3 ), .I1(FIFO_D3_c_3), .I2(n26), 
            .I3(GND_net), .O(n4801));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3713_3_lut (.I0(\REG.mem_39_4 ), .I1(FIFO_D4_c_4), .I2(n26), 
            .I3(GND_net), .O(n4802));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3724_3_lut (.I0(\REG.mem_39_15 ), .I1(FIFO_D15_c_15), .I2(n26), 
            .I3(GND_net), .O(n4813));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3714_3_lut (.I0(\REG.mem_39_5 ), .I1(FIFO_D5_c_5), .I2(n26), 
            .I3(GND_net), .O(n4803));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3715_3_lut (.I0(\REG.mem_39_6 ), .I1(FIFO_D6_c_6), .I2(n26), 
            .I3(GND_net), .O(n4804));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3716_3_lut (.I0(\REG.mem_39_7 ), .I1(FIFO_D7_c_7), .I2(n26), 
            .I3(GND_net), .O(n4805));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3717_3_lut (.I0(\REG.mem_39_8 ), .I1(FIFO_D8_c_8), .I2(n26), 
            .I3(GND_net), .O(n4806));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3718_3_lut (.I0(\REG.mem_39_9 ), .I1(FIFO_D9_c_9), .I2(n26), 
            .I3(GND_net), .O(n4807));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3562_2_lut (.I0(reset_all), .I1(rp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n4651));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3562_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3719_3_lut (.I0(\REG.mem_39_10 ), .I1(FIFO_D10_c_10), .I2(n26), 
            .I3(GND_net), .O(n4808));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3720_3_lut (.I0(\REG.mem_39_11 ), .I1(FIFO_D11_c_11), .I2(n26), 
            .I3(GND_net), .O(n4809));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3721_3_lut (.I0(\REG.mem_39_12 ), .I1(FIFO_D12_c_12), .I2(n26), 
            .I3(GND_net), .O(n4810));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3722_3_lut (.I0(\REG.mem_39_13 ), .I1(FIFO_D13_c_13), .I2(n26), 
            .I3(GND_net), .O(n4811));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3563_2_lut (.I0(reset_all), .I1(rp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4652));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3563_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3564_2_lut (.I0(reset_all), .I1(rp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n4653));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3564_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3565_2_lut (.I0(reset_all), .I1(rp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4654));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3565_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3566_2_lut (.I0(reset_all), .I1(rp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n4655));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3566_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3725_3_lut (.I0(\REG.mem_40_0 ), .I1(FIFO_D0_c_0), .I2(n25), 
            .I3(GND_net), .O(n4814));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3728_3_lut (.I0(\REG.mem_40_1 ), .I1(FIFO_D1_c_1), .I2(n25), 
            .I3(GND_net), .O(n4817));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3729_3_lut (.I0(\REG.mem_40_2 ), .I1(FIFO_D2_c_2), .I2(n25), 
            .I3(GND_net), .O(n4818));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3730_3_lut (.I0(\REG.mem_40_3 ), .I1(FIFO_D3_c_3), .I2(n25), 
            .I3(GND_net), .O(n4819));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3731_3_lut (.I0(\REG.mem_40_4 ), .I1(FIFO_D4_c_4), .I2(n25), 
            .I3(GND_net), .O(n4820));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4103_3_lut (.I0(\REG.mem_61_15 ), .I1(FIFO_D15_c_15), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5192));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3732_3_lut (.I0(\REG.mem_40_5 ), .I1(FIFO_D5_c_5), .I2(n25), 
            .I3(GND_net), .O(n4821));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3733_3_lut (.I0(\REG.mem_40_6 ), .I1(FIFO_D6_c_6), .I2(n25), 
            .I3(GND_net), .O(n4822));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3733_3_lut.LUT_INIT = 16'hcaca;
    SB_IO RST_pad (.PACKAGE_PIN(RST), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RST_pad.PIN_TYPE = 6'b011001;
    defparam RST_pad.PULLUP = 1'b0;
    defparam RST_pad.NEG_TRIGGER = 1'b0;
    defparam RST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i3734_3_lut (.I0(\REG.mem_40_7 ), .I1(FIFO_D7_c_7), .I2(n25), 
            .I3(GND_net), .O(n4823));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3735_3_lut (.I0(\REG.mem_40_8 ), .I1(FIFO_D8_c_8), .I2(n25), 
            .I3(GND_net), .O(n4824));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4104_3_lut (.I0(\REG.mem_62_0 ), .I1(FIFO_D0_c_0), .I2(n3), 
            .I3(GND_net), .O(n5193));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3736_3_lut (.I0(\REG.mem_40_9 ), .I1(FIFO_D9_c_9), .I2(n25), 
            .I3(GND_net), .O(n4825));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3737_3_lut (.I0(\REG.mem_40_10 ), .I1(FIFO_D10_c_10), .I2(n25), 
            .I3(GND_net), .O(n4826));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3738_3_lut (.I0(\REG.mem_40_11 ), .I1(FIFO_D11_c_11), .I2(n25), 
            .I3(GND_net), .O(n4827));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3739_3_lut (.I0(\REG.mem_40_12 ), .I1(FIFO_D12_c_12), .I2(n25), 
            .I3(GND_net), .O(n4828));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3740_3_lut (.I0(\REG.mem_40_13 ), .I1(FIFO_D13_c_13), .I2(n25), 
            .I3(GND_net), .O(n4829));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3741_3_lut (.I0(\REG.mem_40_14 ), .I1(FIFO_D14_c_14), .I2(n25), 
            .I3(GND_net), .O(n4830));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4105_3_lut (.I0(\REG.mem_62_1 ), .I1(FIFO_D1_c_1), .I2(n3), 
            .I3(GND_net), .O(n5194));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4106_3_lut (.I0(\REG.mem_62_2 ), .I1(FIFO_D2_c_2), .I2(n3), 
            .I3(GND_net), .O(n5195));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4107_3_lut (.I0(\REG.mem_62_3 ), .I1(FIFO_D3_c_3), .I2(n3), 
            .I3(GND_net), .O(n5196));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3742_3_lut (.I0(\REG.mem_40_15 ), .I1(FIFO_D15_c_15), .I2(n25), 
            .I3(GND_net), .O(n4831));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3068_3_lut (.I0(\REG.mem_2_3 ), .I1(FIFO_D3_c_3), .I2(n63), 
            .I3(GND_net), .O(n4157));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3743_3_lut (.I0(\REG.mem_41_0 ), .I1(FIFO_D0_c_0), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4832));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4108_3_lut (.I0(\REG.mem_62_4 ), .I1(FIFO_D4_c_4), .I2(n3), 
            .I3(GND_net), .O(n5197));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4109_3_lut (.I0(\REG.mem_62_5 ), .I1(FIFO_D5_c_5), .I2(n3), 
            .I3(GND_net), .O(n5198));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3744_3_lut (.I0(\REG.mem_41_1 ), .I1(FIFO_D1_c_1), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4833));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3745_3_lut (.I0(\REG.mem_41_2 ), .I1(FIFO_D2_c_2), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4834));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4238_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [0]), 
            .I3(fifo_data_out[0]), .O(n5327));
    defparam i4238_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4216_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [15]), 
            .I3(fifo_data_out[15]), .O(n5305));
    defparam i4216_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3746_3_lut (.I0(\REG.mem_41_3 ), .I1(FIFO_D3_c_3), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4835));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3747_3_lut (.I0(\REG.mem_41_4 ), .I1(FIFO_D4_c_4), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4836));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4110_3_lut (.I0(\REG.mem_62_6 ), .I1(FIFO_D6_c_6), .I2(n3), 
            .I3(GND_net), .O(n5199));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3748_3_lut (.I0(\REG.mem_41_5 ), .I1(FIFO_D5_c_5), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4837));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4213_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [14]), 
            .I3(fifo_data_out[14]), .O(n5302));
    defparam i4213_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3749_3_lut (.I0(\REG.mem_41_6 ), .I1(FIFO_D6_c_6), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4838));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3750_3_lut (.I0(\REG.mem_41_7 ), .I1(FIFO_D7_c_7), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4839));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3751_3_lut (.I0(\REG.mem_41_8 ), .I1(FIFO_D8_c_8), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4840));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3752_3_lut (.I0(\REG.mem_41_9 ), .I1(FIFO_D9_c_9), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4841));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3753_3_lut (.I0(\REG.mem_41_10 ), .I1(FIFO_D10_c_10), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4842));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3754_3_lut (.I0(\REG.mem_41_11 ), .I1(FIFO_D11_c_11), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4843));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3755_3_lut (.I0(\REG.mem_41_12 ), .I1(FIFO_D12_c_12), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4844));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3756_3_lut (.I0(\REG.mem_41_13 ), .I1(FIFO_D13_c_13), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4845));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4210_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [13]), 
            .I3(fifo_data_out[13]), .O(n5299));
    defparam i4210_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3757_3_lut (.I0(\REG.mem_41_14 ), .I1(FIFO_D14_c_14), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4846));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4207_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [12]), 
            .I3(fifo_data_out[12]), .O(n5296));
    defparam i4207_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4111_3_lut (.I0(\REG.mem_62_7 ), .I1(FIFO_D7_c_7), .I2(n3), 
            .I3(GND_net), .O(n5200));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 reset_all_w_I_0_1_lut (.I0(reset_all_w), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(RESET_c));   // src/top.v(295[16:28])
    defparam reset_all_w_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4112_3_lut (.I0(\REG.mem_62_8 ), .I1(FIFO_D8_c_8), .I2(n3), 
            .I3(GND_net), .O(n5201));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4113_3_lut (.I0(\REG.mem_62_9 ), .I1(FIFO_D9_c_9), .I2(n3), 
            .I3(GND_net), .O(n5202));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4114_3_lut (.I0(\REG.mem_62_10 ), .I1(FIFO_D10_c_10), .I2(n3), 
            .I3(GND_net), .O(n5203));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4204_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [11]), 
            .I3(fifo_data_out[11]), .O(n5293));
    defparam i4204_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3758_3_lut (.I0(\REG.mem_41_15 ), .I1(FIFO_D15_c_15), .I2(n24_adj_1104), 
            .I3(GND_net), .O(n4847));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3758_3_lut.LUT_INIT = 16'hcaca;
    SB_IO CTS_pad (.PACKAGE_PIN(CTS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CTS_pad.PIN_TYPE = 6'b011001;
    defparam CTS_pad.PULLUP = 1'b0;
    defparam CTS_pad.NEG_TRIGGER = 1'b0;
    defparam CTS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4201_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [10]), 
            .I3(fifo_data_out[10]), .O(n5290));
    defparam i4201_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3759_3_lut (.I0(\REG.mem_42_0 ), .I1(FIFO_D0_c_0), .I2(n23), 
            .I3(GND_net), .O(n4848));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3760_3_lut (.I0(\REG.mem_42_1 ), .I1(FIFO_D1_c_1), .I2(n23), 
            .I3(GND_net), .O(n4849));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3761_3_lut (.I0(\REG.mem_42_2 ), .I1(FIFO_D2_c_2), .I2(n23), 
            .I3(GND_net), .O(n4850));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3762_3_lut (.I0(\REG.mem_42_3 ), .I1(FIFO_D3_c_3), .I2(n23), 
            .I3(GND_net), .O(n4851));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3763_3_lut (.I0(\REG.mem_42_4 ), .I1(FIFO_D4_c_4), .I2(n23), 
            .I3(GND_net), .O(n4852));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3764_3_lut (.I0(\REG.mem_42_5 ), .I1(FIFO_D5_c_5), .I2(n23), 
            .I3(GND_net), .O(n4853));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4115_3_lut (.I0(\REG.mem_62_11 ), .I1(FIFO_D11_c_11), .I2(n3), 
            .I3(GND_net), .O(n5204));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4116_3_lut (.I0(\REG.mem_62_12 ), .I1(FIFO_D12_c_12), .I2(n3), 
            .I3(GND_net), .O(n5205));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3765_3_lut (.I0(\REG.mem_42_6 ), .I1(FIFO_D6_c_6), .I2(n23), 
            .I3(GND_net), .O(n4854));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4166_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [9]), 
            .I3(fifo_data_out[9]), .O(n5255));
    defparam i4166_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3583_2_lut (.I0(reset_all), .I1(rd_addr_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n4672));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3583_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4117_3_lut (.I0(\REG.mem_62_13 ), .I1(FIFO_D13_c_13), .I2(n3), 
            .I3(GND_net), .O(n5206));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4118_3_lut (.I0(\REG.mem_62_14 ), .I1(FIFO_D14_c_14), .I2(n3), 
            .I3(GND_net), .O(n5207));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3766_3_lut (.I0(\REG.mem_42_7 ), .I1(FIFO_D7_c_7), .I2(n23), 
            .I3(GND_net), .O(n4855));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3767_3_lut (.I0(\REG.mem_42_8 ), .I1(FIFO_D8_c_8), .I2(n23), 
            .I3(GND_net), .O(n4856));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3584_2_lut (.I0(reset_all), .I1(rd_grey_sync_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n4673));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3584_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3768_3_lut (.I0(\REG.mem_42_9 ), .I1(FIFO_D9_c_9), .I2(n23), 
            .I3(GND_net), .O(n4857));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3769_3_lut (.I0(\REG.mem_42_10 ), .I1(FIFO_D10_c_10), .I2(n23), 
            .I3(GND_net), .O(n4858));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3770_3_lut (.I0(\REG.mem_42_11 ), .I1(FIFO_D11_c_11), .I2(n23), 
            .I3(GND_net), .O(n4859));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3771_3_lut (.I0(\REG.mem_42_12 ), .I1(FIFO_D12_c_12), .I2(n23), 
            .I3(GND_net), .O(n4860));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3772_3_lut (.I0(\REG.mem_42_13 ), .I1(FIFO_D13_c_13), .I2(n23), 
            .I3(GND_net), .O(n4861));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3773_3_lut (.I0(\REG.mem_42_14 ), .I1(FIFO_D14_c_14), .I2(n23), 
            .I3(GND_net), .O(n4862));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3774_3_lut (.I0(\REG.mem_42_15 ), .I1(FIFO_D15_c_15), .I2(n23), 
            .I3(GND_net), .O(n4863));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3775_3_lut (.I0(\REG.mem_43_0 ), .I1(FIFO_D0_c_0), .I2(n22), 
            .I3(GND_net), .O(n4864));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3776_3_lut (.I0(\REG.mem_43_1 ), .I1(FIFO_D1_c_1), .I2(n22), 
            .I3(GND_net), .O(n4865));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3777_3_lut (.I0(\REG.mem_43_2 ), .I1(FIFO_D2_c_2), .I2(n22), 
            .I3(GND_net), .O(n4866));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4119_3_lut (.I0(\REG.mem_62_15 ), .I1(FIFO_D15_c_15), .I2(n3), 
            .I3(GND_net), .O(n5208));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3778_3_lut (.I0(\REG.mem_43_3 ), .I1(FIFO_D3_c_3), .I2(n22), 
            .I3(GND_net), .O(n4867));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3779_3_lut (.I0(\REG.mem_43_4 ), .I1(FIFO_D4_c_4), .I2(n22), 
            .I3(GND_net), .O(n4868));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3779_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DTR_pad (.PACKAGE_PIN(DTR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DTR_pad.PIN_TYPE = 6'b011001;
    defparam DTR_pad.PULLUP = 1'b0;
    defparam DTR_pad.NEG_TRIGGER = 1'b0;
    defparam DTR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i3780_3_lut (.I0(\REG.mem_43_5 ), .I1(FIFO_D5_c_5), .I2(n22), 
            .I3(GND_net), .O(n4869));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3780_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DSR_pad (.PACKAGE_PIN(DSR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DSR_pad.PIN_TYPE = 6'b011001;
    defparam DSR_pad.PULLUP = 1'b0;
    defparam DSR_pad.NEG_TRIGGER = 1'b0;
    defparam DSR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i3781_3_lut (.I0(\REG.mem_43_6 ), .I1(FIFO_D6_c_6), .I2(n22), 
            .I3(GND_net), .O(n4870));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4163_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [8]), 
            .I3(fifo_data_out[8]), .O(n5252));
    defparam i4163_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_IO DCD_pad (.PACKAGE_PIN(DCD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DCD_pad.PIN_TYPE = 6'b011001;
    defparam DCD_pad.PULLUP = 1'b0;
    defparam DCD_pad.NEG_TRIGGER = 1'b0;
    defparam DCD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i3782_3_lut (.I0(\REG.mem_43_7 ), .I1(FIFO_D7_c_7), .I2(n22), 
            .I3(GND_net), .O(n4871));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3783_3_lut (.I0(\REG.mem_43_8 ), .I1(FIFO_D8_c_8), .I2(n22), 
            .I3(GND_net), .O(n4872));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3585_2_lut (.I0(reset_all), .I1(rd_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4674));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3585_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3784_3_lut (.I0(\REG.mem_43_9 ), .I1(FIFO_D9_c_9), .I2(n22), 
            .I3(GND_net), .O(n4873));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3785_3_lut (.I0(\REG.mem_43_10 ), .I1(FIFO_D10_c_10), .I2(n22), 
            .I3(GND_net), .O(n4874));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4160_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [7]), 
            .I3(fifo_data_out[7]), .O(n5249));
    defparam i4160_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4147_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [6]), 
            .I3(fifo_data_out[6]), .O(n5236));
    defparam i4147_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_IO FIFO_D0_pad (.PACKAGE_PIN(FIFO_D0), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D0_c_0));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D0_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D0_pad.PULLUP = 1'b0;
    defparam FIFO_D0_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i3786_3_lut (.I0(\REG.mem_43_11 ), .I1(FIFO_D11_c_11), .I2(n22), 
            .I3(GND_net), .O(n4875));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3787_3_lut (.I0(\REG.mem_43_12 ), .I1(FIFO_D12_c_12), .I2(n22), 
            .I3(GND_net), .O(n4876));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3788_3_lut (.I0(\REG.mem_43_13 ), .I1(FIFO_D13_c_13), .I2(n22), 
            .I3(GND_net), .O(n4877));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3789_3_lut (.I0(\REG.mem_43_14 ), .I1(FIFO_D14_c_14), .I2(n22), 
            .I3(GND_net), .O(n4878));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3586_2_lut (.I0(reset_all), .I1(rd_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n4675));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3586_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4144_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [5]), 
            .I3(fifo_data_out[5]), .O(n5233));
    defparam i4144_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3790_3_lut (.I0(\REG.mem_43_15 ), .I1(FIFO_D15_c_15), .I2(n22), 
            .I3(GND_net), .O(n4879));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3791_3_lut (.I0(\REG.mem_44_0 ), .I1(FIFO_D0_c_0), .I2(n21), 
            .I3(GND_net), .O(n4880));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4141_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [4]), 
            .I3(fifo_data_out[4]), .O(n5230));
    defparam i4141_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3793_3_lut (.I0(\REG.mem_44_1 ), .I1(FIFO_D1_c_1), .I2(n21), 
            .I3(GND_net), .O(n4882));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3794_3_lut (.I0(\REG.mem_44_2 ), .I1(FIFO_D2_c_2), .I2(n21), 
            .I3(GND_net), .O(n4883));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3795_3_lut (.I0(\REG.mem_44_3 ), .I1(FIFO_D3_c_3), .I2(n21), 
            .I3(GND_net), .O(n4884));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3796_3_lut (.I0(\REG.mem_44_4 ), .I1(FIFO_D4_c_4), .I2(n21), 
            .I3(GND_net), .O(n4885));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3797_3_lut (.I0(\REG.mem_44_5 ), .I1(FIFO_D5_c_5), .I2(n21), 
            .I3(GND_net), .O(n4886));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3798_3_lut (.I0(\REG.mem_44_6 ), .I1(FIFO_D6_c_6), .I2(n21), 
            .I3(GND_net), .O(n4887));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3798_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_936_1013__i0 (.Q(n25_adj_1106), .C(DEBUG_6_c), .D(n130));   // src/top.v(203[20:35])
    SB_LUT4 i3799_3_lut (.I0(\REG.mem_44_7 ), .I1(FIFO_D7_c_7), .I2(n21), 
            .I3(GND_net), .O(n4888));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3800_3_lut (.I0(\REG.mem_44_8 ), .I1(FIFO_D8_c_8), .I2(n21), 
            .I3(GND_net), .O(n4889));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3801_3_lut (.I0(\REG.mem_44_9 ), .I1(FIFO_D9_c_9), .I2(n21), 
            .I3(GND_net), .O(n4890));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3802_3_lut (.I0(\REG.mem_44_10 ), .I1(FIFO_D10_c_10), .I2(n21), 
            .I3(GND_net), .O(n4891));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3803_3_lut (.I0(\REG.mem_44_11 ), .I1(FIFO_D11_c_11), .I2(n21), 
            .I3(GND_net), .O(n4892));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3804_3_lut (.I0(\REG.mem_44_12 ), .I1(FIFO_D12_c_12), .I2(n21), 
            .I3(GND_net), .O(n4893));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3805_3_lut (.I0(\REG.mem_44_13 ), .I1(FIFO_D13_c_13), .I2(n21), 
            .I3(GND_net), .O(n4894));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4123_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [3]), 
            .I3(fifo_data_out[3]), .O(n5212));
    defparam i4123_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3587_2_lut (.I0(reset_all), .I1(rd_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4676));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3587_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3806_3_lut (.I0(\REG.mem_44_14 ), .I1(FIFO_D14_c_14), .I2(n21), 
            .I3(GND_net), .O(n4895));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4024_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [2]), 
            .I3(fifo_data_out[2]), .O(n5113));
    defparam i4024_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4005_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [1]), 
            .I3(fifo_data_out[1]), .O(n5094));
    defparam i4005_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3807_3_lut (.I0(\REG.mem_44_15 ), .I1(FIFO_D15_c_15), .I2(n21), 
            .I3(GND_net), .O(n4896));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3808_3_lut (.I0(\REG.mem_45_0 ), .I1(FIFO_D0_c_0), .I2(n20), 
            .I3(GND_net), .O(n4897));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3809_3_lut (.I0(\REG.mem_45_1 ), .I1(FIFO_D1_c_1), .I2(n20), 
            .I3(GND_net), .O(n4898));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3810_3_lut (.I0(\REG.mem_45_2 ), .I1(FIFO_D2_c_2), .I2(n20), 
            .I3(GND_net), .O(n4899));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3811_3_lut (.I0(\REG.mem_45_3 ), .I1(FIFO_D3_c_3), .I2(n20), 
            .I3(GND_net), .O(n4900));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3812_3_lut (.I0(\REG.mem_45_4 ), .I1(FIFO_D4_c_4), .I2(n20), 
            .I3(GND_net), .O(n4901));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3813_3_lut (.I0(\REG.mem_45_5 ), .I1(FIFO_D5_c_5), .I2(n20), 
            .I3(GND_net), .O(n4902));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3814_3_lut (.I0(\REG.mem_45_6 ), .I1(FIFO_D6_c_6), .I2(n20), 
            .I3(GND_net), .O(n4903));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3815_3_lut (.I0(\REG.mem_45_7 ), .I1(FIFO_D7_c_7), .I2(n20), 
            .I3(GND_net), .O(n4904));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3558_3_lut (.I0(\REG.mem_30_13 ), .I1(FIFO_D13_c_13), .I2(n35), 
            .I3(GND_net), .O(n4647));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3816_3_lut (.I0(\REG.mem_45_8 ), .I1(FIFO_D8_c_8), .I2(n20), 
            .I3(GND_net), .O(n4905));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3817_3_lut (.I0(\REG.mem_45_9 ), .I1(FIFO_D9_c_9), .I2(n20), 
            .I3(GND_net), .O(n4906));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3818_3_lut (.I0(\REG.mem_45_10 ), .I1(FIFO_D10_c_10), .I2(n20), 
            .I3(GND_net), .O(n4907));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3819_3_lut (.I0(\REG.mem_45_11 ), .I1(FIFO_D11_c_11), .I2(n20), 
            .I3(GND_net), .O(n4908));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3820_3_lut (.I0(\REG.mem_45_12 ), .I1(FIFO_D12_c_12), .I2(n20), 
            .I3(GND_net), .O(n4909));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3821_3_lut (.I0(\REG.mem_45_13 ), .I1(FIFO_D13_c_13), .I2(n20), 
            .I3(GND_net), .O(n4910));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3822_3_lut (.I0(\REG.mem_45_14 ), .I1(FIFO_D14_c_14), .I2(n20), 
            .I3(GND_net), .O(n4911));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3823_3_lut (.I0(\REG.mem_45_15 ), .I1(FIFO_D15_c_15), .I2(n20), 
            .I3(GND_net), .O(n4912));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3824_3_lut (.I0(\REG.mem_46_0 ), .I1(FIFO_D0_c_0), .I2(n19), 
            .I3(GND_net), .O(n4913));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3825_3_lut (.I0(\REG.mem_46_1 ), .I1(FIFO_D1_c_1), .I2(n19), 
            .I3(GND_net), .O(n4914));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3826_3_lut (.I0(\REG.mem_46_2 ), .I1(FIFO_D2_c_2), .I2(n19), 
            .I3(GND_net), .O(n4915));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3827_3_lut (.I0(\REG.mem_46_3 ), .I1(FIFO_D3_c_3), .I2(n19), 
            .I3(GND_net), .O(n4916));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3827_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_937__i3 (.Q(reset_clk_counter[3]), .C(DEBUG_6_c), 
           .D(n8863));   // src/top.v(259[27:51])
    SB_LUT4 i3828_3_lut (.I0(\REG.mem_46_4 ), .I1(FIFO_D4_c_4), .I2(n19), 
            .I3(GND_net), .O(n4917));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3829_3_lut (.I0(\REG.mem_46_5 ), .I1(FIFO_D5_c_5), .I2(n19), 
            .I3(GND_net), .O(n4918));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3830_3_lut (.I0(\REG.mem_46_6 ), .I1(FIFO_D6_c_6), .I2(n19), 
            .I3(GND_net), .O(n4919));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3831_3_lut (.I0(\REG.mem_46_7 ), .I1(FIFO_D7_c_7), .I2(n19), 
            .I3(GND_net), .O(n4920));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3832_3_lut (.I0(\REG.mem_46_8 ), .I1(FIFO_D8_c_8), .I2(n19), 
            .I3(GND_net), .O(n4921));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3833_3_lut (.I0(\REG.mem_46_9 ), .I1(FIFO_D9_c_9), .I2(n19), 
            .I3(GND_net), .O(n4922));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3834_3_lut (.I0(\REG.mem_46_10 ), .I1(FIFO_D10_c_10), .I2(n19), 
            .I3(GND_net), .O(n4923));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3835_3_lut (.I0(\REG.mem_46_11 ), .I1(FIFO_D11_c_11), .I2(n19), 
            .I3(GND_net), .O(n4924));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3836_3_lut (.I0(\REG.mem_46_12 ), .I1(FIFO_D12_c_12), .I2(n19), 
            .I3(GND_net), .O(n4925));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3837_3_lut (.I0(\REG.mem_46_13 ), .I1(FIFO_D13_c_13), .I2(n19), 
            .I3(GND_net), .O(n4926));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3838_3_lut (.I0(\REG.mem_46_14 ), .I1(FIFO_D14_c_14), .I2(n19), 
            .I3(GND_net), .O(n4927));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3838_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_937__i2 (.Q(reset_clk_counter[2]), .C(DEBUG_6_c), 
           .D(n8861));   // src/top.v(259[27:51])
    SB_DFF reset_clk_counter_i3_937__i1 (.Q(reset_clk_counter[1]), .C(DEBUG_6_c), 
           .D(n8859));   // src/top.v(259[27:51])
    SB_DFF led_counter_936_1013__i24 (.Q(DEBUG_0_c_24), .C(DEBUG_6_c), .D(n106));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i23 (.Q(n2), .C(DEBUG_6_c), .D(n107));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i22 (.Q(n3_adj_1124), .C(DEBUG_6_c), .D(n108));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i21 (.Q(n4_adj_1123), .C(DEBUG_6_c), .D(n109));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i20 (.Q(n5_adj_1122), .C(DEBUG_6_c), .D(n110));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i19 (.Q(n6), .C(DEBUG_6_c), .D(n111));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i18 (.Q(n7_adj_1121), .C(DEBUG_6_c), .D(n112));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i17 (.Q(n8_adj_1120), .C(DEBUG_6_c), .D(n113));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i16 (.Q(n9_adj_1119), .C(DEBUG_6_c), .D(n114));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i15 (.Q(n10_adj_1118), .C(DEBUG_6_c), .D(n115));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i14 (.Q(n11_adj_1117), .C(DEBUG_6_c), .D(n116));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i13 (.Q(n12_adj_1116), .C(DEBUG_6_c), .D(n117));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i12 (.Q(n13), .C(DEBUG_6_c), .D(n118));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i11 (.Q(n14_adj_1115), .C(DEBUG_6_c), .D(n119));   // src/top.v(203[20:35])
    SB_LUT4 i3054_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[7]), .I2(\mem_LUT.data_raw_r [7]), 
            .I3(n3734), .O(n4143));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3054_4_lut.LUT_INIT = 16'h5044;
    SB_DFF led_counter_936_1013__i10 (.Q(n15_adj_1114), .C(DEBUG_6_c), .D(n120));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i9 (.Q(n16), .C(DEBUG_6_c), .D(n121));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i8 (.Q(n17), .C(DEBUG_6_c), .D(n122));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i7 (.Q(n18_adj_1113), .C(DEBUG_6_c), .D(n123));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i6 (.Q(n19_adj_1112), .C(DEBUG_6_c), .D(n124));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i5 (.Q(n20_adj_1111), .C(DEBUG_6_c), .D(n125));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i4 (.Q(n21_adj_1110), .C(DEBUG_6_c), .D(n126));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i3 (.Q(n22_adj_1109), .C(DEBUG_6_c), .D(n127));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i2 (.Q(n23_adj_1108), .C(DEBUG_6_c), .D(n128));   // src/top.v(203[20:35])
    SB_DFF led_counter_936_1013__i1 (.Q(n24_adj_1107), .C(DEBUG_6_c), .D(n129));   // src/top.v(203[20:35])
    SB_LUT4 i3070_3_lut (.I0(\REG.mem_2_5 ), .I1(FIFO_D5_c_5), .I2(n63), 
            .I3(GND_net), .O(n4159));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3071_3_lut (.I0(\REG.mem_2_6 ), .I1(FIFO_D6_c_6), .I2(n63), 
            .I3(GND_net), .O(n4160));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3839_3_lut (.I0(\REG.mem_46_15 ), .I1(FIFO_D15_c_15), .I2(n19), 
            .I3(GND_net), .O(n4928));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3840_3_lut (.I0(\REG.mem_47_0 ), .I1(FIFO_D0_c_0), .I2(n18), 
            .I3(GND_net), .O(n4929));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3843_3_lut (.I0(\REG.mem_47_1 ), .I1(FIFO_D1_c_1), .I2(n18), 
            .I3(GND_net), .O(n4932));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3844_3_lut (.I0(\REG.mem_47_2 ), .I1(FIFO_D2_c_2), .I2(n18), 
            .I3(GND_net), .O(n4933));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3845_3_lut (.I0(\REG.mem_47_3 ), .I1(FIFO_D3_c_3), .I2(n18), 
            .I3(GND_net), .O(n4934));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3846_3_lut (.I0(\REG.mem_47_4 ), .I1(FIFO_D4_c_4), .I2(n18), 
            .I3(GND_net), .O(n4935));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3847_3_lut (.I0(\REG.mem_47_5 ), .I1(FIFO_D5_c_5), .I2(n18), 
            .I3(GND_net), .O(n4936));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3848_3_lut (.I0(\REG.mem_47_6 ), .I1(FIFO_D6_c_6), .I2(n18), 
            .I3(GND_net), .O(n4937));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3849_3_lut (.I0(\REG.mem_47_7 ), .I1(FIFO_D7_c_7), .I2(n18), 
            .I3(GND_net), .O(n4938));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4176_3_lut (.I0(tx_data_byte[2]), .I1(pc_data_rx[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5265));   // src/top.v(1032[8] 1094[4])
    defparam i4176_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF spi_start_transfer_r_82 (.Q(spi_start_transfer_r), .C(DEBUG_6_c), 
           .D(n2410));   // src/top.v(1032[8] 1094[4])
    SB_LUT4 i3850_3_lut (.I0(\REG.mem_47_8 ), .I1(FIFO_D8_c_8), .I2(n18), 
            .I3(GND_net), .O(n4939));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3851_3_lut (.I0(\REG.mem_47_9 ), .I1(FIFO_D9_c_9), .I2(n18), 
            .I3(GND_net), .O(n4940));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3852_3_lut (.I0(\REG.mem_47_10 ), .I1(FIFO_D10_c_10), .I2(n18), 
            .I3(GND_net), .O(n4941));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3853_3_lut (.I0(\REG.mem_47_11 ), .I1(FIFO_D11_c_11), .I2(n18), 
            .I3(GND_net), .O(n4942));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3854_3_lut (.I0(\REG.mem_47_12 ), .I1(FIFO_D12_c_12), .I2(n18), 
            .I3(GND_net), .O(n4943));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3854_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_data_byte_r_i0_i3 (.Q(tx_data_byte[3]), .C(DEBUG_6_c), .D(n5287));   // src/top.v(1032[8] 1094[4])
    SB_DFF tx_data_byte_r_i0_i4 (.Q(tx_data_byte[4]), .C(DEBUG_6_c), .D(n5286));   // src/top.v(1032[8] 1094[4])
    SB_DFF tx_data_byte_r_i0_i5 (.Q(tx_data_byte[5]), .C(DEBUG_6_c), .D(n5285));   // src/top.v(1032[8] 1094[4])
    SB_DFF tx_data_byte_r_i0_i6 (.Q(tx_data_byte[6]), .C(DEBUG_6_c), .D(n5276));   // src/top.v(1032[8] 1094[4])
    SB_DFF tx_data_byte_r_i0_i7 (.Q(tx_data_byte[7]), .C(DEBUG_6_c), .D(n5275));   // src/top.v(1032[8] 1094[4])
    SB_DFF tx_data_byte_r_i0_i1 (.Q(tx_data_byte[1]), .C(DEBUG_6_c), .D(n5274));   // src/top.v(1032[8] 1094[4])
    SB_LUT4 i4185_3_lut (.I0(tx_data_byte[1]), .I1(pc_data_rx[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5274));   // src/top.v(1032[8] 1094[4])
    defparam i4185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4186_3_lut (.I0(tx_data_byte[7]), .I1(pc_data_rx[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5275));   // src/top.v(1032[8] 1094[4])
    defparam i4186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4187_3_lut (.I0(tx_data_byte[6]), .I1(pc_data_rx[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5276));   // src/top.v(1032[8] 1094[4])
    defparam i4187_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_data_byte_r_i0_i2 (.Q(tx_data_byte[2]), .C(DEBUG_6_c), .D(n5265));   // src/top.v(1032[8] 1094[4])
    SB_LUT4 i3855_3_lut (.I0(\REG.mem_47_13 ), .I1(FIFO_D13_c_13), .I2(n18), 
            .I3(GND_net), .O(n4944));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4196_3_lut (.I0(tx_data_byte[5]), .I1(pc_data_rx[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5285));   // src/top.v(1032[8] 1094[4])
    defparam i4196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3856_3_lut (.I0(\REG.mem_47_14 ), .I1(FIFO_D14_c_14), .I2(n18), 
            .I3(GND_net), .O(n4945));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4197_3_lut (.I0(tx_data_byte[4]), .I1(pc_data_rx[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5286));   // src/top.v(1032[8] 1094[4])
    defparam i4197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4198_3_lut (.I0(tx_data_byte[3]), .I1(pc_data_rx[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5287));   // src/top.v(1032[8] 1094[4])
    defparam i4198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3857_3_lut (.I0(\REG.mem_47_15 ), .I1(FIFO_D15_c_15), .I2(n18), 
            .I3(GND_net), .O(n4946));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3040_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[6]), .I2(\mem_LUT.data_raw_r [6]), 
            .I3(n3734), .O(n4129));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3040_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i3034_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[5]), .I2(\mem_LUT.data_raw_r [5]), 
            .I3(n3734), .O(n4123));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3034_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i3022_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[4]), .I2(\mem_LUT.data_raw_r [4]), 
            .I3(n3734), .O(n4111));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3022_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i1337_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n2410));   // src/top.v(1032[8] 1094[4])
    defparam i1337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7858_4_lut (.I0(n1), .I1(fifo_read_cmd), .I2(wr_addr_r_adj_1162[1]), 
            .I3(rd_addr_r_adj_1165[1]), .O(n9398));
    defparam i7858_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i1_4_lut (.I0(reset_all_w), .I1(n15), .I2(full_nxt_r), .I3(n8824), 
            .O(n8987));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut.LUT_INIT = 16'h5444;
    SB_LUT4 i3878_3_lut (.I0(r_Tx_Data[7]), .I1(fifo_temp_output[7]), .I2(n3151), 
            .I3(GND_net), .O(n4967));   // src/uart_tx.v(38[10] 141[8])
    defparam i3878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4241_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[0]), .I2(\mem_LUT.data_raw_r [0]), 
            .I3(n3734), .O(n5330));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4241_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 led_counter_936_1013_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_1123), .I3(n8773), .O(n109)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3880_3_lut (.I0(r_Tx_Data[6]), .I1(fifo_temp_output[6]), .I2(n3151), 
            .I3(GND_net), .O(n4969));   // src/uart_tx.v(38[10] 141[8])
    defparam i3880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3881_3_lut (.I0(r_Tx_Data[5]), .I1(fifo_temp_output[5]), .I2(n3151), 
            .I3(GND_net), .O(n4970));   // src/uart_tx.v(38[10] 141[8])
    defparam i3881_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_936_1013_add_4_23 (.CI(n8773), .I0(GND_net), .I1(n4_adj_1123), 
            .CO(n8774));
    SB_LUT4 led_counter_936_1013_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_1122), .I3(n8772), .O(n110)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3882_3_lut (.I0(r_Tx_Data[4]), .I1(fifo_temp_output[4]), .I2(n3151), 
            .I3(GND_net), .O(n4971));   // src/uart_tx.v(38[10] 141[8])
    defparam i3882_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_936_1013_add_4_22 (.CI(n8772), .I0(GND_net), .I1(n5_adj_1122), 
            .CO(n8773));
    SB_LUT4 i3883_3_lut (.I0(r_Tx_Data[3]), .I1(fifo_temp_output[3]), .I2(n3151), 
            .I3(GND_net), .O(n4972));   // src/uart_tx.v(38[10] 141[8])
    defparam i3883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3884_3_lut (.I0(r_Tx_Data[2]), .I1(fifo_temp_output[2]), .I2(n3151), 
            .I3(GND_net), .O(n4973));   // src/uart_tx.v(38[10] 141[8])
    defparam i3884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_936_1013_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6), .I3(n8771), .O(n111)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3885_3_lut (.I0(r_Tx_Data[1]), .I1(fifo_temp_output[1]), .I2(n3151), 
            .I3(GND_net), .O(n4974));   // src/uart_tx.v(38[10] 141[8])
    defparam i3885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3072_3_lut (.I0(\REG.mem_2_7 ), .I1(FIFO_D7_c_7), .I2(n63), 
            .I3(GND_net), .O(n4161));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3073_3_lut (.I0(\REG.mem_2_8 ), .I1(FIFO_D8_c_8), .I2(n63), 
            .I3(GND_net), .O(n4162));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3069_3_lut (.I0(\REG.mem_2_4 ), .I1(FIFO_D4_c_4), .I2(n63), 
            .I3(GND_net), .O(n4158));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4248_4_lut (.I0(n3785), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(n131), .O(n5337));   // src/uart_rx.v(49[10] 144[8])
    defparam i4248_4_lut.LUT_INIT = 16'h4464;
    SB_LUT4 i4249_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[1]), .I2(n4), 
            .I3(n3525), .O(n5338));   // src/uart_rx.v(49[10] 144[8])
    defparam i4249_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4250_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[2]), .I2(n4_adj_1098), 
            .I3(n3533), .O(n5339));   // src/uart_rx.v(49[10] 144[8])
    defparam i4250_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY led_counter_936_1013_add_4_21 (.CI(n8771), .I0(GND_net), .I1(n6), 
            .CO(n8772));
    SB_LUT4 led_counter_936_1013_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_1121), .I3(n8770), .O(n112)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_936_1013_add_4_20 (.CI(n8770), .I0(GND_net), .I1(n7_adj_1121), 
            .CO(n8771));
    SB_LUT4 led_counter_936_1013_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_1120), .I3(n8769), .O(n113)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3007_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[3]), .I2(\mem_LUT.data_raw_r [3]), 
            .I3(n3734), .O(n4096));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3007_4_lut.LUT_INIT = 16'h5044;
    SB_CARRY led_counter_936_1013_add_4_19 (.CI(n8769), .I0(GND_net), .I1(n8_adj_1120), 
            .CO(n8770));
    SB_LUT4 led_counter_936_1013_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_1119), .I3(n8768), .O(n114)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_936_1013_add_4_18 (.CI(n8768), .I0(GND_net), .I1(n9_adj_1119), 
            .CO(n8769));
    SB_LUT4 led_counter_936_1013_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_1118), .I3(n8767), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_936_1013_add_4_17 (.CI(n8767), .I0(GND_net), .I1(n10_adj_1118), 
            .CO(n8768));
    SB_LUT4 i4255_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[0]), .I2(n4), 
            .I3(n3533), .O(n5344));   // src/uart_rx.v(49[10] 144[8])
    defparam i4255_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 led_counter_936_1013_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_1117), .I3(n8766), .O(n116)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_936_1013_add_4_16 (.CI(n8766), .I0(GND_net), .I1(n11_adj_1117), 
            .CO(n8767));
    SB_LUT4 i4256_3_lut (.I0(pc_data_rx[3]), .I1(r_Rx_Data), .I2(n9345), 
            .I3(GND_net), .O(n5345));   // src/uart_rx.v(49[10] 144[8])
    defparam i4256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4258_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[4]), .I2(n4_adj_1127), 
            .I3(n3533), .O(n5347));   // src/uart_rx.v(49[10] 144[8])
    defparam i4258_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i3588_2_lut (.I0(reset_all), .I1(rd_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n4677));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3588_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4259_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[5]), .I2(n4_adj_1127), 
            .I3(n3525), .O(n5348));   // src/uart_rx.v(49[10] 144[8])
    defparam i4259_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 led_counter_936_1013_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_1116), .I3(n8765), .O(n117)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_936_1013_add_4_15 (.CI(n8765), .I0(GND_net), .I1(n12_adj_1116), 
            .CO(n8766));
    SB_LUT4 led_counter_936_1013_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13), .I3(n8764), .O(n118)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_936_1013_add_4_14 (.CI(n8764), .I0(GND_net), .I1(n13), 
            .CO(n8765));
    SB_LUT4 led_counter_936_1013_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_1115), .I3(n8763), .O(n119)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_936_1013_add_4_13 (.CI(n8763), .I0(GND_net), .I1(n14_adj_1115), 
            .CO(n8764));
    SB_LUT4 led_counter_936_1013_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_1114), .I3(n8762), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4260_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[6]), .I2(n2414), 
            .I3(n3533), .O(n5349));   // src/uart_rx.v(49[10] 144[8])
    defparam i4260_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY led_counter_936_1013_add_4_12 (.CI(n8762), .I0(GND_net), .I1(n15_adj_1114), 
            .CO(n8763));
    SB_LUT4 led_counter_936_1013_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16), .I3(n8761), .O(n121)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_IO FIFO_D1_pad (.PACKAGE_PIN(FIFO_D1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D1_c_1));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D1_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D1_pad.PULLUP = 1'b0;
    defparam FIFO_D1_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D2_pad (.PACKAGE_PIN(FIFO_D2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D2_c_2));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D2_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D2_pad.PULLUP = 1'b0;
    defparam FIFO_D2_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D3_pad (.PACKAGE_PIN(FIFO_D3), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D3_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D3_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D3_pad.PULLUP = 1'b0;
    defparam FIFO_D3_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D4_pad (.PACKAGE_PIN(FIFO_D4), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D4_c_4));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D4_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D4_pad.PULLUP = 1'b0;
    defparam FIFO_D4_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_936_1013_add_4_11 (.CI(n8761), .I0(GND_net), .I1(n16), 
            .CO(n8762));
    SB_IO FIFO_D5_pad (.PACKAGE_PIN(FIFO_D5), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D5_c_5));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D5_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D5_pad.PULLUP = 1'b0;
    defparam FIFO_D5_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D6_pad (.PACKAGE_PIN(FIFO_D6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D6_c_6));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D6_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D6_pad.PULLUP = 1'b0;
    defparam FIFO_D6_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D7_pad (.PACKAGE_PIN(FIFO_D7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D7_c_7));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D7_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D7_pad.PULLUP = 1'b0;
    defparam FIFO_D7_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D8_pad (.PACKAGE_PIN(FIFO_D8), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D8_c_8));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D8_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D8_pad.PULLUP = 1'b0;
    defparam FIFO_D8_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D9_pad (.PACKAGE_PIN(FIFO_D9), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D9_c_9));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D9_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D9_pad.PULLUP = 1'b0;
    defparam FIFO_D9_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 led_counter_936_1013_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17), .I3(n8760), .O(n122)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_IO FIFO_D10_pad (.PACKAGE_PIN(FIFO_D10), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D10_c_10));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D10_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D10_pad.PULLUP = 1'b0;
    defparam FIFO_D10_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D11_pad (.PACKAGE_PIN(FIFO_D11), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D11_c_11));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D11_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D11_pad.PULLUP = 1'b0;
    defparam FIFO_D11_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D12_pad (.PACKAGE_PIN(FIFO_D12), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D12_c_12));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D12_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D12_pad.PULLUP = 1'b0;
    defparam FIFO_D12_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D13_pad (.PACKAGE_PIN(FIFO_D13), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D13_c_13));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D13_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D13_pad.PULLUP = 1'b0;
    defparam FIFO_D13_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_936_1013_add_4_10 (.CI(n8760), .I0(GND_net), .I1(n17), 
            .CO(n8761));
    SB_IO FIFO_D14_pad (.PACKAGE_PIN(FIFO_D14), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D14_c_14));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D14_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D14_pad.PULLUP = 1'b0;
    defparam FIFO_D14_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D15_pad (.PACKAGE_PIN(FIFO_D15), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D15_c_15));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D15_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D15_pad.PULLUP = 1'b0;
    defparam FIFO_D15_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO FIFO_CLK_pad (.PACKAGE_PIN(FIFO_CLK), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(FIFO_CLK_c));   // src/top.v(84[12:20])
    defparam FIFO_CLK_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_CLK_pad.PULLUP = 1'b0;
    defparam FIFO_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FR_RXF_pad (.PACKAGE_PIN(FR_RXF), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FR_RXF_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FR_RXF_pad.PIN_TYPE = 6'b000001;
    defparam FR_RXF_pad.PULLUP = 1'b0;
    defparam FR_RXF_pad.NEG_TRIGGER = 1'b0;
    defparam FR_RXF_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SOUT_pad (.PACKAGE_PIN(SOUT), .OUTPUT_ENABLE(VCC_net), .D_IN_0(SOUT_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SOUT_pad.PIN_TYPE = 6'b000001;
    defparam SOUT_pad.PULLUP = 1'b0;
    defparam SOUT_pad.NEG_TRIGGER = 1'b0;
    defparam SOUT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UART_RX_pad (.PACKAGE_PIN(UART_RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(UART_RX_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_RX_pad.PIN_TYPE = 6'b000001;
    defparam UART_RX_pad.PULLUP = 1'b0;
    defparam UART_RX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 led_counter_936_1013_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_1113), .I3(n8759), .O(n123)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_IO ICE_SYSCLK_pad (.PACKAGE_PIN(ICE_SYSCLK), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ICE_SYSCLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_SYSCLK_pad.PIN_TYPE = 6'b000001;
    defparam ICE_SYSCLK_pad.PULLUP = 1'b0;
    defparam ICE_SYSCLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_SYSCLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_936_1013_add_4_9 (.CI(n8759), .I0(GND_net), .I1(n18_adj_1113), 
            .CO(n8760));
    SB_IO ICE_CREST_pad (.PACKAGE_PIN(ICE_CREST), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CREST_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CREST_pad.PULLUP = 1'b0;
    defparam ICE_CREST_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CREST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CDONE_pad (.PACKAGE_PIN(ICE_CDONE), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CDONE_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CDONE_pad.PULLUP = 1'b0;
    defparam ICE_CDONE_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CDONE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i12_4_lut (.I0(tx_shift_reg[0]), .I1(n1638), .I2(n3626), .I3(tx_data_byte[0]), 
            .O(n9073));   // src/spi.v(76[8] 221[4])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_IO ICE_CLK_pad (.PACKAGE_PIN(ICE_CLK), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CLK_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CLK_pad.PULLUP = 1'b0;
    defparam ICE_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_9_pad (.PACKAGE_PIN(DEBUG_9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_9_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_9_pad.PULLUP = 1'b0;
    defparam DEBUG_9_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_8_pad (.PACKAGE_PIN(DEBUG_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_8_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_8_pad.PULLUP = 1'b0;
    defparam DEBUG_8_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_6_pad (.PACKAGE_PIN(DEBUG_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_6_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_6_pad.PULLUP = 1'b0;
    defparam DEBUG_6_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_5_pad (.PACKAGE_PIN(DEBUG_5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_5_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_5_pad.PULLUP = 1'b0;
    defparam DEBUG_5_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_3_pad (.PACKAGE_PIN(DEBUG_3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_3_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_3_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_3_pad.PULLUP = 1'b0;
    defparam DEBUG_3_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_2_pad (.PACKAGE_PIN(DEBUG_2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_2_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_2_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_2_pad.PULLUP = 1'b0;
    defparam DEBUG_2_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_1_pad (.PACKAGE_PIN(DEBUG_1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_1_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_1_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_1_pad.PULLUP = 1'b0;
    defparam DEBUG_1_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_0_pad (.PACKAGE_PIN(DEBUG_0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_0_c_24));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_0_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_0_pad.PULLUP = 1'b0;
    defparam DEBUG_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_SIWU_pad (.PACKAGE_PIN(FT_SIWU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_SIWU_pad.PIN_TYPE = 6'b011001;
    defparam FT_SIWU_pad.PULLUP = 1'b0;
    defparam FT_SIWU_pad.NEG_TRIGGER = 1'b0;
    defparam FT_SIWU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_WR_pad (.PACKAGE_PIN(FT_WR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_WR_pad.PIN_TYPE = 6'b011001;
    defparam FT_WR_pad.PULLUP = 1'b0;
    defparam FT_WR_pad.NEG_TRIGGER = 1'b0;
    defparam FT_WR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_RD_pad (.PACKAGE_PIN(FT_RD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_RD_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_RD_pad.PIN_TYPE = 6'b011001;
    defparam FT_RD_pad.PULLUP = 1'b0;
    defparam FT_RD_pad.NEG_TRIGGER = 1'b0;
    defparam FT_RD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_OE_pad (.PACKAGE_PIN(FT_OE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_OE_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_OE_pad.PIN_TYPE = 6'b011001;
    defparam FT_OE_pad.PULLUP = 1'b0;
    defparam FT_OE_pad.NEG_TRIGGER = 1'b0;
    defparam FT_OE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA10_pad (.PACKAGE_PIN(DATA10), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA10_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA10_pad.PIN_TYPE = 6'b011001;
    defparam DATA10_pad.PULLUP = 1'b0;
    defparam DATA10_pad.NEG_TRIGGER = 1'b0;
    defparam DATA10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA9_pad (.PACKAGE_PIN(DATA9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA9_pad.PIN_TYPE = 6'b011001;
    defparam DATA9_pad.PULLUP = 1'b0;
    defparam DATA9_pad.NEG_TRIGGER = 1'b0;
    defparam DATA9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA11_pad (.PACKAGE_PIN(DATA11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA11_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA11_pad.PIN_TYPE = 6'b011001;
    defparam DATA11_pad.PULLUP = 1'b0;
    defparam DATA11_pad.NEG_TRIGGER = 1'b0;
    defparam DATA11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA12_pad (.PACKAGE_PIN(DATA12), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA12_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA12_pad.PIN_TYPE = 6'b011001;
    defparam DATA12_pad.PULLUP = 1'b0;
    defparam DATA12_pad.NEG_TRIGGER = 1'b0;
    defparam DATA12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA13_pad (.PACKAGE_PIN(DATA13), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA13_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA13_pad.PIN_TYPE = 6'b011001;
    defparam DATA13_pad.PULLUP = 1'b0;
    defparam DATA13_pad.NEG_TRIGGER = 1'b0;
    defparam DATA13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4264_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[7]), .I2(n2414), 
            .I3(n3525), .O(n5353));   // src/uart_rx.v(49[10] 144[8])
    defparam i4264_4_lut.LUT_INIT = 16'hccac;
    SB_IO DATA14_pad (.PACKAGE_PIN(DATA14), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA14_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA14_pad.PIN_TYPE = 6'b011001;
    defparam DATA14_pad.PULLUP = 1'b0;
    defparam DATA14_pad.NEG_TRIGGER = 1'b0;
    defparam DATA14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA8_pad (.PACKAGE_PIN(DATA8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA8_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA8_pad.PIN_TYPE = 6'b011001;
    defparam DATA8_pad.PULLUP = 1'b0;
    defparam DATA8_pad.NEG_TRIGGER = 1'b0;
    defparam DATA8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA15_pad (.PACKAGE_PIN(DATA15), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA15_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA15_pad.PIN_TYPE = 6'b011001;
    defparam DATA15_pad.PULLUP = 1'b0;
    defparam DATA15_pad.NEG_TRIGGER = 1'b0;
    defparam DATA15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA16_pad (.PACKAGE_PIN(DATA16), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA16_pad.PIN_TYPE = 6'b011001;
    defparam DATA16_pad.PULLUP = 1'b0;
    defparam DATA16_pad.NEG_TRIGGER = 1'b0;
    defparam DATA16_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA7_pad (.PACKAGE_PIN(DATA7), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA7_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA7_pad.PIN_TYPE = 6'b011001;
    defparam DATA7_pad.PULLUP = 1'b0;
    defparam DATA7_pad.NEG_TRIGGER = 1'b0;
    defparam DATA7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA17_pad (.PACKAGE_PIN(DATA17), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA17_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA17_pad.PIN_TYPE = 6'b011001;
    defparam DATA17_pad.PULLUP = 1'b0;
    defparam DATA17_pad.NEG_TRIGGER = 1'b0;
    defparam DATA17_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA18_pad (.PACKAGE_PIN(DATA18), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA18_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA18_pad.PIN_TYPE = 6'b011001;
    defparam DATA18_pad.PULLUP = 1'b0;
    defparam DATA18_pad.NEG_TRIGGER = 1'b0;
    defparam DATA18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA6_pad (.PACKAGE_PIN(DATA6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA6_pad.PIN_TYPE = 6'b011001;
    defparam DATA6_pad.PULLUP = 1'b0;
    defparam DATA6_pad.NEG_TRIGGER = 1'b0;
    defparam DATA6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA19_pad (.PACKAGE_PIN(DATA19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA19_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA19_pad.PIN_TYPE = 6'b011001;
    defparam DATA19_pad.PULLUP = 1'b0;
    defparam DATA19_pad.NEG_TRIGGER = 1'b0;
    defparam DATA19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA20_pad (.PACKAGE_PIN(DATA20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA20_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA20_pad.PIN_TYPE = 6'b011001;
    defparam DATA20_pad.PULLUP = 1'b0;
    defparam DATA20_pad.NEG_TRIGGER = 1'b0;
    defparam DATA20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 led_counter_936_1013_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_1112), .I3(n8758), .O(n124)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_IO DATA5_pad (.PACKAGE_PIN(DATA5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA5_pad.PIN_TYPE = 6'b011001;
    defparam DATA5_pad.PULLUP = 1'b0;
    defparam DATA5_pad.NEG_TRIGGER = 1'b0;
    defparam DATA5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA21_pad (.PACKAGE_PIN(DATA21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA21_pad.PIN_TYPE = 6'b011001;
    defparam DATA21_pad.PULLUP = 1'b0;
    defparam DATA21_pad.NEG_TRIGGER = 1'b0;
    defparam DATA21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA22_pad (.PACKAGE_PIN(DATA22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA22_pad.PIN_TYPE = 6'b011001;
    defparam DATA22_pad.PULLUP = 1'b0;
    defparam DATA22_pad.NEG_TRIGGER = 1'b0;
    defparam DATA22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA4_pad (.PACKAGE_PIN(DATA4), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA20_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA4_pad.PIN_TYPE = 6'b011001;
    defparam DATA4_pad.PULLUP = 1'b0;
    defparam DATA4_pad.NEG_TRIGGER = 1'b0;
    defparam DATA4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA23_pad (.PACKAGE_PIN(DATA23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA7_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA23_pad.PIN_TYPE = 6'b011001;
    defparam DATA23_pad.PULLUP = 1'b0;
    defparam DATA23_pad.NEG_TRIGGER = 1'b0;
    defparam DATA23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA24_pad (.PACKAGE_PIN(DATA24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA8_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA24_pad.PIN_TYPE = 6'b011001;
    defparam DATA24_pad.PULLUP = 1'b0;
    defparam DATA24_pad.NEG_TRIGGER = 1'b0;
    defparam DATA24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i3000_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[2]), .I2(\mem_LUT.data_raw_r [2]), 
            .I3(n3734), .O(n4089));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i3000_4_lut.LUT_INIT = 16'h5044;
    SB_IO DATA3_pad (.PACKAGE_PIN(DATA3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA19_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA3_pad.PIN_TYPE = 6'b011001;
    defparam DATA3_pad.PULLUP = 1'b0;
    defparam DATA3_pad.NEG_TRIGGER = 1'b0;
    defparam DATA3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA25_pad (.PACKAGE_PIN(DATA25), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA25_pad.PIN_TYPE = 6'b011001;
    defparam DATA25_pad.PULLUP = 1'b0;
    defparam DATA25_pad.NEG_TRIGGER = 1'b0;
    defparam DATA25_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA26_pad (.PACKAGE_PIN(DATA26), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA10_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA26_pad.PIN_TYPE = 6'b011001;
    defparam DATA26_pad.PULLUP = 1'b0;
    defparam DATA26_pad.NEG_TRIGGER = 1'b0;
    defparam DATA26_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA2_pad (.PACKAGE_PIN(DATA2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA18_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA2_pad.PIN_TYPE = 6'b011001;
    defparam DATA2_pad.PULLUP = 1'b0;
    defparam DATA2_pad.NEG_TRIGGER = 1'b0;
    defparam DATA2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i2997_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[1]), .I2(\mem_LUT.data_raw_r [1]), 
            .I3(n3734), .O(n4086));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i2997_4_lut.LUT_INIT = 16'h5044;
    SB_IO DATA27_pad (.PACKAGE_PIN(DATA27), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA11_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA27_pad.PIN_TYPE = 6'b011001;
    defparam DATA27_pad.PULLUP = 1'b0;
    defparam DATA27_pad.NEG_TRIGGER = 1'b0;
    defparam DATA27_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA28_pad (.PACKAGE_PIN(DATA28), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA12_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA28_pad.PIN_TYPE = 6'b011001;
    defparam DATA28_pad.PULLUP = 1'b0;
    defparam DATA28_pad.NEG_TRIGGER = 1'b0;
    defparam DATA28_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA1_pad (.PACKAGE_PIN(DATA1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA17_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA1_pad.PIN_TYPE = 6'b011001;
    defparam DATA1_pad.PULLUP = 1'b0;
    defparam DATA1_pad.NEG_TRIGGER = 1'b0;
    defparam DATA1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA29_pad (.PACKAGE_PIN(DATA29), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA13_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA29_pad.PIN_TYPE = 6'b011001;
    defparam DATA29_pad.PULLUP = 1'b0;
    defparam DATA29_pad.NEG_TRIGGER = 1'b0;
    defparam DATA29_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA30_pad (.PACKAGE_PIN(DATA30), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA14_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA30_pad.PIN_TYPE = 6'b011001;
    defparam DATA30_pad.PULLUP = 1'b0;
    defparam DATA30_pad.NEG_TRIGGER = 1'b0;
    defparam DATA30_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA0_pad (.PACKAGE_PIN(DATA0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA0_pad.PIN_TYPE = 6'b011001;
    defparam DATA0_pad.PULLUP = 1'b0;
    defparam DATA0_pad.NEG_TRIGGER = 1'b0;
    defparam DATA0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA31_pad (.PACKAGE_PIN(DATA31), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA15_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA31_pad.PIN_TYPE = 6'b011001;
    defparam DATA31_pad.PULLUP = 1'b0;
    defparam DATA31_pad.NEG_TRIGGER = 1'b0;
    defparam DATA31_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO VALID_pad (.PACKAGE_PIN(VALID), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam VALID_pad.PIN_TYPE = 6'b011001;
    defparam VALID_pad.PULLUP = 1'b0;
    defparam VALID_pad.NEG_TRIGGER = 1'b0;
    defparam VALID_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SYNC_pad (.PACKAGE_PIN(SYNC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_3_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SYNC_pad.PIN_TYPE = 6'b011001;
    defparam SYNC_pad.PULLUP = 1'b0;
    defparam SYNC_pad.NEG_TRIGGER = 1'b0;
    defparam SYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INVERT_pad (.PACKAGE_PIN(INVERT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INVERT_c_3)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INVERT_pad.PIN_TYPE = 6'b011001;
    defparam INVERT_pad.PULLUP = 1'b0;
    defparam INVERT_pad.NEG_TRIGGER = 1'b0;
    defparam INVERT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SLM_CLK_pad (.PACKAGE_PIN(SLM_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SLM_CLK_pad.PIN_TYPE = 6'b011001;
    defparam SLM_CLK_pad.PULLUP = 1'b0;
    defparam SLM_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam SLM_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO RESET_pad (.PACKAGE_PIN(RESET), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(RESET_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RESET_pad.PIN_TYPE = 6'b011001;
    defparam RESET_pad.PULLUP = 1'b0;
    defparam RESET_pad.NEG_TRIGGER = 1'b0;
    defparam RESET_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UPDATE_pad (.PACKAGE_PIN(UPDATE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UPDATE_c_2));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UPDATE_pad.PIN_TYPE = 6'b011001;
    defparam UPDATE_pad.PULLUP = 1'b0;
    defparam UPDATE_pad.NEG_TRIGGER = 1'b0;
    defparam UPDATE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SDAT_pad (.PACKAGE_PIN(SDAT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SDAT_c_15)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SDAT_pad.PIN_TYPE = 6'b011001;
    defparam SDAT_pad.PULLUP = 1'b0;
    defparam SDAT_pad.NEG_TRIGGER = 1'b0;
    defparam SDAT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SCK_pad (.PACKAGE_PIN(SCK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SCK_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SCK_pad.PIN_TYPE = 6'b011001;
    defparam SCK_pad.PULLUP = 1'b0;
    defparam SCK_pad.NEG_TRIGGER = 1'b0;
    defparam SCK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SEN_pad (.PACKAGE_PIN(SEN), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SEN_c_1)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SEN_pad.PIN_TYPE = 6'b011001;
    defparam SEN_pad.PULLUP = 1'b0;
    defparam SEN_pad.NEG_TRIGGER = 1'b0;
    defparam SEN_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_936_1013_add_4_8 (.CI(n8758), .I0(GND_net), .I1(n19_adj_1112), 
            .CO(n8759));
    SB_LUT4 i3589_3_lut (.I0(rx_buf_byte[7]), .I1(rx_shift_reg[7]), .I2(n2851), 
            .I3(GND_net), .O(n4678));   // src/spi.v(76[8] 221[4])
    defparam i3589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19_4_lut (.I0(n3474), .I1(n10552), .I2(state[3]), .I3(n63_adj_1105), 
            .O(n9057));   // src/timing_controller.v(59[8] 133[4])
    defparam i19_4_lut.LUT_INIT = 16'hfcac;
    SB_LUT4 i3590_3_lut (.I0(rx_buf_byte[6]), .I1(rx_shift_reg[6]), .I2(n2851), 
            .I3(GND_net), .O(n4679));   // src/spi.v(76[8] 221[4])
    defparam i3590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 led_counter_936_1013_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_1111), .I3(n8757), .O(n125)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3591_3_lut (.I0(rx_buf_byte[5]), .I1(rx_shift_reg[5]), .I2(n2851), 
            .I3(GND_net), .O(n4680));   // src/spi.v(76[8] 221[4])
    defparam i3591_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY led_counter_936_1013_add_4_7 (.CI(n8757), .I0(GND_net), .I1(n20_adj_1111), 
            .CO(n8758));
    SB_LUT4 i3_4_lut (.I0(reset_clk_counter[0]), .I1(reset_clk_counter[2]), 
            .I2(reset_clk_counter[3]), .I3(reset_clk_counter[1]), .O(reset_all_w_N_61));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3592_3_lut (.I0(rx_buf_byte[4]), .I1(rx_shift_reg[4]), .I2(n2851), 
            .I3(GND_net), .O(n4681));   // src/spi.v(76[8] 221[4])
    defparam i3592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3903_3_lut (.I0(\REG.mem_50_0 ), .I1(FIFO_D0_c_0), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n4992));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3904_3_lut (.I0(\REG.mem_50_1 ), .I1(FIFO_D1_c_1), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n4993));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(reset_clk_counter[3]), .I1(reset_clk_counter[2]), 
            .I2(n8661), .I3(GND_net), .O(n8863));
    defparam i1_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i3593_3_lut (.I0(rx_buf_byte[3]), .I1(rx_shift_reg[3]), .I2(n2851), 
            .I3(GND_net), .O(n4682));   // src/spi.v(76[8] 221[4])
    defparam i3593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3074_3_lut (.I0(\REG.mem_2_9 ), .I1(FIFO_D9_c_9), .I2(n63), 
            .I3(GND_net), .O(n4163));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3075_3_lut (.I0(\REG.mem_2_10 ), .I1(FIFO_D10_c_10), .I2(n63), 
            .I3(GND_net), .O(n4164));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3594_3_lut (.I0(rx_buf_byte[2]), .I1(rx_shift_reg[2]), .I2(n2851), 
            .I3(GND_net), .O(n4683));   // src/spi.v(76[8] 221[4])
    defparam i3594_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3076_3_lut (.I0(\REG.mem_2_11 ), .I1(FIFO_D11_c_11), .I2(n63), 
            .I3(GND_net), .O(n4165));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3077_3_lut (.I0(\REG.mem_2_12 ), .I1(FIFO_D12_c_12), .I2(n63), 
            .I3(GND_net), .O(n4166));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3078_3_lut (.I0(\REG.mem_2_13 ), .I1(FIFO_D13_c_13), .I2(n63), 
            .I3(GND_net), .O(n4167));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3905_3_lut (.I0(\REG.mem_50_2 ), .I1(FIFO_D2_c_2), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n4994));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3906_3_lut (.I0(\REG.mem_50_3 ), .I1(FIFO_D3_c_3), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n4995));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_936_1013_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_1110), .I3(n8756), .O(n126)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3079_3_lut (.I0(\REG.mem_2_14 ), .I1(FIFO_D14_c_14), .I2(n63), 
            .I3(GND_net), .O(n4168));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3907_3_lut (.I0(\REG.mem_50_4 ), .I1(FIFO_D4_c_4), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n4996));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3908_3_lut (.I0(\REG.mem_50_5 ), .I1(FIFO_D5_c_5), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n4997));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3909_3_lut (.I0(\REG.mem_50_6 ), .I1(FIFO_D6_c_6), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n4998));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3909_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_936_1013_add_4_6 (.CI(n8756), .I0(GND_net), .I1(n21_adj_1110), 
            .CO(n8757));
    SB_LUT4 led_counter_936_1013_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_1109), .I3(n8755), .O(n127)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3910_3_lut (.I0(\REG.mem_50_7 ), .I1(FIFO_D7_c_7), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n4999));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3911_3_lut (.I0(\REG.mem_50_8 ), .I1(FIFO_D8_c_8), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n5000));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3911_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_936_1013_add_4_5 (.CI(n8755), .I0(GND_net), .I1(n22_adj_1109), 
            .CO(n8756));
    SB_LUT4 led_counter_936_1013_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_1108), .I3(n8754), .O(n128)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3080_3_lut (.I0(\REG.mem_2_15 ), .I1(FIFO_D15_c_15), .I2(n63), 
            .I3(GND_net), .O(n4169));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3080_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_936_1013_add_4_4 (.CI(n8754), .I0(GND_net), .I1(n23_adj_1108), 
            .CO(n8755));
    SB_LUT4 led_counter_936_1013_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_1107), .I3(n8753), .O(n129)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3912_3_lut (.I0(\REG.mem_50_9 ), .I1(FIFO_D9_c_9), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n5001));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3913_3_lut (.I0(\REG.mem_50_10 ), .I1(FIFO_D10_c_10), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n5002));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3914_3_lut (.I0(\REG.mem_50_11 ), .I1(FIFO_D11_c_11), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n5003));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3915_3_lut (.I0(\REG.mem_50_12 ), .I1(FIFO_D12_c_12), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n5004));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3916_3_lut (.I0(\REG.mem_50_13 ), .I1(FIFO_D13_c_13), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n5005));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3917_3_lut (.I0(\REG.mem_50_14 ), .I1(FIFO_D14_c_14), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n5006));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3918_3_lut (.I0(\REG.mem_50_15 ), .I1(FIFO_D15_c_15), .I2(n15_adj_1103), 
            .I3(GND_net), .O(n5007));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2783_4_lut (.I0(n63_adj_1105), .I1(n3474), .I2(n6572), .I3(state[3]), 
            .O(n1326));   // src/timing_controller.v(44[11:16])
    defparam i2783_4_lut.LUT_INIT = 16'h0a88;
    SB_CARRY led_counter_936_1013_add_4_3 (.CI(n8753), .I0(GND_net), .I1(n24_adj_1107), 
            .CO(n8754));
    SB_LUT4 led_counter_936_1013_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_1106), .I3(VCC_net), .O(n130)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_936_1013_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_1106), 
            .CO(n8753));
    SB_LUT4 i3610_3_lut (.I0(rx_buf_byte[1]), .I1(rx_shift_reg[1]), .I2(n2851), 
            .I3(GND_net), .O(n4699));   // src/spi.v(76[8] 221[4])
    defparam i3610_3_lut.LUT_INIT = 16'hacac;
    GND i1 (.Y(GND_net));
    SB_LUT4 i3612_3_lut (.I0(rx_shift_reg[1]), .I1(rx_shift_reg[0]), .I2(n3629), 
            .I3(GND_net), .O(n4701));   // src/spi.v(76[8] 221[4])
    defparam i3612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3919_3_lut (.I0(\REG.mem_51_0 ), .I1(FIFO_D0_c_0), .I2(n14), 
            .I3(GND_net), .O(n5008));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3921_3_lut (.I0(\REG.mem_51_1 ), .I1(FIFO_D1_c_1), .I2(n14), 
            .I3(GND_net), .O(n5010));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3922_3_lut (.I0(\REG.mem_51_2 ), .I1(FIFO_D2_c_2), .I2(n14), 
            .I3(GND_net), .O(n5011));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3923_3_lut (.I0(\REG.mem_51_3 ), .I1(FIFO_D3_c_3), .I2(n14), 
            .I3(GND_net), .O(n5012));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3924_3_lut (.I0(\REG.mem_51_4 ), .I1(FIFO_D4_c_4), .I2(n14), 
            .I3(GND_net), .O(n5013));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3925_3_lut (.I0(\REG.mem_51_5 ), .I1(FIFO_D5_c_5), .I2(n14), 
            .I3(GND_net), .O(n5014));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3926_3_lut (.I0(\REG.mem_51_6 ), .I1(FIFO_D6_c_6), .I2(n14), 
            .I3(GND_net), .O(n5015));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3927_3_lut (.I0(\REG.mem_51_7 ), .I1(FIFO_D7_c_7), .I2(n14), 
            .I3(GND_net), .O(n5016));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3928_3_lut (.I0(\REG.mem_51_8 ), .I1(FIFO_D8_c_8), .I2(n14), 
            .I3(GND_net), .O(n5017));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3929_3_lut (.I0(\REG.mem_51_9 ), .I1(FIFO_D9_c_9), .I2(n14), 
            .I3(GND_net), .O(n5018));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3930_3_lut (.I0(\REG.mem_51_10 ), .I1(FIFO_D10_c_10), .I2(n14), 
            .I3(GND_net), .O(n5019));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3931_3_lut (.I0(\REG.mem_51_11 ), .I1(FIFO_D11_c_11), .I2(n14), 
            .I3(GND_net), .O(n5020));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3932_3_lut (.I0(\REG.mem_51_12 ), .I1(FIFO_D12_c_12), .I2(n14), 
            .I3(GND_net), .O(n5021));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3933_3_lut (.I0(\REG.mem_51_13 ), .I1(FIFO_D13_c_13), .I2(n14), 
            .I3(GND_net), .O(n5022));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3934_3_lut (.I0(\REG.mem_51_14 ), .I1(FIFO_D14_c_14), .I2(n14), 
            .I3(GND_net), .O(n5023));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3935_3_lut (.I0(\REG.mem_51_15 ), .I1(FIFO_D15_c_15), .I2(n14), 
            .I3(GND_net), .O(n5024));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3629_3_lut (.I0(\REG.mem_34_0 ), .I1(FIFO_D0_c_0), .I2(n31), 
            .I3(GND_net), .O(n4718));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3630_3_lut (.I0(\REG.mem_34_1 ), .I1(FIFO_D1_c_1), .I2(n31), 
            .I3(GND_net), .O(n4719));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3631_3_lut (.I0(\REG.mem_34_2 ), .I1(FIFO_D2_c_2), .I2(n31), 
            .I3(GND_net), .O(n4720));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3632_3_lut (.I0(\REG.mem_34_3 ), .I1(FIFO_D3_c_3), .I2(n31), 
            .I3(GND_net), .O(n4721));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3633_3_lut (.I0(\REG.mem_34_4 ), .I1(FIFO_D4_c_4), .I2(n31), 
            .I3(GND_net), .O(n4722));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3634_3_lut (.I0(\REG.mem_34_5 ), .I1(FIFO_D5_c_5), .I2(n31), 
            .I3(GND_net), .O(n4723));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3635_3_lut (.I0(\REG.mem_34_6 ), .I1(FIFO_D6_c_6), .I2(n31), 
            .I3(GND_net), .O(n4724));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3635_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_937__i0 (.Q(reset_clk_counter[0]), .C(DEBUG_6_c), 
           .D(n25_adj_1125));   // src/top.v(259[27:51])
    SB_LUT4 i757_4_lut (.I0(n1586), .I1(n6572), .I2(state[3]), .I3(n63_adj_1105), 
            .O(n1431));   // src/timing_controller.v(44[11:16])
    defparam i757_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i3952_3_lut (.I0(\REG.mem_53_0 ), .I1(FIFO_D0_c_0), .I2(n12), 
            .I3(GND_net), .O(n5041));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3953_3_lut (.I0(\REG.mem_53_1 ), .I1(FIFO_D1_c_1), .I2(n12), 
            .I3(GND_net), .O(n5042));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3954_3_lut (.I0(\REG.mem_53_2 ), .I1(FIFO_D2_c_2), .I2(n12), 
            .I3(GND_net), .O(n5043));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3955_3_lut (.I0(\REG.mem_53_3 ), .I1(FIFO_D3_c_3), .I2(n12), 
            .I3(GND_net), .O(n5044));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3956_3_lut (.I0(\REG.mem_53_4 ), .I1(FIFO_D4_c_4), .I2(n12), 
            .I3(GND_net), .O(n5045));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3957_3_lut (.I0(\REG.mem_53_5 ), .I1(FIFO_D5_c_5), .I2(n12), 
            .I3(GND_net), .O(n5046));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3958_3_lut (.I0(\REG.mem_53_6 ), .I1(FIFO_D6_c_6), .I2(n12), 
            .I3(GND_net), .O(n5047));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3959_3_lut (.I0(\REG.mem_53_7 ), .I1(FIFO_D7_c_7), .I2(n12), 
            .I3(GND_net), .O(n5048));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3960_3_lut (.I0(\REG.mem_53_8 ), .I1(FIFO_D8_c_8), .I2(n12), 
            .I3(GND_net), .O(n5049));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3961_3_lut (.I0(\REG.mem_53_9 ), .I1(FIFO_D9_c_9), .I2(n12), 
            .I3(GND_net), .O(n5050));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3962_3_lut (.I0(\REG.mem_53_10 ), .I1(FIFO_D10_c_10), .I2(n12), 
            .I3(GND_net), .O(n5051));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3963_3_lut (.I0(\REG.mem_53_11 ), .I1(FIFO_D11_c_11), .I2(n12), 
            .I3(GND_net), .O(n5052));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3964_3_lut (.I0(\REG.mem_53_12 ), .I1(FIFO_D12_c_12), .I2(n12), 
            .I3(GND_net), .O(n5053));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3965_3_lut (.I0(\REG.mem_53_13 ), .I1(FIFO_D13_c_13), .I2(n12), 
            .I3(GND_net), .O(n5054));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3966_3_lut (.I0(\REG.mem_53_14 ), .I1(FIFO_D14_c_14), .I2(n12), 
            .I3(GND_net), .O(n5055));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3967_3_lut (.I0(\REG.mem_53_15 ), .I1(FIFO_D15_c_15), .I2(n12), 
            .I3(GND_net), .O(n5056));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3968_3_lut (.I0(\REG.mem_54_0 ), .I1(FIFO_D0_c_0), .I2(n11), 
            .I3(GND_net), .O(n5057));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3065_3_lut (.I0(\REG.mem_2_0 ), .I1(FIFO_D0_c_0), .I2(n63), 
            .I3(GND_net), .O(n4154));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3971_3_lut (.I0(\REG.mem_54_1 ), .I1(FIFO_D1_c_1), .I2(n11), 
            .I3(GND_net), .O(n5060));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3066_3_lut (.I0(\REG.mem_2_1 ), .I1(FIFO_D1_c_1), .I2(n63), 
            .I3(GND_net), .O(n4155));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3972_3_lut (.I0(\REG.mem_54_2 ), .I1(FIFO_D2_c_2), .I2(n11), 
            .I3(GND_net), .O(n5061));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3559_3_lut (.I0(\REG.mem_30_14 ), .I1(FIFO_D14_c_14), .I2(n35), 
            .I3(GND_net), .O(n4648));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3973_3_lut (.I0(\REG.mem_54_3 ), .I1(FIFO_D3_c_3), .I2(n11), 
            .I3(GND_net), .O(n5062));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3974_3_lut (.I0(\REG.mem_54_4 ), .I1(FIFO_D4_c_4), .I2(n11), 
            .I3(GND_net), .O(n5063));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3975_3_lut (.I0(\REG.mem_54_5 ), .I1(FIFO_D5_c_5), .I2(n11), 
            .I3(GND_net), .O(n5064));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3976_3_lut (.I0(\REG.mem_54_6 ), .I1(FIFO_D6_c_6), .I2(n11), 
            .I3(GND_net), .O(n5065));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3977_3_lut (.I0(\REG.mem_54_7 ), .I1(FIFO_D7_c_7), .I2(n11), 
            .I3(GND_net), .O(n5066));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3978_3_lut (.I0(\REG.mem_54_8 ), .I1(FIFO_D8_c_8), .I2(n11), 
            .I3(GND_net), .O(n5067));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3979_3_lut (.I0(\REG.mem_54_9 ), .I1(FIFO_D9_c_9), .I2(n11), 
            .I3(GND_net), .O(n5068));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3980_3_lut (.I0(\REG.mem_54_10 ), .I1(FIFO_D10_c_10), .I2(n11), 
            .I3(GND_net), .O(n5069));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3981_3_lut (.I0(\REG.mem_54_11 ), .I1(FIFO_D11_c_11), .I2(n11), 
            .I3(GND_net), .O(n5070));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3982_3_lut (.I0(\REG.mem_54_12 ), .I1(FIFO_D12_c_12), .I2(n11), 
            .I3(GND_net), .O(n5071));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3983_3_lut (.I0(\REG.mem_54_13 ), .I1(FIFO_D13_c_13), .I2(n11), 
            .I3(GND_net), .O(n5072));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3983_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF even_byte_flag_87 (.Q(even_byte_flag), .C(DEBUG_6_c), .D(n2326));   // src/top.v(1032[8] 1094[4])
    SB_LUT4 i3984_3_lut (.I0(\REG.mem_54_14 ), .I1(FIFO_D14_c_14), .I2(n11), 
            .I3(GND_net), .O(n5073));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3636_3_lut (.I0(\REG.mem_34_7 ), .I1(FIFO_D7_c_7), .I2(n31), 
            .I3(GND_net), .O(n4725));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3637_3_lut (.I0(\REG.mem_34_8 ), .I1(FIFO_D8_c_8), .I2(n31), 
            .I3(GND_net), .O(n4726));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3638_3_lut (.I0(\REG.mem_34_9 ), .I1(FIFO_D9_c_9), .I2(n31), 
            .I3(GND_net), .O(n4727));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3639_3_lut (.I0(\REG.mem_34_10 ), .I1(FIFO_D10_c_10), .I2(n31), 
            .I3(GND_net), .O(n4728));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3640_3_lut (.I0(\REG.mem_34_11 ), .I1(FIFO_D11_c_11), .I2(n31), 
            .I3(GND_net), .O(n4729));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3641_3_lut (.I0(\REG.mem_34_12 ), .I1(FIFO_D12_c_12), .I2(n31), 
            .I3(GND_net), .O(n4730));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3642_3_lut (.I0(\REG.mem_34_13 ), .I1(FIFO_D13_c_13), .I2(n31), 
            .I3(GND_net), .O(n4731));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3643_3_lut (.I0(\REG.mem_34_14 ), .I1(FIFO_D14_c_14), .I2(n31), 
            .I3(GND_net), .O(n4732));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3644_3_lut (.I0(\REG.mem_34_15 ), .I1(FIFO_D15_c_15), .I2(n31), 
            .I3(GND_net), .O(n4733));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3644_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF fifo_write_cmd_77 (.Q(fifo_write_cmd), .C(DEBUG_6_c), .D(n4135));   // src/top.v(847[8] 856[4])
    SB_LUT4 i3985_3_lut (.I0(\REG.mem_54_15 ), .I1(FIFO_D15_c_15), .I2(n11), 
            .I3(GND_net), .O(n5074));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3986_3_lut (.I0(\REG.mem_55_0 ), .I1(FIFO_D0_c_0), .I2(n10), 
            .I3(GND_net), .O(n5075));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3987_3_lut (.I0(\REG.mem_55_1 ), .I1(FIFO_D1_c_1), .I2(n10), 
            .I3(GND_net), .O(n5076));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5310_1_lut (.I0(n1326), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n6392));   // src/timing_controller.v(44[11:16])
    defparam i5310_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3988_3_lut (.I0(\REG.mem_55_2 ), .I1(FIFO_D2_c_2), .I2(n10), 
            .I3(GND_net), .O(n5077));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3988_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_all_r_75 (.Q(reset_all_w), .C(DEBUG_6_c), .D(reset_all_w_N_61));   // src/top.v(246[8] 264[4])
    SB_LUT4 i3989_3_lut (.I0(\REG.mem_55_3 ), .I1(FIFO_D3_c_3), .I2(n10), 
            .I3(GND_net), .O(n5078));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3067_3_lut (.I0(\REG.mem_2_2 ), .I1(FIFO_D2_c_2), .I2(n63), 
            .I3(GND_net), .O(n4156));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3990_3_lut (.I0(\REG.mem_55_4 ), .I1(FIFO_D4_c_4), .I2(n10), 
            .I3(GND_net), .O(n5079));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3991_3_lut (.I0(\REG.mem_55_5 ), .I1(FIFO_D5_c_5), .I2(n10), 
            .I3(GND_net), .O(n5080));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3677_3_lut (.I0(\REG.mem_37_0 ), .I1(FIFO_D0_c_0), .I2(n28), 
            .I3(GND_net), .O(n4766));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3992_3_lut (.I0(\REG.mem_55_6 ), .I1(FIFO_D6_c_6), .I2(n10), 
            .I3(GND_net), .O(n5081));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3993_3_lut (.I0(\REG.mem_55_7 ), .I1(FIFO_D7_c_7), .I2(n10), 
            .I3(GND_net), .O(n5082));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3994_3_lut (.I0(\REG.mem_55_8 ), .I1(FIFO_D8_c_8), .I2(n10), 
            .I3(GND_net), .O(n5083));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3995_3_lut (.I0(\REG.mem_55_9 ), .I1(FIFO_D9_c_9), .I2(n10), 
            .I3(GND_net), .O(n5084));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3678_3_lut (.I0(\REG.mem_37_1 ), .I1(FIFO_D1_c_1), .I2(n28), 
            .I3(GND_net), .O(n4767));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3679_3_lut (.I0(\REG.mem_37_2 ), .I1(FIFO_D2_c_2), .I2(n28), 
            .I3(GND_net), .O(n4768));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3680_3_lut (.I0(\REG.mem_37_3 ), .I1(FIFO_D3_c_3), .I2(n28), 
            .I3(GND_net), .O(n4769));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3996_3_lut (.I0(\REG.mem_55_10 ), .I1(FIFO_D10_c_10), .I2(n10), 
            .I3(GND_net), .O(n5085));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3997_3_lut (.I0(\REG.mem_55_11 ), .I1(FIFO_D11_c_11), .I2(n10), 
            .I3(GND_net), .O(n5086));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3998_3_lut (.I0(\REG.mem_55_12 ), .I1(FIFO_D12_c_12), .I2(n10), 
            .I3(GND_net), .O(n5087));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3681_3_lut (.I0(\REG.mem_37_4 ), .I1(FIFO_D4_c_4), .I2(n28), 
            .I3(GND_net), .O(n4770));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3999_3_lut (.I0(\REG.mem_55_13 ), .I1(FIFO_D13_c_13), .I2(n10), 
            .I3(GND_net), .O(n5088));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4000_3_lut (.I0(\REG.mem_55_14 ), .I1(FIFO_D14_c_14), .I2(n10), 
            .I3(GND_net), .O(n5089));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3682_3_lut (.I0(\REG.mem_37_5 ), .I1(FIFO_D5_c_5), .I2(n28), 
            .I3(GND_net), .O(n4771));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4001_3_lut (.I0(\REG.mem_55_15 ), .I1(FIFO_D15_c_15), .I2(n10), 
            .I3(GND_net), .O(n5090));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4002_3_lut (.I0(\REG.mem_56_0 ), .I1(FIFO_D0_c_0), .I2(n9), 
            .I3(GND_net), .O(n5091));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4006_3_lut (.I0(\REG.mem_56_1 ), .I1(FIFO_D1_c_1), .I2(n9), 
            .I3(GND_net), .O(n5095));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4006_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_addr_byte_r_i0_i1 (.Q(tx_addr_byte[1]), .C(DEBUG_6_c), .D(n4295));   // src/top.v(1032[8] 1094[4])
    SB_DFF tx_addr_byte_r_i0_i2 (.Q(tx_addr_byte[2]), .C(DEBUG_6_c), .D(n4294));   // src/top.v(1032[8] 1094[4])
    SB_LUT4 i4007_3_lut (.I0(\REG.mem_56_2 ), .I1(FIFO_D2_c_2), .I2(n9), 
            .I3(GND_net), .O(n5096));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4007_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_addr_byte_r_i0_i3 (.Q(tx_addr_byte[3]), .C(DEBUG_6_c), .D(n4293));   // src/top.v(1032[8] 1094[4])
    SB_DFF tx_addr_byte_r_i0_i4 (.Q(tx_addr_byte[4]), .C(DEBUG_6_c), .D(n4292));   // src/top.v(1032[8] 1094[4])
    SB_LUT4 i4008_3_lut (.I0(\REG.mem_56_3 ), .I1(FIFO_D3_c_3), .I2(n9), 
            .I3(GND_net), .O(n5097));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4008_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_addr_byte_r_i0_i5 (.Q(tx_addr_byte[5]), .C(DEBUG_6_c), .D(n4291));   // src/top.v(1032[8] 1094[4])
    SB_DFF tx_addr_byte_r_i0_i6 (.Q(tx_addr_byte[6]), .C(DEBUG_6_c), .D(n4290));   // src/top.v(1032[8] 1094[4])
    SB_LUT4 i4009_3_lut (.I0(\REG.mem_56_4 ), .I1(FIFO_D4_c_4), .I2(n9), 
            .I3(GND_net), .O(n5098));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4009_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_addr_byte_r_i0_i7 (.Q(tx_addr_byte[7]), .C(DEBUG_6_c), .D(n4289));   // src/top.v(1032[8] 1094[4])
    SB_LUT4 i4010_3_lut (.I0(\REG.mem_56_5 ), .I1(FIFO_D5_c_5), .I2(n9), 
            .I3(GND_net), .O(n5099));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4011_3_lut (.I0(\REG.mem_56_6 ), .I1(FIFO_D6_c_6), .I2(n9), 
            .I3(GND_net), .O(n5100));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4012_3_lut (.I0(\REG.mem_56_7 ), .I1(FIFO_D7_c_7), .I2(n9), 
            .I3(GND_net), .O(n5101));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4013_3_lut (.I0(\REG.mem_56_8 ), .I1(FIFO_D8_c_8), .I2(n9), 
            .I3(GND_net), .O(n5102));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4013_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_addr_byte_r_i0_i0 (.Q(tx_addr_byte[0]), .C(DEBUG_6_c), .D(n4115));   // src/top.v(1032[8] 1094[4])
    SB_LUT4 i3683_3_lut (.I0(\REG.mem_37_6 ), .I1(FIFO_D6_c_6), .I2(n28), 
            .I3(GND_net), .O(n4772));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3684_3_lut (.I0(\REG.mem_37_7 ), .I1(FIFO_D7_c_7), .I2(n28), 
            .I3(GND_net), .O(n4773));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3685_3_lut (.I0(\REG.mem_37_8 ), .I1(FIFO_D8_c_8), .I2(n28), 
            .I3(GND_net), .O(n4774));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3686_3_lut (.I0(\REG.mem_37_9 ), .I1(FIFO_D9_c_9), .I2(n28), 
            .I3(GND_net), .O(n4775));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4014_3_lut (.I0(\REG.mem_56_9 ), .I1(FIFO_D9_c_9), .I2(n9), 
            .I3(GND_net), .O(n5103));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4015_3_lut (.I0(\REG.mem_56_10 ), .I1(FIFO_D10_c_10), .I2(n9), 
            .I3(GND_net), .O(n5104));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4016_3_lut (.I0(\REG.mem_56_11 ), .I1(FIFO_D11_c_11), .I2(n9), 
            .I3(GND_net), .O(n5105));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4017_3_lut (.I0(\REG.mem_56_12 ), .I1(FIFO_D12_c_12), .I2(n9), 
            .I3(GND_net), .O(n5106));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4018_3_lut (.I0(\REG.mem_56_13 ), .I1(FIFO_D13_c_13), .I2(n9), 
            .I3(GND_net), .O(n5107));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4019_3_lut (.I0(\REG.mem_56_14 ), .I1(FIFO_D14_c_14), .I2(n9), 
            .I3(GND_net), .O(n5108));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3687_3_lut (.I0(\REG.mem_37_10 ), .I1(FIFO_D10_c_10), .I2(n28), 
            .I3(GND_net), .O(n4776));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3688_3_lut (.I0(\REG.mem_37_11 ), .I1(FIFO_D11_c_11), .I2(n28), 
            .I3(GND_net), .O(n4777));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3689_3_lut (.I0(\REG.mem_37_12 ), .I1(FIFO_D12_c_12), .I2(n28), 
            .I3(GND_net), .O(n4778));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4020_3_lut (.I0(\REG.mem_56_15 ), .I1(FIFO_D15_c_15), .I2(n9), 
            .I3(GND_net), .O(n5109));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3690_3_lut (.I0(\REG.mem_37_13 ), .I1(FIFO_D13_c_13), .I2(n28), 
            .I3(GND_net), .O(n4779));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4021_3_lut (.I0(\REG.mem_57_0 ), .I1(FIFO_D0_c_0), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5110));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3691_3_lut (.I0(\REG.mem_37_14 ), .I1(FIFO_D14_c_14), .I2(n28), 
            .I3(GND_net), .O(n4780));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3692_3_lut (.I0(\REG.mem_37_15 ), .I1(FIFO_D15_c_15), .I2(n28), 
            .I3(GND_net), .O(n4781));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3693_3_lut (.I0(\REG.mem_38_0 ), .I1(FIFO_D0_c_0), .I2(n27), 
            .I3(GND_net), .O(n4782));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3694_3_lut (.I0(\REG.mem_38_1 ), .I1(FIFO_D1_c_1), .I2(n27), 
            .I3(GND_net), .O(n4783));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3695_3_lut (.I0(\REG.mem_38_2 ), .I1(FIFO_D2_c_2), .I2(n27), 
            .I3(GND_net), .O(n4784));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3696_3_lut (.I0(\REG.mem_38_3 ), .I1(FIFO_D3_c_3), .I2(n27), 
            .I3(GND_net), .O(n4785));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3697_3_lut (.I0(\REG.mem_38_4 ), .I1(FIFO_D4_c_4), .I2(n27), 
            .I3(GND_net), .O(n4786));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3704_3_lut (.I0(\REG.mem_38_11 ), .I1(FIFO_D11_c_11), .I2(n27), 
            .I3(GND_net), .O(n4793));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4025_3_lut (.I0(\REG.mem_57_1 ), .I1(FIFO_D1_c_1), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5114));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4026_3_lut (.I0(\REG.mem_57_2 ), .I1(FIFO_D2_c_2), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5115));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4027_3_lut (.I0(\REG.mem_57_3 ), .I1(FIFO_D3_c_3), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5116));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4028_3_lut (.I0(\REG.mem_57_4 ), .I1(FIFO_D4_c_4), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5117));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4029_3_lut (.I0(\REG.mem_57_5 ), .I1(FIFO_D5_c_5), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5118));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3703_3_lut (.I0(\REG.mem_38_10 ), .I1(FIFO_D10_c_10), .I2(n27), 
            .I3(GND_net), .O(n4792));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3702_3_lut (.I0(\REG.mem_38_9 ), .I1(FIFO_D9_c_9), .I2(n27), 
            .I3(GND_net), .O(n4791));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3701_3_lut (.I0(\REG.mem_38_8 ), .I1(FIFO_D8_c_8), .I2(n27), 
            .I3(GND_net), .O(n4790));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4030_3_lut (.I0(\REG.mem_57_6 ), .I1(FIFO_D6_c_6), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5119));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3700_3_lut (.I0(\REG.mem_38_7 ), .I1(FIFO_D7_c_7), .I2(n27), 
            .I3(GND_net), .O(n4789));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3698_3_lut (.I0(\REG.mem_38_5 ), .I1(FIFO_D5_c_5), .I2(n27), 
            .I3(GND_net), .O(n4787));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4031_3_lut (.I0(\REG.mem_57_7 ), .I1(FIFO_D7_c_7), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5120));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4032_3_lut (.I0(\REG.mem_57_8 ), .I1(FIFO_D8_c_8), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5121));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4033_3_lut (.I0(\REG.mem_57_9 ), .I1(FIFO_D9_c_9), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5122));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4034_3_lut (.I0(\REG.mem_57_10 ), .I1(FIFO_D10_c_10), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5123));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4035_3_lut (.I0(\REG.mem_57_11 ), .I1(FIFO_D11_c_11), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5124));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4036_3_lut (.I0(\REG.mem_57_12 ), .I1(FIFO_D12_c_12), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5125));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4037_3_lut (.I0(\REG.mem_57_13 ), .I1(FIFO_D13_c_13), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5126));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4038_3_lut (.I0(\REG.mem_57_14 ), .I1(FIFO_D14_c_14), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5127));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3699_3_lut (.I0(\REG.mem_38_6 ), .I1(FIFO_D6_c_6), .I2(n27), 
            .I3(GND_net), .O(n4788));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4039_3_lut (.I0(\REG.mem_57_15 ), .I1(FIFO_D15_c_15), .I2(n8_adj_1102), 
            .I3(GND_net), .O(n5128));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4040_3_lut (.I0(\REG.mem_58_0 ), .I1(FIFO_D0_c_0), .I2(n7), 
            .I3(GND_net), .O(n5129));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4041_3_lut (.I0(\REG.mem_58_1 ), .I1(FIFO_D1_c_1), .I2(n7), 
            .I3(GND_net), .O(n5130));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4042_3_lut (.I0(\REG.mem_58_2 ), .I1(FIFO_D2_c_2), .I2(n7), 
            .I3(GND_net), .O(n5131));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4043_3_lut (.I0(\REG.mem_58_3 ), .I1(FIFO_D3_c_3), .I2(n7), 
            .I3(GND_net), .O(n5132));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4044_3_lut (.I0(\REG.mem_58_4 ), .I1(FIFO_D4_c_4), .I2(n7), 
            .I3(GND_net), .O(n5133));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4045_3_lut (.I0(\REG.mem_58_5 ), .I1(FIFO_D5_c_5), .I2(n7), 
            .I3(GND_net), .O(n5134));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4046_3_lut (.I0(\REG.mem_58_6 ), .I1(FIFO_D6_c_6), .I2(n7), 
            .I3(GND_net), .O(n5135));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4047_3_lut (.I0(\REG.mem_58_7 ), .I1(FIFO_D7_c_7), .I2(n7), 
            .I3(GND_net), .O(n5136));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4048_3_lut (.I0(\REG.mem_58_8 ), .I1(FIFO_D8_c_8), .I2(n7), 
            .I3(GND_net), .O(n5137));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4049_3_lut (.I0(\REG.mem_58_9 ), .I1(FIFO_D9_c_9), .I2(n7), 
            .I3(GND_net), .O(n5138));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4050_3_lut (.I0(\REG.mem_58_10 ), .I1(FIFO_D10_c_10), .I2(n7), 
            .I3(GND_net), .O(n5139));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4051_3_lut (.I0(\REG.mem_58_11 ), .I1(FIFO_D11_c_11), .I2(n7), 
            .I3(GND_net), .O(n5140));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4052_3_lut (.I0(\REG.mem_58_12 ), .I1(FIFO_D12_c_12), .I2(n7), 
            .I3(GND_net), .O(n5141));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4053_3_lut (.I0(\REG.mem_58_13 ), .I1(FIFO_D13_c_13), .I2(n7), 
            .I3(GND_net), .O(n5142));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4054_3_lut (.I0(\REG.mem_58_14 ), .I1(FIFO_D14_c_14), .I2(n7), 
            .I3(GND_net), .O(n5143));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4054_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR multi_byte_spi_trans_flag_r_84 (.Q(multi_byte_spi_trans_flag_r), 
            .C(DEBUG_6_c), .D(multi_byte_spi_trans_flag_r_N_72), .R(n3935));   // src/top.v(1032[8] 1094[4])
    SB_LUT4 i4055_3_lut (.I0(\REG.mem_58_15 ), .I1(FIFO_D15_c_15), .I2(n7), 
            .I3(GND_net), .O(n5144));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9065_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(n9355), .O(n10552));
    defparam i9065_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5519_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(n63_adj_1105), 
            .I3(GND_net), .O(n6602));
    defparam i5519_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_DFF uart_rx_complete_rising_edge_80 (.Q(uart_rx_complete_rising_edge), 
           .C(DEBUG_6_c), .D(n4098));   // src/top.v(1023[8] 1029[4])
    SB_LUT4 i4072_3_lut (.I0(\REG.mem_60_0 ), .I1(FIFO_D0_c_0), .I2(n5), 
            .I3(GND_net), .O(n5161));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4073_3_lut (.I0(\REG.mem_60_1 ), .I1(FIFO_D1_c_1), .I2(n5), 
            .I3(GND_net), .O(n5162));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4074_3_lut (.I0(\REG.mem_60_2 ), .I1(FIFO_D2_c_2), .I2(n5), 
            .I3(GND_net), .O(n5163));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4075_3_lut (.I0(\REG.mem_60_3 ), .I1(FIFO_D3_c_3), .I2(n5), 
            .I3(GND_net), .O(n5164));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4076_3_lut (.I0(\REG.mem_60_4 ), .I1(FIFO_D4_c_4), .I2(n5), 
            .I3(GND_net), .O(n5165));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4077_3_lut (.I0(\REG.mem_60_5 ), .I1(FIFO_D5_c_5), .I2(n5), 
            .I3(GND_net), .O(n5166));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4078_3_lut (.I0(\REG.mem_60_6 ), .I1(FIFO_D6_c_6), .I2(n5), 
            .I3(GND_net), .O(n5167));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4079_3_lut (.I0(\REG.mem_60_7 ), .I1(FIFO_D7_c_7), .I2(n5), 
            .I3(GND_net), .O(n5168));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4080_3_lut (.I0(\REG.mem_60_8 ), .I1(FIFO_D8_c_8), .I2(n5), 
            .I3(GND_net), .O(n5169));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4081_3_lut (.I0(\REG.mem_60_9 ), .I1(FIFO_D9_c_9), .I2(n5), 
            .I3(GND_net), .O(n5170));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4082_3_lut (.I0(\REG.mem_60_10 ), .I1(FIFO_D10_c_10), .I2(n5), 
            .I3(GND_net), .O(n5171));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4082_3_lut.LUT_INIT = 16'hcaca;
    FIFO_Quad_Word tx_fifo (.rd_fifo_en_w(rd_fifo_en_w), .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r [0]), 
            .DEBUG_6_c(DEBUG_6_c), .rd_addr_r({rd_addr_r_adj_1165}), .n8(n8_adj_1100), 
            .reset_all_w(reset_all_w), .n8_adj_4(n8), .wr_addr_r({wr_addr_r_adj_1162}), 
            .rx_buf_byte({rx_buf_byte}), .n4086(n4086), .\fifo_temp_output[1] (fifo_temp_output[1]), 
            .n4089(n4089), .\fifo_temp_output[2] (fifo_temp_output[2]), 
            .n4096(n4096), .\fifo_temp_output[3] (fifo_temp_output[3]), 
            .n5330(n5330), .VCC_net(VCC_net), .\fifo_temp_output[0] (fifo_temp_output[0]), 
            .n8987(n8987), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .n4111(n4111), .\fifo_temp_output[4] (fifo_temp_output[4]), 
            .n4123(n4123), .\fifo_temp_output[5] (fifo_temp_output[5]), 
            .n4129(n4129), .\fifo_temp_output[6] (fifo_temp_output[6]), 
            .n5317(n5317), .n5314(n5314), .n5311(n5311), .n5308(n5308), 
            .n4143(n4143), .\fifo_temp_output[7] (fifo_temp_output[7]), 
            .\rd_addr_p1_w[1] (rd_addr_p1_w_adj_1167[1]), .GND_net(GND_net), 
            .\rd_addr_p1_w[2] (rd_addr_p1_w_adj_1167[2]), .\wr_addr_p1_w[1] (wr_addr_p1_w_adj_1164[1]), 
            .n1(n1), .\wr_addr_p1_w[2] (wr_addr_p1_w_adj_1164[2]), .n8824(n8824), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r [7]), .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r [6]), 
            .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r [5]), .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r [4]), 
            .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r [3]), .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r [2]), 
            .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r [1]), .fifo_write_cmd(fifo_write_cmd), 
            .full_nxt_r(full_nxt_r), .fifo_read_cmd(fifo_read_cmd), .is_fifo_empty_flag(is_fifo_empty_flag), 
            .n9299(n9299), .n4093(n4093), .rd_fifo_en_prev_r(rd_fifo_en_prev_r)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(891[16] 907[2])
    SB_LUT4 i4083_3_lut (.I0(\REG.mem_60_11 ), .I1(FIFO_D11_c_11), .I2(n5), 
            .I3(GND_net), .O(n5172));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4084_3_lut (.I0(\REG.mem_60_12 ), .I1(FIFO_D12_c_12), .I2(n5), 
            .I3(GND_net), .O(n5173));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4219_4_lut_4_lut (.I0(rd_fifo_en_w), .I1(reset_all_w), .I2(rd_addr_p1_w_adj_1167[1]), 
            .I3(rd_addr_r_adj_1165[1]), .O(n5308));
    defparam i4219_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_DFF start_tx_79 (.Q(r_SM_Main_2__N_728[0]), .C(DEBUG_6_c), .D(n4082));   // src/top.v(868[8] 886[4])
    SB_LUT4 i4222_4_lut_4_lut (.I0(rd_fifo_en_w), .I1(reset_all_w), .I2(rd_addr_p1_w_adj_1167[2]), 
            .I3(rd_addr_r_adj_1165[2]), .O(n5311));
    defparam i4222_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4085_3_lut (.I0(\REG.mem_60_13 ), .I1(FIFO_D13_c_13), .I2(n5), 
            .I3(GND_net), .O(n5174));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4086_3_lut (.I0(\REG.mem_60_14 ), .I1(FIFO_D14_c_14), .I2(n5), 
            .I3(GND_net), .O(n5175));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4086_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF fifo_read_cmd_78 (.Q(fifo_read_cmd), .C(DEBUG_6_c), .D(start_tx_N_64));   // src/top.v(868[8] 886[4])
    SB_DFF tx_data_byte_r_i0_i0 (.Q(tx_data_byte[0]), .C(DEBUG_6_c), .D(n4073));   // src/top.v(1032[8] 1094[4])
    SB_LUT4 i3557_3_lut (.I0(\REG.mem_30_12 ), .I1(FIFO_D12_c_12), .I2(n35), 
            .I3(GND_net), .O(n4646));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4087_3_lut (.I0(\REG.mem_60_15 ), .I1(FIFO_D15_c_15), .I2(n5), 
            .I3(GND_net), .O(n5176));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4088_3_lut (.I0(\REG.mem_61_0 ), .I1(FIFO_D0_c_0), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5177));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4225_4_lut_4_lut (.I0(full_nxt_r), .I1(reset_all_w), .I2(wr_addr_p1_w_adj_1164[1]), 
            .I3(wr_addr_r_adj_1162[1]), .O(n5314));
    defparam i4225_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4228_4_lut_4_lut (.I0(full_nxt_r), .I1(reset_all_w), .I2(wr_addr_p1_w_adj_1164[2]), 
            .I3(wr_addr_r_adj_1162[2]), .O(n5317));
    defparam i4228_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i4089_3_lut (.I0(\REG.mem_61_1 ), .I1(FIFO_D1_c_1), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5178));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4090_3_lut (.I0(\REG.mem_61_2 ), .I1(FIFO_D2_c_2), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5179));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4091_3_lut (.I0(\REG.mem_61_3 ), .I1(FIFO_D3_c_3), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5180));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4092_3_lut (.I0(\REG.mem_61_4 ), .I1(FIFO_D4_c_4), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5181));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4093_3_lut (.I0(\REG.mem_61_5 ), .I1(FIFO_D5_c_5), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5182));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4094_3_lut (.I0(\REG.mem_61_6 ), .I1(FIFO_D6_c_6), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5183));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4095_3_lut (.I0(\REG.mem_61_7 ), .I1(FIFO_D7_c_7), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5184));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4096_3_lut (.I0(\REG.mem_61_8 ), .I1(FIFO_D8_c_8), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5185));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_936_1013_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(DEBUG_0_c_24), .I3(n8776), .O(n106)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 led_counter_936_1013_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n2), .I3(n8775), .O(n107)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4097_3_lut (.I0(\REG.mem_61_9 ), .I1(FIFO_D9_c_9), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5186));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4098_3_lut (.I0(\REG.mem_61_10 ), .I1(FIFO_D10_c_10), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5187));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4098_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_936_1013_add_4_25 (.CI(n8775), .I0(GND_net), .I1(n2), 
            .CO(n8776));
    SB_LUT4 i4099_3_lut (.I0(\REG.mem_61_11 ), .I1(FIFO_D11_c_11), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5188));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_936_1013_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_1124), .I3(n8774), .O(n108)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_936_1013_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_936_1013_add_4_24 (.CI(n8774), .I0(GND_net), .I1(n3_adj_1124), 
            .CO(n8775));
    SB_LUT4 i4100_3_lut (.I0(\REG.mem_61_12 ), .I1(FIFO_D12_c_12), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5189));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4101_3_lut (.I0(\REG.mem_61_13 ), .I1(FIFO_D13_c_13), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5190));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4102_3_lut (.I0(\REG.mem_61_14 ), .I1(FIFO_D14_c_14), .I2(n4_adj_1101), 
            .I3(GND_net), .O(n5191));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i4102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3723_3_lut (.I0(\REG.mem_39_14 ), .I1(FIFO_D14_c_14), .I2(n26), 
            .I3(GND_net), .O(n4812));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3556_3_lut (.I0(\REG.mem_30_11 ), .I1(FIFO_D11_c_11), .I2(n35), 
            .I3(GND_net), .O(n4645));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3555_3_lut (.I0(\REG.mem_30_10 ), .I1(FIFO_D10_c_10), .I2(n35), 
            .I3(GND_net), .O(n4644));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3554_3_lut (.I0(\REG.mem_30_9 ), .I1(FIFO_D9_c_9), .I2(n35), 
            .I3(GND_net), .O(n4643));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3553_3_lut (.I0(\REG.mem_30_8 ), .I1(FIFO_D8_c_8), .I2(n35), 
            .I3(GND_net), .O(n4642));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3552_3_lut (.I0(\REG.mem_30_7 ), .I1(FIFO_D7_c_7), .I2(n35), 
            .I3(GND_net), .O(n4641));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3551_3_lut (.I0(\REG.mem_30_6 ), .I1(FIFO_D6_c_6), .I2(n35), 
            .I3(GND_net), .O(n4640));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3550_3_lut (.I0(\REG.mem_30_5 ), .I1(FIFO_D5_c_5), .I2(n35), 
            .I3(GND_net), .O(n4639));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3549_3_lut (.I0(\REG.mem_30_4 ), .I1(FIFO_D4_c_4), .I2(n35), 
            .I3(GND_net), .O(n4638));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3548_3_lut (.I0(\REG.mem_30_3 ), .I1(FIFO_D3_c_3), .I2(n35), 
            .I3(GND_net), .O(n4637));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3547_3_lut (.I0(\REG.mem_30_2 ), .I1(FIFO_D2_c_2), .I2(n35), 
            .I3(GND_net), .O(n4636));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3546_3_lut (.I0(\REG.mem_30_1 ), .I1(FIFO_D1_c_1), .I2(n35), 
            .I3(GND_net), .O(n4635));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3545_3_lut (.I0(\REG.mem_30_0 ), .I1(FIFO_D0_c_0), .I2(n35), 
            .I3(GND_net), .O(n4634));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3544_2_lut (.I0(reset_all), .I1(rd_addr_nxt_c_6__N_176[1]), 
            .I2(GND_net), .I3(GND_net), .O(n4633));   // src/fifo_dc_32_lut_gen.v(558[21] 574[24])
    defparam i3544_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3542_2_lut (.I0(reset_all), .I1(rd_addr_nxt_c_6__N_176[3]), 
            .I2(GND_net), .I3(GND_net), .O(n4631));   // src/fifo_dc_32_lut_gen.v(558[21] 574[24])
    defparam i3542_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3540_2_lut (.I0(reset_all), .I1(rd_addr_nxt_c_6__N_176[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4629));   // src/fifo_dc_32_lut_gen.v(558[21] 574[24])
    defparam i3540_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3538_3_lut (.I0(\REG.mem_29_15 ), .I1(FIFO_D15_c_15), .I2(n36), 
            .I3(GND_net), .O(n4627));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3537_3_lut (.I0(\REG.mem_29_14 ), .I1(FIFO_D14_c_14), .I2(n36), 
            .I3(GND_net), .O(n4626));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3536_3_lut (.I0(\REG.mem_29_13 ), .I1(FIFO_D13_c_13), .I2(n36), 
            .I3(GND_net), .O(n4625));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3535_3_lut (.I0(\REG.mem_29_12 ), .I1(FIFO_D12_c_12), .I2(n36), 
            .I3(GND_net), .O(n4624));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3534_3_lut (.I0(\REG.mem_29_11 ), .I1(FIFO_D11_c_11), .I2(n36), 
            .I3(GND_net), .O(n4623));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3533_3_lut (.I0(\REG.mem_29_10 ), .I1(FIFO_D10_c_10), .I2(n36), 
            .I3(GND_net), .O(n4622));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3532_3_lut (.I0(\REG.mem_29_9 ), .I1(FIFO_D9_c_9), .I2(n36), 
            .I3(GND_net), .O(n4621));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3531_3_lut (.I0(\REG.mem_29_8 ), .I1(FIFO_D8_c_8), .I2(n36), 
            .I3(GND_net), .O(n4620));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3530_3_lut (.I0(\REG.mem_29_7 ), .I1(FIFO_D7_c_7), .I2(n36), 
            .I3(GND_net), .O(n4619));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3529_3_lut (.I0(\REG.mem_29_6 ), .I1(FIFO_D6_c_6), .I2(n36), 
            .I3(GND_net), .O(n4618));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3528_3_lut (.I0(\REG.mem_29_5 ), .I1(FIFO_D5_c_5), .I2(n36), 
            .I3(GND_net), .O(n4617));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3527_3_lut (.I0(\REG.mem_29_4 ), .I1(FIFO_D4_c_4), .I2(n36), 
            .I3(GND_net), .O(n4616));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3526_3_lut (.I0(\REG.mem_29_3 ), .I1(FIFO_D3_c_3), .I2(n36), 
            .I3(GND_net), .O(n4615));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3525_3_lut (.I0(\REG.mem_29_2 ), .I1(FIFO_D2_c_2), .I2(n36), 
            .I3(GND_net), .O(n4614));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3524_3_lut (.I0(\REG.mem_29_1 ), .I1(FIFO_D1_c_1), .I2(n36), 
            .I3(GND_net), .O(n4613));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3523_3_lut (.I0(\REG.mem_29_0 ), .I1(FIFO_D0_c_0), .I2(n36), 
            .I3(GND_net), .O(n4612));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3522_3_lut (.I0(\REG.mem_28_15 ), .I1(FIFO_D15_c_15), .I2(n37), 
            .I3(GND_net), .O(n4611));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3521_3_lut (.I0(\REG.mem_28_14 ), .I1(FIFO_D14_c_14), .I2(n37), 
            .I3(GND_net), .O(n4610));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3520_3_lut (.I0(\REG.mem_28_13 ), .I1(FIFO_D13_c_13), .I2(n37), 
            .I3(GND_net), .O(n4609));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3519_3_lut (.I0(\REG.mem_28_12 ), .I1(FIFO_D12_c_12), .I2(n37), 
            .I3(GND_net), .O(n4608));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3518_3_lut (.I0(\REG.mem_28_11 ), .I1(FIFO_D11_c_11), .I2(n37), 
            .I3(GND_net), .O(n4607));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3517_3_lut (.I0(\REG.mem_28_10 ), .I1(FIFO_D10_c_10), .I2(n37), 
            .I3(GND_net), .O(n4606));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3516_3_lut (.I0(\REG.mem_28_9 ), .I1(FIFO_D9_c_9), .I2(n37), 
            .I3(GND_net), .O(n4605));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3515_3_lut (.I0(\REG.mem_28_8 ), .I1(FIFO_D8_c_8), .I2(n37), 
            .I3(GND_net), .O(n4604));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3514_3_lut (.I0(\REG.mem_28_7 ), .I1(FIFO_D7_c_7), .I2(n37), 
            .I3(GND_net), .O(n4603));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3513_3_lut (.I0(\REG.mem_28_6 ), .I1(FIFO_D6_c_6), .I2(n37), 
            .I3(GND_net), .O(n4602));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3512_3_lut (.I0(\REG.mem_28_5 ), .I1(FIFO_D5_c_5), .I2(n37), 
            .I3(GND_net), .O(n4601));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3511_3_lut (.I0(\REG.mem_28_4 ), .I1(FIFO_D4_c_4), .I2(n37), 
            .I3(GND_net), .O(n4600));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3510_3_lut (.I0(\REG.mem_28_3 ), .I1(FIFO_D3_c_3), .I2(n37), 
            .I3(GND_net), .O(n4599));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3509_3_lut (.I0(\REG.mem_28_2 ), .I1(FIFO_D2_c_2), .I2(n37), 
            .I3(GND_net), .O(n4598));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3508_3_lut (.I0(\REG.mem_28_1 ), .I1(FIFO_D1_c_1), .I2(n37), 
            .I3(GND_net), .O(n4597));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3507_3_lut (.I0(\REG.mem_28_0 ), .I1(FIFO_D0_c_0), .I2(n37), 
            .I3(GND_net), .O(n4596));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3490_3_lut (.I0(\REG.mem_26_15 ), .I1(FIFO_D15_c_15), .I2(n39), 
            .I3(GND_net), .O(n4579));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3489_3_lut (.I0(\REG.mem_26_14 ), .I1(FIFO_D14_c_14), .I2(n39), 
            .I3(GND_net), .O(n4578));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3488_3_lut (.I0(\REG.mem_26_13 ), .I1(FIFO_D13_c_13), .I2(n39), 
            .I3(GND_net), .O(n4577));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3487_3_lut (.I0(\REG.mem_26_12 ), .I1(FIFO_D12_c_12), .I2(n39), 
            .I3(GND_net), .O(n4576));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3486_3_lut (.I0(\REG.mem_26_11 ), .I1(FIFO_D11_c_11), .I2(n39), 
            .I3(GND_net), .O(n4575));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3485_3_lut (.I0(\REG.mem_26_10 ), .I1(FIFO_D10_c_10), .I2(n39), 
            .I3(GND_net), .O(n4574));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3484_3_lut (.I0(\REG.mem_26_9 ), .I1(FIFO_D9_c_9), .I2(n39), 
            .I3(GND_net), .O(n4573));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3483_3_lut (.I0(\REG.mem_26_8 ), .I1(FIFO_D8_c_8), .I2(n39), 
            .I3(GND_net), .O(n4572));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3482_3_lut (.I0(\REG.mem_26_7 ), .I1(FIFO_D7_c_7), .I2(n39), 
            .I3(GND_net), .O(n4571));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3481_3_lut (.I0(\REG.mem_26_6 ), .I1(FIFO_D6_c_6), .I2(n39), 
            .I3(GND_net), .O(n4570));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3480_3_lut (.I0(\REG.mem_26_5 ), .I1(FIFO_D5_c_5), .I2(n39), 
            .I3(GND_net), .O(n4569));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3479_3_lut (.I0(\REG.mem_26_4 ), .I1(FIFO_D4_c_4), .I2(n39), 
            .I3(GND_net), .O(n4568));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3478_3_lut (.I0(\REG.mem_26_3 ), .I1(FIFO_D3_c_3), .I2(n39), 
            .I3(GND_net), .O(n4567));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3477_3_lut (.I0(\REG.mem_26_2 ), .I1(FIFO_D2_c_2), .I2(n39), 
            .I3(GND_net), .O(n4566));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3476_3_lut (.I0(\REG.mem_26_1 ), .I1(FIFO_D1_c_1), .I2(n39), 
            .I3(GND_net), .O(n4565));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3475_3_lut (.I0(\REG.mem_26_0 ), .I1(FIFO_D0_c_0), .I2(n39), 
            .I3(GND_net), .O(n4564));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3474_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n4563));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3474_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3473_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4562));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3473_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3472_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n4561));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3472_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3471_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4560));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3471_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3470_3_lut (.I0(\REG.mem_25_15 ), .I1(FIFO_D15_c_15), .I2(n40), 
            .I3(GND_net), .O(n4559));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3469_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n4558));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3469_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3468_3_lut (.I0(\REG.mem_25_14 ), .I1(FIFO_D14_c_14), .I2(n40), 
            .I3(GND_net), .O(n4557));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3467_3_lut (.I0(\REG.mem_25_13 ), .I1(FIFO_D13_c_13), .I2(n40), 
            .I3(GND_net), .O(n4556));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3466_3_lut (.I0(\REG.mem_25_12 ), .I1(FIFO_D12_c_12), .I2(n40), 
            .I3(GND_net), .O(n4555));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3465_3_lut (.I0(\REG.mem_25_11 ), .I1(FIFO_D11_c_11), .I2(n40), 
            .I3(GND_net), .O(n4554));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3464_3_lut (.I0(\REG.mem_25_10 ), .I1(FIFO_D10_c_10), .I2(n40), 
            .I3(GND_net), .O(n4553));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3463_3_lut (.I0(\REG.mem_25_9 ), .I1(FIFO_D9_c_9), .I2(n40), 
            .I3(GND_net), .O(n4552));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3462_3_lut (.I0(\REG.mem_25_8 ), .I1(FIFO_D8_c_8), .I2(n40), 
            .I3(GND_net), .O(n4551));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3461_3_lut (.I0(\REG.mem_25_7 ), .I1(FIFO_D7_c_7), .I2(n40), 
            .I3(GND_net), .O(n4550));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3460_3_lut (.I0(\REG.mem_25_6 ), .I1(FIFO_D6_c_6), .I2(n40), 
            .I3(GND_net), .O(n4549));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3459_3_lut (.I0(\REG.mem_25_5 ), .I1(FIFO_D5_c_5), .I2(n40), 
            .I3(GND_net), .O(n4548));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3458_3_lut (.I0(\REG.mem_25_4 ), .I1(FIFO_D4_c_4), .I2(n40), 
            .I3(GND_net), .O(n4547));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3457_3_lut (.I0(\REG.mem_25_3 ), .I1(FIFO_D3_c_3), .I2(n40), 
            .I3(GND_net), .O(n4546));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3456_3_lut (.I0(\REG.mem_25_2 ), .I1(FIFO_D2_c_2), .I2(n40), 
            .I3(GND_net), .O(n4545));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3455_3_lut (.I0(\REG.mem_25_1 ), .I1(FIFO_D1_c_1), .I2(n40), 
            .I3(GND_net), .O(n4544));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3454_3_lut (.I0(\REG.mem_25_0 ), .I1(FIFO_D0_c_0), .I2(n40), 
            .I3(GND_net), .O(n4543));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3453_2_lut (.I0(reset_all), .I1(wr_addr_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n4542));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3453_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3452_2_lut (.I0(reset_all), .I1(wp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n4541));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3452_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3451_2_lut (.I0(reset_all), .I1(wp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4540));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3451_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3450_2_lut (.I0(reset_all), .I1(wp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n4539));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3450_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3449_2_lut (.I0(reset_all), .I1(wp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4538));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3449_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3448_2_lut (.I0(reset_all), .I1(wp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n4537));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3448_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3447_2_lut (.I0(reset_all), .I1(wp_sync1_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n4536));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3447_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3446_3_lut (.I0(\REG.mem_24_15 ), .I1(FIFO_D15_c_15), .I2(n41), 
            .I3(GND_net), .O(n4535));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3445_3_lut (.I0(\REG.mem_24_14 ), .I1(FIFO_D14_c_14), .I2(n41), 
            .I3(GND_net), .O(n4534));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3444_3_lut (.I0(\REG.mem_24_13 ), .I1(FIFO_D13_c_13), .I2(n41), 
            .I3(GND_net), .O(n4533));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3443_3_lut (.I0(\REG.mem_24_12 ), .I1(FIFO_D12_c_12), .I2(n41), 
            .I3(GND_net), .O(n4532));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3442_3_lut (.I0(\REG.mem_24_11 ), .I1(FIFO_D11_c_11), .I2(n41), 
            .I3(GND_net), .O(n4531));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3441_3_lut (.I0(\REG.mem_24_10 ), .I1(FIFO_D10_c_10), .I2(n41), 
            .I3(GND_net), .O(n4530));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3440_3_lut (.I0(\REG.mem_24_9 ), .I1(FIFO_D9_c_9), .I2(n41), 
            .I3(GND_net), .O(n4529));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3439_3_lut (.I0(\REG.mem_24_8 ), .I1(FIFO_D8_c_8), .I2(n41), 
            .I3(GND_net), .O(n4528));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3438_3_lut (.I0(\REG.mem_24_7 ), .I1(FIFO_D7_c_7), .I2(n41), 
            .I3(GND_net), .O(n4527));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3437_3_lut (.I0(\REG.mem_24_6 ), .I1(FIFO_D6_c_6), .I2(n41), 
            .I3(GND_net), .O(n4526));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3436_3_lut (.I0(\REG.mem_24_5 ), .I1(FIFO_D5_c_5), .I2(n41), 
            .I3(GND_net), .O(n4525));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3435_3_lut (.I0(\REG.mem_24_4 ), .I1(FIFO_D4_c_4), .I2(n41), 
            .I3(GND_net), .O(n4524));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3434_3_lut (.I0(\REG.mem_24_3 ), .I1(FIFO_D3_c_3), .I2(n41), 
            .I3(GND_net), .O(n4523));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3433_3_lut (.I0(\REG.mem_24_2 ), .I1(FIFO_D2_c_2), .I2(n41), 
            .I3(GND_net), .O(n4522));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3432_3_lut (.I0(\REG.mem_24_1 ), .I1(FIFO_D1_c_1), .I2(n41), 
            .I3(GND_net), .O(n4521));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3431_3_lut (.I0(\REG.mem_24_0 ), .I1(FIFO_D0_c_0), .I2(n41), 
            .I3(GND_net), .O(n4520));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3430_3_lut (.I0(\REG.mem_23_15 ), .I1(FIFO_D15_c_15), .I2(n42), 
            .I3(GND_net), .O(n4519));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7245_2_lut_3_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(reset_clk_counter[1]), .I3(GND_net), .O(n8661));   // src/top.v(259[27:51])
    defparam i7245_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i3429_3_lut (.I0(\REG.mem_23_14 ), .I1(FIFO_D14_c_14), .I2(n42), 
            .I3(GND_net), .O(n4518));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3428_3_lut (.I0(\REG.mem_23_13 ), .I1(FIFO_D13_c_13), .I2(n42), 
            .I3(GND_net), .O(n4517));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3427_3_lut (.I0(\REG.mem_23_12 ), .I1(FIFO_D12_c_12), .I2(n42), 
            .I3(GND_net), .O(n4516));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3426_3_lut (.I0(\REG.mem_23_11 ), .I1(FIFO_D11_c_11), .I2(n42), 
            .I3(GND_net), .O(n4515));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3425_3_lut (.I0(\REG.mem_23_10 ), .I1(FIFO_D10_c_10), .I2(n42), 
            .I3(GND_net), .O(n4514));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3424_3_lut (.I0(\REG.mem_23_9 ), .I1(FIFO_D9_c_9), .I2(n42), 
            .I3(GND_net), .O(n4513));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3423_3_lut (.I0(\REG.mem_23_8 ), .I1(FIFO_D8_c_8), .I2(n42), 
            .I3(GND_net), .O(n4512));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3422_3_lut (.I0(\REG.mem_23_7 ), .I1(FIFO_D7_c_7), .I2(n42), 
            .I3(GND_net), .O(n4511));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3421_3_lut (.I0(\REG.mem_23_6 ), .I1(FIFO_D6_c_6), .I2(n42), 
            .I3(GND_net), .O(n4510));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3420_3_lut (.I0(\REG.mem_23_5 ), .I1(FIFO_D5_c_5), .I2(n42), 
            .I3(GND_net), .O(n4509));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3419_3_lut (.I0(\REG.mem_23_4 ), .I1(FIFO_D4_c_4), .I2(n42), 
            .I3(GND_net), .O(n4508));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3418_3_lut (.I0(\REG.mem_23_3 ), .I1(FIFO_D3_c_3), .I2(n42), 
            .I3(GND_net), .O(n4507));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3417_3_lut (.I0(\REG.mem_23_2 ), .I1(FIFO_D2_c_2), .I2(n42), 
            .I3(GND_net), .O(n4506));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3416_3_lut (.I0(\REG.mem_23_1 ), .I1(FIFO_D1_c_1), .I2(n42), 
            .I3(GND_net), .O(n4505));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3415_3_lut (.I0(\REG.mem_23_0 ), .I1(FIFO_D0_c_0), .I2(n42), 
            .I3(GND_net), .O(n4504));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3414_3_lut (.I0(\REG.mem_22_15 ), .I1(FIFO_D15_c_15), .I2(n43), 
            .I3(GND_net), .O(n4503));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(reset_clk_counter[1]), .I3(GND_net), .O(n8859));   // src/top.v(259[27:51])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i3413_3_lut (.I0(\REG.mem_22_14 ), .I1(FIFO_D14_c_14), .I2(n43), 
            .I3(GND_net), .O(n4502));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3412_3_lut (.I0(\REG.mem_22_13 ), .I1(FIFO_D13_c_13), .I2(n43), 
            .I3(GND_net), .O(n4501));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3411_3_lut (.I0(\REG.mem_22_12 ), .I1(FIFO_D12_c_12), .I2(n43), 
            .I3(GND_net), .O(n4500));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3410_3_lut (.I0(\REG.mem_22_11 ), .I1(FIFO_D11_c_11), .I2(n43), 
            .I3(GND_net), .O(n4499));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3409_3_lut (.I0(\REG.mem_22_10 ), .I1(FIFO_D10_c_10), .I2(n43), 
            .I3(GND_net), .O(n4498));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3408_3_lut (.I0(\REG.mem_22_9 ), .I1(FIFO_D9_c_9), .I2(n43), 
            .I3(GND_net), .O(n4497));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3407_3_lut (.I0(\REG.mem_22_8 ), .I1(FIFO_D8_c_8), .I2(n43), 
            .I3(GND_net), .O(n4496));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3406_3_lut (.I0(\REG.mem_22_7 ), .I1(FIFO_D7_c_7), .I2(n43), 
            .I3(GND_net), .O(n4495));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3405_3_lut (.I0(\REG.mem_22_6 ), .I1(FIFO_D6_c_6), .I2(n43), 
            .I3(GND_net), .O(n4494));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3404_3_lut (.I0(\REG.mem_22_5 ), .I1(FIFO_D5_c_5), .I2(n43), 
            .I3(GND_net), .O(n4493));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3403_3_lut (.I0(\REG.mem_22_4 ), .I1(FIFO_D4_c_4), .I2(n43), 
            .I3(GND_net), .O(n4492));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3402_3_lut (.I0(\REG.mem_22_3 ), .I1(FIFO_D3_c_3), .I2(n43), 
            .I3(GND_net), .O(n4491));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3401_3_lut (.I0(\REG.mem_22_2 ), .I1(FIFO_D2_c_2), .I2(n43), 
            .I3(GND_net), .O(n4490));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3400_3_lut (.I0(\REG.mem_22_1 ), .I1(FIFO_D1_c_1), .I2(n43), 
            .I3(GND_net), .O(n4489));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3399_3_lut (.I0(\REG.mem_22_0 ), .I1(FIFO_D0_c_0), .I2(n43), 
            .I3(GND_net), .O(n4488));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3398_3_lut (.I0(\REG.mem_21_15 ), .I1(FIFO_D15_c_15), .I2(n44), 
            .I3(GND_net), .O(n4487));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3397_3_lut (.I0(\REG.mem_21_14 ), .I1(FIFO_D14_c_14), .I2(n44), 
            .I3(GND_net), .O(n4486));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3396_3_lut (.I0(\REG.mem_21_13 ), .I1(FIFO_D13_c_13), .I2(n44), 
            .I3(GND_net), .O(n4485));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3395_3_lut (.I0(\REG.mem_21_12 ), .I1(FIFO_D12_c_12), .I2(n44), 
            .I3(GND_net), .O(n4484));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3394_3_lut (.I0(\REG.mem_21_11 ), .I1(FIFO_D11_c_11), .I2(n44), 
            .I3(GND_net), .O(n4483));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3393_3_lut (.I0(\REG.mem_21_10 ), .I1(FIFO_D10_c_10), .I2(n44), 
            .I3(GND_net), .O(n4482));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3392_3_lut (.I0(\REG.mem_21_9 ), .I1(FIFO_D9_c_9), .I2(n44), 
            .I3(GND_net), .O(n4481));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3391_3_lut (.I0(\REG.mem_21_8 ), .I1(FIFO_D8_c_8), .I2(n44), 
            .I3(GND_net), .O(n4480));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3390_3_lut (.I0(\REG.mem_21_7 ), .I1(FIFO_D7_c_7), .I2(n44), 
            .I3(GND_net), .O(n4479));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3389_3_lut (.I0(\REG.mem_21_6 ), .I1(FIFO_D6_c_6), .I2(n44), 
            .I3(GND_net), .O(n4478));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3388_3_lut (.I0(\REG.mem_21_5 ), .I1(FIFO_D5_c_5), .I2(n44), 
            .I3(GND_net), .O(n4477));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3387_3_lut (.I0(\REG.mem_21_4 ), .I1(FIFO_D4_c_4), .I2(n44), 
            .I3(GND_net), .O(n4476));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3386_3_lut (.I0(\REG.mem_21_3 ), .I1(FIFO_D3_c_3), .I2(n44), 
            .I3(GND_net), .O(n4475));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3385_3_lut (.I0(\REG.mem_21_2 ), .I1(FIFO_D2_c_2), .I2(n44), 
            .I3(GND_net), .O(n4474));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_1125));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3384_3_lut (.I0(\REG.mem_21_1 ), .I1(FIFO_D1_c_1), .I2(n44), 
            .I3(GND_net), .O(n4473));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3383_3_lut (.I0(\REG.mem_21_0 ), .I1(FIFO_D0_c_0), .I2(n44), 
            .I3(GND_net), .O(n4472));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3366_3_lut (.I0(\REG.mem_19_15 ), .I1(FIFO_D15_c_15), .I2(n46), 
            .I3(GND_net), .O(n4455));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3365_3_lut (.I0(\REG.mem_19_14 ), .I1(FIFO_D14_c_14), .I2(n46), 
            .I3(GND_net), .O(n4454));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3364_3_lut (.I0(\REG.mem_19_13 ), .I1(FIFO_D13_c_13), .I2(n46), 
            .I3(GND_net), .O(n4453));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3363_3_lut (.I0(\REG.mem_19_12 ), .I1(FIFO_D12_c_12), .I2(n46), 
            .I3(GND_net), .O(n4452));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3362_3_lut (.I0(\REG.mem_19_11 ), .I1(FIFO_D11_c_11), .I2(n46), 
            .I3(GND_net), .O(n4451));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3361_3_lut (.I0(\REG.mem_19_10 ), .I1(FIFO_D10_c_10), .I2(n46), 
            .I3(GND_net), .O(n4450));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3360_3_lut (.I0(\REG.mem_19_9 ), .I1(FIFO_D9_c_9), .I2(n46), 
            .I3(GND_net), .O(n4449));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3359_3_lut (.I0(\REG.mem_19_8 ), .I1(FIFO_D8_c_8), .I2(n46), 
            .I3(GND_net), .O(n4448));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3358_3_lut (.I0(\REG.mem_19_7 ), .I1(FIFO_D7_c_7), .I2(n46), 
            .I3(GND_net), .O(n4447));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3357_3_lut (.I0(\REG.mem_19_6 ), .I1(FIFO_D6_c_6), .I2(n46), 
            .I3(GND_net), .O(n4446));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3356_3_lut (.I0(\REG.mem_19_5 ), .I1(FIFO_D5_c_5), .I2(n46), 
            .I3(GND_net), .O(n4445));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3355_3_lut (.I0(\REG.mem_19_4 ), .I1(FIFO_D4_c_4), .I2(n46), 
            .I3(GND_net), .O(n4444));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3354_3_lut (.I0(\REG.mem_19_3 ), .I1(FIFO_D3_c_3), .I2(n46), 
            .I3(GND_net), .O(n4443));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3353_3_lut (.I0(\REG.mem_19_2 ), .I1(FIFO_D2_c_2), .I2(n46), 
            .I3(GND_net), .O(n4442));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3352_3_lut (.I0(\REG.mem_19_1 ), .I1(FIFO_D1_c_1), .I2(n46), 
            .I3(GND_net), .O(n4441));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3351_3_lut (.I0(\REG.mem_19_0 ), .I1(FIFO_D0_c_0), .I2(n46), 
            .I3(GND_net), .O(n4440));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3350_3_lut (.I0(\REG.mem_18_15 ), .I1(FIFO_D15_c_15), .I2(n47), 
            .I3(GND_net), .O(n4439));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3056_3_lut (.I0(rx_shift_reg[2]), .I1(rx_shift_reg[1]), .I2(n3629), 
            .I3(GND_net), .O(n4145));   // src/spi.v(76[8] 221[4])
    defparam i3056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3349_3_lut (.I0(\REG.mem_18_14 ), .I1(FIFO_D14_c_14), .I2(n47), 
            .I3(GND_net), .O(n4438));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3348_3_lut (.I0(\REG.mem_18_13 ), .I1(FIFO_D13_c_13), .I2(n47), 
            .I3(GND_net), .O(n4437));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3347_3_lut (.I0(\REG.mem_18_12 ), .I1(FIFO_D12_c_12), .I2(n47), 
            .I3(GND_net), .O(n4436));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3346_3_lut (.I0(\REG.mem_18_11 ), .I1(FIFO_D11_c_11), .I2(n47), 
            .I3(GND_net), .O(n4435));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3345_3_lut (.I0(\REG.mem_18_10 ), .I1(FIFO_D10_c_10), .I2(n47), 
            .I3(GND_net), .O(n4434));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3344_3_lut (.I0(\REG.mem_18_9 ), .I1(FIFO_D9_c_9), .I2(n47), 
            .I3(GND_net), .O(n4433));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3343_3_lut (.I0(\REG.mem_18_8 ), .I1(FIFO_D8_c_8), .I2(n47), 
            .I3(GND_net), .O(n4432));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3342_3_lut (.I0(\REG.mem_18_7 ), .I1(FIFO_D7_c_7), .I2(n47), 
            .I3(GND_net), .O(n4431));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3341_3_lut (.I0(\REG.mem_18_6 ), .I1(FIFO_D6_c_6), .I2(n47), 
            .I3(GND_net), .O(n4430));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3340_3_lut (.I0(\REG.mem_18_5 ), .I1(FIFO_D5_c_5), .I2(n47), 
            .I3(GND_net), .O(n4429));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3339_3_lut (.I0(\REG.mem_18_4 ), .I1(FIFO_D4_c_4), .I2(n47), 
            .I3(GND_net), .O(n4428));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3338_3_lut (.I0(\REG.mem_18_3 ), .I1(FIFO_D3_c_3), .I2(n47), 
            .I3(GND_net), .O(n4427));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3337_3_lut (.I0(\REG.mem_18_2 ), .I1(FIFO_D2_c_2), .I2(n47), 
            .I3(GND_net), .O(n4426));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3336_3_lut (.I0(\REG.mem_18_1 ), .I1(FIFO_D1_c_1), .I2(n47), 
            .I3(GND_net), .O(n4425));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3335_3_lut (.I0(\REG.mem_18_0 ), .I1(FIFO_D0_c_0), .I2(n47), 
            .I3(GND_net), .O(n4424));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3302_3_lut (.I0(\REG.mem_15_15 ), .I1(FIFO_D15_c_15), .I2(n50), 
            .I3(GND_net), .O(n4391));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3301_3_lut (.I0(\REG.mem_15_14 ), .I1(FIFO_D14_c_14), .I2(n50), 
            .I3(GND_net), .O(n4390));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3300_3_lut (.I0(\REG.mem_15_13 ), .I1(FIFO_D13_c_13), .I2(n50), 
            .I3(GND_net), .O(n4389));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3299_3_lut (.I0(\REG.mem_15_12 ), .I1(FIFO_D12_c_12), .I2(n50), 
            .I3(GND_net), .O(n4388));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3298_3_lut (.I0(\REG.mem_15_11 ), .I1(FIFO_D11_c_11), .I2(n50), 
            .I3(GND_net), .O(n4387));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3297_3_lut (.I0(\REG.mem_15_10 ), .I1(FIFO_D10_c_10), .I2(n50), 
            .I3(GND_net), .O(n4386));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3296_3_lut (.I0(\REG.mem_15_9 ), .I1(FIFO_D9_c_9), .I2(n50), 
            .I3(GND_net), .O(n4385));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3295_3_lut (.I0(\REG.mem_15_8 ), .I1(FIFO_D8_c_8), .I2(n50), 
            .I3(GND_net), .O(n4384));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3294_3_lut (.I0(\REG.mem_15_7 ), .I1(FIFO_D7_c_7), .I2(n50), 
            .I3(GND_net), .O(n4383));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3293_3_lut (.I0(\REG.mem_15_6 ), .I1(FIFO_D6_c_6), .I2(n50), 
            .I3(GND_net), .O(n4382));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3292_3_lut (.I0(\REG.mem_15_5 ), .I1(FIFO_D5_c_5), .I2(n50), 
            .I3(GND_net), .O(n4381));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3291_3_lut (.I0(\REG.mem_15_4 ), .I1(FIFO_D4_c_4), .I2(n50), 
            .I3(GND_net), .O(n4380));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3290_3_lut (.I0(\REG.mem_15_3 ), .I1(FIFO_D3_c_3), .I2(n50), 
            .I3(GND_net), .O(n4379));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3289_3_lut (.I0(\REG.mem_15_2 ), .I1(FIFO_D2_c_2), .I2(n50), 
            .I3(GND_net), .O(n4378));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3288_3_lut (.I0(\REG.mem_15_1 ), .I1(FIFO_D1_c_1), .I2(n50), 
            .I3(GND_net), .O(n4377));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3287_3_lut (.I0(\REG.mem_15_0 ), .I1(FIFO_D0_c_0), .I2(n50), 
            .I3(GND_net), .O(n4376));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3286_3_lut (.I0(\REG.mem_14_15 ), .I1(FIFO_D15_c_15), .I2(n51), 
            .I3(GND_net), .O(n4375));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3285_3_lut (.I0(\REG.mem_14_14 ), .I1(FIFO_D14_c_14), .I2(n51), 
            .I3(GND_net), .O(n4374));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3055_3_lut (.I0(rx_shift_reg[3]), .I1(rx_shift_reg[2]), .I2(n3629), 
            .I3(GND_net), .O(n4144));   // src/spi.v(76[8] 221[4])
    defparam i3055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3284_3_lut (.I0(\REG.mem_14_13 ), .I1(FIFO_D13_c_13), .I2(n51), 
            .I3(GND_net), .O(n4373));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1266_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n2326));   // src/top.v(1032[8] 1094[4])
    defparam i1266_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3283_3_lut (.I0(\REG.mem_14_12 ), .I1(FIFO_D12_c_12), .I2(n51), 
            .I3(GND_net), .O(n4372));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3282_3_lut (.I0(\REG.mem_14_11 ), .I1(FIFO_D11_c_11), .I2(n51), 
            .I3(GND_net), .O(n4371));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3281_3_lut (.I0(\REG.mem_14_10 ), .I1(FIFO_D10_c_10), .I2(n51), 
            .I3(GND_net), .O(n4370));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3280_3_lut (.I0(\REG.mem_14_9 ), .I1(FIFO_D9_c_9), .I2(n51), 
            .I3(GND_net), .O(n4369));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3279_3_lut (.I0(\REG.mem_14_8 ), .I1(FIFO_D8_c_8), .I2(n51), 
            .I3(GND_net), .O(n4368));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3278_3_lut (.I0(\REG.mem_14_7 ), .I1(FIFO_D7_c_7), .I2(n51), 
            .I3(GND_net), .O(n4367));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3277_3_lut (.I0(\REG.mem_14_6 ), .I1(FIFO_D6_c_6), .I2(n51), 
            .I3(GND_net), .O(n4366));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3276_3_lut (.I0(\REG.mem_14_5 ), .I1(FIFO_D5_c_5), .I2(n51), 
            .I3(GND_net), .O(n4365));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3275_3_lut (.I0(\REG.mem_14_4 ), .I1(FIFO_D4_c_4), .I2(n51), 
            .I3(GND_net), .O(n4364));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3274_3_lut (.I0(\REG.mem_14_3 ), .I1(FIFO_D3_c_3), .I2(n51), 
            .I3(GND_net), .O(n4363));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3273_3_lut (.I0(\REG.mem_14_2 ), .I1(FIFO_D2_c_2), .I2(n51), 
            .I3(GND_net), .O(n4362));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3272_3_lut (.I0(\REG.mem_14_1 ), .I1(FIFO_D1_c_1), .I2(n51), 
            .I3(GND_net), .O(n4361));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3271_3_lut (.I0(\REG.mem_14_0 ), .I1(FIFO_D0_c_0), .I2(n51), 
            .I3(GND_net), .O(n4360));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3270_3_lut (.I0(\REG.mem_13_15 ), .I1(FIFO_D15_c_15), .I2(n52), 
            .I3(GND_net), .O(n4359));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3269_3_lut (.I0(\REG.mem_13_14 ), .I1(FIFO_D14_c_14), .I2(n52), 
            .I3(GND_net), .O(n4358));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3268_3_lut (.I0(\REG.mem_13_13 ), .I1(FIFO_D13_c_13), .I2(n52), 
            .I3(GND_net), .O(n4357));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3267_3_lut (.I0(\REG.mem_13_12 ), .I1(FIFO_D12_c_12), .I2(n52), 
            .I3(GND_net), .O(n4356));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3266_3_lut (.I0(\REG.mem_13_11 ), .I1(FIFO_D11_c_11), .I2(n52), 
            .I3(GND_net), .O(n4355));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3265_3_lut (.I0(\REG.mem_13_10 ), .I1(FIFO_D10_c_10), .I2(n52), 
            .I3(GND_net), .O(n4354));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3264_3_lut (.I0(\REG.mem_13_9 ), .I1(FIFO_D9_c_9), .I2(n52), 
            .I3(GND_net), .O(n4353));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3263_3_lut (.I0(\REG.mem_13_8 ), .I1(FIFO_D8_c_8), .I2(n52), 
            .I3(GND_net), .O(n4352));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3262_3_lut (.I0(\REG.mem_13_7 ), .I1(FIFO_D7_c_7), .I2(n52), 
            .I3(GND_net), .O(n4351));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3048_3_lut (.I0(rx_shift_reg[4]), .I1(rx_shift_reg[3]), .I2(n3629), 
            .I3(GND_net), .O(n4137));   // src/spi.v(76[8] 221[4])
    defparam i3048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3261_3_lut (.I0(\REG.mem_13_6 ), .I1(FIFO_D6_c_6), .I2(n52), 
            .I3(GND_net), .O(n4350));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3046_2_lut (.I0(is_tx_fifo_full_flag), .I1(spi_rx_byte_ready), 
            .I2(GND_net), .I3(GND_net), .O(n4135));   // src/top.v(847[8] 856[4])
    defparam i3046_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3260_3_lut (.I0(\REG.mem_13_5 ), .I1(FIFO_D5_c_5), .I2(n52), 
            .I3(GND_net), .O(n4349));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3259_3_lut (.I0(\REG.mem_13_4 ), .I1(FIFO_D4_c_4), .I2(n52), 
            .I3(GND_net), .O(n4348));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3258_3_lut (.I0(\REG.mem_13_3 ), .I1(FIFO_D3_c_3), .I2(n52), 
            .I3(GND_net), .O(n4347));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3257_3_lut (.I0(\REG.mem_13_2 ), .I1(FIFO_D2_c_2), .I2(n52), 
            .I3(GND_net), .O(n4346));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3256_3_lut (.I0(\REG.mem_13_1 ), .I1(FIFO_D1_c_1), .I2(n52), 
            .I3(GND_net), .O(n4345));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3255_3_lut (.I0(\REG.mem_13_0 ), .I1(FIFO_D0_c_0), .I2(n52), 
            .I3(GND_net), .O(n4344));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3254_3_lut (.I0(\REG.mem_12_15 ), .I1(FIFO_D15_c_15), .I2(n53), 
            .I3(GND_net), .O(n4343));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3253_3_lut (.I0(\REG.mem_12_14 ), .I1(FIFO_D14_c_14), .I2(n53), 
            .I3(GND_net), .O(n4342));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3252_3_lut (.I0(\REG.mem_12_13 ), .I1(FIFO_D13_c_13), .I2(n53), 
            .I3(GND_net), .O(n4341));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3251_3_lut (.I0(\REG.mem_12_12 ), .I1(FIFO_D12_c_12), .I2(n53), 
            .I3(GND_net), .O(n4340));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3250_3_lut (.I0(\REG.mem_12_11 ), .I1(FIFO_D11_c_11), .I2(n53), 
            .I3(GND_net), .O(n4339));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3249_3_lut (.I0(\REG.mem_12_10 ), .I1(FIFO_D10_c_10), .I2(n53), 
            .I3(GND_net), .O(n4338));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3248_3_lut (.I0(\REG.mem_12_9 ), .I1(FIFO_D9_c_9), .I2(n53), 
            .I3(GND_net), .O(n4337));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3247_3_lut (.I0(\REG.mem_12_8 ), .I1(FIFO_D8_c_8), .I2(n53), 
            .I3(GND_net), .O(n4336));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3246_3_lut (.I0(\REG.mem_12_7 ), .I1(FIFO_D7_c_7), .I2(n53), 
            .I3(GND_net), .O(n4335));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3245_3_lut (.I0(\REG.mem_12_6 ), .I1(FIFO_D6_c_6), .I2(n53), 
            .I3(GND_net), .O(n4334));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3244_3_lut (.I0(\REG.mem_12_5 ), .I1(FIFO_D5_c_5), .I2(n53), 
            .I3(GND_net), .O(n4333));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3243_3_lut (.I0(\REG.mem_12_4 ), .I1(FIFO_D4_c_4), .I2(n53), 
            .I3(GND_net), .O(n4332));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3242_3_lut (.I0(\REG.mem_12_3 ), .I1(FIFO_D3_c_3), .I2(n53), 
            .I3(GND_net), .O(n4331));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3241_3_lut (.I0(\REG.mem_12_2 ), .I1(FIFO_D2_c_2), .I2(n53), 
            .I3(GND_net), .O(n4330));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3240_3_lut (.I0(\REG.mem_12_1 ), .I1(FIFO_D1_c_1), .I2(n53), 
            .I3(GND_net), .O(n4329));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3239_3_lut (.I0(\REG.mem_12_0 ), .I1(FIFO_D0_c_0), .I2(n53), 
            .I3(GND_net), .O(n4328));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3238_3_lut (.I0(\REG.mem_11_15 ), .I1(FIFO_D15_c_15), .I2(n54), 
            .I3(GND_net), .O(n4327));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3237_3_lut (.I0(\REG.mem_11_14 ), .I1(FIFO_D14_c_14), .I2(n54), 
            .I3(GND_net), .O(n4326));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3236_3_lut (.I0(\REG.mem_11_13 ), .I1(FIFO_D13_c_13), .I2(n54), 
            .I3(GND_net), .O(n4325));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3235_3_lut (.I0(\REG.mem_11_12 ), .I1(FIFO_D12_c_12), .I2(n54), 
            .I3(GND_net), .O(n4324));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2993_3_lut_4_lut (.I0(fifo_read_cmd), .I1(r_SM_Main_2__N_728[0]), 
            .I2(is_fifo_empty_flag), .I3(tx_uart_active_flag), .O(n4082));   // src/top.v(868[8] 886[4])
    defparam i2993_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i3234_3_lut (.I0(\REG.mem_11_11 ), .I1(FIFO_D11_c_11), .I2(n54), 
            .I3(GND_net), .O(n4323));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3233_3_lut (.I0(\REG.mem_11_10 ), .I1(FIFO_D10_c_10), .I2(n54), 
            .I3(GND_net), .O(n4322));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3232_3_lut (.I0(\REG.mem_11_9 ), .I1(FIFO_D9_c_9), .I2(n54), 
            .I3(GND_net), .O(n4321));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_1138[1]), .I1(r_SM_Main_2__N_725[1]), 
            .I2(r_SM_Main_adj_1138[0]), .I3(r_SM_Main_adj_1138[2]), .O(n12410));   // src/uart_tx.v(38[10] 141[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i3231_3_lut (.I0(\REG.mem_11_8 ), .I1(FIFO_D8_c_8), .I2(n54), 
            .I3(GND_net), .O(n4320));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3230_3_lut (.I0(\REG.mem_11_7 ), .I1(FIFO_D7_c_7), .I2(n54), 
            .I3(GND_net), .O(n4319));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3001_4_lut_4_lut (.I0(tx_uart_active_flag), .I1(r_SM_Main_adj_1138[1]), 
            .I2(r_SM_Main_adj_1138[2]), .I3(n4_adj_1099), .O(n4090));   // src/uart_tx.v(38[10] 141[8])
    defparam i3001_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i3229_3_lut (.I0(\REG.mem_11_6 ), .I1(FIFO_D6_c_6), .I2(n54), 
            .I3(GND_net), .O(n4318));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3228_3_lut (.I0(\REG.mem_11_5 ), .I1(FIFO_D5_c_5), .I2(n54), 
            .I3(GND_net), .O(n4317));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3227_3_lut (.I0(\REG.mem_11_4 ), .I1(FIFO_D4_c_4), .I2(n54), 
            .I3(GND_net), .O(n4316));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3226_3_lut (.I0(\REG.mem_11_3 ), .I1(FIFO_D3_c_3), .I2(n54), 
            .I3(GND_net), .O(n4315));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3225_3_lut (.I0(\REG.mem_11_2 ), .I1(FIFO_D2_c_2), .I2(n54), 
            .I3(GND_net), .O(n4314));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3224_3_lut (.I0(\REG.mem_11_1 ), .I1(FIFO_D1_c_1), .I2(n54), 
            .I3(GND_net), .O(n4313));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3223_3_lut (.I0(\REG.mem_11_0 ), .I1(FIFO_D0_c_0), .I2(n54), 
            .I3(GND_net), .O(n4312));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3222_3_lut (.I0(\REG.mem_10_15 ), .I1(FIFO_D15_c_15), .I2(n55), 
            .I3(GND_net), .O(n4311));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3004_2_lut_3_lut (.I0(reset_all_w), .I1(fifo_read_cmd), .I2(is_fifo_empty_flag), 
            .I3(GND_net), .O(n4093));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    defparam i3004_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i3221_3_lut (.I0(\REG.mem_10_14 ), .I1(FIFO_D14_c_14), .I2(n55), 
            .I3(GND_net), .O(n4310));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3220_3_lut (.I0(\REG.mem_10_13 ), .I1(FIFO_D13_c_13), .I2(n55), 
            .I3(GND_net), .O(n4309));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3219_3_lut (.I0(\REG.mem_10_12 ), .I1(FIFO_D12_c_12), .I2(n55), 
            .I3(GND_net), .O(n4308));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3218_3_lut (.I0(\REG.mem_10_11 ), .I1(FIFO_D11_c_11), .I2(n55), 
            .I3(GND_net), .O(n4307));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3217_3_lut (.I0(\REG.mem_10_10 ), .I1(FIFO_D10_c_10), .I2(n55), 
            .I3(GND_net), .O(n4306));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3216_3_lut (.I0(\REG.mem_10_9 ), .I1(FIFO_D9_c_9), .I2(n55), 
            .I3(GND_net), .O(n4305));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3215_3_lut (.I0(\REG.mem_10_8 ), .I1(FIFO_D8_c_8), .I2(n55), 
            .I3(GND_net), .O(n4304));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3214_3_lut (.I0(\REG.mem_10_7 ), .I1(FIFO_D7_c_7), .I2(n55), 
            .I3(GND_net), .O(n4303));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3213_3_lut (.I0(\REG.mem_10_6 ), .I1(FIFO_D6_c_6), .I2(n55), 
            .I3(GND_net), .O(n4302));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3212_3_lut (.I0(\REG.mem_10_5 ), .I1(FIFO_D5_c_5), .I2(n55), 
            .I3(GND_net), .O(n4301));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3211_3_lut (.I0(\REG.mem_10_4 ), .I1(FIFO_D4_c_4), .I2(n55), 
            .I3(GND_net), .O(n4300));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3210_3_lut (.I0(\REG.mem_10_3 ), .I1(FIFO_D3_c_3), .I2(n55), 
            .I3(GND_net), .O(n4299));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3209_3_lut (.I0(\REG.mem_10_2 ), .I1(FIFO_D2_c_2), .I2(n55), 
            .I3(GND_net), .O(n4298));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3208_3_lut (.I0(\REG.mem_10_1 ), .I1(FIFO_D1_c_1), .I2(n55), 
            .I3(GND_net), .O(n4297));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3207_3_lut (.I0(\REG.mem_10_0 ), .I1(FIFO_D0_c_0), .I2(n55), 
            .I3(GND_net), .O(n4296));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3206_3_lut (.I0(tx_addr_byte[1]), .I1(tx_data_byte[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4295));   // src/top.v(1032[8] 1094[4])
    defparam i3206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3205_3_lut (.I0(tx_addr_byte[2]), .I1(tx_data_byte[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4294));   // src/top.v(1032[8] 1094[4])
    defparam i3205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3204_3_lut (.I0(tx_addr_byte[3]), .I1(tx_data_byte[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4293));   // src/top.v(1032[8] 1094[4])
    defparam i3204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3203_3_lut (.I0(tx_addr_byte[4]), .I1(tx_data_byte[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4292));   // src/top.v(1032[8] 1094[4])
    defparam i3203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3202_3_lut (.I0(tx_addr_byte[5]), .I1(tx_data_byte[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4291));   // src/top.v(1032[8] 1094[4])
    defparam i3202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3201_3_lut (.I0(tx_addr_byte[6]), .I1(tx_data_byte[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4290));   // src/top.v(1032[8] 1094[4])
    defparam i3201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2846_1_lut_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n3935));   // src/top.v(1032[8] 1094[4])
    defparam i2846_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1_2_lut_4_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(wr_addr_r_adj_1162[0]), .I3(rd_addr_r_adj_1165[0]), .O(n4_adj_1126));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0220;
    SB_LUT4 i3200_3_lut (.I0(tx_addr_byte[7]), .I1(tx_data_byte[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4289));   // src/top.v(1032[8] 1094[4])
    defparam i3200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3199_3_lut (.I0(\REG.mem_9_15 ), .I1(FIFO_D15_c_15), .I2(n56), 
            .I3(GND_net), .O(n4288));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3041_2_lut_3_lut (.I0(reset_all), .I1(DEBUG_9_c), .I2(DEBUG_1_c), 
            .I3(GND_net), .O(n4130));   // src/fifo_dc_32_lut_gen.v(749[29] 759[32])
    defparam i3041_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i3198_2_lut (.I0(reset_all), .I1(wr_addr_nxt_c[1]), .I2(GND_net), 
            .I3(GND_net), .O(n4287));   // src/fifo_dc_32_lut_gen.v(308[21] 324[24])
    defparam i3198_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3197_3_lut (.I0(\REG.mem_9_14 ), .I1(FIFO_D14_c_14), .I2(n56), 
            .I3(GND_net), .O(n4286));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3196_3_lut (.I0(\REG.mem_9_13 ), .I1(FIFO_D13_c_13), .I2(n56), 
            .I3(GND_net), .O(n4285));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3195_3_lut (.I0(\REG.mem_9_12 ), .I1(FIFO_D12_c_12), .I2(n56), 
            .I3(GND_net), .O(n4284));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3194_3_lut (.I0(\REG.mem_9_11 ), .I1(FIFO_D11_c_11), .I2(n56), 
            .I3(GND_net), .O(n4283));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3193_3_lut (.I0(\REG.mem_9_10 ), .I1(FIFO_D10_c_10), .I2(n56), 
            .I3(GND_net), .O(n4282));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3192_3_lut (.I0(\REG.mem_9_9 ), .I1(FIFO_D9_c_9), .I2(n56), 
            .I3(GND_net), .O(n4281));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1275_2_lut_3_lut_4_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(reset_all_w), .I3(wr_addr_r_adj_1162[0]), .O(n8));
    defparam i1275_2_lut_3_lut_4_lut.LUT_INIT = 16'h0df2;
    SB_LUT4 i1274_2_lut_3_lut_4_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(reset_all_w), .I3(rd_addr_r_adj_1165[0]), .O(n8_adj_1100));
    defparam i1274_2_lut_3_lut_4_lut.LUT_INIT = 16'h0df2;
    SB_LUT4 i1_4_lut_adj_62 (.I0(reset_all_w), .I1(n9406), .I2(n24), .I3(n4_adj_1126), 
            .O(n9299));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_62.LUT_INIT = 16'hfbfa;
    SB_LUT4 i7866_4_lut (.I0(rd_addr_p1_w_adj_1167[2]), .I1(rd_addr_p1_w_adj_1167[1]), 
            .I2(wr_addr_r_adj_1162[2]), .I3(wr_addr_r_adj_1162[1]), .O(n9406));
    defparam i7866_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_3_lut_adj_63 (.I0(is_fifo_empty_flag), .I1(fifo_write_cmd), 
            .I2(n32), .I3(GND_net), .O(n24));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_3_lut_adj_63.LUT_INIT = 16'h2020;
    SB_LUT4 i1_4_lut_adj_64 (.I0(rd_addr_r_adj_1165[1]), .I1(rd_addr_r_adj_1165[0]), 
            .I2(wr_addr_r_adj_1162[1]), .I3(wr_addr_r_adj_1162[0]), .O(n32));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_64.LUT_INIT = 16'h8421;
    SB_LUT4 i3026_3_lut (.I0(tx_addr_byte[0]), .I1(tx_data_byte[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4115));   // src/top.v(1032[8] 1094[4])
    defparam i3026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(reset_all_w), .I3(rd_fifo_en_prev_r), .O(n3734));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff2;
    SB_LUT4 i3191_3_lut (.I0(\REG.mem_9_8 ), .I1(FIFO_D8_c_8), .I2(n56), 
            .I3(GND_net), .O(n4280));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3190_3_lut (.I0(\REG.mem_9_7 ), .I1(FIFO_D7_c_7), .I2(n56), 
            .I3(GND_net), .O(n4279));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3189_3_lut (.I0(\REG.mem_9_6 ), .I1(FIFO_D6_c_6), .I2(n56), 
            .I3(GND_net), .O(n4278));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3188_3_lut (.I0(\REG.mem_9_5 ), .I1(FIFO_D5_c_5), .I2(n56), 
            .I3(GND_net), .O(n4277));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3019_2_lut (.I0(reset_all), .I1(wp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4108));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3019_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3187_3_lut (.I0(\REG.mem_9_4 ), .I1(FIFO_D4_c_4), .I2(n56), 
            .I3(GND_net), .O(n4276));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3186_3_lut (.I0(\REG.mem_9_3 ), .I1(FIFO_D3_c_3), .I2(n56), 
            .I3(GND_net), .O(n4275));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3185_3_lut (.I0(\REG.mem_9_2 ), .I1(FIFO_D2_c_2), .I2(n56), 
            .I3(GND_net), .O(n4274));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3184_3_lut (.I0(\REG.mem_9_1 ), .I1(FIFO_D1_c_1), .I2(n56), 
            .I3(GND_net), .O(n4273));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3183_3_lut (.I0(\REG.mem_9_0 ), .I1(FIFO_D0_c_0), .I2(n56), 
            .I3(GND_net), .O(n4272));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3181_2_lut (.I0(reset_all), .I1(wr_addr_nxt_c[3]), .I2(GND_net), 
            .I3(GND_net), .O(n4270));   // src/fifo_dc_32_lut_gen.v(308[21] 324[24])
    defparam i3181_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3179_2_lut (.I0(reset_all), .I1(wr_addr_nxt_c[5]), .I2(GND_net), 
            .I3(GND_net), .O(n4268));   // src/fifo_dc_32_lut_gen.v(308[21] 324[24])
    defparam i3179_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3018_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4107));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    defparam i3018_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3176_3_lut (.I0(\REG.mem_8_15 ), .I1(FIFO_D15_c_15), .I2(n57), 
            .I3(GND_net), .O(n4265));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3175_3_lut (.I0(\REG.mem_8_14 ), .I1(FIFO_D14_c_14), .I2(n57), 
            .I3(GND_net), .O(n4264));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3174_3_lut (.I0(\REG.mem_8_13 ), .I1(FIFO_D13_c_13), .I2(n57), 
            .I3(GND_net), .O(n4263));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3173_3_lut (.I0(\REG.mem_8_12 ), .I1(FIFO_D12_c_12), .I2(n57), 
            .I3(GND_net), .O(n4262));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9123_4_lut (.I0(tx_data_byte[0]), .I1(tx_data_byte[1]), .I2(tx_data_byte[6]), 
            .I3(n9482), .O(multi_byte_spi_trans_flag_r_N_72));   // src/top.v(1081[10:31])
    defparam i9123_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i7940_4_lut (.I0(tx_data_byte[3]), .I1(tx_data_byte[2]), .I2(tx_data_byte[4]), 
            .I3(n9440), .O(n9482));
    defparam i7940_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i7899_2_lut (.I0(tx_data_byte[5]), .I1(tx_data_byte[7]), .I2(GND_net), 
            .I3(GND_net), .O(n9440));
    defparam i7899_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3172_3_lut (.I0(\REG.mem_8_11 ), .I1(FIFO_D11_c_11), .I2(n57), 
            .I3(GND_net), .O(n4261));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3171_3_lut (.I0(\REG.mem_8_10 ), .I1(FIFO_D10_c_10), .I2(n57), 
            .I3(GND_net), .O(n4260));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3170_3_lut (.I0(\REG.mem_8_9 ), .I1(FIFO_D9_c_9), .I2(n57), 
            .I3(GND_net), .O(n4259));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3169_3_lut (.I0(\REG.mem_8_8 ), .I1(FIFO_D8_c_8), .I2(n57), 
            .I3(GND_net), .O(n4258));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3168_3_lut (.I0(\REG.mem_8_7 ), .I1(FIFO_D7_c_7), .I2(n57), 
            .I3(GND_net), .O(n4257));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3167_3_lut (.I0(\REG.mem_8_6 ), .I1(FIFO_D6_c_6), .I2(n57), 
            .I3(GND_net), .O(n4256));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3166_3_lut (.I0(\REG.mem_8_5 ), .I1(FIFO_D5_c_5), .I2(n57), 
            .I3(GND_net), .O(n4255));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3165_3_lut (.I0(\REG.mem_8_4 ), .I1(FIFO_D4_c_4), .I2(n57), 
            .I3(GND_net), .O(n4254));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3164_3_lut (.I0(\REG.mem_8_3 ), .I1(FIFO_D3_c_3), .I2(n57), 
            .I3(GND_net), .O(n4253));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3163_3_lut (.I0(\REG.mem_8_2 ), .I1(FIFO_D2_c_2), .I2(n57), 
            .I3(GND_net), .O(n4252));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3162_3_lut (.I0(\REG.mem_8_1 ), .I1(FIFO_D1_c_1), .I2(n57), 
            .I3(GND_net), .O(n4251));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3161_3_lut (.I0(\REG.mem_8_0 ), .I1(FIFO_D0_c_0), .I2(n57), 
            .I3(GND_net), .O(n4250));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3160_3_lut (.I0(\REG.mem_7_15 ), .I1(FIFO_D15_c_15), .I2(n58), 
            .I3(GND_net), .O(n4249));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3159_3_lut (.I0(\REG.mem_7_14 ), .I1(FIFO_D14_c_14), .I2(n58), 
            .I3(GND_net), .O(n4248));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3158_3_lut (.I0(\REG.mem_7_13 ), .I1(FIFO_D13_c_13), .I2(n58), 
            .I3(GND_net), .O(n4247));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3157_3_lut (.I0(\REG.mem_7_12 ), .I1(FIFO_D12_c_12), .I2(n58), 
            .I3(GND_net), .O(n4246));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3156_3_lut (.I0(\REG.mem_7_11 ), .I1(FIFO_D11_c_11), .I2(n58), 
            .I3(GND_net), .O(n4245));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3155_3_lut (.I0(\REG.mem_7_10 ), .I1(FIFO_D10_c_10), .I2(n58), 
            .I3(GND_net), .O(n4244));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3154_3_lut (.I0(\REG.mem_7_9 ), .I1(FIFO_D9_c_9), .I2(n58), 
            .I3(GND_net), .O(n4243));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3153_3_lut (.I0(\REG.mem_7_8 ), .I1(FIFO_D8_c_8), .I2(n58), 
            .I3(GND_net), .O(n4242));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3152_3_lut (.I0(\REG.mem_7_7 ), .I1(FIFO_D7_c_7), .I2(n58), 
            .I3(GND_net), .O(n4241));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3151_3_lut (.I0(\REG.mem_7_6 ), .I1(FIFO_D6_c_6), .I2(n58), 
            .I3(GND_net), .O(n4240));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3150_3_lut (.I0(\REG.mem_7_5 ), .I1(FIFO_D5_c_5), .I2(n58), 
            .I3(GND_net), .O(n4239));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3149_3_lut (.I0(\REG.mem_7_4 ), .I1(FIFO_D4_c_4), .I2(n58), 
            .I3(GND_net), .O(n4238));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3148_3_lut (.I0(\REG.mem_7_3 ), .I1(FIFO_D3_c_3), .I2(n58), 
            .I3(GND_net), .O(n4237));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3147_3_lut (.I0(\REG.mem_7_2 ), .I1(FIFO_D2_c_2), .I2(n58), 
            .I3(GND_net), .O(n4236));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3146_3_lut (.I0(\REG.mem_7_1 ), .I1(FIFO_D1_c_1), .I2(n58), 
            .I3(GND_net), .O(n4235));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3145_3_lut (.I0(\REG.mem_7_0 ), .I1(FIFO_D0_c_0), .I2(n58), 
            .I3(GND_net), .O(n4234));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3144_3_lut (.I0(\REG.mem_6_15 ), .I1(FIFO_D15_c_15), .I2(n59), 
            .I3(GND_net), .O(n4233));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3143_3_lut (.I0(\REG.mem_6_14 ), .I1(FIFO_D14_c_14), .I2(n59), 
            .I3(GND_net), .O(n4232));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3142_3_lut (.I0(\REG.mem_6_13 ), .I1(FIFO_D13_c_13), .I2(n59), 
            .I3(GND_net), .O(n4231));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3141_3_lut (.I0(\REG.mem_6_12 ), .I1(FIFO_D12_c_12), .I2(n59), 
            .I3(GND_net), .O(n4230));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3140_3_lut (.I0(\REG.mem_6_11 ), .I1(FIFO_D11_c_11), .I2(n59), 
            .I3(GND_net), .O(n4229));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3139_3_lut (.I0(\REG.mem_6_10 ), .I1(FIFO_D10_c_10), .I2(n59), 
            .I3(GND_net), .O(n4228));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3138_3_lut (.I0(\REG.mem_6_9 ), .I1(FIFO_D9_c_9), .I2(n59), 
            .I3(GND_net), .O(n4227));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3137_3_lut (.I0(\REG.mem_6_8 ), .I1(FIFO_D8_c_8), .I2(n59), 
            .I3(GND_net), .O(n4226));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3136_3_lut (.I0(\REG.mem_6_7 ), .I1(FIFO_D7_c_7), .I2(n59), 
            .I3(GND_net), .O(n4225));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3135_3_lut (.I0(\REG.mem_6_6 ), .I1(FIFO_D6_c_6), .I2(n59), 
            .I3(GND_net), .O(n4224));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3134_3_lut (.I0(\REG.mem_6_5 ), .I1(FIFO_D5_c_5), .I2(n59), 
            .I3(GND_net), .O(n4223));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3133_3_lut (.I0(\REG.mem_6_4 ), .I1(FIFO_D4_c_4), .I2(n59), 
            .I3(GND_net), .O(n4222));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3132_3_lut (.I0(\REG.mem_6_3 ), .I1(FIFO_D3_c_3), .I2(n59), 
            .I3(GND_net), .O(n4221));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3131_3_lut (.I0(\REG.mem_6_2 ), .I1(FIFO_D2_c_2), .I2(n59), 
            .I3(GND_net), .O(n4220));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3130_3_lut (.I0(\REG.mem_6_1 ), .I1(FIFO_D1_c_1), .I2(n59), 
            .I3(GND_net), .O(n4219));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3129_3_lut (.I0(\REG.mem_6_0 ), .I1(FIFO_D0_c_0), .I2(n59), 
            .I3(GND_net), .O(n4218));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3128_3_lut (.I0(\REG.mem_5_15 ), .I1(FIFO_D15_c_15), .I2(n60), 
            .I3(GND_net), .O(n4217));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3127_3_lut (.I0(\REG.mem_5_14 ), .I1(FIFO_D14_c_14), .I2(n60), 
            .I3(GND_net), .O(n4216));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3126_3_lut (.I0(\REG.mem_5_13 ), .I1(FIFO_D13_c_13), .I2(n60), 
            .I3(GND_net), .O(n4215));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3125_3_lut (.I0(\REG.mem_5_12 ), .I1(FIFO_D12_c_12), .I2(n60), 
            .I3(GND_net), .O(n4214));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3124_3_lut (.I0(\REG.mem_5_11 ), .I1(FIFO_D11_c_11), .I2(n60), 
            .I3(GND_net), .O(n4213));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3123_3_lut (.I0(\REG.mem_5_10 ), .I1(FIFO_D10_c_10), .I2(n60), 
            .I3(GND_net), .O(n4212));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3122_3_lut (.I0(\REG.mem_5_9 ), .I1(FIFO_D9_c_9), .I2(n60), 
            .I3(GND_net), .O(n4211));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3121_3_lut (.I0(\REG.mem_5_8 ), .I1(FIFO_D8_c_8), .I2(n60), 
            .I3(GND_net), .O(n4210));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3120_3_lut (.I0(\REG.mem_5_7 ), .I1(FIFO_D7_c_7), .I2(n60), 
            .I3(GND_net), .O(n4209));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3119_3_lut (.I0(\REG.mem_5_6 ), .I1(FIFO_D6_c_6), .I2(n60), 
            .I3(GND_net), .O(n4208));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3118_3_lut (.I0(\REG.mem_5_5 ), .I1(FIFO_D5_c_5), .I2(n60), 
            .I3(GND_net), .O(n4207));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3117_3_lut (.I0(\REG.mem_5_4 ), .I1(FIFO_D4_c_4), .I2(n60), 
            .I3(GND_net), .O(n4206));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3116_3_lut (.I0(\REG.mem_5_3 ), .I1(FIFO_D3_c_3), .I2(n60), 
            .I3(GND_net), .O(n4205));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3115_3_lut (.I0(\REG.mem_5_2 ), .I1(FIFO_D2_c_2), .I2(n60), 
            .I3(GND_net), .O(n4204));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3114_3_lut (.I0(\REG.mem_5_1 ), .I1(FIFO_D1_c_1), .I2(n60), 
            .I3(GND_net), .O(n4203));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3113_3_lut (.I0(\REG.mem_5_0 ), .I1(FIFO_D0_c_0), .I2(n60), 
            .I3(GND_net), .O(n4202));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    defparam i3113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3014_2_lut (.I0(reset_all), .I1(rp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4103));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3014_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i752_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(n63_adj_1105), 
            .I3(state[2]), .O(n1586));   // src/timing_controller.v(44[11:16])
    defparam i752_4_lut_4_lut.LUT_INIT = 16'h0806;
    SB_LUT4 i3012_2_lut (.I0(reset_all), .I1(rd_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4101));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    defparam i3012_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3010_3_lut (.I0(rx_buf_byte[0]), .I1(rx_shift_reg[0]), .I2(n2851), 
            .I3(GND_net), .O(n4099));   // src/spi.v(76[8] 221[4])
    defparam i3010_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3009_2_lut (.I0(uart_rx_complete_prev), .I1(debug_led3), .I2(GND_net), 
            .I3(GND_net), .O(n4098));   // src/top.v(1023[8] 1029[4])
    defparam i3009_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3002_3_lut (.I0(r_Tx_Data[0]), .I1(fifo_temp_output[0]), .I2(n3151), 
            .I3(GND_net), .O(n4091));   // src/uart_tx.v(38[10] 141[8])
    defparam i3002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_65 (.I0(reset_clk_counter[2]), .I1(reset_all_w_N_61), 
            .I2(reset_clk_counter[0]), .I3(reset_clk_counter[1]), .O(n8861));
    defparam i1_2_lut_4_lut_adj_65.LUT_INIT = 16'haaa6;
    SB_LUT4 i9120_2_lut (.I0(is_fifo_empty_flag), .I1(tx_uart_active_flag), 
            .I2(GND_net), .I3(GND_net), .O(start_tx_N_64));
    defparam i9120_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2992_3_lut (.I0(rx_shift_reg[5]), .I1(rx_shift_reg[4]), .I2(n3629), 
            .I3(GND_net), .O(n4081));   // src/spi.v(76[8] 221[4])
    defparam i2992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2991_3_lut (.I0(rx_shift_reg[6]), .I1(rx_shift_reg[5]), .I2(n3629), 
            .I3(GND_net), .O(n4080));   // src/spi.v(76[8] 221[4])
    defparam i2991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2990_3_lut (.I0(rx_shift_reg[7]), .I1(rx_shift_reg[6]), .I2(n3629), 
            .I3(GND_net), .O(n4079));   // src/spi.v(76[8] 221[4])
    defparam i2990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2984_3_lut (.I0(tx_data_byte[0]), .I1(pc_data_rx[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4073));   // src/top.v(1032[8] 1094[4])
    defparam i2984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut_4_lut (.I0(debug_led3), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n3642), .O(n8963));   // src/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    usb3_if usb3_if_inst (.VCC_net(VCC_net), .FIFO_CLK_c(FIFO_CLK_c), .FT_OE_c(FT_OE_c), 
            .GND_net(GND_net), .FT_RD_c(FT_RD_c), .dc32_fifo_is_full(dc32_fifo_is_full), 
            .FR_RXF_c(FR_RXF_c), .write_to_dc32_fifo(write_to_dc32_fifo)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(447[9] 458[3])
    \uart_rx(CLKS_PER_BIT=20)  pc_rx (.DEBUG_6_c(DEBUG_6_c), .\r_SM_Main[2] (r_SM_Main[2]), 
            .r_Rx_Data(r_Rx_Data), .n5353(n5353), .pc_data_rx({pc_data_rx}), 
            .n5349(n5349), .n5348(n5348), .n5347(n5347), .n5345(n5345), 
            .n5344(n5344), .n8963(n8963), .VCC_net(VCC_net), .debug_led3(debug_led3), 
            .n5339(n5339), .n5338(n5338), .n5337(n5337), .r_Bit_Index({Open_0, 
            Open_1, r_Bit_Index[0]}), .GND_net(GND_net), .n4(n4), .\r_SM_Main[1] (r_SM_Main[1]), 
            .n4_adj_1(n4_adj_1098), .n9345(n9345), .n4_adj_2(n4_adj_1127), 
            .UART_RX_c(UART_RX_c), .n2414(n2414), .n3785(n3785), .n3533(n3533), 
            .n3525(n3525), .n3642(n3642), .n131(n131)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(657[42] 662[3])
    fifo_dc_32_lut_gen fifo_dc_32_lut_gen_inst (.FIFO_D6_c_6(FIFO_D6_c_6), 
            .\REG.mem_42_15 (\REG.mem_42_15 ), .\REG.mem_43_15 (\REG.mem_43_15 ), 
            .FIFO_D5_c_5(FIFO_D5_c_5), .\REG.mem_29_14 (\REG.mem_29_14 ), 
            .\REG.mem_28_14 (\REG.mem_28_14 ), .FIFO_CLK_c(FIFO_CLK_c), 
            .\REG.mem_41_15 (\REG.mem_41_15 ), .\REG.mem_40_15 (\REG.mem_40_15 ), 
            .GND_net(GND_net), .\REG.mem_2_0 (\REG.mem_2_0 ), .\REG.mem_2_2 (\REG.mem_2_2 ), 
            .FIFO_D4_c_4(FIFO_D4_c_4), .\REG.mem_18_5 (\REG.mem_18_5 ), 
            .\REG.mem_19_5 (\REG.mem_19_5 ), .FIFO_D3_c_3(FIFO_D3_c_3), 
            .\REG.mem_62_5 (\REG.mem_62_5 ), .\REG.mem_61_5 (\REG.mem_61_5 ), 
            .\REG.mem_60_5 (\REG.mem_60_5 ), .FIFO_D2_c_2(FIFO_D2_c_2), 
            .t_rd_fifo_en_w(t_rd_fifo_en_w), .\REG.out_raw[0] (\REG.out_raw [0]), 
            .DEBUG_6_c(DEBUG_6_c), .\REG.mem_30_10 (\REG.mem_30_10 ), .\REG.mem_29_10 (\REG.mem_29_10 ), 
            .\REG.mem_28_10 (\REG.mem_28_10 ), .\REG.mem_58_8 (\REG.mem_58_8 ), 
            .\REG.mem_57_8 (\REG.mem_57_8 ), .\REG.mem_56_8 (\REG.mem_56_8 ), 
            .FIFO_D1_c_1(FIFO_D1_c_1), .\REG.mem_2_14 (\REG.mem_2_14 ), 
            .FIFO_D0_c_0(FIFO_D0_c_0), .\REG.mem_14_15 (\REG.mem_14_15 ), 
            .\REG.mem_15_15 (\REG.mem_15_15 ), .\REG.mem_13_15 (\REG.mem_13_15 ), 
            .\REG.mem_12_15 (\REG.mem_12_15 ), .\REG.mem_10_15 (\REG.mem_10_15 ), 
            .\REG.mem_11_15 (\REG.mem_11_15 ), .n56(n56), .\REG.mem_62_8 (\REG.mem_62_8 ), 
            .\REG.mem_61_8 (\REG.mem_61_8 ), .\REG.mem_60_8 (\REG.mem_60_8 ), 
            .\REG.mem_46_6 (\REG.mem_46_6 ), .\REG.mem_47_6 (\REG.mem_47_6 ), 
            .n24(n24_adj_1104), .write_to_dc32_fifo(write_to_dc32_fifo), 
            .reset_all(reset_all), .\wr_addr_nxt_c[1] (wr_addr_nxt_c[1]), 
            .\REG.mem_45_6 (\REG.mem_45_6 ), .\REG.mem_44_6 (\REG.mem_44_6 ), 
            .dc32_fifo_is_full(dc32_fifo_is_full), .\REG.mem_34_10 (\REG.mem_34_10 ), 
            .\REG.mem_18_8 (\REG.mem_18_8 ), .\REG.mem_19_8 (\REG.mem_19_8 ), 
            .\REG.mem_58_11 (\REG.mem_58_11 ), .\rd_grey_sync_r[0] (rd_grey_sync_r[0]), 
            .\REG.mem_57_11 (\REG.mem_57_11 ), .\REG.mem_56_11 (\REG.mem_56_11 ), 
            .\REG.mem_6_14 (\REG.mem_6_14 ), .\REG.mem_7_14 (\REG.mem_7_14 ), 
            .\REG.mem_5_14 (\REG.mem_5_14 ), .\REG.mem_10_12 (\REG.mem_10_12 ), 
            .\REG.mem_11_12 (\REG.mem_11_12 ), .\REG.mem_9_12 (\REG.mem_9_12 ), 
            .\REG.mem_8_12 (\REG.mem_8_12 ), .\REG.mem_6_10 (\REG.mem_6_10 ), 
            .\REG.mem_7_10 (\REG.mem_7_10 ), .\REG.mem_26_9 (\REG.mem_26_9 ), 
            .DEBUG_1_c(DEBUG_1_c), .\REG.mem_6_0 (\REG.mem_6_0 ), .\REG.mem_7_0 (\REG.mem_7_0 ), 
            .\REG.mem_5_0 (\REG.mem_5_0 ), .\REG.mem_5_10 (\REG.mem_5_10 ), 
            .\REG.mem_25_9 (\REG.mem_25_9 ), .\REG.mem_24_9 (\REG.mem_24_9 ), 
            .\REG.mem_56_7 (\REG.mem_56_7 ), .\REG.mem_57_7 (\REG.mem_57_7 ), 
            .\REG.mem_58_7 (\REG.mem_58_7 ), .\num_words_in_buffer[3] (num_words_in_buffer[3]), 
            .\wr_grey_sync_r[0] (wr_grey_sync_r[0]), .\REG.mem_10_14 (\REG.mem_10_14 ), 
            .\REG.mem_11_14 (\REG.mem_11_14 ), .\REG.mem_9_14 (\REG.mem_9_14 ), 
            .\REG.mem_8_14 (\REG.mem_8_14 ), .\REG.mem_14_14 (\REG.mem_14_14 ), 
            .\REG.mem_15_14 (\REG.mem_15_14 ), .\REG.mem_13_14 (\REG.mem_13_14 ), 
            .\REG.mem_12_14 (\REG.mem_12_14 ), .\REG.mem_38_9 (\REG.mem_38_9 ), 
            .\REG.mem_39_9 (\REG.mem_39_9 ), .\REG.mem_37_9 (\REG.mem_37_9 ), 
            .\REG.mem_34_7 (\REG.mem_34_7 ), .\REG.mem_42_9 (\REG.mem_42_9 ), 
            .\REG.mem_43_9 (\REG.mem_43_9 ), .\REG.mem_10_10 (\REG.mem_10_10 ), 
            .\REG.mem_11_10 (\REG.mem_11_10 ), .\REG.mem_9_10 (\REG.mem_9_10 ), 
            .\REG.mem_8_10 (\REG.mem_8_10 ), .\REG.mem_41_9 (\REG.mem_41_9 ), 
            .\REG.mem_40_9 (\REG.mem_40_9 ), .\REG.mem_9_15 (\REG.mem_9_15 ), 
            .\REG.mem_8_15 (\REG.mem_8_15 ), .\REG.mem_18_6 (\REG.mem_18_6 ), 
            .\REG.mem_19_6 (\REG.mem_19_6 ), .\wr_addr_nxt_c[3] (wr_addr_nxt_c[3]), 
            .FIFO_D15_c_15(FIFO_D15_c_15), .\REG.mem_22_5 (\REG.mem_22_5 ), 
            .\REG.mem_23_5 (\REG.mem_23_5 ), .\REG.mem_21_5 (\REG.mem_21_5 ), 
            .\REG.mem_38_10 (\REG.mem_38_10 ), .\REG.mem_39_10 (\REG.mem_39_10 ), 
            .\REG.mem_37_10 (\REG.mem_37_10 ), .\REG.mem_18_10 (\REG.mem_18_10 ), 
            .\REG.mem_19_10 (\REG.mem_19_10 ), .FIFO_D14_c_14(FIFO_D14_c_14), 
            .\REG.mem_34_12 (\REG.mem_34_12 ), .\REG.mem_22_6 (\REG.mem_22_6 ), 
            .\REG.mem_23_6 (\REG.mem_23_6 ), .\REG.mem_26_14 (\REG.mem_26_14 ), 
            .\REG.mem_25_14 (\REG.mem_25_14 ), .\REG.mem_24_14 (\REG.mem_24_14 ), 
            .\REG.mem_18_13 (\REG.mem_18_13 ), .\REG.mem_19_13 (\REG.mem_19_13 ), 
            .\REG.mem_62_7 (\REG.mem_62_7 ), .\REG.mem_21_6 (\REG.mem_21_6 ), 
            .\REG.mem_60_7 (\REG.mem_60_7 ), .\REG.mem_61_7 (\REG.mem_61_7 ), 
            .\REG.mem_30_14 (\REG.mem_30_14 ), .\REG.mem_50_3 (\REG.mem_50_3 ), 
            .\REG.mem_51_3 (\REG.mem_51_3 ), .\REG.mem_38_12 (\REG.mem_38_12 ), 
            .\REG.mem_39_12 (\REG.mem_39_12 ), .\REG.mem_37_12 (\REG.mem_37_12 ), 
            .\REG.mem_46_8 (\REG.mem_46_8 ), .\REG.mem_47_8 (\REG.mem_47_8 ), 
            .\REG.mem_45_8 (\REG.mem_45_8 ), .\REG.mem_44_8 (\REG.mem_44_8 ), 
            .\REG.mem_58_10 (\REG.mem_58_10 ), .\REG.mem_2_3 (\REG.mem_2_3 ), 
            .\REG.mem_57_10 (\REG.mem_57_10 ), .\REG.mem_56_10 (\REG.mem_56_10 ), 
            .\REG.mem_62_2 (\REG.mem_62_2 ), .\REG.mem_61_2 (\REG.mem_61_2 ), 
            .\REG.mem_60_2 (\REG.mem_60_2 ), .\REG.mem_58_15 (\REG.mem_58_15 ), 
            .\REG.mem_10_0 (\REG.mem_10_0 ), .\REG.mem_11_0 (\REG.mem_11_0 ), 
            .\REG.mem_9_0 (\REG.mem_9_0 ), .\REG.mem_8_0 (\REG.mem_8_0 ), 
            .\REG.mem_57_15 (\REG.mem_57_15 ), .\REG.mem_56_15 (\REG.mem_56_15 ), 
            .\REG.mem_30_0 (\REG.mem_30_0 ), .\REG.mem_29_0 (\REG.mem_29_0 ), 
            .\REG.mem_28_0 (\REG.mem_28_0 ), .\REG.mem_38_7 (\REG.mem_38_7 ), 
            .\REG.mem_39_7 (\REG.mem_39_7 ), .FIFO_D13_c_13(FIFO_D13_c_13), 
            .\REG.mem_37_7 (\REG.mem_37_7 ), .n58(n58), .FIFO_D12_c_12(FIFO_D12_c_12), 
            .\REG.mem_26_5 (\REG.mem_26_5 ), .\REG.mem_25_5 (\REG.mem_25_5 ), 
            .\REG.mem_24_5 (\REG.mem_24_5 ), .n50(n50), .\REG.mem_46_0 (\REG.mem_46_0 ), 
            .\REG.mem_47_0 (\REG.mem_47_0 ), .\REG.mem_6_3 (\REG.mem_6_3 ), 
            .\REG.mem_7_3 (\REG.mem_7_3 ), .\REG.mem_5_3 (\REG.mem_5_3 ), 
            .\REG.mem_45_0 (\REG.mem_45_0 ), .\REG.mem_44_0 (\REG.mem_44_0 ), 
            .\REG.mem_50_8 (\REG.mem_50_8 ), .\REG.mem_51_8 (\REG.mem_51_8 ), 
            .n18(n18), .\REG.mem_10_3 (\REG.mem_10_3 ), .\REG.mem_11_3 (\REG.mem_11_3 ), 
            .\REG.mem_6_2 (\REG.mem_6_2 ), .\REG.mem_7_2 (\REG.mem_7_2 ), 
            .\REG.mem_5_2 (\REG.mem_5_2 ), .\REG.mem_9_3 (\REG.mem_9_3 ), 
            .\REG.mem_8_3 (\REG.mem_8_3 ), .\wr_addr_nxt_c[5] (wr_addr_nxt_c[5]), 
            .\REG.mem_42_12 (\REG.mem_42_12 ), .\REG.mem_43_12 (\REG.mem_43_12 ), 
            .\REG.mem_41_12 (\REG.mem_41_12 ), .\REG.mem_40_12 (\REG.mem_40_12 ), 
            .\REG.mem_10_2 (\REG.mem_10_2 ), .\REG.mem_11_2 (\REG.mem_11_2 ), 
            .n4169(n4169), .\REG.mem_2_15 (\REG.mem_2_15 ), .\REG.mem_9_2 (\REG.mem_9_2 ), 
            .\REG.mem_8_2 (\REG.mem_8_2 ), .n4168(n4168), .n4167(n4167), 
            .\REG.mem_2_13 (\REG.mem_2_13 ), .n4166(n4166), .\REG.mem_2_12 (\REG.mem_2_12 ), 
            .n4165(n4165), .\REG.mem_2_11 (\REG.mem_2_11 ), .n4164(n4164), 
            .\REG.mem_2_10 (\REG.mem_2_10 ), .\REG.mem_6_6 (\REG.mem_6_6 ), 
            .\REG.mem_7_6 (\REG.mem_7_6 ), .n4163(n4163), .\REG.mem_2_9 (\REG.mem_2_9 ), 
            .\REG.mem_5_6 (\REG.mem_5_6 ), .\REG.mem_30_3 (\REG.mem_30_3 ), 
            .\REG.mem_29_3 (\REG.mem_29_3 ), .\REG.mem_28_3 (\REG.mem_28_3 ), 
            .\REG.mem_22_13 (\REG.mem_22_13 ), .\REG.mem_23_13 (\REG.mem_23_13 ), 
            .\REG.mem_21_13 (\REG.mem_21_13 ), .\REG.mem_54_3 (\REG.mem_54_3 ), 
            .\REG.mem_55_3 (\REG.mem_55_3 ), .\REG.mem_53_3 (\REG.mem_53_3 ), 
            .\REG.mem_42_10 (\REG.mem_42_10 ), .\REG.mem_43_10 (\REG.mem_43_10 ), 
            .\REG.mem_41_10 (\REG.mem_41_10 ), .\REG.mem_40_10 (\REG.mem_40_10 ), 
            .\REG.mem_56_4 (\REG.mem_56_4 ), .\REG.mem_57_4 (\REG.mem_57_4 ), 
            .\REG.mem_6_15 (\REG.mem_6_15 ), .\REG.mem_7_15 (\REG.mem_7_15 ), 
            .\REG.mem_58_4 (\REG.mem_58_4 ), .\REG.mem_26_15 (\REG.mem_26_15 ), 
            .\REG.mem_5_15 (\REG.mem_5_15 ), .\REG.mem_25_15 (\REG.mem_25_15 ), 
            .\REG.mem_24_15 (\REG.mem_24_15 ), .\REG.mem_58_3 (\REG.mem_58_3 ), 
            .\REG.mem_57_3 (\REG.mem_57_3 ), .\REG.mem_56_3 (\REG.mem_56_3 ), 
            .\REG.mem_62_3 (\REG.mem_62_3 ), .\REG.mem_62_4 (\REG.mem_62_4 ), 
            .\REG.mem_60_4 (\REG.mem_60_4 ), .\REG.mem_61_4 (\REG.mem_61_4 ), 
            .\REG.mem_61_3 (\REG.mem_61_3 ), .\REG.mem_60_3 (\REG.mem_60_3 ), 
            .\rd_addr_r[6] (rd_addr_r[6]), .\rd_addr_nxt_c_6__N_176[5] (rd_addr_nxt_c_6__N_176[5]), 
            .\REG.mem_22_8 (\REG.mem_22_8 ), .\REG.mem_23_8 (\REG.mem_23_8 ), 
            .\rd_addr_nxt_c_6__N_176[3] (rd_addr_nxt_c_6__N_176[3]), .\REG.mem_21_8 (\REG.mem_21_8 ), 
            .\REG.mem_54_8 (\REG.mem_54_8 ), .\REG.mem_55_8 (\REG.mem_55_8 ), 
            .FIFO_D11_c_11(FIFO_D11_c_11), .\REG.mem_14_3 (\REG.mem_14_3 ), 
            .\REG.mem_15_3 (\REG.mem_15_3 ), .\REG.mem_53_8 (\REG.mem_53_8 ), 
            .\REG.mem_14_2 (\REG.mem_14_2 ), .\REG.mem_15_2 (\REG.mem_15_2 ), 
            .\REG.mem_13_3 (\REG.mem_13_3 ), .\REG.mem_12_3 (\REG.mem_12_3 ), 
            .\REG.mem_13_2 (\REG.mem_13_2 ), .\REG.mem_12_2 (\REG.mem_12_2 ), 
            .\REG.mem_30_5 (\REG.mem_30_5 ), .\REG.mem_58_13 (\REG.mem_58_13 ), 
            .\REG.mem_29_5 (\REG.mem_29_5 ), .\REG.mem_28_5 (\REG.mem_28_5 ), 
            .\REG.mem_34_5 (\REG.mem_34_5 ), .\REG.mem_57_13 (\REG.mem_57_13 ), 
            .\REG.mem_56_13 (\REG.mem_56_13 ), .\REG.mem_14_6 (\REG.mem_14_6 ), 
            .\REG.mem_15_6 (\REG.mem_15_6 ), .\REG.mem_13_6 (\REG.mem_13_6 ), 
            .\REG.mem_12_6 (\REG.mem_12_6 ), .\REG.mem_54_9 (\REG.mem_54_9 ), 
            .\REG.mem_55_9 (\REG.mem_55_9 ), .\REG.mem_53_9 (\REG.mem_53_9 ), 
            .\REG.mem_34_0 (\REG.mem_34_0 ), .\REG.mem_14_0 (\REG.mem_14_0 ), 
            .\REG.mem_15_0 (\REG.mem_15_0 ), .\REG.mem_13_0 (\REG.mem_13_0 ), 
            .\REG.mem_12_0 (\REG.mem_12_0 ), .FIFO_D10_c_10(FIFO_D10_c_10), 
            .\REG.mem_42_14 (\REG.mem_42_14 ), .\REG.mem_43_14 (\REG.mem_43_14 ), 
            .\REG.mem_41_14 (\REG.mem_41_14 ), .\REG.mem_40_14 (\REG.mem_40_14 ), 
            .n4162(n4162), .\REG.mem_2_8 (\REG.mem_2_8 ), .n4161(n4161), 
            .\REG.mem_2_7 (\REG.mem_2_7 ), .FIFO_D9_c_9(FIFO_D9_c_9), .n5327(n5327), 
            .VCC_net(VCC_net), .\fifo_data_out[0] (fifo_data_out[0]), .\REG.mem_10_11 (\REG.mem_10_11 ), 
            .\REG.mem_11_11 (\REG.mem_11_11 ), .FIFO_D8_c_8(FIFO_D8_c_8), 
            .FIFO_D7_c_7(FIFO_D7_c_7), .\REG.mem_9_11 (\REG.mem_9_11 ), 
            .\REG.mem_8_11 (\REG.mem_8_11 ), .\REG.mem_62_15 (\REG.mem_62_15 ), 
            .\REG.mem_62_10 (\REG.mem_62_10 ), .n5305(n5305), .\fifo_data_out[15] (fifo_data_out[15]), 
            .\REG.mem_46_12 (\REG.mem_46_12 ), .\REG.mem_47_12 (\REG.mem_47_12 ), 
            .n5302(n5302), .\fifo_data_out[14] (fifo_data_out[14]), .\REG.mem_61_10 (\REG.mem_61_10 ), 
            .\REG.mem_60_10 (\REG.mem_60_10 ), .\REG.mem_61_15 (\REG.mem_61_15 ), 
            .\REG.mem_60_15 (\REG.mem_60_15 ), .n5299(n5299), .\fifo_data_out[13] (fifo_data_out[13]), 
            .n5296(n5296), .\fifo_data_out[12] (fifo_data_out[12]), .n5293(n5293), 
            .\fifo_data_out[11] (fifo_data_out[11]), .n5290(n5290), .\fifo_data_out[10] (fifo_data_out[10]), 
            .\REG.mem_45_12 (\REG.mem_45_12 ), .\REG.mem_44_12 (\REG.mem_44_12 ), 
            .\REG.mem_46_15 (\REG.mem_46_15 ), .\REG.mem_47_15 (\REG.mem_47_15 ), 
            .\REG.mem_18_3 (\REG.mem_18_3 ), .\REG.mem_19_3 (\REG.mem_19_3 ), 
            .n5255(n5255), .\fifo_data_out[9] (fifo_data_out[9]), .n5252(n5252), 
            .\fifo_data_out[8] (fifo_data_out[8]), .n5249(n5249), .\fifo_data_out[7] (fifo_data_out[7]), 
            .\REG.mem_45_15 (\REG.mem_45_15 ), .\REG.mem_44_15 (\REG.mem_44_15 ), 
            .n4160(n4160), .\REG.mem_2_6 (\REG.mem_2_6 ), .\REG.mem_14_11 (\REG.mem_14_11 ), 
            .\REG.mem_15_11 (\REG.mem_15_11 ), .n4159(n4159), .\REG.mem_2_5 (\REG.mem_2_5 ), 
            .n5236(n5236), .\fifo_data_out[6] (fifo_data_out[6]), .n5233(n5233), 
            .\fifo_data_out[5] (fifo_data_out[5]), .\REG.mem_13_11 (\REG.mem_13_11 ), 
            .\REG.mem_12_11 (\REG.mem_12_11 ), .n5230(n5230), .\fifo_data_out[4] (fifo_data_out[4]), 
            .\wr_grey_sync_r[5] (wr_grey_sync_r[5]), .\wr_grey_sync_r[4] (wr_grey_sync_r[4]), 
            .\wr_grey_sync_r[3] (wr_grey_sync_r[3]), .n5212(n5212), .\fifo_data_out[3] (fifo_data_out[3]), 
            .\REG.mem_18_2 (\REG.mem_18_2 ), .\REG.mem_19_2 (\REG.mem_19_2 ), 
            .n5208(n5208), .n5207(n5207), .\REG.mem_62_14 (\REG.mem_62_14 ), 
            .n5206(n5206), .\REG.mem_62_13 (\REG.mem_62_13 ), .n5205(n5205), 
            .\REG.mem_62_12 (\REG.mem_62_12 ), .n5204(n5204), .\REG.mem_62_11 (\REG.mem_62_11 ), 
            .n5203(n5203), .n5202(n5202), .\REG.mem_62_9 (\REG.mem_62_9 ), 
            .n5201(n5201), .n5200(n5200), .\wr_grey_sync_r[2] (wr_grey_sync_r[2]), 
            .\wr_grey_sync_r[1] (wr_grey_sync_r[1]), .n5199(n5199), .\REG.mem_62_6 (\REG.mem_62_6 ), 
            .n5198(n5198), .n5197(n5197), .n5196(n5196), .n5195(n5195), 
            .n5194(n5194), .\REG.mem_62_1 (\REG.mem_62_1 ), .n5193(n5193), 
            .\REG.mem_62_0 (\REG.mem_62_0 ), .n5192(n5192), .n5191(n5191), 
            .\REG.mem_61_14 (\REG.mem_61_14 ), .n5190(n5190), .\REG.mem_61_13 (\REG.mem_61_13 ), 
            .n5189(n5189), .\REG.mem_61_12 (\REG.mem_61_12 ), .n5188(n5188), 
            .\REG.mem_61_11 (\REG.mem_61_11 ), .n5187(n5187), .n5186(n5186), 
            .\REG.mem_61_9 (\REG.mem_61_9 ), .n5185(n5185), .n5184(n5184), 
            .n5183(n5183), .\REG.mem_61_6 (\REG.mem_61_6 ), .\REG.mem_22_3 (\REG.mem_22_3 ), 
            .\REG.mem_23_3 (\REG.mem_23_3 ), .\REG.mem_26_8 (\REG.mem_26_8 ), 
            .n5182(n5182), .\REG.mem_21_3 (\REG.mem_21_3 ), .n5181(n5181), 
            .n5180(n5180), .n5179(n5179), .n5178(n5178), .\REG.mem_61_1 (\REG.mem_61_1 ), 
            .n5177(n5177), .\REG.mem_61_0 (\REG.mem_61_0 ), .n5176(n5176), 
            .n5175(n5175), .\REG.mem_60_14 (\REG.mem_60_14 ), .n5174(n5174), 
            .\REG.mem_60_13 (\REG.mem_60_13 ), .n5173(n5173), .\REG.mem_60_12 (\REG.mem_60_12 ), 
            .n5172(n5172), .\REG.mem_60_11 (\REG.mem_60_11 ), .n5171(n5171), 
            .n5170(n5170), .\REG.mem_60_9 (\REG.mem_60_9 ), .n5169(n5169), 
            .n5168(n5168), .n5167(n5167), .\REG.mem_60_6 (\REG.mem_60_6 ), 
            .\REG.mem_25_8 (\REG.mem_25_8 ), .\REG.mem_24_8 (\REG.mem_24_8 ), 
            .\REG.mem_46_9 (\REG.mem_46_9 ), .\REG.mem_47_9 (\REG.mem_47_9 ), 
            .\REG.mem_45_9 (\REG.mem_45_9 ), .\REG.mem_44_9 (\REG.mem_44_9 ), 
            .\REG.mem_30_7 (\REG.mem_30_7 ), .n5166(n5166), .n5165(n5165), 
            .n5164(n5164), .n5163(n5163), .n5162(n5162), .\REG.mem_60_1 (\REG.mem_60_1 ), 
            .n5161(n5161), .\REG.mem_60_0 (\REG.mem_60_0 ), .\REG.mem_29_7 (\REG.mem_29_7 ), 
            .\REG.mem_28_7 (\REG.mem_28_7 ), .n5144(n5144), .n5143(n5143), 
            .\REG.mem_58_14 (\REG.mem_58_14 ), .n5142(n5142), .n5141(n5141), 
            .\REG.mem_58_12 (\REG.mem_58_12 ), .n5140(n5140), .n5139(n5139), 
            .n5138(n5138), .\REG.mem_58_9 (\REG.mem_58_9 ), .n5137(n5137), 
            .n5136(n5136), .n5135(n5135), .\REG.mem_58_6 (\REG.mem_58_6 ), 
            .\REG.mem_46_10 (\REG.mem_46_10 ), .\REG.mem_47_10 (\REG.mem_47_10 ), 
            .\REG.mem_45_10 (\REG.mem_45_10 ), .\REG.mem_44_10 (\REG.mem_44_10 ), 
            .n5134(n5134), .\REG.mem_58_5 (\REG.mem_58_5 ), .\REG.mem_30_9 (\REG.mem_30_9 ), 
            .n5133(n5133), .n5132(n5132), .n5131(n5131), .\REG.mem_58_2 (\REG.mem_58_2 ), 
            .n5130(n5130), .\REG.mem_58_1 (\REG.mem_58_1 ), .n5129(n5129), 
            .\REG.mem_58_0 (\REG.mem_58_0 ), .n5128(n5128), .n5127(n5127), 
            .\REG.mem_57_14 (\REG.mem_57_14 ), .n5126(n5126), .n5125(n5125), 
            .\REG.mem_57_12 (\REG.mem_57_12 ), .n5124(n5124), .n5123(n5123), 
            .n5122(n5122), .\REG.mem_57_9 (\REG.mem_57_9 ), .n5121(n5121), 
            .n5120(n5120), .n5119(n5119), .\REG.mem_57_6 (\REG.mem_57_6 ), 
            .\REG.mem_29_9 (\REG.mem_29_9 ), .\REG.mem_28_9 (\REG.mem_28_9 ), 
            .n5118(n5118), .\REG.mem_57_5 (\REG.mem_57_5 ), .n5117(n5117), 
            .n5116(n5116), .n5115(n5115), .\REG.mem_57_2 (\REG.mem_57_2 ), 
            .n5114(n5114), .\REG.mem_57_1 (\REG.mem_57_1 ), .n5113(n5113), 
            .\fifo_data_out[2] (fifo_data_out[2]), .n5110(n5110), .\REG.mem_57_0 (\REG.mem_57_0 ), 
            .n5109(n5109), .n5108(n5108), .\REG.mem_56_14 (\REG.mem_56_14 ), 
            .n5107(n5107), .n5106(n5106), .\REG.mem_56_12 (\REG.mem_56_12 ), 
            .n5105(n5105), .n5104(n5104), .n5103(n5103), .\REG.mem_56_9 (\REG.mem_56_9 ), 
            .\REG.mem_10_6 (\REG.mem_10_6 ), .\REG.mem_11_6 (\REG.mem_11_6 ), 
            .n5102(n5102), .\REG.mem_9_6 (\REG.mem_9_6 ), .\REG.mem_8_6 (\REG.mem_8_6 ), 
            .n5101(n5101), .n5100(n5100), .\REG.mem_56_6 (\REG.mem_56_6 ), 
            .n5099(n5099), .\REG.mem_56_5 (\REG.mem_56_5 ), .n5098(n5098), 
            .n5097(n5097), .n5096(n5096), .\REG.mem_56_2 (\REG.mem_56_2 ), 
            .n5095(n5095), .\REG.mem_56_1 (\REG.mem_56_1 ), .n5094(n5094), 
            .\fifo_data_out[1] (fifo_data_out[1]), .n5091(n5091), .\REG.mem_56_0 (\REG.mem_56_0 ), 
            .n5090(n5090), .\REG.mem_55_15 (\REG.mem_55_15 ), .n5089(n5089), 
            .\REG.mem_55_14 (\REG.mem_55_14 ), .n5088(n5088), .\REG.mem_55_13 (\REG.mem_55_13 ), 
            .n5087(n5087), .\REG.mem_55_12 (\REG.mem_55_12 ), .\REG.mem_22_2 (\REG.mem_22_2 ), 
            .\REG.mem_23_2 (\REG.mem_23_2 ), .\REG.mem_21_2 (\REG.mem_21_2 ), 
            .n5086(n5086), .\REG.mem_55_11 (\REG.mem_55_11 ), .n5085(n5085), 
            .\REG.mem_55_10 (\REG.mem_55_10 ), .n5084(n5084), .n5083(n5083), 
            .n5082(n5082), .\REG.mem_55_7 (\REG.mem_55_7 ), .n5081(n5081), 
            .\REG.mem_55_6 (\REG.mem_55_6 ), .n5080(n5080), .\REG.mem_55_5 (\REG.mem_55_5 ), 
            .n5079(n5079), .\REG.mem_55_4 (\REG.mem_55_4 ), .n5078(n5078), 
            .n5077(n5077), .\REG.mem_55_2 (\REG.mem_55_2 ), .n5076(n5076), 
            .\REG.mem_55_1 (\REG.mem_55_1 ), .n5075(n5075), .\REG.mem_55_0 (\REG.mem_55_0 ), 
            .n5074(n5074), .\REG.mem_54_15 (\REG.mem_54_15 ), .n5073(n5073), 
            .\REG.mem_54_14 (\REG.mem_54_14 ), .n5072(n5072), .\REG.mem_54_13 (\REG.mem_54_13 ), 
            .\num_words_in_buffer[6] (num_words_in_buffer[6]), .\num_words_in_buffer[5] (num_words_in_buffer[5]), 
            .\num_words_in_buffer[4] (num_words_in_buffer[4]), .n5071(n5071), 
            .\REG.mem_54_12 (\REG.mem_54_12 ), .n5070(n5070), .\REG.mem_54_11 (\REG.mem_54_11 ), 
            .n5069(n5069), .\REG.mem_54_10 (\REG.mem_54_10 ), .n5068(n5068), 
            .n5067(n5067), .n5066(n5066), .\REG.mem_54_7 (\REG.mem_54_7 ), 
            .n5065(n5065), .\REG.mem_54_6 (\REG.mem_54_6 ), .n5064(n5064), 
            .\REG.mem_54_5 (\REG.mem_54_5 ), .n5063(n5063), .\REG.mem_54_4 (\REG.mem_54_4 ), 
            .n5062(n5062), .n5061(n5061), .\REG.mem_54_2 (\REG.mem_54_2 ), 
            .n5060(n5060), .\REG.mem_54_1 (\REG.mem_54_1 ), .n5057(n5057), 
            .\REG.mem_54_0 (\REG.mem_54_0 ), .n5056(n5056), .\REG.mem_53_15 (\REG.mem_53_15 ), 
            .n5055(n5055), .\REG.mem_53_14 (\REG.mem_53_14 ), .\REG.mem_50_12 (\REG.mem_50_12 ), 
            .\REG.mem_51_12 (\REG.mem_51_12 ), .\REG.mem_38_5 (\REG.mem_38_5 ), 
            .\REG.mem_39_5 (\REG.mem_39_5 ), .\REG.mem_37_5 (\REG.mem_37_5 ), 
            .n5054(n5054), .\REG.mem_53_13 (\REG.mem_53_13 ), .n5053(n5053), 
            .\REG.mem_53_12 (\REG.mem_53_12 ), .n5052(n5052), .\REG.mem_53_11 (\REG.mem_53_11 ), 
            .n5051(n5051), .\REG.mem_53_10 (\REG.mem_53_10 ), .n5050(n5050), 
            .n5049(n5049), .n5048(n5048), .\REG.mem_53_7 (\REG.mem_53_7 ), 
            .n5047(n5047), .\REG.mem_53_6 (\REG.mem_53_6 ), .n5046(n5046), 
            .\REG.mem_53_5 (\REG.mem_53_5 ), .n5045(n5045), .\REG.mem_53_4 (\REG.mem_53_4 ), 
            .n5044(n5044), .n5043(n5043), .\REG.mem_53_2 (\REG.mem_53_2 ), 
            .n5042(n5042), .\REG.mem_53_1 (\REG.mem_53_1 ), .n5041(n5041), 
            .\REG.mem_53_0 (\REG.mem_53_0 ), .\REG.mem_26_2 (\REG.mem_26_2 ), 
            .\REG.mem_18_11 (\REG.mem_18_11 ), .\REG.mem_19_11 (\REG.mem_19_11 ), 
            .\REG.mem_25_2 (\REG.mem_25_2 ), .\REG.mem_24_2 (\REG.mem_24_2 ), 
            .n5024(n5024), .\REG.mem_51_15 (\REG.mem_51_15 ), .n5023(n5023), 
            .\REG.mem_51_14 (\REG.mem_51_14 ), .n26(n26), .\REG.mem_26_3 (\REG.mem_26_3 ), 
            .\REG.mem_25_3 (\REG.mem_25_3 ), .\REG.mem_24_3 (\REG.mem_24_3 ), 
            .\REG.mem_40_4 (\REG.mem_40_4 ), .\REG.mem_41_4 (\REG.mem_41_4 ), 
            .n5022(n5022), .\REG.mem_51_13 (\REG.mem_51_13 ), .n5021(n5021), 
            .n5020(n5020), .\REG.mem_51_11 (\REG.mem_51_11 ), .n5019(n5019), 
            .\REG.mem_51_10 (\REG.mem_51_10 ), .n5018(n5018), .\REG.mem_51_9 (\REG.mem_51_9 ), 
            .n5017(n5017), .n5016(n5016), .\REG.mem_51_7 (\REG.mem_51_7 ), 
            .n5015(n5015), .\REG.mem_51_6 (\REG.mem_51_6 ), .n5014(n5014), 
            .\REG.mem_51_5 (\REG.mem_51_5 ), .n5013(n5013), .\REG.mem_51_4 (\REG.mem_51_4 ), 
            .n5012(n5012), .n5011(n5011), .\REG.mem_51_2 (\REG.mem_51_2 ), 
            .n5010(n5010), .\REG.mem_51_1 (\REG.mem_51_1 ), .n5008(n5008), 
            .\REG.mem_51_0 (\REG.mem_51_0 ), .\REG.mem_42_4 (\REG.mem_42_4 ), 
            .\REG.mem_43_4 (\REG.mem_43_4 ), .\REG.mem_22_11 (\REG.mem_22_11 ), 
            .\REG.mem_23_11 (\REG.mem_23_11 ), .n5007(n5007), .\REG.mem_50_15 (\REG.mem_50_15 ), 
            .n5006(n5006), .\REG.mem_50_14 (\REG.mem_50_14 ), .n5005(n5005), 
            .\REG.mem_50_13 (\REG.mem_50_13 ), .n5004(n5004), .n5003(n5003), 
            .\REG.mem_50_11 (\REG.mem_50_11 ), .n5002(n5002), .\REG.mem_50_10 (\REG.mem_50_10 ), 
            .n5001(n5001), .\REG.mem_50_9 (\REG.mem_50_9 ), .n5000(n5000), 
            .n4999(n4999), .\REG.mem_50_7 (\REG.mem_50_7 ), .n4998(n4998), 
            .\REG.mem_50_6 (\REG.mem_50_6 ), .n4997(n4997), .\REG.mem_50_5 (\REG.mem_50_5 ), 
            .n4996(n4996), .\REG.mem_50_4 (\REG.mem_50_4 ), .n4995(n4995), 
            .n4994(n4994), .\REG.mem_50_2 (\REG.mem_50_2 ), .n4993(n4993), 
            .\REG.mem_50_1 (\REG.mem_50_1 ), .n4992(n4992), .\REG.mem_50_0 (\REG.mem_50_0 ), 
            .\REG.mem_21_11 (\REG.mem_21_11 ), .\rd_addr_nxt_c_6__N_176[1] (rd_addr_nxt_c_6__N_176[1]), 
            .n4158(n4158), .\REG.mem_2_4 (\REG.mem_2_4 ), .\REG.mem_30_15 (\REG.mem_30_15 ), 
            .\REG.mem_29_15 (\REG.mem_29_15 ), .\REG.mem_28_15 (\REG.mem_28_15 ), 
            .\REG.mem_30_8 (\REG.mem_30_8 ), .\REG.mem_29_8 (\REG.mem_29_8 ), 
            .\REG.mem_28_8 (\REG.mem_28_8 ), .\REG.mem_46_4 (\REG.mem_46_4 ), 
            .\REG.mem_47_4 (\REG.mem_47_4 ), .n4946(n4946), .n4945(n4945), 
            .\REG.mem_47_14 (\REG.mem_47_14 ), .n4944(n4944), .\REG.mem_47_13 (\REG.mem_47_13 ), 
            .\rd_grey_sync_r[5] (rd_grey_sync_r[5]), .\rd_grey_sync_r[4] (rd_grey_sync_r[4]), 
            .\rd_grey_sync_r[3] (rd_grey_sync_r[3]), .\rd_grey_sync_r[2] (rd_grey_sync_r[2]), 
            .\rd_grey_sync_r[1] (rd_grey_sync_r[1]), .n4943(n4943), .\REG.mem_44_4 (\REG.mem_44_4 ), 
            .\REG.mem_45_4 (\REG.mem_45_4 ), .n4942(n4942), .\REG.mem_47_11 (\REG.mem_47_11 ), 
            .n4941(n4941), .n4940(n4940), .n4939(n4939), .n4938(n4938), 
            .\REG.mem_47_7 (\REG.mem_47_7 ), .n4937(n4937), .n4936(n4936), 
            .\REG.mem_47_5 (\REG.mem_47_5 ), .n4935(n4935), .n4934(n4934), 
            .\REG.mem_47_3 (\REG.mem_47_3 ), .n4933(n4933), .\REG.mem_47_2 (\REG.mem_47_2 ), 
            .n4932(n4932), .\REG.mem_47_1 (\REG.mem_47_1 ), .n4929(n4929), 
            .n4928(n4928), .n4927(n4927), .\REG.mem_46_14 (\REG.mem_46_14 ), 
            .\wr_addr_r[6] (wr_addr_r[6]), .n4926(n4926), .\REG.mem_46_13 (\REG.mem_46_13 ), 
            .n4925(n4925), .n4924(n4924), .\REG.mem_46_11 (\REG.mem_46_11 ), 
            .n4923(n4923), .n4922(n4922), .n4921(n4921), .n4920(n4920), 
            .\REG.mem_46_7 (\REG.mem_46_7 ), .n4919(n4919), .n4918(n4918), 
            .\REG.mem_46_5 (\REG.mem_46_5 ), .n4917(n4917), .n4916(n4916), 
            .\REG.mem_46_3 (\REG.mem_46_3 ), .n4915(n4915), .\REG.mem_46_2 (\REG.mem_46_2 ), 
            .n4914(n4914), .\REG.mem_46_1 (\REG.mem_46_1 ), .n4913(n4913), 
            .n4912(n4912), .n4911(n4911), .\REG.mem_45_14 (\REG.mem_45_14 ), 
            .n59(n59), .n4910(n4910), .\REG.mem_45_13 (\REG.mem_45_13 ), 
            .n4909(n4909), .n4908(n4908), .\REG.mem_45_11 (\REG.mem_45_11 ), 
            .n4907(n4907), .n4906(n4906), .n4905(n4905), .n4904(n4904), 
            .\REG.mem_45_7 (\REG.mem_45_7 ), .n4903(n4903), .n4902(n4902), 
            .\REG.mem_45_5 (\REG.mem_45_5 ), .n4901(n4901), .n4900(n4900), 
            .\REG.mem_45_3 (\REG.mem_45_3 ), .n4899(n4899), .\REG.mem_45_2 (\REG.mem_45_2 ), 
            .n4898(n4898), .\REG.mem_45_1 (\REG.mem_45_1 ), .n4897(n4897), 
            .n4896(n4896), .n27(n27), .n4895(n4895), .\REG.mem_44_14 (\REG.mem_44_14 ), 
            .n4894(n4894), .\REG.mem_44_13 (\REG.mem_44_13 ), .n4893(n4893), 
            .n4892(n4892), .\REG.mem_44_11 (\REG.mem_44_11 ), .n4891(n4891), 
            .n4890(n4890), .n4889(n4889), .n4888(n4888), .\REG.mem_44_7 (\REG.mem_44_7 ), 
            .n4887(n4887), .n4886(n4886), .\REG.mem_44_5 (\REG.mem_44_5 ), 
            .n4885(n4885), .n4884(n4884), .\REG.mem_44_3 (\REG.mem_44_3 ), 
            .n4883(n4883), .\REG.mem_44_2 (\REG.mem_44_2 ), .n4882(n4882), 
            .\REG.mem_44_1 (\REG.mem_44_1 ), .n4880(n4880), .n4879(n4879), 
            .n4878(n4878), .n4877(n4877), .\REG.mem_43_13 (\REG.mem_43_13 ), 
            .n4876(n4876), .n4875(n4875), .\REG.mem_43_11 (\REG.mem_43_11 ), 
            .n4874(n4874), .n4873(n4873), .n4872(n4872), .\REG.mem_43_8 (\REG.mem_43_8 ), 
            .n4871(n4871), .\REG.mem_43_7 (\REG.mem_43_7 ), .n4870(n4870), 
            .\REG.mem_43_6 (\REG.mem_43_6 ), .n4869(n4869), .\REG.mem_43_5 (\REG.mem_43_5 ), 
            .n4868(n4868), .n4867(n4867), .\REG.mem_43_3 (\REG.mem_43_3 ), 
            .n4866(n4866), .\REG.mem_43_2 (\REG.mem_43_2 ), .n4865(n4865), 
            .\REG.mem_43_1 (\REG.mem_43_1 ), .n4864(n4864), .\REG.mem_43_0 (\REG.mem_43_0 ), 
            .n4863(n4863), .\REG.mem_30_2 (\REG.mem_30_2 ), .n4862(n4862), 
            .n4861(n4861), .\REG.mem_42_13 (\REG.mem_42_13 ), .n4860(n4860), 
            .n4859(n4859), .\REG.mem_42_11 (\REG.mem_42_11 ), .n4858(n4858), 
            .n4857(n4857), .n4856(n4856), .\REG.mem_42_8 (\REG.mem_42_8 ), 
            .n4855(n4855), .\REG.mem_42_7 (\REG.mem_42_7 ), .n4854(n4854), 
            .\REG.mem_42_6 (\REG.mem_42_6 ), .n4853(n4853), .\REG.mem_42_5 (\REG.mem_42_5 ), 
            .n4852(n4852), .n4851(n4851), .\REG.mem_42_3 (\REG.mem_42_3 ), 
            .n4850(n4850), .\REG.mem_42_2 (\REG.mem_42_2 ), .n4849(n4849), 
            .\REG.mem_42_1 (\REG.mem_42_1 ), .n4848(n4848), .\REG.mem_42_0 (\REG.mem_42_0 ), 
            .n4847(n4847), .\REG.mem_29_2 (\REG.mem_29_2 ), .\REG.mem_28_2 (\REG.mem_28_2 ), 
            .\REG.mem_26_11 (\REG.mem_26_11 ), .\REG.mem_6_7 (\REG.mem_6_7 ), 
            .\REG.mem_7_7 (\REG.mem_7_7 ), .\REG.mem_5_7 (\REG.mem_5_7 ), 
            .n4846(n4846), .n4845(n4845), .\REG.mem_41_13 (\REG.mem_41_13 ), 
            .n4844(n4844), .n4843(n4843), .\REG.mem_41_11 (\REG.mem_41_11 ), 
            .n4842(n4842), .n4841(n4841), .n4840(n4840), .\REG.mem_41_8 (\REG.mem_41_8 ), 
            .n4839(n4839), .\REG.mem_41_7 (\REG.mem_41_7 ), .n4838(n4838), 
            .\REG.mem_41_6 (\REG.mem_41_6 ), .n4837(n4837), .\REG.mem_41_5 (\REG.mem_41_5 ), 
            .n4836(n4836), .n4835(n4835), .\REG.mem_41_3 (\REG.mem_41_3 ), 
            .n4834(n4834), .\REG.mem_41_2 (\REG.mem_41_2 ), .n4833(n4833), 
            .\REG.mem_41_1 (\REG.mem_41_1 ), .n4832(n4832), .\REG.mem_41_0 (\REG.mem_41_0 ), 
            .\REG.mem_18_7 (\REG.mem_18_7 ), .\REG.mem_19_7 (\REG.mem_19_7 ), 
            .\REG.mem_25_11 (\REG.mem_25_11 ), .\REG.mem_24_11 (\REG.mem_24_11 ), 
            .n4157(n4157), .n4831(n4831), .n4830(n4830), .n4829(n4829), 
            .\REG.mem_40_13 (\REG.mem_40_13 ), .n4828(n4828), .n4827(n4827), 
            .\REG.mem_40_11 (\REG.mem_40_11 ), .n4826(n4826), .n4825(n4825), 
            .n4824(n4824), .\REG.mem_40_8 (\REG.mem_40_8 ), .n4823(n4823), 
            .\REG.mem_40_7 (\REG.mem_40_7 ), .n4822(n4822), .\REG.mem_40_6 (\REG.mem_40_6 ), 
            .n4821(n4821), .\REG.mem_40_5 (\REG.mem_40_5 ), .n4820(n4820), 
            .n4819(n4819), .\REG.mem_40_3 (\REG.mem_40_3 ), .n4818(n4818), 
            .\REG.mem_40_2 (\REG.mem_40_2 ), .n4817(n4817), .\REG.mem_40_1 (\REG.mem_40_1 ), 
            .n4814(n4814), .\REG.mem_40_0 (\REG.mem_40_0 ), .n4813(n4813), 
            .\REG.mem_39_15 (\REG.mem_39_15 ), .n4812(n4812), .\REG.mem_39_14 (\REG.mem_39_14 ), 
            .\REG.mem_22_7 (\REG.mem_22_7 ), .\REG.mem_23_7 (\REG.mem_23_7 ), 
            .n4811(n4811), .\REG.mem_39_13 (\REG.mem_39_13 ), .n4810(n4810), 
            .n4809(n4809), .\REG.mem_39_11 (\REG.mem_39_11 ), .\REG.mem_21_7 (\REG.mem_21_7 ), 
            .n4808(n4808), .\REG.mem_30_11 (\REG.mem_30_11 ), .n4807(n4807), 
            .n4806(n4806), .\REG.mem_39_8 (\REG.mem_39_8 ), .n4805(n4805), 
            .n4804(n4804), .\REG.mem_39_6 (\REG.mem_39_6 ), .n4803(n4803), 
            .n4802(n4802), .\REG.mem_39_4 (\REG.mem_39_4 ), .n4801(n4801), 
            .\REG.mem_39_3 (\REG.mem_39_3 ), .n4800(n4800), .\REG.mem_39_2 (\REG.mem_39_2 ), 
            .n4799(n4799), .\REG.mem_39_1 (\REG.mem_39_1 ), .n4798(n4798), 
            .\REG.mem_39_0 (\REG.mem_39_0 ), .n4797(n4797), .\REG.mem_38_15 (\REG.mem_38_15 ), 
            .n4796(n4796), .\REG.mem_38_14 (\REG.mem_38_14 ), .n4795(n4795), 
            .\REG.mem_38_13 (\REG.mem_38_13 ), .n4794(n4794), .n4793(n4793), 
            .\REG.mem_38_11 (\REG.mem_38_11 ), .\REG.mem_29_11 (\REG.mem_29_11 ), 
            .\REG.mem_28_11 (\REG.mem_28_11 ), .n4792(n4792), .\REG.mem_34_2 (\REG.mem_34_2 ), 
            .n4791(n4791), .n4790(n4790), .\REG.mem_38_8 (\REG.mem_38_8 ), 
            .n4789(n4789), .n4788(n4788), .\REG.mem_38_6 (\REG.mem_38_6 ), 
            .n4787(n4787), .n4786(n4786), .\REG.mem_38_4 (\REG.mem_38_4 ), 
            .n4785(n4785), .\REG.mem_38_3 (\REG.mem_38_3 ), .n4784(n4784), 
            .\REG.mem_38_2 (\REG.mem_38_2 ), .n4783(n4783), .\REG.mem_38_1 (\REG.mem_38_1 ), 
            .n4782(n4782), .\REG.mem_38_0 (\REG.mem_38_0 ), .n4781(n4781), 
            .\REG.mem_37_15 (\REG.mem_37_15 ), .n4780(n4780), .\REG.mem_37_14 (\REG.mem_37_14 ), 
            .n4779(n4779), .\REG.mem_37_13 (\REG.mem_37_13 ), .n4778(n4778), 
            .n4777(n4777), .\REG.mem_37_11 (\REG.mem_37_11 ), .n4776(n4776), 
            .n4775(n4775), .n4774(n4774), .\REG.mem_37_8 (\REG.mem_37_8 ), 
            .n4773(n4773), .n4772(n4772), .\REG.mem_37_6 (\REG.mem_37_6 ), 
            .n4771(n4771), .n4770(n4770), .\REG.mem_37_4 (\REG.mem_37_4 ), 
            .n4769(n4769), .\REG.mem_37_3 (\REG.mem_37_3 ), .n4768(n4768), 
            .\REG.mem_37_2 (\REG.mem_37_2 ), .n4767(n4767), .\REG.mem_37_1 (\REG.mem_37_1 ), 
            .n4766(n4766), .\REG.mem_37_0 (\REG.mem_37_0 ), .n4156(n4156), 
            .\REG.mem_26_6 (\REG.mem_26_6 ), .\REG.mem_25_6 (\REG.mem_25_6 ), 
            .\REG.mem_24_6 (\REG.mem_24_6 ), .\REG.mem_34_9 (\REG.mem_34_9 ), 
            .n4733(n4733), .\REG.mem_34_15 (\REG.mem_34_15 ), .n4732(n4732), 
            .\REG.mem_34_14 (\REG.mem_34_14 ), .n4731(n4731), .\REG.mem_34_13 (\REG.mem_34_13 ), 
            .n4730(n4730), .n4729(n4729), .\REG.mem_34_11 (\REG.mem_34_11 ), 
            .n4728(n4728), .n4727(n4727), .n4726(n4726), .\REG.mem_34_8 (\REG.mem_34_8 ), 
            .n4725(n4725), .n4155(n4155), .\REG.mem_2_1 (\REG.mem_2_1 ), 
            .n4154(n4154), .\REG.mem_24_4 (\REG.mem_24_4 ), .\REG.mem_25_4 (\REG.mem_25_4 ), 
            .\REG.mem_26_4 (\REG.mem_26_4 ), .n4724(n4724), .\REG.mem_34_6 (\REG.mem_34_6 ), 
            .\REG.mem_30_4 (\REG.mem_30_4 ), .\REG.mem_28_4 (\REG.mem_28_4 ), 
            .\REG.mem_29_4 (\REG.mem_29_4 ), .n4723(n4723), .n4722(n4722), 
            .\REG.mem_34_4 (\REG.mem_34_4 ), .n4721(n4721), .\REG.mem_34_3 (\REG.mem_34_3 ), 
            .n4720(n4720), .n4719(n4719), .\REG.mem_34_1 (\REG.mem_34_1 ), 
            .n4718(n4718), .\REG.mem_8_4 (\REG.mem_8_4 ), .\REG.mem_9_4 (\REG.mem_9_4 ), 
            .\REG.mem_10_4 (\REG.mem_10_4 ), .\REG.mem_11_4 (\REG.mem_11_4 ), 
            .\REG.mem_14_4 (\REG.mem_14_4 ), .\REG.mem_15_4 (\REG.mem_15_4 ), 
            .\REG.mem_12_4 (\REG.mem_12_4 ), .\REG.mem_13_4 (\REG.mem_13_4 ), 
            .\REG.mem_6_1 (\REG.mem_6_1 ), .\REG.mem_7_1 (\REG.mem_7_1 ), 
            .\REG.mem_5_1 (\REG.mem_5_1 ), .n4677(n4677), .rp_sync1_r({rp_sync1_r}), 
            .\REG.mem_26_10 (\REG.mem_26_10 ), .\REG.mem_18_1 (\REG.mem_18_1 ), 
            .\REG.mem_19_1 (\REG.mem_19_1 ), .n4676(n4676), .n4675(n4675), 
            .n4674(n4674), .n4673(n4673), .n4672(n4672), .\REG.mem_25_10 (\REG.mem_25_10 ), 
            .\REG.mem_24_10 (\REG.mem_24_10 ), .\REG.mem_22_1 (\REG.mem_22_1 ), 
            .\REG.mem_23_1 (\REG.mem_23_1 ), .\REG.mem_21_1 (\REG.mem_21_1 ), 
            .n46(n46), .n14(n14), .n4655(n4655), .n4654(n4654), .n4653(n4653), 
            .n4652(n4652), .n4651(n4651), .n4650(n4650), .n4649(n4649), 
            .n4648(n4648), .n4647(n4647), .\REG.mem_30_13 (\REG.mem_30_13 ), 
            .n4646(n4646), .\REG.mem_30_12 (\REG.mem_30_12 ), .n4645(n4645), 
            .n37(n37), .n5(n5), .n4644(n4644), .n4643(n4643), .n4642(n4642), 
            .n4641(n4641), .n4640(n4640), .\REG.mem_30_6 (\REG.mem_30_6 ), 
            .n4639(n4639), .n4638(n4638), .n4637(n4637), .n4636(n4636), 
            .n4635(n4635), .\REG.mem_30_1 (\REG.mem_30_1 ), .n4634(n4634), 
            .n4633(n4633), .n4631(n4631), .n4629(n4629), .\REG.mem_18_14 (\REG.mem_18_14 ), 
            .\REG.mem_19_14 (\REG.mem_19_14 ), .n4627(n4627), .n51(n51), 
            .n4626(n4626), .n4625(n4625), .\REG.mem_29_13 (\REG.mem_29_13 ), 
            .\REG.mem_22_14 (\REG.mem_22_14 ), .\REG.mem_23_14 (\REG.mem_23_14 ), 
            .\REG.mem_21_14 (\REG.mem_21_14 ), .n4624(n4624), .\REG.mem_29_12 (\REG.mem_29_12 ), 
            .n4623(n4623), .n4622(n4622), .n4621(n4621), .n4620(n4620), 
            .n4619(n4619), .n4618(n4618), .\REG.mem_29_6 (\REG.mem_29_6 ), 
            .n4617(n4617), .n4616(n4616), .n4615(n4615), .n4614(n4614), 
            .n4613(n4613), .\REG.mem_29_1 (\REG.mem_29_1 ), .n4612(n4612), 
            .n4611(n4611), .n4610(n4610), .n4609(n4609), .\REG.mem_28_13 (\REG.mem_28_13 ), 
            .n19(n19), .n4608(n4608), .\REG.mem_28_12 (\REG.mem_28_12 ), 
            .n4607(n4607), .\REG.mem_18_12 (\REG.mem_18_12 ), .\REG.mem_19_12 (\REG.mem_19_12 ), 
            .\REG.mem_22_12 (\REG.mem_22_12 ), .\REG.mem_23_12 (\REG.mem_23_12 ), 
            .n4606(n4606), .n4605(n4605), .n4604(n4604), .n4603(n4603), 
            .n4602(n4602), .\REG.mem_28_6 (\REG.mem_28_6 ), .n4601(n4601), 
            .n4600(n4600), .n4599(n4599), .n4598(n4598), .n4597(n4597), 
            .\REG.mem_28_1 (\REG.mem_28_1 ), .n4596(n4596), .\REG.mem_21_12 (\REG.mem_21_12 ), 
            .n4579(n4579), .n4578(n4578), .n4577(n4577), .\REG.mem_26_13 (\REG.mem_26_13 ), 
            .n4576(n4576), .\REG.mem_26_12 (\REG.mem_26_12 ), .n4575(n4575), 
            .n4574(n4574), .n4573(n4573), .n4572(n4572), .n4571(n4571), 
            .\REG.mem_26_7 (\REG.mem_26_7 ), .n4570(n4570), .n4569(n4569), 
            .n4568(n4568), .n4567(n4567), .\REG.mem_6_13 (\REG.mem_6_13 ), 
            .\REG.mem_7_13 (\REG.mem_7_13 ), .n4566(n4566), .n4565(n4565), 
            .\REG.mem_26_1 (\REG.mem_26_1 ), .n4564(n4564), .\REG.mem_26_0 (\REG.mem_26_0 ), 
            .n4563(n4563), .wp_sync1_r({wp_sync1_r}), .n4562(n4562), .n4561(n4561), 
            .n4560(n4560), .n4559(n4559), .n4558(n4558), .n4557(n4557), 
            .n4556(n4556), .\REG.mem_25_13 (\REG.mem_25_13 ), .n4555(n4555), 
            .\REG.mem_25_12 (\REG.mem_25_12 ), .n4554(n4554), .n4553(n4553), 
            .n4552(n4552), .n4551(n4551), .\REG.mem_5_13 (\REG.mem_5_13 ), 
            .n4550(n4550), .\REG.mem_25_7 (\REG.mem_25_7 ), .n4549(n4549), 
            .n4548(n4548), .n4547(n4547), .n4546(n4546), .n4545(n4545), 
            .n4544(n4544), .\REG.mem_25_1 (\REG.mem_25_1 ), .n4543(n4543), 
            .\REG.mem_25_0 (\REG.mem_25_0 ), .n4542(n4542), .n4541(n4541), 
            .n4540(n4540), .n4539(n4539), .n4538(n4538), .n4537(n4537), 
            .n4536(n4536), .n4535(n4535), .n4534(n4534), .\REG.mem_18_0 (\REG.mem_18_0 ), 
            .\REG.mem_19_0 (\REG.mem_19_0 ), .\REG.mem_22_0 (\REG.mem_22_0 ), 
            .\REG.mem_23_0 (\REG.mem_23_0 ), .\REG.mem_21_0 (\REG.mem_21_0 ), 
            .DEBUG_9_c(DEBUG_9_c), .n4533(n4533), .\REG.mem_24_13 (\REG.mem_24_13 ), 
            .n4532(n4532), .\REG.mem_24_12 (\REG.mem_24_12 ), .n4531(n4531), 
            .n4530(n4530), .n4529(n4529), .n4528(n4528), .n4527(n4527), 
            .\REG.mem_24_7 (\REG.mem_24_7 ), .n4526(n4526), .n4525(n4525), 
            .n4524(n4524), .n4523(n4523), .n4522(n4522), .n4521(n4521), 
            .\REG.mem_24_1 (\REG.mem_24_1 ), .n4520(n4520), .\REG.mem_24_0 (\REG.mem_24_0 ), 
            .n4519(n4519), .\REG.mem_23_15 (\REG.mem_23_15 ), .n4518(n4518), 
            .n4517(n4517), .n4516(n4516), .n4515(n4515), .n4514(n4514), 
            .\REG.mem_23_10 (\REG.mem_23_10 ), .n4513(n4513), .\REG.mem_23_9 (\REG.mem_23_9 ), 
            .n4512(n4512), .n4511(n4511), .n4510(n4510), .n4509(n4509), 
            .n4508(n4508), .\REG.mem_23_4 (\REG.mem_23_4 ), .n4507(n4507), 
            .n4506(n4506), .n4505(n4505), .n4504(n4504), .n4503(n4503), 
            .\REG.mem_22_15 (\REG.mem_22_15 ), .n4502(n4502), .n4501(n4501), 
            .n4500(n4500), .n4499(n4499), .n4498(n4498), .\REG.mem_22_10 (\REG.mem_22_10 ), 
            .n4497(n4497), .\REG.mem_22_9 (\REG.mem_22_9 ), .n4496(n4496), 
            .n4495(n4495), .n4494(n4494), .n4493(n4493), .n4492(n4492), 
            .\REG.mem_22_4 (\REG.mem_22_4 ), .n4491(n4491), .n4490(n4490), 
            .n4489(n4489), .n4488(n4488), .n4487(n4487), .\REG.mem_21_15 (\REG.mem_21_15 ), 
            .n4486(n4486), .n4485(n4485), .n4484(n4484), .n4483(n4483), 
            .n4482(n4482), .\REG.mem_21_10 (\REG.mem_21_10 ), .n4481(n4481), 
            .\REG.mem_21_9 (\REG.mem_21_9 ), .n4480(n4480), .n4479(n4479), 
            .n4478(n4478), .n4477(n4477), .n4476(n4476), .\REG.mem_21_4 (\REG.mem_21_4 ), 
            .n4475(n4475), .n4474(n4474), .n4473(n4473), .\REG.mem_6_12 (\REG.mem_6_12 ), 
            .\REG.mem_7_12 (\REG.mem_7_12 ), .n4472(n4472), .\REG.out_raw[15] (\REG.out_raw [15]), 
            .\REG.out_raw[14] (\REG.out_raw [14]), .\REG.out_raw[13] (\REG.out_raw [13]), 
            .\REG.mem_5_12 (\REG.mem_5_12 ), .\REG.out_raw[12] (\REG.out_raw [12]), 
            .\REG.out_raw[11] (\REG.out_raw [11]), .\REG.out_raw[10] (\REG.out_raw [10]), 
            .n4455(n4455), .\REG.mem_19_15 (\REG.mem_19_15 ), .n4454(n4454), 
            .n4453(n4453), .n4452(n4452), .n4451(n4451), .n4450(n4450), 
            .n4449(n4449), .\REG.mem_19_9 (\REG.mem_19_9 ), .n4448(n4448), 
            .n4447(n4447), .n4446(n4446), .n4445(n4445), .n4444(n4444), 
            .\REG.mem_19_4 (\REG.mem_19_4 ), .n4443(n4443), .n4442(n4442), 
            .n4441(n4441), .n4440(n4440), .\REG.out_raw[9] (\REG.out_raw [9]), 
            .\REG.out_raw[8] (\REG.out_raw [8]), .n4439(n4439), .\REG.mem_18_15 (\REG.mem_18_15 ), 
            .\REG.out_raw[7] (\REG.out_raw [7]), .\REG.out_raw[6] (\REG.out_raw [6]), 
            .\REG.out_raw[5] (\REG.out_raw [5]), .\REG.out_raw[4] (\REG.out_raw [4]), 
            .\REG.out_raw[3] (\REG.out_raw [3]), .n4438(n4438), .\REG.mem_6_9 (\REG.mem_6_9 ), 
            .\REG.mem_7_9 (\REG.mem_7_9 ), .n54(n54), .\REG.mem_5_9 (\REG.mem_5_9 ), 
            .n4437(n4437), .n4436(n4436), .n4435(n4435), .n4434(n4434), 
            .n4433(n4433), .\REG.mem_18_9 (\REG.mem_18_9 ), .n4432(n4432), 
            .n4431(n4431), .n4430(n4430), .n4429(n4429), .n4428(n4428), 
            .\REG.mem_18_4 (\REG.mem_18_4 ), .n4427(n4427), .n4426(n4426), 
            .n4425(n4425), .n4424(n4424), .\REG.out_raw[2] (\REG.out_raw [2]), 
            .n22(n22), .n39(n39), .\REG.mem_10_9 (\REG.mem_10_9 ), .\REG.mem_11_9 (\REG.mem_11_9 ), 
            .\REG.mem_10_13 (\REG.mem_10_13 ), .\REG.mem_11_13 (\REG.mem_11_13 ), 
            .n7(n7), .n40(n40), .\REG.mem_9_9 (\REG.mem_9_9 ), .\REG.mem_8_9 (\REG.mem_8_9 ), 
            .\REG.mem_9_13 (\REG.mem_9_13 ), .\REG.mem_8_13 (\REG.mem_8_13 ), 
            .n8(n8_adj_1102), .\REG.mem_14_12 (\REG.mem_14_12 ), .\REG.mem_15_12 (\REG.mem_15_12 ), 
            .n4391(n4391), .\REG.out_raw[1] (\REG.out_raw [1]), .n4390(n4390), 
            .\REG.mem_13_12 (\REG.mem_13_12 ), .\REG.mem_12_12 (\REG.mem_12_12 ), 
            .n4389(n4389), .\REG.mem_15_13 (\REG.mem_15_13 ), .n4388(n4388), 
            .n4387(n4387), .n4386(n4386), .\REG.mem_15_10 (\REG.mem_15_10 ), 
            .n4385(n4385), .\REG.mem_15_9 (\REG.mem_15_9 ), .n4384(n4384), 
            .\REG.mem_15_8 (\REG.mem_15_8 ), .n4383(n4383), .\REG.mem_15_7 (\REG.mem_15_7 ), 
            .n4382(n4382), .n4381(n4381), .\REG.mem_15_5 (\REG.mem_15_5 ), 
            .n4380(n4380), .n4379(n4379), .n4378(n4378), .n4377(n4377), 
            .\REG.mem_15_1 (\REG.mem_15_1 ), .n4376(n4376), .n4375(n4375), 
            .n4374(n4374), .\REG.mem_6_8 (\REG.mem_6_8 ), .\REG.mem_7_8 (\REG.mem_7_8 ), 
            .\REG.mem_5_8 (\REG.mem_5_8 ), .\REG.mem_14_9 (\REG.mem_14_9 ), 
            .\REG.mem_13_9 (\REG.mem_13_9 ), .\REG.mem_12_9 (\REG.mem_12_9 ), 
            .\REG.mem_6_5 (\REG.mem_6_5 ), .\REG.mem_7_5 (\REG.mem_7_5 ), 
            .n4373(n4373), .\REG.mem_14_13 (\REG.mem_14_13 ), .n4372(n4372), 
            .n4371(n4371), .n4370(n4370), .\REG.mem_14_10 (\REG.mem_14_10 ), 
            .n4369(n4369), .n4368(n4368), .\REG.mem_14_8 (\REG.mem_14_8 ), 
            .n4367(n4367), .\REG.mem_14_7 (\REG.mem_14_7 ), .\REG.mem_5_5 (\REG.mem_5_5 ), 
            .n4366(n4366), .n4365(n4365), .\REG.mem_14_5 (\REG.mem_14_5 ), 
            .n4364(n4364), .n4363(n4363), .n4362(n4362), .n4361(n4361), 
            .\REG.mem_14_1 (\REG.mem_14_1 ), .n4360(n4360), .n4359(n4359), 
            .n4358(n4358), .n4357(n4357), .\REG.mem_13_13 (\REG.mem_13_13 ), 
            .n4356(n4356), .n4355(n4355), .n4354(n4354), .\REG.mem_13_10 (\REG.mem_13_10 ), 
            .n4353(n4353), .n4352(n4352), .\REG.mem_13_8 (\REG.mem_13_8 ), 
            .n4351(n4351), .\REG.mem_13_7 (\REG.mem_13_7 ), .n4350(n4350), 
            .n4349(n4349), .\REG.mem_13_5 (\REG.mem_13_5 ), .n4348(n4348), 
            .n4347(n4347), .n4346(n4346), .n4345(n4345), .\REG.mem_13_1 (\REG.mem_13_1 ), 
            .n4344(n4344), .n4343(n4343), .n4342(n4342), .n4341(n4341), 
            .\REG.mem_12_13 (\REG.mem_12_13 ), .n4340(n4340), .n4339(n4339), 
            .n4338(n4338), .\REG.mem_12_10 (\REG.mem_12_10 ), .n4337(n4337), 
            .n4336(n4336), .\REG.mem_12_8 (\REG.mem_12_8 ), .n4335(n4335), 
            .\REG.mem_12_7 (\REG.mem_12_7 ), .n4334(n4334), .n4333(n4333), 
            .\REG.mem_12_5 (\REG.mem_12_5 ), .n4332(n4332), .n4331(n4331), 
            .n4330(n4330), .n4329(n4329), .\REG.mem_12_1 (\REG.mem_12_1 ), 
            .n4328(n4328), .n4327(n4327), .n4326(n4326), .n4325(n4325), 
            .n4324(n4324), .n4323(n4323), .n60(n60), .n4322(n4322), 
            .n28(n28), .n41(n41), .n9(n9), .n4321(n4321), .n4320(n4320), 
            .\REG.mem_11_8 (\REG.mem_11_8 ), .n4319(n4319), .\REG.mem_11_7 (\REG.mem_11_7 ), 
            .n4318(n4318), .n4317(n4317), .\REG.mem_11_5 (\REG.mem_11_5 ), 
            .n4316(n4316), .n4315(n4315), .n4314(n4314), .n4313(n4313), 
            .\REG.mem_11_1 (\REG.mem_11_1 ), .n4312(n4312), .n4311(n4311), 
            .n42(n42), .n4310(n4310), .n4309(n4309), .n4308(n4308), 
            .n10(n10), .n4307(n4307), .n4306(n4306), .n4305(n4305), 
            .n4304(n4304), .\REG.mem_10_8 (\REG.mem_10_8 ), .n4303(n4303), 
            .\REG.mem_10_7 (\REG.mem_10_7 ), .n4302(n4302), .n4301(n4301), 
            .\REG.mem_10_5 (\REG.mem_10_5 ), .n4300(n4300), .n4299(n4299), 
            .n4298(n4298), .n4297(n4297), .\REG.mem_10_1 (\REG.mem_10_1 ), 
            .n4296(n4296), .n4130(n4130), .n57(n57), .\REG.mem_9_5 (\REG.mem_9_5 ), 
            .\REG.mem_8_5 (\REG.mem_8_5 ), .n4288(n4288), .n4287(n4287), 
            .n4286(n4286), .n4285(n4285), .n4284(n4284), .n4283(n4283), 
            .n4282(n4282), .n4281(n4281), .n4280(n4280), .\REG.mem_9_8 (\REG.mem_9_8 ), 
            .n4279(n4279), .\REG.mem_9_7 (\REG.mem_9_7 ), .n4278(n4278), 
            .n4277(n4277), .n4108(n4108), .n25(n25), .n4276(n4276), 
            .n43(n43), .n11(n11), .n44(n44), .n12(n12), .n4275(n4275), 
            .n4274(n4274), .n4273(n4273), .\REG.mem_9_1 (\REG.mem_9_1 ), 
            .n4272(n4272), .n4270(n4270), .n4268(n4268), .n4107(n4107), 
            .\REG.mem_8_7 (\REG.mem_8_7 ), .n4265(n4265), .n4264(n4264), 
            .n4263(n4263), .n4262(n4262), .n4261(n4261), .n52(n52), 
            .n4260(n4260), .\REG.mem_8_8 (\REG.mem_8_8 ), .n4259(n4259), 
            .n4258(n4258), .n4257(n4257), .n4256(n4256), .n4255(n4255), 
            .n4254(n4254), .n4253(n4253), .n4252(n4252), .n4251(n4251), 
            .\REG.mem_8_1 (\REG.mem_8_1 ), .n4250(n4250), .n4249(n4249), 
            .n4248(n4248), .n4247(n4247), .n4246(n4246), .n4245(n4245), 
            .\REG.mem_7_11 (\REG.mem_7_11 ), .n4244(n4244), .n4243(n4243), 
            .n4242(n4242), .n4241(n4241), .n4240(n4240), .n4239(n4239), 
            .n4238(n4238), .\REG.mem_7_4 (\REG.mem_7_4 ), .n4237(n4237), 
            .n4236(n4236), .n4235(n4235), .n4234(n4234), .n4233(n4233), 
            .n4232(n4232), .n4231(n4231), .n4230(n4230), .n4229(n4229), 
            .\REG.mem_6_11 (\REG.mem_6_11 ), .n4228(n4228), .n4227(n4227), 
            .n4226(n4226), .n4225(n4225), .n4224(n4224), .n4223(n4223), 
            .n4222(n4222), .\REG.mem_6_4 (\REG.mem_6_4 ), .n4221(n4221), 
            .n4220(n4220), .n4219(n4219), .n4218(n4218), .n4217(n4217), 
            .n4216(n4216), .n4215(n4215), .n4214(n4214), .n4213(n4213), 
            .\REG.mem_5_11 (\REG.mem_5_11 ), .n4212(n4212), .n4211(n4211), 
            .n4210(n4210), .n4209(n4209), .n4208(n4208), .n4207(n4207), 
            .n4206(n4206), .\REG.mem_5_4 (\REG.mem_5_4 ), .n4205(n4205), 
            .n4204(n4204), .n4203(n4203), .n4202(n4202), .n4103(n4103), 
            .n20(n20), .n53(n53), .n4101(n4101), .n21(n21), .n35(n35), 
            .n3(n3), .n36(n36), .n55(n55), .n23(n23), .n4(n4_adj_1101), 
            .n47(n47), .n15(n15_adj_1103), .n31(n31), .n63(n63)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(476[20] 491[2])
    SB_LUT4 i1_4_lut_4_lut (.I0(is_tx_fifo_full_flag), .I1(n9398), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h2222;
    spi spi0 (.SEN_c_1(SEN_c_1), .DEBUG_6_c(DEBUG_6_c), .SOUT_c(SOUT_c), 
        .n3629(n3629), .\rx_shift_reg[0] (rx_shift_reg[0]), .GND_net(GND_net), 
        .multi_byte_spi_trans_flag_r(multi_byte_spi_trans_flag_r), .n9073(n9073), 
        .VCC_net(VCC_net), .\tx_shift_reg[0] (tx_shift_reg[0]), .spi_start_transfer_r(spi_start_transfer_r), 
        .n1638(n1638), .spi_rx_byte_ready(spi_rx_byte_ready), .n4701(n4701), 
        .\rx_shift_reg[1] (rx_shift_reg[1]), .n4699(n4699), .rx_buf_byte({rx_buf_byte}), 
        .n4683(n4683), .n4682(n4682), .n4681(n4681), .n4680(n4680), 
        .n4679(n4679), .n4678(n4678), .n4145(n4145), .\rx_shift_reg[2] (rx_shift_reg[2]), 
        .n4144(n4144), .\rx_shift_reg[3] (rx_shift_reg[3]), .n4137(n4137), 
        .\rx_shift_reg[4] (rx_shift_reg[4]), .n3626(n3626), .SCK_c_0(SCK_c_0), 
        .SDAT_c_15(SDAT_c_15), .n4099(n4099), .n4081(n4081), .\rx_shift_reg[5] (rx_shift_reg[5]), 
        .n4080(n4080), .\rx_shift_reg[6] (rx_shift_reg[6]), .n4079(n4079), 
        .\rx_shift_reg[7] (rx_shift_reg[7]), .tx_addr_byte({tx_addr_byte}), 
        .\tx_data_byte[7] (tx_data_byte[7]), .\tx_data_byte[6] (tx_data_byte[6]), 
        .\tx_data_byte[5] (tx_data_byte[5]), .\tx_data_byte[4] (tx_data_byte[4]), 
        .\tx_data_byte[3] (tx_data_byte[3]), .\tx_data_byte[2] (tx_data_byte[2]), 
        .\tx_data_byte[1] (tx_data_byte[1]), .n2851(n2851)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(791[5] 815[2])
    clock clock_inst (.GND_net(GND_net), .VCC_net(VCC_net), .ICE_SYSCLK_c(ICE_SYSCLK_c), 
          .pll_clk_unbuf(pll_clk_unbuf)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(222[7] 228[3])
    \uart_tx(CLKS_PER_BIT=20)  pc_tx (.DEBUG_6_c(DEBUG_6_c), .UART_TX_c(UART_TX_c), 
            .r_SM_Main({r_SM_Main_adj_1138}), .VCC_net(VCC_net), .n4974(n4974), 
            .r_Tx_Data({r_Tx_Data}), .n4973(n4973), .n4972(n4972), .n4971(n4971), 
            .n4970(n4970), .n4969(n4969), .n4967(n4967), .GND_net(GND_net), 
            .\r_SM_Main_2__N_728[0] (r_SM_Main_2__N_728[0]), .\r_SM_Main_2__N_725[1] (r_SM_Main_2__N_725[1]), 
            .n3151(n3151), .n4091(n4091), .n4090(n4090), .tx_uart_active_flag(tx_uart_active_flag), 
            .n12410(n12410), .n4(n4_adj_1099)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(726[42] 735[3])
    
endmodule
//
// Verilog Description of module timing_controller
//

module timing_controller (state, DEBUG_6_c, \num_words_in_buffer[4] , 
            \num_words_in_buffer[6] , \num_words_in_buffer[5] , \num_words_in_buffer[3] , 
            DEBUG_2_c, n9057, buffer_switch_done, n63, GND_net, n9355, 
            VCC_net, n1326, n1431, n6392, n6602, n6572, n3474, 
            INVERT_c_3, reset_all, UPDATE_c_2) /* synthesis syn_module_defined=1 */ ;
    output [3:0]state;
    input DEBUG_6_c;
    input \num_words_in_buffer[4] ;
    input \num_words_in_buffer[6] ;
    input \num_words_in_buffer[5] ;
    input \num_words_in_buffer[3] ;
    output DEBUG_2_c;
    input n9057;
    output buffer_switch_done;
    output n63;
    input GND_net;
    output n9355;
    input VCC_net;
    input n1326;
    input n1431;
    input n6392;
    input n6602;
    output n6572;
    output n3474;
    output INVERT_c_3;
    output reset_all;
    output UPDATE_c_2;
    
    wire DEBUG_6_c /* synthesis SET_AS_NETWORK=DEBUG_6_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [3:0]state_3__N_313;
    
    wire n9356;
    wire [31:0]n1504;
    
    wire n3668;
    wire [31:0]state_timeout_counter;   // src/timing_controller.v(45[12:33])
    wire [31:0]n1432;
    
    wire n3998;
    wire [31:0]n507;
    
    wire n3984, n9330, n9361;
    wire [3:0]n596;
    
    wire n3830, n10561, n8699, n8700, n10562, n8698, n8710, n8709, 
        n8690, n8691, n8683, n8684, n10567, n8689, n10563, n8697, 
        n10569, n8682, n8696, n8708, n10568, n8688, n8707, n8706, 
        n10571, n8680, n9329, n8695, n8685, n8687, n10582, n1503, 
        n10572, n8705, n8704, n8686, n9338, n10558, n8703, n10564, 
        n8694, n10559, n8702, n10560, n8701, n10570, n8681, n10565, 
        n8693, n10530, n8692, n10566, n5, n1585, n9350, n38, 
        n52, n56, n54, n55, n53, n50, n58, n62, n49, n6606, 
        n7, n10656;
    
    SB_DFFE state_i0 (.Q(state[0]), .C(DEBUG_6_c), .E(n9356), .D(state_3__N_313[0]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[0]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1432[1]), .R(n3998));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1432[2]), .R(n3998));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(DEBUG_6_c), 
            .E(n3668), .D(n507[6]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(DEBUG_6_c), 
            .E(n3668), .D(n507[7]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i8 (.Q(state_timeout_counter[8]), .C(DEBUG_6_c), 
            .E(n3668), .D(n507[8]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i11 (.Q(state_timeout_counter[11]), 
            .C(DEBUG_6_c), .E(n3668), .D(n507[11]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i13 (.Q(state_timeout_counter[13]), 
            .C(DEBUG_6_c), .E(n3668), .D(n507[13]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i16 (.Q(state_timeout_counter[16]), 
            .C(DEBUG_6_c), .E(n3668), .D(n507[16]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i17 (.Q(state_timeout_counter[17]), 
            .C(DEBUG_6_c), .E(n3668), .D(n507[17]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i21 (.Q(state_timeout_counter[21]), 
            .C(DEBUG_6_c), .E(n3668), .D(n507[21]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i25 (.Q(state_timeout_counter[25]), 
            .C(DEBUG_6_c), .E(n3668), .D(n507[25]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_LUT4 i1017_4_lut (.I0(\num_words_in_buffer[4] ), .I1(\num_words_in_buffer[6] ), 
            .I2(\num_words_in_buffer[5] ), .I3(\num_words_in_buffer[3] ), 
            .O(DEBUG_2_c));
    defparam i1017_4_lut.LUT_INIT = 16'hfcec;
    SB_DFF state_i3 (.Q(state[3]), .C(DEBUG_6_c), .D(n9057));   // src/timing_controller.v(59[8] 133[4])
    SB_DFF invert_52_i1 (.Q(buffer_switch_done), .C(DEBUG_6_c), .D(n9330));   // src/timing_controller.v(64[5] 132[12])
    SB_LUT4 i1_2_lut_3_lut (.I0(state[2]), .I1(state[0]), .I2(n63), .I3(GND_net), 
            .O(n9361));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_187_Mux_3_i15_4_lut_4_lut_4_lut (.I0(state[2]), .I1(state[0]), 
            .I2(state[3]), .I3(state[1]), .O(n596[3]));
    defparam mux_187_Mux_3_i15_4_lut_4_lut_4_lut.LUT_INIT = 16'h0a10;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[2]), .I1(state[0]), .I2(n9355), 
            .I3(state[1]), .O(n3830));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hf0f1;
    SB_LUT4 sub_32_add_2_22_lut (.I0(n1326), .I1(state_timeout_counter[20]), 
            .I2(VCC_net), .I3(n8699), .O(n10561)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_32_add_2_22 (.CI(n8699), .I0(state_timeout_counter[20]), 
            .I1(VCC_net), .CO(n8700));
    SB_LUT4 sub_32_add_2_21_lut (.I0(n1326), .I1(state_timeout_counter[19]), 
            .I2(VCC_net), .I3(n8698), .O(n10562)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_32_add_2_21 (.CI(n8698), .I0(state_timeout_counter[19]), 
            .I1(VCC_net), .CO(n8699));
    SB_DFFE state_timeout_counter_i0_i24 (.Q(state_timeout_counter[24]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[24]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i23 (.Q(state_timeout_counter[23]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[23]));   // src/timing_controller.v(59[8] 133[4])
    SB_LUT4 sub_32_add_2_33_lut (.I0(GND_net), .I1(state_timeout_counter[31]), 
            .I2(VCC_net), .I3(n8710), .O(n507[31])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_33_lut.LUT_INIT = 16'hC33C;
    SB_DFFE state_timeout_counter_i0_i22 (.Q(state_timeout_counter[22]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[22]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i20 (.Q(state_timeout_counter[20]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[20]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i19 (.Q(state_timeout_counter[19]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[19]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i18 (.Q(state_timeout_counter[18]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[18]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i15 (.Q(state_timeout_counter[15]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[15]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i14 (.Q(state_timeout_counter[14]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[14]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i12 (.Q(state_timeout_counter[12]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[12]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i10 (.Q(state_timeout_counter[10]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[10]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i9 (.Q(state_timeout_counter[9]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[9]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[5]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[4]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(DEBUG_6_c), 
            .E(n3668), .D(n1504[3]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i26 (.Q(state_timeout_counter[26]), 
            .C(DEBUG_6_c), .E(n3668), .D(n507[26]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_LUT4 sub_32_add_2_32_lut (.I0(GND_net), .I1(state_timeout_counter[30]), 
            .I2(VCC_net), .I3(n8709), .O(n507[30])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_32_add_2_13_lut (.I0(GND_net), .I1(state_timeout_counter[11]), 
            .I2(VCC_net), .I3(n8690), .O(n507[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_32_add_2_13 (.CI(n8690), .I0(state_timeout_counter[11]), 
            .I1(VCC_net), .CO(n8691));
    SB_DFFESR state_timeout_counter_i0_i27 (.Q(state_timeout_counter[27]), 
            .C(DEBUG_6_c), .E(n3668), .D(n507[27]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_CARRY sub_32_add_2_6 (.CI(n8683), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n8684));
    SB_CARRY sub_32_add_2_32 (.CI(n8709), .I0(state_timeout_counter[30]), 
            .I1(VCC_net), .CO(n8710));
    SB_LUT4 sub_32_add_2_12_lut (.I0(n1326), .I1(state_timeout_counter[10]), 
            .I2(VCC_net), .I3(n8689), .O(n10567)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_32_add_2_20_lut (.I0(n1326), .I1(state_timeout_counter[18]), 
            .I2(VCC_net), .I3(n8697), .O(n10563)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_32_add_2_12 (.CI(n8689), .I0(state_timeout_counter[10]), 
            .I1(VCC_net), .CO(n8690));
    SB_CARRY sub_32_add_2_20 (.CI(n8697), .I0(state_timeout_counter[18]), 
            .I1(VCC_net), .CO(n8698));
    SB_LUT4 sub_32_add_2_5_lut (.I0(n1326), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n8682), .O(n10569)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_32_add_2_19_lut (.I0(GND_net), .I1(state_timeout_counter[17]), 
            .I2(VCC_net), .I3(n8696), .O(n507[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_32_add_2_31_lut (.I0(GND_net), .I1(state_timeout_counter[29]), 
            .I2(VCC_net), .I3(n8708), .O(n507[29])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_32_add_2_31 (.CI(n8708), .I0(state_timeout_counter[29]), 
            .I1(VCC_net), .CO(n8709));
    SB_LUT4 sub_32_add_2_11_lut (.I0(n1326), .I1(state_timeout_counter[9]), 
            .I2(VCC_net), .I3(n8688), .O(n10568)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_32_add_2_19 (.CI(n8696), .I0(state_timeout_counter[17]), 
            .I1(VCC_net), .CO(n8697));
    SB_LUT4 sub_32_add_2_30_lut (.I0(GND_net), .I1(state_timeout_counter[28]), 
            .I2(VCC_net), .I3(n8707), .O(n507[28])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_32_add_2_30 (.CI(n8707), .I0(state_timeout_counter[28]), 
            .I1(VCC_net), .CO(n8708));
    SB_CARRY sub_32_add_2_11 (.CI(n8688), .I0(state_timeout_counter[9]), 
            .I1(VCC_net), .CO(n8689));
    SB_LUT4 sub_32_add_2_29_lut (.I0(GND_net), .I1(state_timeout_counter[27]), 
            .I2(VCC_net), .I3(n8706), .O(n507[27])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_32_add_2_3_lut (.I0(n1326), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n8680), .O(n10571)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(state[3]), 
            .I3(state[2]), .O(n9329));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 sub_32_add_2_18_lut (.I0(GND_net), .I1(state_timeout_counter[16]), 
            .I2(VCC_net), .I3(n8695), .O(n507[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_32_add_2_7 (.CI(n8684), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n8685));
    SB_LUT4 i1_2_lut_4_lut_adj_59 (.I0(state[0]), .I1(state[1]), .I2(state[3]), 
            .I3(state[2]), .O(n9330));
    defparam i1_2_lut_4_lut_adj_59.LUT_INIT = 16'h0200;
    SB_LUT4 sub_32_add_2_10_lut (.I0(GND_net), .I1(state_timeout_counter[8]), 
            .I2(VCC_net), .I3(n8687), .O(n507[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_32_add_2_29 (.CI(n8706), .I0(state_timeout_counter[27]), 
            .I1(VCC_net), .CO(n8707));
    SB_CARRY sub_32_add_2_18 (.CI(n8695), .I0(state_timeout_counter[16]), 
            .I1(VCC_net), .CO(n8696));
    SB_LUT4 mux_693_i4_3_lut (.I0(n10569), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[3]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7890_4_lut (.I0(n10582), .I1(state[1]), .I2(n1431), .I3(n1503), 
            .O(n1504[4]));   // src/timing_controller.v(64[5] 132[12])
    defparam i7890_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_701_i6_3_lut (.I0(n10572), .I1(state[1]), .I2(n1503), 
            .I3(GND_net), .O(n1504[5]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_701_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_693_i10_3_lut (.I0(n10568), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[9]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 sub_32_add_2_28_lut (.I0(GND_net), .I1(state_timeout_counter[26]), 
            .I2(VCC_net), .I3(n8705), .O(n507[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_693_i11_3_lut (.I0(n10567), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[10]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i11_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFESR state_timeout_counter_i0_i28 (.Q(state_timeout_counter[28]), 
            .C(DEBUG_6_c), .E(n3668), .D(n507[28]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_CARRY sub_32_add_2_28 (.CI(n8705), .I0(state_timeout_counter[26]), 
            .I1(VCC_net), .CO(n8706));
    SB_CARRY sub_32_add_2_10 (.CI(n8687), .I0(state_timeout_counter[8]), 
            .I1(VCC_net), .CO(n8688));
    SB_LUT4 sub_32_add_2_27_lut (.I0(GND_net), .I1(state_timeout_counter[25]), 
            .I2(VCC_net), .I3(n8704), .O(n507[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_32_add_2_27 (.CI(n8704), .I0(state_timeout_counter[25]), 
            .I1(VCC_net), .CO(n8705));
    SB_LUT4 sub_32_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n8686), .O(n507[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_32_add_2_9 (.CI(n8686), .I0(state_timeout_counter[7]), 
            .I1(VCC_net), .CO(n8687));
    SB_LUT4 sub_32_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n8685), .O(n507[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_32_add_2_7_lut (.I0(n9338), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n8684), .O(n10572)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_32_add_2_26_lut (.I0(n1326), .I1(state_timeout_counter[24]), 
            .I2(VCC_net), .I3(n8703), .O(n10558)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_32_add_2_5 (.CI(n8682), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n8683));
    SB_LUT4 sub_32_add_2_17_lut (.I0(n1326), .I1(state_timeout_counter[15]), 
            .I2(VCC_net), .I3(n8694), .O(n10564)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_32_add_2_17 (.CI(n8694), .I0(state_timeout_counter[15]), 
            .I1(VCC_net), .CO(n8695));
    SB_CARRY sub_32_add_2_26 (.CI(n8703), .I0(state_timeout_counter[24]), 
            .I1(VCC_net), .CO(n8704));
    SB_CARRY sub_32_add_2_8 (.CI(n8685), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n8686));
    SB_DFFESR state_timeout_counter_i0_i29 (.Q(state_timeout_counter[29]), 
            .C(DEBUG_6_c), .E(n3668), .D(n507[29]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFESR state_timeout_counter_i0_i30 (.Q(state_timeout_counter[30]), 
            .C(DEBUG_6_c), .E(n3668), .D(n507[30]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_LUT4 sub_32_add_2_25_lut (.I0(n1326), .I1(state_timeout_counter[23]), 
            .I2(VCC_net), .I3(n8702), .O(n10559)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_32_add_2_25 (.CI(n8702), .I0(state_timeout_counter[23]), 
            .I1(VCC_net), .CO(n8703));
    SB_LUT4 sub_32_add_2_24_lut (.I0(n1326), .I1(state_timeout_counter[22]), 
            .I2(VCC_net), .I3(n8701), .O(n10560)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_32_add_2_4_lut (.I0(n6392), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n8681), .O(n10570)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_32_add_2_16_lut (.I0(n1326), .I1(state_timeout_counter[14]), 
            .I2(VCC_net), .I3(n8693), .O(n10565)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_32_add_2_24 (.CI(n8701), .I0(state_timeout_counter[22]), 
            .I1(VCC_net), .CO(n8702));
    SB_CARRY sub_32_add_2_3 (.CI(n8680), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n8681));
    SB_DFFESR state_timeout_counter_i0_i31 (.Q(state_timeout_counter[31]), 
            .C(DEBUG_6_c), .E(n3668), .D(n507[31]), .R(n3984));   // src/timing_controller.v(59[8] 133[4])
    SB_LUT4 sub_32_add_2_2_lut (.I0(n6392), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n10530)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_32_add_2_16 (.CI(n8693), .I0(state_timeout_counter[14]), 
            .I1(VCC_net), .CO(n8694));
    SB_LUT4 sub_32_add_2_15_lut (.I0(GND_net), .I1(state_timeout_counter[13]), 
            .I2(VCC_net), .I3(n8692), .O(n507[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_32_add_2_6_lut (.I0(n1326), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n8683), .O(n10582)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_32_add_2_15 (.CI(n8692), .I0(state_timeout_counter[13]), 
            .I1(VCC_net), .CO(n8693));
    SB_CARRY sub_32_add_2_4 (.CI(n8681), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n8682));
    SB_CARRY sub_32_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n8680));
    SB_LUT4 sub_32_add_2_14_lut (.I0(n1326), .I1(state_timeout_counter[12]), 
            .I2(VCC_net), .I3(n8691), .O(n10566)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_32_add_2_14 (.CI(n8691), .I0(state_timeout_counter[12]), 
            .I1(VCC_net), .CO(n8692));
    SB_LUT4 mux_693_i13_3_lut (.I0(n10566), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[12]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i13_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 sub_32_add_2_23_lut (.I0(GND_net), .I1(state_timeout_counter[21]), 
            .I2(VCC_net), .I3(n8700), .O(n507[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_32_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_693_i15_3_lut (.I0(n10565), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[14]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i15_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_2_lut (.I0(n1326), .I1(n1431), .I2(GND_net), .I3(GND_net), 
            .O(n9338));   // src/timing_controller.v(64[5] 132[12])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_693_i3_3_lut (.I0(n10570), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[2]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY sub_32_add_2_23 (.CI(n8700), .I0(state_timeout_counter[21]), 
            .I1(VCC_net), .CO(n8701));
    SB_LUT4 mux_693_i2_3_lut (.I0(n10571), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[1]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_693_i16_3_lut (.I0(n10564), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[15]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_693_i19_3_lut (.I0(n10563), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[18]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i19_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_693_i20_3_lut (.I0(n10562), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[19]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_693_i21_3_lut (.I0(n10561), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[20]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i21_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_693_i23_3_lut (.I0(n10560), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[22]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i23_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_693_i24_3_lut (.I0(n10559), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[23]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_693_i25_3_lut (.I0(n10558), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[24]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i25_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i9149_2_lut (.I0(state[3]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n5));   // src/timing_controller.v(59[8] 133[4])
    defparam i9149_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i762_4_lut (.I0(state[3]), .I1(n1585), .I2(n6602), .I3(state[2]), 
            .O(n1503));   // src/timing_controller.v(59[8] 133[4])
    defparam i762_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i5489_3_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n6572));
    defparam i5489_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut (.I0(state[2]), .I1(state[1]), .I2(state[0]), .I3(GND_net), 
            .O(n3474));   // src/timing_controller.v(64[5] 132[12])
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9153_2_lut (.I0(state[3]), .I1(n3474), .I2(GND_net), .I3(GND_net), 
            .O(n3668));   // src/timing_controller.v(64[5] 132[12])
    defparam i9153_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 mux_693_i1_3_lut (.I0(n10530), .I1(state[1]), .I2(n1431), 
            .I3(GND_net), .O(n1432[0]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_693_i1_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_701_i1_4_lut (.I0(n1432[0]), .I1(state[1]), .I2(n1503), 
            .I3(n9350), .O(n1504[0]));   // src/timing_controller.v(64[5] 132[12])
    defparam mux_701_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 state_3__I_0_56_Mux_1_i15_4_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[3]), .I3(n9361), .O(state_3__N_313[1]));   // src/timing_controller.v(64[5] 132[12])
    defparam state_3__I_0_56_Mux_1_i15_4_lut_4_lut.LUT_INIT = 16'hc6f6;
    SB_DFFE state_i2 (.Q(state[2]), .C(DEBUG_6_c), .E(n3830), .D(state_3__N_313[2]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(DEBUG_6_c), .E(n3830), .D(state_3__N_313[1]));   // src/timing_controller.v(59[8] 133[4])
    SB_DFF invert_52_i3 (.Q(INVERT_c_3), .C(DEBUG_6_c), .D(n596[3]));   // src/timing_controller.v(64[5] 132[12])
    SB_LUT4 i1_2_lut_adj_60 (.I0(state[3]), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n9355));
    defparam i1_2_lut_adj_60.LUT_INIT = 16'hbbbb;
    SB_LUT4 i751_2_lut_3_lut (.I0(state[0]), .I1(n63), .I2(state[1]), 
            .I3(GND_net), .O(n1585));   // src/timing_controller.v(59[8] 133[4])
    defparam i751_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i6_2_lut (.I0(state_timeout_counter[19]), .I1(state_timeout_counter[21]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // src/timing_controller.v(59[8] 133[4])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut (.I0(state_timeout_counter[22]), .I1(state_timeout_counter[26]), 
            .I2(state_timeout_counter[25]), .I3(state_timeout_counter[28]), 
            .O(n52));   // src/timing_controller.v(59[8] 133[4])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(state_timeout_counter[4]), .I1(state_timeout_counter[16]), 
            .I2(state_timeout_counter[8]), .I3(state_timeout_counter[0]), 
            .O(n56));   // src/timing_controller.v(59[8] 133[4])
    defparam i24_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i22_4_lut (.I0(state_timeout_counter[10]), .I1(state_timeout_counter[17]), 
            .I2(state_timeout_counter[12]), .I3(state_timeout_counter[18]), 
            .O(n54));   // src/timing_controller.v(59[8] 133[4])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(state_timeout_counter[20]), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[24]), .I3(state_timeout_counter[2]), 
            .O(n55));   // src/timing_controller.v(59[8] 133[4])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[6]), 
            .I2(state_timeout_counter[5]), .I3(state_timeout_counter[9]), 
            .O(n53));   // src/timing_controller.v(59[8] 133[4])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(state_timeout_counter[29]), .I1(state_timeout_counter[7]), 
            .I2(state_timeout_counter[30]), .I3(state_timeout_counter[11]), 
            .O(n50));   // src/timing_controller.v(59[8] 133[4])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(state_timeout_counter[13]), .I1(n52), .I2(n38), 
            .I3(state_timeout_counter[14]), .O(n58));   // src/timing_controller.v(59[8] 133[4])
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30_4_lut (.I0(n53), .I1(n55), .I2(n54), .I3(n56), .O(n62));   // src/timing_controller.v(59[8] 133[4])
    defparam i30_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(state_timeout_counter[31]), .I1(state_timeout_counter[23]), 
            .I2(state_timeout_counter[15]), .I3(state_timeout_counter[27]), 
            .O(n49));   // src/timing_controller.v(59[8] 133[4])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31_4_lut (.I0(n49), .I1(n62), .I2(n58), .I3(n50), .O(n63));   // src/timing_controller.v(59[8] 133[4])
    defparam i31_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5523_3_lut (.I0(n63), .I1(state[1]), .I2(state[2]), .I3(GND_net), 
            .O(n6606));
    defparam i5523_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 state_3__I_0_56_Mux_0_i7_4_lut (.I0(state[1]), .I1(n63), .I2(state[2]), 
            .I3(state[0]), .O(n7));   // src/timing_controller.v(64[5] 132[12])
    defparam state_3__I_0_56_Mux_0_i7_4_lut.LUT_INIT = 16'hc535;
    SB_LUT4 state_3__I_0_56_Mux_0_i15_4_lut (.I0(n7), .I1(n6606), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_313[0]));   // src/timing_controller.v(64[5] 132[12])
    defparam state_3__I_0_56_Mux_0_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_DFF invert_52_i0 (.Q(reset_all), .C(DEBUG_6_c), .D(n9329));   // src/timing_controller.v(64[5] 132[12])
    SB_LUT4 mux_701_i4_3_lut_4_lut (.I0(state[1]), .I1(n9350), .I2(n1503), 
            .I3(n1432[3]), .O(n1504[3]));   // src/timing_controller.v(59[8] 133[4])
    defparam mux_701_i4_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_701_i10_3_lut_4_lut (.I0(state[1]), .I1(n9350), .I2(n1503), 
            .I3(n1432[9]), .O(n1504[9]));   // src/timing_controller.v(59[8] 133[4])
    defparam mux_701_i10_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_701_i11_3_lut_4_lut (.I0(state[1]), .I1(n9350), .I2(n1503), 
            .I3(n1432[10]), .O(n1504[10]));   // src/timing_controller.v(59[8] 133[4])
    defparam mux_701_i11_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_701_i13_3_lut_4_lut (.I0(state[1]), .I1(n9350), .I2(n1503), 
            .I3(n1432[12]), .O(n1504[12]));   // src/timing_controller.v(59[8] 133[4])
    defparam mux_701_i13_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_701_i15_3_lut_4_lut (.I0(state[1]), .I1(n9350), .I2(n1503), 
            .I3(n1432[14]), .O(n1504[14]));   // src/timing_controller.v(59[8] 133[4])
    defparam mux_701_i15_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_701_i16_3_lut_4_lut (.I0(state[1]), .I1(n9350), .I2(n1503), 
            .I3(n1432[15]), .O(n1504[15]));   // src/timing_controller.v(59[8] 133[4])
    defparam mux_701_i16_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_DFFESR invert_52_i2 (.Q(UPDATE_c_2), .C(DEBUG_6_c), .E(VCC_net), 
            .D(n10656), .R(n5));   // src/timing_controller.v(64[5] 132[12])
    SB_LUT4 mux_701_i19_3_lut_4_lut (.I0(state[1]), .I1(n9350), .I2(n1503), 
            .I3(n1432[18]), .O(n1504[18]));   // src/timing_controller.v(59[8] 133[4])
    defparam mux_701_i19_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_701_i20_3_lut_4_lut (.I0(state[1]), .I1(n9350), .I2(n1503), 
            .I3(n1432[19]), .O(n1504[19]));   // src/timing_controller.v(59[8] 133[4])
    defparam mux_701_i20_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_701_i21_3_lut_4_lut (.I0(state[1]), .I1(n9350), .I2(n1503), 
            .I3(n1432[20]), .O(n1504[20]));   // src/timing_controller.v(59[8] 133[4])
    defparam mux_701_i21_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_701_i24_3_lut_4_lut (.I0(state[1]), .I1(n9350), .I2(n1503), 
            .I3(n1432[23]), .O(n1504[23]));   // src/timing_controller.v(59[8] 133[4])
    defparam mux_701_i24_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_701_i25_3_lut_4_lut (.I0(state[1]), .I1(n9350), .I2(n1503), 
            .I3(n1432[24]), .O(n1504[24]));   // src/timing_controller.v(59[8] 133[4])
    defparam mux_701_i25_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_701_i23_3_lut_4_lut (.I0(state[1]), .I1(n9350), .I2(n1503), 
            .I3(n1432[22]), .O(n1504[22]));   // src/timing_controller.v(59[8] 133[4])
    defparam mux_701_i23_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 state_3__I_0_56_Mux_2_i15_4_lut (.I0(state[1]), .I1(state[2]), 
            .I2(state[3]), .I3(state[0]), .O(state_3__N_313[2]));   // src/timing_controller.v(64[5] 132[12])
    defparam state_3__I_0_56_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[3]), .I1(n63), .I2(state[1]), .I3(state[2]), 
            .O(n9356));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_61 (.I0(state[0]), .I1(n63), .I2(state[3]), 
            .I3(state[2]), .O(n9350));   // src/timing_controller.v(59[8] 133[4])
    defparam i1_2_lut_3_lut_4_lut_adj_61.LUT_INIT = 16'h0200;
    SB_LUT4 i2909_2_lut_3_lut (.I0(state[3]), .I1(n3474), .I2(n1503), 
            .I3(GND_net), .O(n3998));   // src/timing_controller.v(59[8] 133[4])
    defparam i2909_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i9139_3_lut_4_lut (.I0(state[3]), .I1(n3474), .I2(n1503), 
            .I3(n9338), .O(n3984));
    defparam i9139_3_lut_4_lut.LUT_INIT = 16'h7077;
    SB_LUT4 i9114_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n10656));   // src/timing_controller.v(64[5] 132[12])
    defparam i9114_2_lut.LUT_INIT = 16'h9999;
    
endmodule
//
// Verilog Description of module bluejay_data
//

module bluejay_data (DEBUG_6_c, GND_net, DEBUG_9_c, DEBUG_3_c, buffer_switch_done, 
            DEBUG_2_c, DEBUG_5_c, VCC_net, DATA15_c, DATA14_c, DATA13_c, 
            DATA12_c, DATA11_c, DATA10_c, DATA9_c, DATA8_c, DATA7_c, 
            DATA6_c, DATA5_c, DATA20_c, DATA19_c, DATA18_c, \fifo_data_out[1] , 
            \fifo_data_out[2] , \fifo_data_out[0] , \fifo_data_out[5] , 
            \fifo_data_out[6] , \fifo_data_out[7] , \fifo_data_out[8] , 
            \fifo_data_out[9] , \fifo_data_out[10] , \fifo_data_out[11] , 
            \fifo_data_out[12] , \fifo_data_out[13] , \fifo_data_out[14] , 
            \fifo_data_out[15] , \fifo_data_out[3] , \fifo_data_out[4] , 
            DATA17_c) /* synthesis syn_module_defined=1 */ ;
    input DEBUG_6_c;
    input GND_net;
    output DEBUG_9_c;
    output DEBUG_3_c;
    input buffer_switch_done;
    input DEBUG_2_c;
    output DEBUG_5_c;
    input VCC_net;
    output DATA15_c;
    output DATA14_c;
    output DATA13_c;
    output DATA12_c;
    output DATA11_c;
    output DATA10_c;
    output DATA9_c;
    output DATA8_c;
    output DATA7_c;
    output DATA6_c;
    output DATA5_c;
    output DATA20_c;
    output DATA19_c;
    output DATA18_c;
    input \fifo_data_out[1] ;
    input \fifo_data_out[2] ;
    input \fifo_data_out[0] ;
    input \fifo_data_out[5] ;
    input \fifo_data_out[6] ;
    input \fifo_data_out[7] ;
    input \fifo_data_out[8] ;
    input \fifo_data_out[9] ;
    input \fifo_data_out[10] ;
    input \fifo_data_out[11] ;
    input \fifo_data_out[12] ;
    input \fifo_data_out[13] ;
    input \fifo_data_out[14] ;
    input \fifo_data_out[15] ;
    input \fifo_data_out[3] ;
    input \fifo_data_out[4] ;
    output DATA17_c;
    
    wire DEBUG_6_c /* synthesis SET_AS_NETWORK=DEBUG_6_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [8:0]n47;
    
    wire n3625;
    wire [7:0]state_timeout_counter;   // src/bluejay_data.v(52[11:32])
    
    wire n6151, data_o_31__N_619, n73, data_o_31__N_620;
    wire [7:0]n1791;
    
    wire n2401, n3927;
    wire [7:0]n1771;
    
    wire n4056, get_next_word_N_623;
    wire [10:0]v_counter_10__N_600;
    
    wire n3809;
    wire [10:0]v_counter;   // src/bluejay_data.v(50[12:21])
    wire [7:0]n520;
    
    wire n9362, n10, n9288, n9388, n8903, n9303, n544, n6, n10_adj_1095, 
        n4, n6185, n2389, n9, n9474, n9484, n553, n5346, n2367, 
        n2377, data_o_31__N_621, n2397, n8750, n8751, n8749, n8712, 
        n8713, n8711, n6154, n8748, n8747, n2422, n5059, n5058, 
        n8746, n8745, n8744, n5009, n8743, n4991, n4951, n4950, 
        n4949, n4948, n4947, n4931, n4930, n4881, n4816, n4815, 
        n8717, n8716, n8715, n82, n8714, n74, n8752, n6148, 
        n4267, n9448, n7;
    
    SB_DFFESR state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(DEBUG_6_c), 
            .E(n3625), .D(n47[7]), .R(n6151));   // src/bluejay_data.v(56[8] 114[4])
    SB_LUT4 i1_3_lut (.I0(data_o_31__N_619), .I1(n73), .I2(data_o_31__N_620), 
            .I3(GND_net), .O(n1791[5]));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_DFFESS state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(DEBUG_6_c), 
            .E(n3625), .D(n2401), .S(n3927));   // src/bluejay_data.v(56[8] 114[4])
    SB_DFFESR state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(DEBUG_6_c), 
            .E(n3625), .D(n1771[2]), .R(n4056));   // src/bluejay_data.v(56[8] 114[4])
    SB_DFFN get_next_word_54 (.Q(DEBUG_9_c), .C(DEBUG_6_c), .D(get_next_word_N_623));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFN sync_55 (.Q(DEBUG_3_c), .C(DEBUG_6_c), .D(data_o_31__N_619));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFESR v_counter_i1 (.Q(v_counter[1]), .C(DEBUG_6_c), .E(n3809), 
            .D(v_counter_10__N_600[1]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 114[4])
    SB_DFFESR v_counter_i2 (.Q(v_counter[2]), .C(DEBUG_6_c), .E(n3809), 
            .D(v_counter_10__N_600[2]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 114[4])
    SB_DFFESR v_counter_i3 (.Q(v_counter[3]), .C(DEBUG_6_c), .E(n3809), 
            .D(v_counter_10__N_600[3]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 114[4])
    SB_DFF state_FSM_i0 (.Q(n520[0]), .C(DEBUG_6_c), .D(buffer_switch_done));   // src/bluejay_data.v(62[9] 112[16])
    SB_DFFESR v_counter_i4 (.Q(v_counter[4]), .C(DEBUG_6_c), .E(n3809), 
            .D(v_counter_10__N_600[4]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 114[4])
    SB_DFFESR v_counter_i5 (.Q(v_counter[5]), .C(DEBUG_6_c), .E(n3809), 
            .D(v_counter_10__N_600[5]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 114[4])
    SB_DFFESR v_counter_i6 (.Q(v_counter[6]), .C(DEBUG_6_c), .E(n3809), 
            .D(v_counter_10__N_600[6]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 114[4])
    SB_DFFESR v_counter_i7 (.Q(v_counter[7]), .C(DEBUG_6_c), .E(n3809), 
            .D(v_counter_10__N_600[7]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 114[4])
    SB_DFFESS v_counter_i8 (.Q(v_counter[8]), .C(DEBUG_6_c), .E(n3809), 
            .D(v_counter_10__N_600[8]), .S(buffer_switch_done));   // src/bluejay_data.v(56[8] 114[4])
    SB_DFFESR v_counter_i9 (.Q(v_counter[9]), .C(DEBUG_6_c), .E(n3809), 
            .D(v_counter_10__N_600[9]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 114[4])
    SB_DFFESS v_counter_i10 (.Q(v_counter[10]), .C(DEBUG_6_c), .E(n3809), 
            .D(v_counter_10__N_600[10]), .S(buffer_switch_done));   // src/bluejay_data.v(56[8] 114[4])
    SB_LUT4 i7848_4_lut (.I0(n9362), .I1(n10), .I2(n9288), .I3(state_timeout_counter[4]), 
            .O(n9388));
    defparam i7848_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut (.I0(v_counter[0]), .I1(n520[7]), .I2(state_timeout_counter[0]), 
            .I3(n9388), .O(n8903));
    defparam i3_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i1_4_lut (.I0(n520[1]), .I1(n8903), .I2(n520[0]), .I3(DEBUG_2_c), 
            .O(n9303));
    defparam i1_4_lut.LUT_INIT = 16'heefe;
    SB_LUT4 i166_2_lut (.I0(DEBUG_2_c), .I1(n520[0]), .I2(GND_net), .I3(GND_net), 
            .O(n544));   // src/bluejay_data.v(62[9] 112[16])
    defparam i166_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut (.I0(v_counter[8]), .I1(v_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // src/bluejay_data.v(56[8] 114[4])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(v_counter[0]), .I1(v_counter[3]), .I2(v_counter[6]), 
            .I3(n6), .O(n9288));   // src/bluejay_data.v(56[8] 114[4])
    defparam i4_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_4_lut_adj_47 (.I0(v_counter[10]), .I1(v_counter[9]), .I2(v_counter[7]), 
            .I3(v_counter[1]), .O(n10_adj_1095));
    defparam i4_4_lut_adj_47.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(v_counter[2]), .I1(n10_adj_1095), .I2(v_counter[5]), 
            .I3(GND_net), .O(n10));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_adj_48 (.I0(n10), .I1(n520[7]), .I2(n9288), .I3(GND_net), 
            .O(n4));   // src/bluejay_data.v(62[9] 112[16])
    defparam i1_3_lut_adj_48.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1316_4_lut (.I0(n520[4]), .I1(n6185), .I2(DEBUG_2_c), .I3(n4), 
            .O(n2389));   // src/bluejay_data.v(62[9] 112[16])
    defparam i1316_4_lut.LUT_INIT = 16'h3b0a;
    SB_LUT4 i7942_4_lut (.I0(n9), .I1(n9474), .I2(state_timeout_counter[3]), 
            .I3(state_timeout_counter[2]), .O(n9484));
    defparam i7942_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 reduce_or_174_i1_4_lut (.I0(DEBUG_2_c), .I1(n520[3]), .I2(n520[4]), 
            .I3(n9484), .O(n553));   // src/bluejay_data.v(62[9] 112[16])
    defparam reduce_or_174_i1_4_lut.LUT_INIT = 16'ha0ec;
    SB_DFFN data_o_i1 (.Q(DEBUG_5_c), .C(DEBUG_6_c), .D(n5346));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFSR state_FSM_i7 (.Q(n520[7]), .C(DEBUG_6_c), .D(n2367), .R(buffer_switch_done));   // src/bluejay_data.v(62[9] 112[16])
    SB_DFFSR state_FSM_i6 (.Q(data_o_31__N_621), .C(DEBUG_6_c), .D(n2377), 
            .R(buffer_switch_done));   // src/bluejay_data.v(62[9] 112[16])
    SB_DFFSR state_FSM_i5 (.Q(data_o_31__N_620), .C(DEBUG_6_c), .D(n553), 
            .R(buffer_switch_done));   // src/bluejay_data.v(62[9] 112[16])
    SB_DFFSR state_FSM_i4 (.Q(n520[4]), .C(DEBUG_6_c), .D(n2389), .R(buffer_switch_done));   // src/bluejay_data.v(62[9] 112[16])
    SB_DFFSR state_FSM_i3 (.Q(n520[3]), .C(DEBUG_6_c), .D(n2397), .R(buffer_switch_done));   // src/bluejay_data.v(62[9] 112[16])
    SB_DFFSR state_FSM_i2 (.Q(data_o_31__N_619), .C(DEBUG_6_c), .D(n544), 
            .R(buffer_switch_done));   // src/bluejay_data.v(62[9] 112[16])
    SB_DFFSR state_FSM_i1 (.Q(n520[1]), .C(DEBUG_6_c), .D(n9303), .R(buffer_switch_done));   // src/bluejay_data.v(62[9] 112[16])
    SB_CARRY sub_110_add_2_10 (.CI(n8750), .I0(v_counter[8]), .I1(VCC_net), 
            .CO(n8751));
    SB_LUT4 sub_110_add_2_9_lut (.I0(GND_net), .I1(v_counter[7]), .I2(VCC_net), 
            .I3(n8749), .O(v_counter_10__N_600[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_110_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_110_add_2_9 (.CI(n8749), .I0(v_counter[7]), .I1(VCC_net), 
            .CO(n8750));
    SB_CARRY sub_108_add_2_4 (.CI(n8712), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n8713));
    SB_LUT4 sub_108_add_2_3_lut (.I0(n6154), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n8711), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_108_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_110_add_2_8_lut (.I0(GND_net), .I1(v_counter[6]), .I2(VCC_net), 
            .I3(n8748), .O(v_counter_10__N_600[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_110_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_110_add_2_8 (.CI(n8748), .I0(v_counter[6]), .I1(VCC_net), 
            .CO(n8749));
    SB_CARRY sub_108_add_2_3 (.CI(n8711), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n8712));
    SB_LUT4 sub_110_add_2_7_lut (.I0(GND_net), .I1(v_counter[5]), .I2(VCC_net), 
            .I3(n8747), .O(v_counter_10__N_600[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_110_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_108_add_2_2_lut (.I0(n6154), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n2422)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_108_add_2_2_lut.LUT_INIT = 16'h8228;
    SB_DFFN data_o_i16 (.Q(DATA15_c), .C(DEBUG_6_c), .D(n5059));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFN data_o_i15 (.Q(DATA14_c), .C(DEBUG_6_c), .D(n5058));   // src/bluejay_data.v(117[8] 137[4])
    SB_CARRY sub_110_add_2_7 (.CI(n8747), .I0(v_counter[5]), .I1(VCC_net), 
            .CO(n8748));
    SB_LUT4 sub_110_add_2_6_lut (.I0(GND_net), .I1(v_counter[4]), .I2(VCC_net), 
            .I3(n8746), .O(v_counter_10__N_600[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_110_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_110_add_2_6 (.CI(n8746), .I0(v_counter[4]), .I1(VCC_net), 
            .CO(n8747));
    SB_LUT4 sub_110_add_2_5_lut (.I0(GND_net), .I1(v_counter[3]), .I2(VCC_net), 
            .I3(n8745), .O(v_counter_10__N_600[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_110_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_110_add_2_5 (.CI(n8745), .I0(v_counter[3]), .I1(VCC_net), 
            .CO(n8746));
    SB_LUT4 sub_110_add_2_4_lut (.I0(GND_net), .I1(v_counter[2]), .I2(VCC_net), 
            .I3(n8744), .O(v_counter_10__N_600[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_110_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_108_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n8711));
    SB_DFFN data_o_i14 (.Q(DATA13_c), .C(DEBUG_6_c), .D(n5009));   // src/bluejay_data.v(117[8] 137[4])
    SB_CARRY sub_110_add_2_4 (.CI(n8744), .I0(v_counter[2]), .I1(VCC_net), 
            .CO(n8745));
    SB_LUT4 sub_110_add_2_3_lut (.I0(GND_net), .I1(v_counter[1]), .I2(VCC_net), 
            .I3(n8743), .O(v_counter_10__N_600[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_110_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_110_add_2_3 (.CI(n8743), .I0(v_counter[1]), .I1(VCC_net), 
            .CO(n8744));
    SB_LUT4 sub_110_add_2_2_lut (.I0(GND_net), .I1(v_counter[0]), .I2(n6185), 
            .I3(VCC_net), .O(v_counter_10__N_600[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_110_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_110_add_2_2 (.CI(VCC_net), .I0(v_counter[0]), .I1(n6185), 
            .CO(n8743));
    SB_DFFN data_o_i13 (.Q(DATA12_c), .C(DEBUG_6_c), .D(n4991));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFN data_o_i12 (.Q(DATA11_c), .C(DEBUG_6_c), .D(n4951));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFN data_o_i11 (.Q(DATA10_c), .C(DEBUG_6_c), .D(n4950));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFN data_o_i10 (.Q(DATA9_c), .C(DEBUG_6_c), .D(n4949));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFN data_o_i9 (.Q(DATA8_c), .C(DEBUG_6_c), .D(n4948));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFN data_o_i8 (.Q(DATA7_c), .C(DEBUG_6_c), .D(n4947));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFN data_o_i7 (.Q(DATA6_c), .C(DEBUG_6_c), .D(n4931));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFN data_o_i6 (.Q(DATA5_c), .C(DEBUG_6_c), .D(n4930));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFN data_o_i5 (.Q(DATA20_c), .C(DEBUG_6_c), .D(n4881));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFN data_o_i4 (.Q(DATA19_c), .C(DEBUG_6_c), .D(n4816));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFN data_o_i3 (.Q(DATA18_c), .C(DEBUG_6_c), .D(n4815));   // src/bluejay_data.v(117[8] 137[4])
    SB_DFFE state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(DEBUG_6_c), 
            .E(n3625), .D(n1791[5]));   // src/bluejay_data.v(56[8] 114[4])
    SB_LUT4 sub_108_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n8717), .O(n47[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_108_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_108_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n8716), .O(n47[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_108_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_108_add_2_8 (.CI(n8716), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n8717));
    SB_LUT4 sub_108_add_2_7_lut (.I0(n82), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n8715), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_108_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_108_add_2_7 (.CI(n8715), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n8716));
    SB_LUT4 sub_108_add_2_6_lut (.I0(GND_net), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n8714), .O(n47[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_108_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_108_add_2_6 (.CI(n8714), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n8715));
    SB_LUT4 sub_108_add_2_5_lut (.I0(n82), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n8713), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_108_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_110_add_2_12_lut (.I0(GND_net), .I1(v_counter[10]), .I2(VCC_net), 
            .I3(n8752), .O(v_counter_10__N_600[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_110_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_110_add_2_11_lut (.I0(GND_net), .I1(v_counter[9]), .I2(VCC_net), 
            .I3(n8751), .O(v_counter_10__N_600[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_110_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_108_add_2_5 (.CI(n8713), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n8714));
    SB_LUT4 sub_108_add_2_4_lut (.I0(n6148), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n8712), .O(n1771[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_108_add_2_4_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_110_add_2_11 (.CI(n8751), .I0(v_counter[9]), .I1(VCC_net), 
            .CO(n8752));
    SB_LUT4 sub_110_add_2_10_lut (.I0(GND_net), .I1(v_counter[8]), .I2(VCC_net), 
            .I3(n8750), .O(v_counter_10__N_600[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_110_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut (.I0(data_o_31__N_620), .I1(n6148), .I2(data_o_31__N_619), 
            .I3(n3625), .O(n6151));   // src/bluejay_data.v(62[9] 112[16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_DFFESR state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(DEBUG_6_c), 
            .E(n3625), .D(n47[4]), .R(n6151));   // src/bluejay_data.v(56[8] 114[4])
    SB_DFFESR state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(DEBUG_6_c), 
            .E(n3625), .D(n47[6]), .R(n6151));   // src/bluejay_data.v(56[8] 114[4])
    SB_LUT4 i3178_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[1] ), .I3(GND_net), .O(n4267));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3178_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3726_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[2] ), .I3(GND_net), .O(n4815));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3726_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i4257_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[0] ), .I3(GND_net), .O(n5346));   // src/bluejay_data.v(62[9] 112[16])
    defparam i4257_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3841_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[5] ), .I3(GND_net), .O(n4930));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3841_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3842_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[6] ), .I3(GND_net), .O(n4931));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3842_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3858_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[7] ), .I3(GND_net), .O(n4947));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3858_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3859_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[8] ), .I3(GND_net), .O(n4948));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3859_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3860_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[9] ), .I3(GND_net), .O(n4949));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3860_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3861_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[10] ), .I3(GND_net), .O(n4950));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3861_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3862_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[11] ), .I3(GND_net), .O(n4951));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3862_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3902_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[12] ), .I3(GND_net), .O(n4991));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3902_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3920_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[13] ), .I3(GND_net), .O(n5009));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3920_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3969_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[14] ), .I3(GND_net), .O(n5058));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3969_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_DFFE state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(DEBUG_6_c), 
            .E(n3625), .D(n1791[3]));   // src/bluejay_data.v(56[8] 114[4])
    SB_LUT4 i3970_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[15] ), .I3(GND_net), .O(n5059));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3970_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(data_o_31__N_619), .I3(GND_net), .O(get_next_word_N_623));   // src/bluejay_data.v(62[9] 112[16])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i3727_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[3] ), .I3(GND_net), .O(n4816));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3727_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3792_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(\fifo_data_out[4] ), .I3(GND_net), .O(n4881));   // src/bluejay_data.v(62[9] 112[16])
    defparam i3792_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_49 (.I0(n520[7]), .I1(buffer_switch_done), .I2(GND_net), 
            .I3(GND_net), .O(n3809));
    defparam i1_2_lut_adj_49.LUT_INIT = 16'heeee;
    SB_DFFN data_o_i2 (.Q(DATA17_c), .C(DEBUG_6_c), .D(n4267));   // src/bluejay_data.v(117[8] 137[4])
    SB_LUT4 i1_3_lut_adj_50 (.I0(n3625), .I1(data_o_31__N_619), .I2(data_o_31__N_620), 
            .I3(GND_net), .O(n4056));   // src/bluejay_data.v(61[10] 113[8])
    defparam i1_3_lut_adj_50.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_2_lut_adj_51 (.I0(n3625), .I1(data_o_31__N_619), .I2(GND_net), 
            .I3(GND_net), .O(n3927));   // src/bluejay_data.v(61[10] 113[8])
    defparam i1_2_lut_adj_51.LUT_INIT = 16'h8888;
    SB_LUT4 i7907_2_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[7]), 
            .I2(GND_net), .I3(GND_net), .O(n9448));
    defparam i7907_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_52 (.I0(state_timeout_counter[2]), .I1(state_timeout_counter[6]), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // src/bluejay_data.v(43[15:21])
    defparam i1_2_lut_adj_52.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(state_timeout_counter[5]), .I1(n7), .I2(state_timeout_counter[3]), 
            .I3(n9448), .O(n9362));   // src/bluejay_data.v(43[15:21])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_53 (.I0(state_timeout_counter[0]), .I1(state_timeout_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // src/bluejay_data.v(97[21:49])
    defparam i1_2_lut_adj_53.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_54 (.I0(data_o_31__N_621), .I1(n6185), .I2(GND_net), 
            .I3(GND_net), .O(n6148));   // src/bluejay_data.v(62[9] 112[16])
    defparam i1_2_lut_adj_54.LUT_INIT = 16'h2222;
    SB_DFFESR v_counter_i0 (.Q(v_counter[0]), .C(DEBUG_6_c), .E(n3809), 
            .D(v_counter_10__N_600[0]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 114[4])
    SB_LUT4 i9165_4_lut (.I0(n520[0]), .I1(buffer_switch_done), .I2(n520[4]), 
            .I3(n520[1]), .O(n3625));   // src/bluejay_data.v(61[10] 113[8])
    defparam i9165_4_lut.LUT_INIT = 16'h0001;
    SB_DFFESS state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(DEBUG_6_c), 
            .E(n3625), .D(n2422), .S(n3927));   // src/bluejay_data.v(56[8] 114[4])
    SB_LUT4 i1_3_lut_adj_55 (.I0(data_o_31__N_619), .I1(n74), .I2(data_o_31__N_620), 
            .I3(GND_net), .O(n1791[3]));
    defparam i1_3_lut_adj_55.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(data_o_31__N_621), .I1(state_timeout_counter[0]), 
            .I2(state_timeout_counter[4]), .I3(n9362), .O(n82));   // src/bluejay_data.v(43[15:21])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_adj_56 (.I0(state_timeout_counter[0]), .I1(state_timeout_counter[4]), 
            .I2(n9362), .I3(GND_net), .O(n6185));   // src/bluejay_data.v(43[15:21])
    defparam i1_2_lut_3_lut_adj_56.LUT_INIT = 16'hfdfd;
    SB_LUT4 i5067_1_lut_2_lut_3_lut (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(n6185), .I3(GND_net), .O(n6154));   // src/bluejay_data.v(62[9] 112[16])
    defparam i5067_1_lut_2_lut_3_lut.LUT_INIT = 16'h5151;
    SB_LUT4 i1_3_lut_3_lut (.I0(n520[7]), .I1(data_o_31__N_621), .I2(n6185), 
            .I3(GND_net), .O(n2367));
    defparam i1_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_4_lut_adj_57 (.I0(data_o_31__N_620), .I1(data_o_31__N_621), 
            .I2(n9), .I3(n9362), .O(n2377));   // src/bluejay_data.v(62[9] 112[16])
    defparam i1_3_lut_4_lut_adj_57.LUT_INIT = 16'heeea;
    SB_LUT4 i7933_3_lut_4_lut (.I0(state_timeout_counter[6]), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[7]), .I3(state_timeout_counter[5]), 
            .O(n9474));
    defparam i7933_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_58 (.I0(data_o_31__N_619), .I1(n9), .I2(n9362), 
            .I3(n520[3]), .O(n2397));   // src/bluejay_data.v(62[9] 112[16])
    defparam i1_3_lut_4_lut_adj_58.LUT_INIT = 16'hfeaa;
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word
//

module FIFO_Quad_Word (rd_fifo_en_w, \mem_LUT.data_raw_r[0] , DEBUG_6_c, 
            rd_addr_r, n8, reset_all_w, n8_adj_4, wr_addr_r, rx_buf_byte, 
            n4086, \fifo_temp_output[1] , n4089, \fifo_temp_output[2] , 
            n4096, \fifo_temp_output[3] , n5330, VCC_net, \fifo_temp_output[0] , 
            n8987, is_tx_fifo_full_flag, n4111, \fifo_temp_output[4] , 
            n4123, \fifo_temp_output[5] , n4129, \fifo_temp_output[6] , 
            n5317, n5314, n5311, n5308, n4143, \fifo_temp_output[7] , 
            \rd_addr_p1_w[1] , GND_net, \rd_addr_p1_w[2] , \wr_addr_p1_w[1] , 
            n1, \wr_addr_p1_w[2] , n8824, \mem_LUT.data_raw_r[7] , \mem_LUT.data_raw_r[6] , 
            \mem_LUT.data_raw_r[5] , \mem_LUT.data_raw_r[4] , \mem_LUT.data_raw_r[3] , 
            \mem_LUT.data_raw_r[2] , \mem_LUT.data_raw_r[1] , fifo_write_cmd, 
            full_nxt_r, fifo_read_cmd, is_fifo_empty_flag, n9299, n4093, 
            rd_fifo_en_prev_r) /* synthesis syn_module_defined=1 */ ;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[0] ;
    input DEBUG_6_c;
    output [2:0]rd_addr_r;
    input n8;
    input reset_all_w;
    input n8_adj_4;
    output [2:0]wr_addr_r;
    input [7:0]rx_buf_byte;
    input n4086;
    output \fifo_temp_output[1] ;
    input n4089;
    output \fifo_temp_output[2] ;
    input n4096;
    output \fifo_temp_output[3] ;
    input n5330;
    input VCC_net;
    output \fifo_temp_output[0] ;
    input n8987;
    output is_tx_fifo_full_flag;
    input n4111;
    output \fifo_temp_output[4] ;
    input n4123;
    output \fifo_temp_output[5] ;
    input n4129;
    output \fifo_temp_output[6] ;
    input n5317;
    input n5314;
    input n5311;
    input n5308;
    input n4143;
    output \fifo_temp_output[7] ;
    output \rd_addr_p1_w[1] ;
    input GND_net;
    output \rd_addr_p1_w[2] ;
    output \wr_addr_p1_w[1] ;
    output n1;
    output \wr_addr_p1_w[2] ;
    output n8824;
    output \mem_LUT.data_raw_r[7] ;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[3] ;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[1] ;
    input fifo_write_cmd;
    output full_nxt_r;
    input fifo_read_cmd;
    output is_fifo_empty_flag;
    input n9299;
    input n4093;
    output rd_fifo_en_prev_r;
    
    wire DEBUG_6_c /* synthesis SET_AS_NETWORK=DEBUG_6_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2 lscc_fifo_inst (.rd_fifo_en_w(rd_fifo_en_w), 
            .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r[0] ), .DEBUG_6_c(DEBUG_6_c), 
            .rd_addr_r({rd_addr_r}), .n8(n8), .reset_all_w(reset_all_w), 
            .n8_adj_3(n8_adj_4), .wr_addr_r({wr_addr_r}), .rx_buf_byte({rx_buf_byte}), 
            .n4086(n4086), .\fifo_temp_output[1] (\fifo_temp_output[1] ), 
            .n4089(n4089), .\fifo_temp_output[2] (\fifo_temp_output[2] ), 
            .n4096(n4096), .\fifo_temp_output[3] (\fifo_temp_output[3] ), 
            .n5330(n5330), .VCC_net(VCC_net), .\fifo_temp_output[0] (\fifo_temp_output[0] ), 
            .n8987(n8987), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .n4111(n4111), .\fifo_temp_output[4] (\fifo_temp_output[4] ), 
            .n4123(n4123), .\fifo_temp_output[5] (\fifo_temp_output[5] ), 
            .n4129(n4129), .\fifo_temp_output[6] (\fifo_temp_output[6] ), 
            .n5317(n5317), .n5314(n5314), .n5311(n5311), .n5308(n5308), 
            .n4143(n4143), .\fifo_temp_output[7] (\fifo_temp_output[7] ), 
            .\rd_addr_p1_w[1] (\rd_addr_p1_w[1] ), .GND_net(GND_net), .\rd_addr_p1_w[2] (\rd_addr_p1_w[2] ), 
            .\wr_addr_p1_w[1] (\wr_addr_p1_w[1] ), .n1(n1), .\wr_addr_p1_w[2] (\wr_addr_p1_w[2] ), 
            .n8824(n8824), .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r[7] ), 
            .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r[6] ), .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r[5] ), 
            .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r[4] ), .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r[3] ), 
            .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r[2] ), .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r[1] ), 
            .fifo_write_cmd(fifo_write_cmd), .full_nxt_r(full_nxt_r), .fifo_read_cmd(fifo_read_cmd), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .n9299(n9299), .n4093(n4093), 
            .rd_fifo_en_prev_r(rd_fifo_en_prev_r)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_quad_word_mod.v(20[37:380])
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2
//

module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2 (rd_fifo_en_w, 
            \mem_LUT.data_raw_r[0] , DEBUG_6_c, rd_addr_r, n8, reset_all_w, 
            n8_adj_3, wr_addr_r, rx_buf_byte, n4086, \fifo_temp_output[1] , 
            n4089, \fifo_temp_output[2] , n4096, \fifo_temp_output[3] , 
            n5330, VCC_net, \fifo_temp_output[0] , n8987, is_tx_fifo_full_flag, 
            n4111, \fifo_temp_output[4] , n4123, \fifo_temp_output[5] , 
            n4129, \fifo_temp_output[6] , n5317, n5314, n5311, n5308, 
            n4143, \fifo_temp_output[7] , \rd_addr_p1_w[1] , GND_net, 
            \rd_addr_p1_w[2] , \wr_addr_p1_w[1] , n1, \wr_addr_p1_w[2] , 
            n8824, \mem_LUT.data_raw_r[7] , \mem_LUT.data_raw_r[6] , \mem_LUT.data_raw_r[5] , 
            \mem_LUT.data_raw_r[4] , \mem_LUT.data_raw_r[3] , \mem_LUT.data_raw_r[2] , 
            \mem_LUT.data_raw_r[1] , fifo_write_cmd, full_nxt_r, fifo_read_cmd, 
            is_fifo_empty_flag, n9299, n4093, rd_fifo_en_prev_r) /* synthesis syn_module_defined=1 */ ;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[0] ;
    input DEBUG_6_c;
    output [2:0]rd_addr_r;
    input n8;
    input reset_all_w;
    input n8_adj_3;
    output [2:0]wr_addr_r;
    input [7:0]rx_buf_byte;
    input n4086;
    output \fifo_temp_output[1] ;
    input n4089;
    output \fifo_temp_output[2] ;
    input n4096;
    output \fifo_temp_output[3] ;
    input n5330;
    input VCC_net;
    output \fifo_temp_output[0] ;
    input n8987;
    output is_tx_fifo_full_flag;
    input n4111;
    output \fifo_temp_output[4] ;
    input n4123;
    output \fifo_temp_output[5] ;
    input n4129;
    output \fifo_temp_output[6] ;
    input n5317;
    input n5314;
    input n5311;
    input n5308;
    input n4143;
    output \fifo_temp_output[7] ;
    output \rd_addr_p1_w[1] ;
    input GND_net;
    output \rd_addr_p1_w[2] ;
    output \wr_addr_p1_w[1] ;
    output n1;
    output \wr_addr_p1_w[2] ;
    output n8824;
    output \mem_LUT.data_raw_r[7] ;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[3] ;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[1] ;
    input fifo_write_cmd;
    output full_nxt_r;
    input fifo_read_cmd;
    output is_fifo_empty_flag;
    input n9299;
    input n4093;
    output rd_fifo_en_prev_r;
    
    wire DEBUG_6_c /* synthesis SET_AS_NETWORK=DEBUG_6_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [31:0]\mem_LUT.data_raw_r_31__N_968 ;
    
    wire \mem_LUT.mem_2_7 , \mem_LUT.mem_3_7 , n12204, \mem_LUT.mem_1_7 , 
        \mem_LUT.mem_0_7 , \mem_LUT.mem_2_6 , \mem_LUT.mem_3_6 , n12150, 
        \mem_LUT.mem_1_6 , \mem_LUT.mem_0_6 , \mem_LUT.mem_2_5 , \mem_LUT.mem_3_5 , 
        n12126, \mem_LUT.mem_1_5 , \mem_LUT.mem_0_5 , n3, n5284, n5283, 
        \mem_LUT.mem_2_4 , \mem_LUT.mem_3_4 , n12114, \mem_LUT.mem_1_4 , 
        \mem_LUT.mem_0_4 , n5282, n5281, \mem_LUT.mem_2_3 , \mem_LUT.mem_3_3 , 
        n12096, \mem_LUT.mem_1_3 , \mem_LUT.mem_0_3 , n5280, \mem_LUT.mem_3_2 , 
        n5279, \mem_LUT.mem_3_1 , n5278, \mem_LUT.mem_3_0 , n5277, 
        n4, n5273, n5272, n5271, n5270, n5269, n5268, \mem_LUT.mem_2_2 , 
        n5267, \mem_LUT.mem_2_1 , n5266, \mem_LUT.mem_2_0 , n5262, 
        n5261, n5260, n5259, n5258, n5257, \mem_LUT.mem_1_2 , n5256, 
        \mem_LUT.mem_1_1 , n5246, \mem_LUT.mem_1_0 , n5245, n5244, 
        n5243, n5242, n5241, n5240, \mem_LUT.mem_0_2 , n5239, \mem_LUT.mem_0_1 , 
        n5238, \mem_LUT.mem_0_0 , n3_adj_1093, n11850, n11844, n11832;
    
    SB_DFFE \mem_LUT.data_raw_r__i1  (.Q(\mem_LUT.data_raw_r[0] ), .C(DEBUG_6_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_968 [0]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_7 ), 
            .I2(\mem_LUT.mem_3_7 ), .I3(rd_addr_r[1]), .O(n12204));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n12204_bdd_4_lut (.I0(n12204), .I1(\mem_LUT.mem_1_7 ), .I2(\mem_LUT.mem_0_7 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_968 [7]));
    defparam n12204_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(DEBUG_6_c), .D(n8), .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFSR wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(DEBUG_6_c), .D(n8_adj_3), 
            .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10409 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_6 ), 
            .I2(\mem_LUT.mem_3_6 ), .I3(rd_addr_r[1]), .O(n12150));
    defparam rd_addr_r_0__bdd_4_lut_10409.LUT_INIT = 16'he4aa;
    SB_LUT4 n12150_bdd_4_lut (.I0(n12150), .I1(\mem_LUT.mem_1_6 ), .I2(\mem_LUT.mem_0_6 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_968 [6]));
    defparam n12150_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10364 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_5 ), 
            .I2(\mem_LUT.mem_3_5 ), .I3(rd_addr_r[1]), .O(n12126));
    defparam rd_addr_r_0__bdd_4_lut_10364.LUT_INIT = 16'he4aa;
    SB_LUT4 n12126_bdd_4_lut (.I0(n12126), .I1(\mem_LUT.mem_1_5 ), .I2(\mem_LUT.mem_0_5 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_968 [5]));
    defparam n12126_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4195_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_3_7 ), .O(n5284));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4195_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4194_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_3_6 ), .O(n5283));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4194_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10344 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_4 ), 
            .I2(\mem_LUT.mem_3_4 ), .I3(rd_addr_r[1]), .O(n12114));
    defparam rd_addr_r_0__bdd_4_lut_10344.LUT_INIT = 16'he4aa;
    SB_LUT4 n12114_bdd_4_lut (.I0(n12114), .I1(\mem_LUT.mem_1_4 ), .I2(\mem_LUT.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_968 [4]));
    defparam n12114_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4193_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_3_5 ), .O(n5282));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4193_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4192_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_3_4 ), .O(n5281));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4192_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10334 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_3 ), 
            .I2(\mem_LUT.mem_3_3 ), .I3(rd_addr_r[1]), .O(n12096));
    defparam rd_addr_r_0__bdd_4_lut_10334.LUT_INIT = 16'he4aa;
    SB_LUT4 n12096_bdd_4_lut (.I0(n12096), .I1(\mem_LUT.mem_1_3 ), .I2(\mem_LUT.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_968 [3]));
    defparam n12096_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4191_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_3_3 ), .O(n5280));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4191_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4190_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_3_2 ), .O(n5279));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4190_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4189_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_3_1 ), .O(n5278));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4189_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4188_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_3_0 ), .O(n5277));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4188_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4184_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_2_7 ), .O(n5273));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4184_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF \mem_LUT.data_buff_r__i1  (.Q(\fifo_temp_output[1] ), .C(DEBUG_6_c), 
           .D(n4086));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i2  (.Q(\fifo_temp_output[2] ), .C(DEBUG_6_c), 
           .D(n4089));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i3  (.Q(\fifo_temp_output[3] ), .C(DEBUG_6_c), 
           .D(n4096));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 i4183_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_2_6 ), .O(n5272));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4183_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE \mem_LUT.data_buff_r__i0  (.Q(\fifo_temp_output[0] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5330));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE full_r_84 (.Q(is_tx_fifo_full_flag), .C(DEBUG_6_c), .E(VCC_net), 
            .D(n8987));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF \mem_LUT.data_buff_r__i4  (.Q(\fifo_temp_output[4] ), .C(DEBUG_6_c), 
           .D(n4111));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i5  (.Q(\fifo_temp_output[5] ), .C(DEBUG_6_c), 
           .D(n4123));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFF \mem_LUT.data_buff_r__i6  (.Q(\fifo_temp_output[6] ), .C(DEBUG_6_c), 
           .D(n4129));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(DEBUG_6_c), .E(VCC_net), 
            .D(n5317));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFE wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(DEBUG_6_c), .E(VCC_net), 
            .D(n5314));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFE rd_addr_r__i2 (.Q(rd_addr_r[2]), .C(DEBUG_6_c), .E(VCC_net), 
            .D(n5311));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFE rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(DEBUG_6_c), .E(VCC_net), 
            .D(n5308));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF i347_348 (.Q(\mem_LUT.mem_3_7 ), .C(DEBUG_6_c), .D(n5284));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i344_345 (.Q(\mem_LUT.mem_3_6 ), .C(DEBUG_6_c), .D(n5283));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i341_342 (.Q(\mem_LUT.mem_3_5 ), .C(DEBUG_6_c), .D(n5282));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i338_339 (.Q(\mem_LUT.mem_3_4 ), .C(DEBUG_6_c), .D(n5281));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i335_336 (.Q(\mem_LUT.mem_3_3 ), .C(DEBUG_6_c), .D(n5280));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i332_333 (.Q(\mem_LUT.mem_3_2 ), .C(DEBUG_6_c), .D(n5279));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i329_330 (.Q(\mem_LUT.mem_3_1 ), .C(DEBUG_6_c), .D(n5278));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i326_327 (.Q(\mem_LUT.mem_3_0 ), .C(DEBUG_6_c), .D(n5277));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i251_252 (.Q(\mem_LUT.mem_2_7 ), .C(DEBUG_6_c), .D(n5273));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i248_249 (.Q(\mem_LUT.mem_2_6 ), .C(DEBUG_6_c), .D(n5272));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i245_246 (.Q(\mem_LUT.mem_2_5 ), .C(DEBUG_6_c), .D(n5271));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i242_243 (.Q(\mem_LUT.mem_2_4 ), .C(DEBUG_6_c), .D(n5270));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i239_240 (.Q(\mem_LUT.mem_2_3 ), .C(DEBUG_6_c), .D(n5269));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i236_237 (.Q(\mem_LUT.mem_2_2 ), .C(DEBUG_6_c), .D(n5268));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i233_234 (.Q(\mem_LUT.mem_2_1 ), .C(DEBUG_6_c), .D(n5267));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i230_231 (.Q(\mem_LUT.mem_2_0 ), .C(DEBUG_6_c), .D(n5266));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i155_156 (.Q(\mem_LUT.mem_1_7 ), .C(DEBUG_6_c), .D(n5262));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i152_153 (.Q(\mem_LUT.mem_1_6 ), .C(DEBUG_6_c), .D(n5261));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i149_150 (.Q(\mem_LUT.mem_1_5 ), .C(DEBUG_6_c), .D(n5260));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i146_147 (.Q(\mem_LUT.mem_1_4 ), .C(DEBUG_6_c), .D(n5259));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i143_144 (.Q(\mem_LUT.mem_1_3 ), .C(DEBUG_6_c), .D(n5258));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i140_141 (.Q(\mem_LUT.mem_1_2 ), .C(DEBUG_6_c), .D(n5257));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i137_138 (.Q(\mem_LUT.mem_1_1 ), .C(DEBUG_6_c), .D(n5256));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i134_135 (.Q(\mem_LUT.mem_1_0 ), .C(DEBUG_6_c), .D(n5246));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i59_60 (.Q(\mem_LUT.mem_0_7 ), .C(DEBUG_6_c), .D(n5245));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i56_57 (.Q(\mem_LUT.mem_0_6 ), .C(DEBUG_6_c), .D(n5244));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i53_54 (.Q(\mem_LUT.mem_0_5 ), .C(DEBUG_6_c), .D(n5243));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i50_51 (.Q(\mem_LUT.mem_0_4 ), .C(DEBUG_6_c), .D(n5242));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i47_48 (.Q(\mem_LUT.mem_0_3 ), .C(DEBUG_6_c), .D(n5241));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i44_45 (.Q(\mem_LUT.mem_0_2 ), .C(DEBUG_6_c), .D(n5240));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i41_42 (.Q(\mem_LUT.mem_0_1 ), .C(DEBUG_6_c), .D(n5239));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i38_39 (.Q(\mem_LUT.mem_0_0 ), .C(DEBUG_6_c), .D(n5238));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF \mem_LUT.data_buff_r__i7  (.Q(\fifo_temp_output[7] ), .C(DEBUG_6_c), 
           .D(n4143));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 i4182_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_2_5 ), .O(n5271));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4182_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4181_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_2_4 ), .O(n5270));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4181_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1127_2_lut (.I0(rd_addr_r[1]), .I1(rd_addr_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(\rd_addr_p1_w[1] ));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1127_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1134_3_lut (.I0(rd_addr_r[2]), .I1(rd_addr_r[1]), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(\rd_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1134_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1105_2_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(\wr_addr_p1_w[1] ));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam i1105_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 wr_addr_r_1__I_0_i1_2_lut (.I0(wr_addr_r[0]), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(GND_net), .O(n1));   // src/fifo_quad_word_mod.v(115[26:58])
    defparam wr_addr_r_1__I_0_i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1112_3_lut (.I0(wr_addr_r[2]), .I1(wr_addr_r[1]), .I2(wr_addr_r[0]), 
            .I3(GND_net), .O(\wr_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam i1112_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_4_lut (.I0(n1), .I1(\wr_addr_p1_w[1] ), .I2(n3_adj_1093), 
            .I3(rd_addr_r[1]), .O(n8824));
    defparam i1_4_lut.LUT_INIT = 16'h8020;
    SB_LUT4 i4180_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_2_3 ), .O(n5269));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4180_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4179_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_2_2 ), .O(n5268));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4179_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4178_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_2_1 ), .O(n5267));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4178_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4177_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_2_0 ), .O(n5266));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4177_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE \mem_LUT.data_raw_r__i8  (.Q(\mem_LUT.data_raw_r[7] ), .C(DEBUG_6_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_968 [7]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i7  (.Q(\mem_LUT.data_raw_r[6] ), .C(DEBUG_6_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_968 [6]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i6  (.Q(\mem_LUT.data_raw_r[5] ), .C(DEBUG_6_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_968 [5]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 i4173_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_1_7 ), .O(n5262));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4173_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4172_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_1_6 ), .O(n5261));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4172_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4171_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_1_5 ), .O(n5260));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4171_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \mem_LUT.data_raw_r__i5  (.Q(\mem_LUT.data_raw_r[4] ), .C(DEBUG_6_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_968 [4]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i4  (.Q(\mem_LUT.data_raw_r[3] ), .C(DEBUG_6_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_968 [3]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i3  (.Q(\mem_LUT.data_raw_r[2] ), .C(DEBUG_6_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_968 [2]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i2  (.Q(\mem_LUT.data_raw_r[1] ), .C(DEBUG_6_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_968 [1]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_LUT4 i4170_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_1_4 ), .O(n5259));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4170_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4169_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_1_3 ), .O(n5258));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4169_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4168_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_1_2 ), .O(n5257));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4168_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4167_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_1_1 ), .O(n5256));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4167_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4157_3_lut_4_lut (.I0(n3), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_1_0 ), .O(n5246));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4157_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_en_i_I_0_2_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(GND_net), .I3(GND_net), .O(full_nxt_r));   // src/fifo_quad_word_mod.v(103[21:60])
    defparam wr_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10319 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_2 ), 
            .I2(\mem_LUT.mem_3_2 ), .I3(rd_addr_r[1]), .O(n11850));
    defparam rd_addr_r_0__bdd_4_lut_10319.LUT_INIT = 16'he4aa;
    SB_LUT4 n11850_bdd_4_lut (.I0(n11850), .I1(\mem_LUT.mem_1_2 ), .I2(\mem_LUT.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_968 [2]));
    defparam n11850_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10114 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_1 ), 
            .I2(\mem_LUT.mem_3_1 ), .I3(rd_addr_r[1]), .O(n11844));
    defparam rd_addr_r_0__bdd_4_lut_10114.LUT_INIT = 16'he4aa;
    SB_LUT4 n11844_bdd_4_lut (.I0(n11844), .I1(\mem_LUT.mem_1_1 ), .I2(\mem_LUT.mem_0_1 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_968 [1]));
    defparam n11844_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10109 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_0 ), 
            .I2(\mem_LUT.mem_3_0 ), .I3(rd_addr_r[1]), .O(n11832));
    defparam rd_addr_r_0__bdd_4_lut_10109.LUT_INIT = 16'he4aa;
    SB_LUT4 n11832_bdd_4_lut (.I0(n11832), .I1(\mem_LUT.mem_1_0 ), .I2(\mem_LUT.mem_0_0 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_968 [0]));
    defparam n11832_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4156_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_0_7 ), .O(n5245));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4156_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4155_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_0_6 ), .O(n5244));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4155_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4154_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_0_5 ), .O(n5243));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4154_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4153_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_0_4 ), .O(n5242));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4153_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4152_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_0_3 ), .O(n5241));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4152_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_en_i_I_0_2_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(GND_net), .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_quad_word_mod.v(62[29:51])
    defparam rd_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4151_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_0_2 ), .O(n5240));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4151_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4150_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_0_1 ), .O(n5239));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4150_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4149_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_0_0 ), .O(n5238));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4149_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF empty_r_85 (.Q(is_fifo_empty_flag), .C(DEBUG_6_c), .D(n9299));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF rd_fifo_en_prev_r_86 (.Q(rd_fifo_en_prev_r), .C(DEBUG_6_c), .D(n4093));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    SB_LUT4 wr_addr_p1_w_2__I_0_i3_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[0]), .I3(rd_addr_r[2]), .O(n3_adj_1093));   // src/fifo_quad_word_mod.v(107[37:64])
    defparam wr_addr_p1_w_2__I_0_i3_2_lut_4_lut.LUT_INIT = 16'h956a;
    SB_LUT4 EnabledDecoder_2_i3_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n3));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i3_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i4_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n4));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i4_2_lut_3_lut.LUT_INIT = 16'h0202;
    
endmodule
//
// Verilog Description of module usb3_if
//

module usb3_if (VCC_net, FIFO_CLK_c, FT_OE_c, GND_net, FT_RD_c, dc32_fifo_is_full, 
            FR_RXF_c, write_to_dc32_fifo) /* synthesis syn_module_defined=1 */ ;
    input VCC_net;
    input FIFO_CLK_c;
    output FT_OE_c;
    input GND_net;
    output FT_RD_c;
    input dc32_fifo_is_full;
    input FR_RXF_c;
    output write_to_dc32_fifo;
    
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    
    wire OE_N_N_90, OE_N, n2094, RD_N;
    
    SB_DFFNE OE_N_36 (.Q(OE_N), .C(FIFO_CLK_c), .E(VCC_net), .D(OE_N_N_90));   // src/usb3_if.v(57[8] 70[4])
    SB_DFFNE RD_N_37 (.Q(RD_N), .C(FIFO_CLK_c), .E(VCC_net), .D(n2094));   // src/usb3_if.v(57[8] 70[4])
    SB_LUT4 OE_N_I_0_1_lut (.I0(OE_N), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(FT_OE_c));   // src/usb3_if.v(53[16:23])
    defparam OE_N_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 RD_N_I_0_1_lut (.I0(RD_N), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(FT_RD_c));   // src/usb3_if.v(54[16:23])
    defparam RD_N_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut (.I0(dc32_fifo_is_full), .I1(OE_N), .I2(FR_RXF_c), 
            .I3(GND_net), .O(n2094));   // src/usb3_if.v(57[8] 70[4])
    defparam i2_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i9130_2_lut (.I0(FR_RXF_c), .I1(dc32_fifo_is_full), .I2(GND_net), 
            .I3(GND_net), .O(OE_N_N_90));   // src/usb3_if.v(58[9:57])
    defparam i9130_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2_4_lut (.I0(dc32_fifo_is_full), .I1(RD_N), .I2(FR_RXF_c), 
            .I3(OE_N), .O(write_to_dc32_fifo));   // src/usb3_if.v(74[9:93])
    defparam i2_4_lut.LUT_INIT = 16'h0400;
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=20) 
//

module \uart_rx(CLKS_PER_BIT=20)  (DEBUG_6_c, \r_SM_Main[2] , r_Rx_Data, 
            n5353, pc_data_rx, n5349, n5348, n5347, n5345, n5344, 
            n8963, VCC_net, debug_led3, n5339, n5338, n5337, r_Bit_Index, 
            GND_net, n4, \r_SM_Main[1] , n4_adj_1, n9345, n4_adj_2, 
            UART_RX_c, n2414, n3785, n3533, n3525, n3642, n131) /* synthesis syn_module_defined=1 */ ;
    input DEBUG_6_c;
    output \r_SM_Main[2] ;
    output r_Rx_Data;
    input n5353;
    output [7:0]pc_data_rx;
    input n5349;
    input n5348;
    input n5347;
    input n5345;
    input n5344;
    input n8963;
    input VCC_net;
    output debug_led3;
    input n5339;
    input n5338;
    input n5337;
    output [2:0]r_Bit_Index;
    input GND_net;
    output n4;
    output \r_SM_Main[1] ;
    output n4_adj_1;
    output n9345;
    output n4_adj_2;
    input UART_RX_c;
    output n2414;
    output n3785;
    output n3533;
    output n3525;
    output n3642;
    output n131;
    
    wire DEBUG_6_c /* synthesis SET_AS_NETWORK=DEBUG_6_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n3;
    wire [2:0]r_SM_Main;   // src/uart_rx.v(36[17:26])
    
    wire r_Rx_Data_R, n8813, n4_c, n9418;
    wire [2:0]r_Bit_Index_c;   // src/uart_rx.v(33[17:28])
    wire [9:0]n45;
    
    wire n5932;
    wire [9:0]r_Clock_Count;   // src/uart_rx.v(32[17:30])
    
    wire n5919, n9344, n154, n13, n9374, n33, n9027, n8794, 
        n8793, n8792, n8791, n8790, n8789, n8788, n8787, n8786, 
        n6, n147, n8, n4_adj_1090;
    wire [2:0]r_SM_Main_2__N_649;
    
    wire n55_adj_1091, n5950;
    wire [2:0]n340;
    
    wire n4016, n132;
    
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(DEBUG_6_c), .D(n3), .R(\r_SM_Main[2] ));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(DEBUG_6_c), .D(r_Rx_Data_R));   // src/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Byte_i7 (.Q(pc_data_rx[7]), .C(DEBUG_6_c), .D(n5353));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(pc_data_rx[6]), .C(DEBUG_6_c), .D(n5349));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(pc_data_rx[5]), .C(DEBUG_6_c), .D(n5348));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(pc_data_rx[4]), .C(DEBUG_6_c), .D(n5347));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(pc_data_rx[3]), .C(DEBUG_6_c), .D(n5345));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(pc_data_rx[0]), .C(DEBUG_6_c), .D(n5344));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Rx_DV_52 (.Q(debug_led3), .C(DEBUG_6_c), .E(VCC_net), .D(n8963));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(pc_data_rx[2]), .C(DEBUG_6_c), .D(n5339));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(pc_data_rx[1]), .C(DEBUG_6_c), .D(n5338));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(DEBUG_6_c), .E(VCC_net), 
            .D(n5337));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(DEBUG_6_c), .D(n8813));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(n4_c), .I2(GND_net), .I3(GND_net), 
            .O(n8813));   // src/uart_rx.v(49[10] 144[8])
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7877_2_lut (.I0(\r_SM_Main[2] ), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n9418));
    defparam i7877_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_132_i4_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // src/uart_rx.v(97[17:39])
    defparam equal_132_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESR r_Clock_Count_941__i0 (.Q(r_Clock_Count[0]), .C(DEBUG_6_c), 
            .E(n5932), .D(n45[0]), .R(n5919));   // src/uart_rx.v(120[34:51])
    SB_LUT4 i1_2_lut (.I0(\r_SM_Main[1] ), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n9344));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 equal_131_i4_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // src/uart_rx.v(97[17:39])
    defparam equal_131_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i3_4_lut (.I0(n154), .I1(n4_adj_1), .I2(r_SM_Main[0]), .I3(n9344), 
            .O(n9345));
    defparam i3_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 equal_128_i4_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // src/uart_rx.v(97[17:39])
    defparam equal_128_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i7834_2_lut (.I0(r_Rx_Data), .I1(n13), .I2(GND_net), .I3(GND_net), 
            .O(n9374));
    defparam i7834_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9127_4_lut (.I0(\r_SM_Main[1] ), .I1(\r_SM_Main[2] ), .I2(n33), 
            .I3(r_Rx_Data), .O(n5932));
    defparam i9127_4_lut.LUT_INIT = 16'h2333;
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(DEBUG_6_c), .D(UART_RX_c));   // src/uart_rx.v(41[10] 45[8])
    SB_DFFSR r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(DEBUG_6_c), .D(n9027), 
            .R(\r_SM_Main[2] ));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_941_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n8794), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_941_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_941_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n8793), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_941_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_941_add_4_10 (.CI(n8793), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n8794));
    SB_LUT4 r_Clock_Count_941_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[7]), 
            .I3(n8792), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_941_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_941_add_4_9 (.CI(n8792), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n8793));
    SB_LUT4 r_Clock_Count_941_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[6]), 
            .I3(n8791), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_941_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_941_add_4_8 (.CI(n8791), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n8792));
    SB_LUT4 r_Clock_Count_941_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[5]), 
            .I3(n8790), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_941_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_941_add_4_7 (.CI(n8790), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n8791));
    SB_LUT4 r_Clock_Count_941_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[4]), 
            .I3(n8789), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_941_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_941_add_4_6 (.CI(n8789), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n8790));
    SB_LUT4 r_Clock_Count_941_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[3]), 
            .I3(n8788), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_941_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_941_add_4_5 (.CI(n8788), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n8789));
    SB_LUT4 r_Clock_Count_941_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[2]), 
            .I3(n8787), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_941_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_941_add_4_4 (.CI(n8787), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n8788));
    SB_LUT4 r_Clock_Count_941_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[1]), 
            .I3(n8786), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_941_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_941_add_4_3 (.CI(n8786), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n8787));
    SB_LUT4 r_Clock_Count_941_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_941_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_941_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n8786));
    SB_DFFESR r_Clock_Count_941__i1 (.Q(r_Clock_Count[1]), .C(DEBUG_6_c), 
            .E(n5932), .D(n45[1]), .R(n5919));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_941__i2 (.Q(r_Clock_Count[2]), .C(DEBUG_6_c), 
            .E(n5932), .D(n45[2]), .R(n5919));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_941__i3 (.Q(r_Clock_Count[3]), .C(DEBUG_6_c), 
            .E(n5932), .D(n45[3]), .R(n5919));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_941__i4 (.Q(r_Clock_Count[4]), .C(DEBUG_6_c), 
            .E(n5932), .D(n45[4]), .R(n5919));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_941__i5 (.Q(r_Clock_Count[5]), .C(DEBUG_6_c), 
            .E(n5932), .D(n45[5]), .R(n5919));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_941__i6 (.Q(r_Clock_Count[6]), .C(DEBUG_6_c), 
            .E(n5932), .D(n45[6]), .R(n5919));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_941__i7 (.Q(r_Clock_Count[7]), .C(DEBUG_6_c), 
            .E(n5932), .D(n45[7]), .R(n5919));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_941__i8 (.Q(r_Clock_Count[8]), .C(DEBUG_6_c), 
            .E(n5932), .D(n45[8]), .R(n5919));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_941__i9 (.Q(r_Clock_Count[9]), .C(DEBUG_6_c), 
            .E(n5932), .D(n45[9]), .R(n5919));   // src/uart_rx.v(120[34:51])
    SB_LUT4 i1_2_lut_adj_38 (.I0(r_Clock_Count[9]), .I1(r_Clock_Count[7]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // src/uart_rx.v(32[17:30])
    defparam i1_2_lut_adj_38.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[5]), 
            .I3(n6), .O(n147));   // src/uart_rx.v(32[17:30])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_39 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), 
            .I2(r_Clock_Count[3]), .I3(r_Clock_Count[4]), .O(n8));
    defparam i3_4_lut_adj_39.LUT_INIT = 16'hffdf;
    SB_LUT4 i4_3_lut (.I0(n147), .I1(n8), .I2(r_Clock_Count[2]), .I3(GND_net), 
            .O(n13));
    defparam i4_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_40 (.I0(r_SM_Main[0]), .I1(n13), .I2(GND_net), 
            .I3(GND_net), .O(n33));
    defparam i1_2_lut_adj_40.LUT_INIT = 16'h2222;
    SB_LUT4 i1341_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), .I2(GND_net), 
            .I3(GND_net), .O(n2414));   // src/uart_rx.v(100[21:36])
    defparam i1341_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[0]), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n4_adj_1090));   // src/uart_rx.v(118[17:47])
    defparam i1_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[4]), .I1(n147), .I2(r_Clock_Count[3]), 
            .I3(n4_adj_1090), .O(r_SM_Main_2__N_649[2]));   // src/uart_rx.v(32[17:30])
    defparam i1_4_lut.LUT_INIT = 16'heeec;
    SB_LUT4 i1_2_lut_adj_41 (.I0(r_SM_Main_2__N_649[2]), .I1(r_Bit_Index[0]), 
            .I2(GND_net), .I3(GND_net), .O(n154));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_41.LUT_INIT = 16'h8888;
    SB_LUT4 i54_3_lut (.I0(n55_adj_1091), .I1(n5950), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n3));   // src/uart_rx.v(30[17:26])
    defparam i54_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index_c[1]), .C(DEBUG_6_c), .E(n3785), 
            .D(n340[1]), .R(n4016));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index_c[2]), .C(DEBUG_6_c), .E(n3785), 
            .D(n340[2]), .R(n4016));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i20_4_lut (.I0(n9374), .I1(r_SM_Main_2__N_649[2]), .I2(\r_SM_Main[1] ), 
            .I3(r_SM_Main[0]), .O(n9027));   // src/uart_rx.v(30[17:26])
    defparam i20_4_lut.LUT_INIT = 16'h35f0;
    SB_LUT4 i1_2_lut_3_lut (.I0(r_SM_Main[0]), .I1(n4_c), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n3533));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_42 (.I0(r_SM_Main[0]), .I1(n4_c), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n3525));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_adj_42.LUT_INIT = 16'hbfbf;
    SB_LUT4 i26_4_lut_4_lut (.I0(\r_SM_Main[2] ), .I1(r_SM_Main_2__N_649[2]), 
            .I2(n132), .I3(\r_SM_Main[1] ), .O(n5919));   // src/uart_rx.v(49[10] 144[8])
    defparam i26_4_lut_4_lut.LUT_INIT = 16'h4405;
    SB_LUT4 i1_2_lut_3_lut_adj_43 (.I0(\r_SM_Main[2] ), .I1(r_SM_Main_2__N_649[2]), 
            .I2(\r_SM_Main[1] ), .I3(GND_net), .O(n4_c));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_adj_43.LUT_INIT = 16'h4040;
    SB_LUT4 i53_4_lut_3_lut (.I0(r_SM_Main[0]), .I1(n13), .I2(r_Rx_Data), 
            .I3(GND_net), .O(n55_adj_1091));   // src/uart_rx.v(30[17:26])
    defparam i53_4_lut_3_lut.LUT_INIT = 16'h8d8d;
    SB_LUT4 i4861_4_lut_4_lut (.I0(r_SM_Main_2__N_649[2]), .I1(r_Bit_Index[0]), 
            .I2(r_SM_Main[0]), .I3(n2414), .O(n5950));   // src/uart_rx.v(36[17:26])
    defparam i4861_4_lut_4_lut.LUT_INIT = 16'h5850;
    SB_LUT4 i1_2_lut_3_lut_adj_44 (.I0(r_Rx_Data), .I1(n13), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n132));   // src/uart_rx.v(30[17:26])
    defparam i1_2_lut_3_lut_adj_44.LUT_INIT = 16'he0e0;
    SB_LUT4 i13_4_lut_4_lut (.I0(\r_SM_Main[1] ), .I1(\r_SM_Main[2] ), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main_2__N_649[2]), .O(n3642));
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2505;
    SB_LUT4 i1061_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n340[1]));   // src/uart_rx.v(102[36:51])
    defparam i1061_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_45 (.I0(r_SM_Main_2__N_649[2]), .I1(n9418), .I2(\r_SM_Main[1] ), 
            .I3(n131), .O(n4016));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_4_lut_adj_45.LUT_INIT = 16'h2303;
    SB_LUT4 i1068_3_lut (.I0(r_Bit_Index_c[2]), .I1(r_Bit_Index_c[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n340[2]));   // src/uart_rx.v(102[36:51])
    defparam i1068_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main_2__N_649[2]), .I1(\r_SM_Main[2] ), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main[1] ), .O(n3785));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0203;
    SB_LUT4 i1_2_lut_3_lut_adj_46 (.I0(r_Bit_Index[0]), .I1(r_Bit_Index_c[1]), 
            .I2(r_Bit_Index_c[2]), .I3(GND_net), .O(n131));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_adj_46.LUT_INIT = 16'h8080;
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen
//

module fifo_dc_32_lut_gen (FIFO_D6_c_6, \REG.mem_42_15 , \REG.mem_43_15 , 
            FIFO_D5_c_5, \REG.mem_29_14 , \REG.mem_28_14 , FIFO_CLK_c, 
            \REG.mem_41_15 , \REG.mem_40_15 , GND_net, \REG.mem_2_0 , 
            \REG.mem_2_2 , FIFO_D4_c_4, \REG.mem_18_5 , \REG.mem_19_5 , 
            FIFO_D3_c_3, \REG.mem_62_5 , \REG.mem_61_5 , \REG.mem_60_5 , 
            FIFO_D2_c_2, t_rd_fifo_en_w, \REG.out_raw[0] , DEBUG_6_c, 
            \REG.mem_30_10 , \REG.mem_29_10 , \REG.mem_28_10 , \REG.mem_58_8 , 
            \REG.mem_57_8 , \REG.mem_56_8 , FIFO_D1_c_1, \REG.mem_2_14 , 
            FIFO_D0_c_0, \REG.mem_14_15 , \REG.mem_15_15 , \REG.mem_13_15 , 
            \REG.mem_12_15 , \REG.mem_10_15 , \REG.mem_11_15 , n56, 
            \REG.mem_62_8 , \REG.mem_61_8 , \REG.mem_60_8 , \REG.mem_46_6 , 
            \REG.mem_47_6 , n24, write_to_dc32_fifo, reset_all, \wr_addr_nxt_c[1] , 
            \REG.mem_45_6 , \REG.mem_44_6 , dc32_fifo_is_full, \REG.mem_34_10 , 
            \REG.mem_18_8 , \REG.mem_19_8 , \REG.mem_58_11 , \rd_grey_sync_r[0] , 
            \REG.mem_57_11 , \REG.mem_56_11 , \REG.mem_6_14 , \REG.mem_7_14 , 
            \REG.mem_5_14 , \REG.mem_10_12 , \REG.mem_11_12 , \REG.mem_9_12 , 
            \REG.mem_8_12 , \REG.mem_6_10 , \REG.mem_7_10 , \REG.mem_26_9 , 
            DEBUG_1_c, \REG.mem_6_0 , \REG.mem_7_0 , \REG.mem_5_0 , 
            \REG.mem_5_10 , \REG.mem_25_9 , \REG.mem_24_9 , \REG.mem_56_7 , 
            \REG.mem_57_7 , \REG.mem_58_7 , \num_words_in_buffer[3] , 
            \wr_grey_sync_r[0] , \REG.mem_10_14 , \REG.mem_11_14 , \REG.mem_9_14 , 
            \REG.mem_8_14 , \REG.mem_14_14 , \REG.mem_15_14 , \REG.mem_13_14 , 
            \REG.mem_12_14 , \REG.mem_38_9 , \REG.mem_39_9 , \REG.mem_37_9 , 
            \REG.mem_34_7 , \REG.mem_42_9 , \REG.mem_43_9 , \REG.mem_10_10 , 
            \REG.mem_11_10 , \REG.mem_9_10 , \REG.mem_8_10 , \REG.mem_41_9 , 
            \REG.mem_40_9 , \REG.mem_9_15 , \REG.mem_8_15 , \REG.mem_18_6 , 
            \REG.mem_19_6 , \wr_addr_nxt_c[3] , FIFO_D15_c_15, \REG.mem_22_5 , 
            \REG.mem_23_5 , \REG.mem_21_5 , \REG.mem_38_10 , \REG.mem_39_10 , 
            \REG.mem_37_10 , \REG.mem_18_10 , \REG.mem_19_10 , FIFO_D14_c_14, 
            \REG.mem_34_12 , \REG.mem_22_6 , \REG.mem_23_6 , \REG.mem_26_14 , 
            \REG.mem_25_14 , \REG.mem_24_14 , \REG.mem_18_13 , \REG.mem_19_13 , 
            \REG.mem_62_7 , \REG.mem_21_6 , \REG.mem_60_7 , \REG.mem_61_7 , 
            \REG.mem_30_14 , \REG.mem_50_3 , \REG.mem_51_3 , \REG.mem_38_12 , 
            \REG.mem_39_12 , \REG.mem_37_12 , \REG.mem_46_8 , \REG.mem_47_8 , 
            \REG.mem_45_8 , \REG.mem_44_8 , \REG.mem_58_10 , \REG.mem_2_3 , 
            \REG.mem_57_10 , \REG.mem_56_10 , \REG.mem_62_2 , \REG.mem_61_2 , 
            \REG.mem_60_2 , \REG.mem_58_15 , \REG.mem_10_0 , \REG.mem_11_0 , 
            \REG.mem_9_0 , \REG.mem_8_0 , \REG.mem_57_15 , \REG.mem_56_15 , 
            \REG.mem_30_0 , \REG.mem_29_0 , \REG.mem_28_0 , \REG.mem_38_7 , 
            \REG.mem_39_7 , FIFO_D13_c_13, \REG.mem_37_7 , n58, FIFO_D12_c_12, 
            \REG.mem_26_5 , \REG.mem_25_5 , \REG.mem_24_5 , n50, \REG.mem_46_0 , 
            \REG.mem_47_0 , \REG.mem_6_3 , \REG.mem_7_3 , \REG.mem_5_3 , 
            \REG.mem_45_0 , \REG.mem_44_0 , \REG.mem_50_8 , \REG.mem_51_8 , 
            n18, \REG.mem_10_3 , \REG.mem_11_3 , \REG.mem_6_2 , \REG.mem_7_2 , 
            \REG.mem_5_2 , \REG.mem_9_3 , \REG.mem_8_3 , \wr_addr_nxt_c[5] , 
            \REG.mem_42_12 , \REG.mem_43_12 , \REG.mem_41_12 , \REG.mem_40_12 , 
            \REG.mem_10_2 , \REG.mem_11_2 , n4169, \REG.mem_2_15 , \REG.mem_9_2 , 
            \REG.mem_8_2 , n4168, n4167, \REG.mem_2_13 , n4166, \REG.mem_2_12 , 
            n4165, \REG.mem_2_11 , n4164, \REG.mem_2_10 , \REG.mem_6_6 , 
            \REG.mem_7_6 , n4163, \REG.mem_2_9 , \REG.mem_5_6 , \REG.mem_30_3 , 
            \REG.mem_29_3 , \REG.mem_28_3 , \REG.mem_22_13 , \REG.mem_23_13 , 
            \REG.mem_21_13 , \REG.mem_54_3 , \REG.mem_55_3 , \REG.mem_53_3 , 
            \REG.mem_42_10 , \REG.mem_43_10 , \REG.mem_41_10 , \REG.mem_40_10 , 
            \REG.mem_56_4 , \REG.mem_57_4 , \REG.mem_6_15 , \REG.mem_7_15 , 
            \REG.mem_58_4 , \REG.mem_26_15 , \REG.mem_5_15 , \REG.mem_25_15 , 
            \REG.mem_24_15 , \REG.mem_58_3 , \REG.mem_57_3 , \REG.mem_56_3 , 
            \REG.mem_62_3 , \REG.mem_62_4 , \REG.mem_60_4 , \REG.mem_61_4 , 
            \REG.mem_61_3 , \REG.mem_60_3 , \rd_addr_r[6] , \rd_addr_nxt_c_6__N_176[5] , 
            \REG.mem_22_8 , \REG.mem_23_8 , \rd_addr_nxt_c_6__N_176[3] , 
            \REG.mem_21_8 , \REG.mem_54_8 , \REG.mem_55_8 , FIFO_D11_c_11, 
            \REG.mem_14_3 , \REG.mem_15_3 , \REG.mem_53_8 , \REG.mem_14_2 , 
            \REG.mem_15_2 , \REG.mem_13_3 , \REG.mem_12_3 , \REG.mem_13_2 , 
            \REG.mem_12_2 , \REG.mem_30_5 , \REG.mem_58_13 , \REG.mem_29_5 , 
            \REG.mem_28_5 , \REG.mem_34_5 , \REG.mem_57_13 , \REG.mem_56_13 , 
            \REG.mem_14_6 , \REG.mem_15_6 , \REG.mem_13_6 , \REG.mem_12_6 , 
            \REG.mem_54_9 , \REG.mem_55_9 , \REG.mem_53_9 , \REG.mem_34_0 , 
            \REG.mem_14_0 , \REG.mem_15_0 , \REG.mem_13_0 , \REG.mem_12_0 , 
            FIFO_D10_c_10, \REG.mem_42_14 , \REG.mem_43_14 , \REG.mem_41_14 , 
            \REG.mem_40_14 , n4162, \REG.mem_2_8 , n4161, \REG.mem_2_7 , 
            FIFO_D9_c_9, n5327, VCC_net, \fifo_data_out[0] , \REG.mem_10_11 , 
            \REG.mem_11_11 , FIFO_D8_c_8, FIFO_D7_c_7, \REG.mem_9_11 , 
            \REG.mem_8_11 , \REG.mem_62_15 , \REG.mem_62_10 , n5305, 
            \fifo_data_out[15] , \REG.mem_46_12 , \REG.mem_47_12 , n5302, 
            \fifo_data_out[14] , \REG.mem_61_10 , \REG.mem_60_10 , \REG.mem_61_15 , 
            \REG.mem_60_15 , n5299, \fifo_data_out[13] , n5296, \fifo_data_out[12] , 
            n5293, \fifo_data_out[11] , n5290, \fifo_data_out[10] , 
            \REG.mem_45_12 , \REG.mem_44_12 , \REG.mem_46_15 , \REG.mem_47_15 , 
            \REG.mem_18_3 , \REG.mem_19_3 , n5255, \fifo_data_out[9] , 
            n5252, \fifo_data_out[8] , n5249, \fifo_data_out[7] , \REG.mem_45_15 , 
            \REG.mem_44_15 , n4160, \REG.mem_2_6 , \REG.mem_14_11 , 
            \REG.mem_15_11 , n4159, \REG.mem_2_5 , n5236, \fifo_data_out[6] , 
            n5233, \fifo_data_out[5] , \REG.mem_13_11 , \REG.mem_12_11 , 
            n5230, \fifo_data_out[4] , \wr_grey_sync_r[5] , \wr_grey_sync_r[4] , 
            \wr_grey_sync_r[3] , n5212, \fifo_data_out[3] , \REG.mem_18_2 , 
            \REG.mem_19_2 , n5208, n5207, \REG.mem_62_14 , n5206, 
            \REG.mem_62_13 , n5205, \REG.mem_62_12 , n5204, \REG.mem_62_11 , 
            n5203, n5202, \REG.mem_62_9 , n5201, n5200, \wr_grey_sync_r[2] , 
            \wr_grey_sync_r[1] , n5199, \REG.mem_62_6 , n5198, n5197, 
            n5196, n5195, n5194, \REG.mem_62_1 , n5193, \REG.mem_62_0 , 
            n5192, n5191, \REG.mem_61_14 , n5190, \REG.mem_61_13 , 
            n5189, \REG.mem_61_12 , n5188, \REG.mem_61_11 , n5187, 
            n5186, \REG.mem_61_9 , n5185, n5184, n5183, \REG.mem_61_6 , 
            \REG.mem_22_3 , \REG.mem_23_3 , \REG.mem_26_8 , n5182, \REG.mem_21_3 , 
            n5181, n5180, n5179, n5178, \REG.mem_61_1 , n5177, \REG.mem_61_0 , 
            n5176, n5175, \REG.mem_60_14 , n5174, \REG.mem_60_13 , 
            n5173, \REG.mem_60_12 , n5172, \REG.mem_60_11 , n5171, 
            n5170, \REG.mem_60_9 , n5169, n5168, n5167, \REG.mem_60_6 , 
            \REG.mem_25_8 , \REG.mem_24_8 , \REG.mem_46_9 , \REG.mem_47_9 , 
            \REG.mem_45_9 , \REG.mem_44_9 , \REG.mem_30_7 , n5166, n5165, 
            n5164, n5163, n5162, \REG.mem_60_1 , n5161, \REG.mem_60_0 , 
            \REG.mem_29_7 , \REG.mem_28_7 , n5144, n5143, \REG.mem_58_14 , 
            n5142, n5141, \REG.mem_58_12 , n5140, n5139, n5138, 
            \REG.mem_58_9 , n5137, n5136, n5135, \REG.mem_58_6 , \REG.mem_46_10 , 
            \REG.mem_47_10 , \REG.mem_45_10 , \REG.mem_44_10 , n5134, 
            \REG.mem_58_5 , \REG.mem_30_9 , n5133, n5132, n5131, \REG.mem_58_2 , 
            n5130, \REG.mem_58_1 , n5129, \REG.mem_58_0 , n5128, n5127, 
            \REG.mem_57_14 , n5126, n5125, \REG.mem_57_12 , n5124, 
            n5123, n5122, \REG.mem_57_9 , n5121, n5120, n5119, \REG.mem_57_6 , 
            \REG.mem_29_9 , \REG.mem_28_9 , n5118, \REG.mem_57_5 , n5117, 
            n5116, n5115, \REG.mem_57_2 , n5114, \REG.mem_57_1 , n5113, 
            \fifo_data_out[2] , n5110, \REG.mem_57_0 , n5109, n5108, 
            \REG.mem_56_14 , n5107, n5106, \REG.mem_56_12 , n5105, 
            n5104, n5103, \REG.mem_56_9 , \REG.mem_10_6 , \REG.mem_11_6 , 
            n5102, \REG.mem_9_6 , \REG.mem_8_6 , n5101, n5100, \REG.mem_56_6 , 
            n5099, \REG.mem_56_5 , n5098, n5097, n5096, \REG.mem_56_2 , 
            n5095, \REG.mem_56_1 , n5094, \fifo_data_out[1] , n5091, 
            \REG.mem_56_0 , n5090, \REG.mem_55_15 , n5089, \REG.mem_55_14 , 
            n5088, \REG.mem_55_13 , n5087, \REG.mem_55_12 , \REG.mem_22_2 , 
            \REG.mem_23_2 , \REG.mem_21_2 , n5086, \REG.mem_55_11 , 
            n5085, \REG.mem_55_10 , n5084, n5083, n5082, \REG.mem_55_7 , 
            n5081, \REG.mem_55_6 , n5080, \REG.mem_55_5 , n5079, \REG.mem_55_4 , 
            n5078, n5077, \REG.mem_55_2 , n5076, \REG.mem_55_1 , n5075, 
            \REG.mem_55_0 , n5074, \REG.mem_54_15 , n5073, \REG.mem_54_14 , 
            n5072, \REG.mem_54_13 , \num_words_in_buffer[6] , \num_words_in_buffer[5] , 
            \num_words_in_buffer[4] , n5071, \REG.mem_54_12 , n5070, 
            \REG.mem_54_11 , n5069, \REG.mem_54_10 , n5068, n5067, 
            n5066, \REG.mem_54_7 , n5065, \REG.mem_54_6 , n5064, \REG.mem_54_5 , 
            n5063, \REG.mem_54_4 , n5062, n5061, \REG.mem_54_2 , n5060, 
            \REG.mem_54_1 , n5057, \REG.mem_54_0 , n5056, \REG.mem_53_15 , 
            n5055, \REG.mem_53_14 , \REG.mem_50_12 , \REG.mem_51_12 , 
            \REG.mem_38_5 , \REG.mem_39_5 , \REG.mem_37_5 , n5054, \REG.mem_53_13 , 
            n5053, \REG.mem_53_12 , n5052, \REG.mem_53_11 , n5051, 
            \REG.mem_53_10 , n5050, n5049, n5048, \REG.mem_53_7 , 
            n5047, \REG.mem_53_6 , n5046, \REG.mem_53_5 , n5045, \REG.mem_53_4 , 
            n5044, n5043, \REG.mem_53_2 , n5042, \REG.mem_53_1 , n5041, 
            \REG.mem_53_0 , \REG.mem_26_2 , \REG.mem_18_11 , \REG.mem_19_11 , 
            \REG.mem_25_2 , \REG.mem_24_2 , n5024, \REG.mem_51_15 , 
            n5023, \REG.mem_51_14 , n26, \REG.mem_26_3 , \REG.mem_25_3 , 
            \REG.mem_24_3 , \REG.mem_40_4 , \REG.mem_41_4 , n5022, \REG.mem_51_13 , 
            n5021, n5020, \REG.mem_51_11 , n5019, \REG.mem_51_10 , 
            n5018, \REG.mem_51_9 , n5017, n5016, \REG.mem_51_7 , n5015, 
            \REG.mem_51_6 , n5014, \REG.mem_51_5 , n5013, \REG.mem_51_4 , 
            n5012, n5011, \REG.mem_51_2 , n5010, \REG.mem_51_1 , n5008, 
            \REG.mem_51_0 , \REG.mem_42_4 , \REG.mem_43_4 , \REG.mem_22_11 , 
            \REG.mem_23_11 , n5007, \REG.mem_50_15 , n5006, \REG.mem_50_14 , 
            n5005, \REG.mem_50_13 , n5004, n5003, \REG.mem_50_11 , 
            n5002, \REG.mem_50_10 , n5001, \REG.mem_50_9 , n5000, 
            n4999, \REG.mem_50_7 , n4998, \REG.mem_50_6 , n4997, \REG.mem_50_5 , 
            n4996, \REG.mem_50_4 , n4995, n4994, \REG.mem_50_2 , n4993, 
            \REG.mem_50_1 , n4992, \REG.mem_50_0 , \REG.mem_21_11 , 
            \rd_addr_nxt_c_6__N_176[1] , n4158, \REG.mem_2_4 , \REG.mem_30_15 , 
            \REG.mem_29_15 , \REG.mem_28_15 , \REG.mem_30_8 , \REG.mem_29_8 , 
            \REG.mem_28_8 , \REG.mem_46_4 , \REG.mem_47_4 , n4946, n4945, 
            \REG.mem_47_14 , n4944, \REG.mem_47_13 , \rd_grey_sync_r[5] , 
            \rd_grey_sync_r[4] , \rd_grey_sync_r[3] , \rd_grey_sync_r[2] , 
            \rd_grey_sync_r[1] , n4943, \REG.mem_44_4 , \REG.mem_45_4 , 
            n4942, \REG.mem_47_11 , n4941, n4940, n4939, n4938, 
            \REG.mem_47_7 , n4937, n4936, \REG.mem_47_5 , n4935, n4934, 
            \REG.mem_47_3 , n4933, \REG.mem_47_2 , n4932, \REG.mem_47_1 , 
            n4929, n4928, n4927, \REG.mem_46_14 , \wr_addr_r[6] , 
            n4926, \REG.mem_46_13 , n4925, n4924, \REG.mem_46_11 , 
            n4923, n4922, n4921, n4920, \REG.mem_46_7 , n4919, n4918, 
            \REG.mem_46_5 , n4917, n4916, \REG.mem_46_3 , n4915, \REG.mem_46_2 , 
            n4914, \REG.mem_46_1 , n4913, n4912, n4911, \REG.mem_45_14 , 
            n59, n4910, \REG.mem_45_13 , n4909, n4908, \REG.mem_45_11 , 
            n4907, n4906, n4905, n4904, \REG.mem_45_7 , n4903, n4902, 
            \REG.mem_45_5 , n4901, n4900, \REG.mem_45_3 , n4899, \REG.mem_45_2 , 
            n4898, \REG.mem_45_1 , n4897, n4896, n27, n4895, \REG.mem_44_14 , 
            n4894, \REG.mem_44_13 , n4893, n4892, \REG.mem_44_11 , 
            n4891, n4890, n4889, n4888, \REG.mem_44_7 , n4887, n4886, 
            \REG.mem_44_5 , n4885, n4884, \REG.mem_44_3 , n4883, \REG.mem_44_2 , 
            n4882, \REG.mem_44_1 , n4880, n4879, n4878, n4877, \REG.mem_43_13 , 
            n4876, n4875, \REG.mem_43_11 , n4874, n4873, n4872, 
            \REG.mem_43_8 , n4871, \REG.mem_43_7 , n4870, \REG.mem_43_6 , 
            n4869, \REG.mem_43_5 , n4868, n4867, \REG.mem_43_3 , n4866, 
            \REG.mem_43_2 , n4865, \REG.mem_43_1 , n4864, \REG.mem_43_0 , 
            n4863, \REG.mem_30_2 , n4862, n4861, \REG.mem_42_13 , 
            n4860, n4859, \REG.mem_42_11 , n4858, n4857, n4856, 
            \REG.mem_42_8 , n4855, \REG.mem_42_7 , n4854, \REG.mem_42_6 , 
            n4853, \REG.mem_42_5 , n4852, n4851, \REG.mem_42_3 , n4850, 
            \REG.mem_42_2 , n4849, \REG.mem_42_1 , n4848, \REG.mem_42_0 , 
            n4847, \REG.mem_29_2 , \REG.mem_28_2 , \REG.mem_26_11 , 
            \REG.mem_6_7 , \REG.mem_7_7 , \REG.mem_5_7 , n4846, n4845, 
            \REG.mem_41_13 , n4844, n4843, \REG.mem_41_11 , n4842, 
            n4841, n4840, \REG.mem_41_8 , n4839, \REG.mem_41_7 , n4838, 
            \REG.mem_41_6 , n4837, \REG.mem_41_5 , n4836, n4835, \REG.mem_41_3 , 
            n4834, \REG.mem_41_2 , n4833, \REG.mem_41_1 , n4832, \REG.mem_41_0 , 
            \REG.mem_18_7 , \REG.mem_19_7 , \REG.mem_25_11 , \REG.mem_24_11 , 
            n4157, n4831, n4830, n4829, \REG.mem_40_13 , n4828, 
            n4827, \REG.mem_40_11 , n4826, n4825, n4824, \REG.mem_40_8 , 
            n4823, \REG.mem_40_7 , n4822, \REG.mem_40_6 , n4821, \REG.mem_40_5 , 
            n4820, n4819, \REG.mem_40_3 , n4818, \REG.mem_40_2 , n4817, 
            \REG.mem_40_1 , n4814, \REG.mem_40_0 , n4813, \REG.mem_39_15 , 
            n4812, \REG.mem_39_14 , \REG.mem_22_7 , \REG.mem_23_7 , 
            n4811, \REG.mem_39_13 , n4810, n4809, \REG.mem_39_11 , 
            \REG.mem_21_7 , n4808, \REG.mem_30_11 , n4807, n4806, 
            \REG.mem_39_8 , n4805, n4804, \REG.mem_39_6 , n4803, n4802, 
            \REG.mem_39_4 , n4801, \REG.mem_39_3 , n4800, \REG.mem_39_2 , 
            n4799, \REG.mem_39_1 , n4798, \REG.mem_39_0 , n4797, \REG.mem_38_15 , 
            n4796, \REG.mem_38_14 , n4795, \REG.mem_38_13 , n4794, 
            n4793, \REG.mem_38_11 , \REG.mem_29_11 , \REG.mem_28_11 , 
            n4792, \REG.mem_34_2 , n4791, n4790, \REG.mem_38_8 , n4789, 
            n4788, \REG.mem_38_6 , n4787, n4786, \REG.mem_38_4 , n4785, 
            \REG.mem_38_3 , n4784, \REG.mem_38_2 , n4783, \REG.mem_38_1 , 
            n4782, \REG.mem_38_0 , n4781, \REG.mem_37_15 , n4780, 
            \REG.mem_37_14 , n4779, \REG.mem_37_13 , n4778, n4777, 
            \REG.mem_37_11 , n4776, n4775, n4774, \REG.mem_37_8 , 
            n4773, n4772, \REG.mem_37_6 , n4771, n4770, \REG.mem_37_4 , 
            n4769, \REG.mem_37_3 , n4768, \REG.mem_37_2 , n4767, \REG.mem_37_1 , 
            n4766, \REG.mem_37_0 , n4156, \REG.mem_26_6 , \REG.mem_25_6 , 
            \REG.mem_24_6 , \REG.mem_34_9 , n4733, \REG.mem_34_15 , 
            n4732, \REG.mem_34_14 , n4731, \REG.mem_34_13 , n4730, 
            n4729, \REG.mem_34_11 , n4728, n4727, n4726, \REG.mem_34_8 , 
            n4725, n4155, \REG.mem_2_1 , n4154, \REG.mem_24_4 , \REG.mem_25_4 , 
            \REG.mem_26_4 , n4724, \REG.mem_34_6 , \REG.mem_30_4 , \REG.mem_28_4 , 
            \REG.mem_29_4 , n4723, n4722, \REG.mem_34_4 , n4721, \REG.mem_34_3 , 
            n4720, n4719, \REG.mem_34_1 , n4718, \REG.mem_8_4 , \REG.mem_9_4 , 
            \REG.mem_10_4 , \REG.mem_11_4 , \REG.mem_14_4 , \REG.mem_15_4 , 
            \REG.mem_12_4 , \REG.mem_13_4 , \REG.mem_6_1 , \REG.mem_7_1 , 
            \REG.mem_5_1 , n4677, rp_sync1_r, \REG.mem_26_10 , \REG.mem_18_1 , 
            \REG.mem_19_1 , n4676, n4675, n4674, n4673, n4672, \REG.mem_25_10 , 
            \REG.mem_24_10 , \REG.mem_22_1 , \REG.mem_23_1 , \REG.mem_21_1 , 
            n46, n14, n4655, n4654, n4653, n4652, n4651, n4650, 
            n4649, n4648, n4647, \REG.mem_30_13 , n4646, \REG.mem_30_12 , 
            n4645, n37, n5, n4644, n4643, n4642, n4641, n4640, 
            \REG.mem_30_6 , n4639, n4638, n4637, n4636, n4635, \REG.mem_30_1 , 
            n4634, n4633, n4631, n4629, \REG.mem_18_14 , \REG.mem_19_14 , 
            n4627, n51, n4626, n4625, \REG.mem_29_13 , \REG.mem_22_14 , 
            \REG.mem_23_14 , \REG.mem_21_14 , n4624, \REG.mem_29_12 , 
            n4623, n4622, n4621, n4620, n4619, n4618, \REG.mem_29_6 , 
            n4617, n4616, n4615, n4614, n4613, \REG.mem_29_1 , n4612, 
            n4611, n4610, n4609, \REG.mem_28_13 , n19, n4608, \REG.mem_28_12 , 
            n4607, \REG.mem_18_12 , \REG.mem_19_12 , \REG.mem_22_12 , 
            \REG.mem_23_12 , n4606, n4605, n4604, n4603, n4602, 
            \REG.mem_28_6 , n4601, n4600, n4599, n4598, n4597, \REG.mem_28_1 , 
            n4596, \REG.mem_21_12 , n4579, n4578, n4577, \REG.mem_26_13 , 
            n4576, \REG.mem_26_12 , n4575, n4574, n4573, n4572, 
            n4571, \REG.mem_26_7 , n4570, n4569, n4568, n4567, \REG.mem_6_13 , 
            \REG.mem_7_13 , n4566, n4565, \REG.mem_26_1 , n4564, \REG.mem_26_0 , 
            n4563, wp_sync1_r, n4562, n4561, n4560, n4559, n4558, 
            n4557, n4556, \REG.mem_25_13 , n4555, \REG.mem_25_12 , 
            n4554, n4553, n4552, n4551, \REG.mem_5_13 , n4550, \REG.mem_25_7 , 
            n4549, n4548, n4547, n4546, n4545, n4544, \REG.mem_25_1 , 
            n4543, \REG.mem_25_0 , n4542, n4541, n4540, n4539, n4538, 
            n4537, n4536, n4535, n4534, \REG.mem_18_0 , \REG.mem_19_0 , 
            \REG.mem_22_0 , \REG.mem_23_0 , \REG.mem_21_0 , DEBUG_9_c, 
            n4533, \REG.mem_24_13 , n4532, \REG.mem_24_12 , n4531, 
            n4530, n4529, n4528, n4527, \REG.mem_24_7 , n4526, n4525, 
            n4524, n4523, n4522, n4521, \REG.mem_24_1 , n4520, \REG.mem_24_0 , 
            n4519, \REG.mem_23_15 , n4518, n4517, n4516, n4515, 
            n4514, \REG.mem_23_10 , n4513, \REG.mem_23_9 , n4512, 
            n4511, n4510, n4509, n4508, \REG.mem_23_4 , n4507, n4506, 
            n4505, n4504, n4503, \REG.mem_22_15 , n4502, n4501, 
            n4500, n4499, n4498, \REG.mem_22_10 , n4497, \REG.mem_22_9 , 
            n4496, n4495, n4494, n4493, n4492, \REG.mem_22_4 , n4491, 
            n4490, n4489, n4488, n4487, \REG.mem_21_15 , n4486, 
            n4485, n4484, n4483, n4482, \REG.mem_21_10 , n4481, 
            \REG.mem_21_9 , n4480, n4479, n4478, n4477, n4476, \REG.mem_21_4 , 
            n4475, n4474, n4473, \REG.mem_6_12 , \REG.mem_7_12 , n4472, 
            \REG.out_raw[15] , \REG.out_raw[14] , \REG.out_raw[13] , \REG.mem_5_12 , 
            \REG.out_raw[12] , \REG.out_raw[11] , \REG.out_raw[10] , n4455, 
            \REG.mem_19_15 , n4454, n4453, n4452, n4451, n4450, 
            n4449, \REG.mem_19_9 , n4448, n4447, n4446, n4445, n4444, 
            \REG.mem_19_4 , n4443, n4442, n4441, n4440, \REG.out_raw[9] , 
            \REG.out_raw[8] , n4439, \REG.mem_18_15 , \REG.out_raw[7] , 
            \REG.out_raw[6] , \REG.out_raw[5] , \REG.out_raw[4] , \REG.out_raw[3] , 
            n4438, \REG.mem_6_9 , \REG.mem_7_9 , n54, \REG.mem_5_9 , 
            n4437, n4436, n4435, n4434, n4433, \REG.mem_18_9 , n4432, 
            n4431, n4430, n4429, n4428, \REG.mem_18_4 , n4427, n4426, 
            n4425, n4424, \REG.out_raw[2] , n22, n39, \REG.mem_10_9 , 
            \REG.mem_11_9 , \REG.mem_10_13 , \REG.mem_11_13 , n7, n40, 
            \REG.mem_9_9 , \REG.mem_8_9 , \REG.mem_9_13 , \REG.mem_8_13 , 
            n8, \REG.mem_14_12 , \REG.mem_15_12 , n4391, \REG.out_raw[1] , 
            n4390, \REG.mem_13_12 , \REG.mem_12_12 , n4389, \REG.mem_15_13 , 
            n4388, n4387, n4386, \REG.mem_15_10 , n4385, \REG.mem_15_9 , 
            n4384, \REG.mem_15_8 , n4383, \REG.mem_15_7 , n4382, n4381, 
            \REG.mem_15_5 , n4380, n4379, n4378, n4377, \REG.mem_15_1 , 
            n4376, n4375, n4374, \REG.mem_6_8 , \REG.mem_7_8 , \REG.mem_5_8 , 
            \REG.mem_14_9 , \REG.mem_13_9 , \REG.mem_12_9 , \REG.mem_6_5 , 
            \REG.mem_7_5 , n4373, \REG.mem_14_13 , n4372, n4371, n4370, 
            \REG.mem_14_10 , n4369, n4368, \REG.mem_14_8 , n4367, 
            \REG.mem_14_7 , \REG.mem_5_5 , n4366, n4365, \REG.mem_14_5 , 
            n4364, n4363, n4362, n4361, \REG.mem_14_1 , n4360, n4359, 
            n4358, n4357, \REG.mem_13_13 , n4356, n4355, n4354, 
            \REG.mem_13_10 , n4353, n4352, \REG.mem_13_8 , n4351, 
            \REG.mem_13_7 , n4350, n4349, \REG.mem_13_5 , n4348, n4347, 
            n4346, n4345, \REG.mem_13_1 , n4344, n4343, n4342, n4341, 
            \REG.mem_12_13 , n4340, n4339, n4338, \REG.mem_12_10 , 
            n4337, n4336, \REG.mem_12_8 , n4335, \REG.mem_12_7 , n4334, 
            n4333, \REG.mem_12_5 , n4332, n4331, n4330, n4329, \REG.mem_12_1 , 
            n4328, n4327, n4326, n4325, n4324, n4323, n60, n4322, 
            n28, n41, n9, n4321, n4320, \REG.mem_11_8 , n4319, 
            \REG.mem_11_7 , n4318, n4317, \REG.mem_11_5 , n4316, n4315, 
            n4314, n4313, \REG.mem_11_1 , n4312, n4311, n42, n4310, 
            n4309, n4308, n10, n4307, n4306, n4305, n4304, \REG.mem_10_8 , 
            n4303, \REG.mem_10_7 , n4302, n4301, \REG.mem_10_5 , n4300, 
            n4299, n4298, n4297, \REG.mem_10_1 , n4296, n4130, n57, 
            \REG.mem_9_5 , \REG.mem_8_5 , n4288, n4287, n4286, n4285, 
            n4284, n4283, n4282, n4281, n4280, \REG.mem_9_8 , n4279, 
            \REG.mem_9_7 , n4278, n4277, n4108, n25, n4276, n43, 
            n11, n44, n12, n4275, n4274, n4273, \REG.mem_9_1 , 
            n4272, n4270, n4268, n4107, \REG.mem_8_7 , n4265, n4264, 
            n4263, n4262, n4261, n52, n4260, \REG.mem_8_8 , n4259, 
            n4258, n4257, n4256, n4255, n4254, n4253, n4252, n4251, 
            \REG.mem_8_1 , n4250, n4249, n4248, n4247, n4246, n4245, 
            \REG.mem_7_11 , n4244, n4243, n4242, n4241, n4240, n4239, 
            n4238, \REG.mem_7_4 , n4237, n4236, n4235, n4234, n4233, 
            n4232, n4231, n4230, n4229, \REG.mem_6_11 , n4228, n4227, 
            n4226, n4225, n4224, n4223, n4222, \REG.mem_6_4 , n4221, 
            n4220, n4219, n4218, n4217, n4216, n4215, n4214, n4213, 
            \REG.mem_5_11 , n4212, n4211, n4210, n4209, n4208, n4207, 
            n4206, \REG.mem_5_4 , n4205, n4204, n4203, n4202, n4103, 
            n20, n53, n4101, n21, n35, n3, n36, n55, n23, 
            n4, n47, n15, n31, n63) /* synthesis syn_module_defined=1 */ ;
    input FIFO_D6_c_6;
    output \REG.mem_42_15 ;
    output \REG.mem_43_15 ;
    input FIFO_D5_c_5;
    output \REG.mem_29_14 ;
    output \REG.mem_28_14 ;
    input FIFO_CLK_c;
    output \REG.mem_41_15 ;
    output \REG.mem_40_15 ;
    input GND_net;
    output \REG.mem_2_0 ;
    output \REG.mem_2_2 ;
    input FIFO_D4_c_4;
    output \REG.mem_18_5 ;
    output \REG.mem_19_5 ;
    input FIFO_D3_c_3;
    output \REG.mem_62_5 ;
    output \REG.mem_61_5 ;
    output \REG.mem_60_5 ;
    input FIFO_D2_c_2;
    output t_rd_fifo_en_w;
    output \REG.out_raw[0] ;
    input DEBUG_6_c;
    output \REG.mem_30_10 ;
    output \REG.mem_29_10 ;
    output \REG.mem_28_10 ;
    output \REG.mem_58_8 ;
    output \REG.mem_57_8 ;
    output \REG.mem_56_8 ;
    input FIFO_D1_c_1;
    output \REG.mem_2_14 ;
    input FIFO_D0_c_0;
    output \REG.mem_14_15 ;
    output \REG.mem_15_15 ;
    output \REG.mem_13_15 ;
    output \REG.mem_12_15 ;
    output \REG.mem_10_15 ;
    output \REG.mem_11_15 ;
    output n56;
    output \REG.mem_62_8 ;
    output \REG.mem_61_8 ;
    output \REG.mem_60_8 ;
    output \REG.mem_46_6 ;
    output \REG.mem_47_6 ;
    output n24;
    input write_to_dc32_fifo;
    input reset_all;
    output \wr_addr_nxt_c[1] ;
    output \REG.mem_45_6 ;
    output \REG.mem_44_6 ;
    output dc32_fifo_is_full;
    output \REG.mem_34_10 ;
    output \REG.mem_18_8 ;
    output \REG.mem_19_8 ;
    output \REG.mem_58_11 ;
    output \rd_grey_sync_r[0] ;
    output \REG.mem_57_11 ;
    output \REG.mem_56_11 ;
    output \REG.mem_6_14 ;
    output \REG.mem_7_14 ;
    output \REG.mem_5_14 ;
    output \REG.mem_10_12 ;
    output \REG.mem_11_12 ;
    output \REG.mem_9_12 ;
    output \REG.mem_8_12 ;
    output \REG.mem_6_10 ;
    output \REG.mem_7_10 ;
    output \REG.mem_26_9 ;
    output DEBUG_1_c;
    output \REG.mem_6_0 ;
    output \REG.mem_7_0 ;
    output \REG.mem_5_0 ;
    output \REG.mem_5_10 ;
    output \REG.mem_25_9 ;
    output \REG.mem_24_9 ;
    output \REG.mem_56_7 ;
    output \REG.mem_57_7 ;
    output \REG.mem_58_7 ;
    output \num_words_in_buffer[3] ;
    output \wr_grey_sync_r[0] ;
    output \REG.mem_10_14 ;
    output \REG.mem_11_14 ;
    output \REG.mem_9_14 ;
    output \REG.mem_8_14 ;
    output \REG.mem_14_14 ;
    output \REG.mem_15_14 ;
    output \REG.mem_13_14 ;
    output \REG.mem_12_14 ;
    output \REG.mem_38_9 ;
    output \REG.mem_39_9 ;
    output \REG.mem_37_9 ;
    output \REG.mem_34_7 ;
    output \REG.mem_42_9 ;
    output \REG.mem_43_9 ;
    output \REG.mem_10_10 ;
    output \REG.mem_11_10 ;
    output \REG.mem_9_10 ;
    output \REG.mem_8_10 ;
    output \REG.mem_41_9 ;
    output \REG.mem_40_9 ;
    output \REG.mem_9_15 ;
    output \REG.mem_8_15 ;
    output \REG.mem_18_6 ;
    output \REG.mem_19_6 ;
    output \wr_addr_nxt_c[3] ;
    input FIFO_D15_c_15;
    output \REG.mem_22_5 ;
    output \REG.mem_23_5 ;
    output \REG.mem_21_5 ;
    output \REG.mem_38_10 ;
    output \REG.mem_39_10 ;
    output \REG.mem_37_10 ;
    output \REG.mem_18_10 ;
    output \REG.mem_19_10 ;
    input FIFO_D14_c_14;
    output \REG.mem_34_12 ;
    output \REG.mem_22_6 ;
    output \REG.mem_23_6 ;
    output \REG.mem_26_14 ;
    output \REG.mem_25_14 ;
    output \REG.mem_24_14 ;
    output \REG.mem_18_13 ;
    output \REG.mem_19_13 ;
    output \REG.mem_62_7 ;
    output \REG.mem_21_6 ;
    output \REG.mem_60_7 ;
    output \REG.mem_61_7 ;
    output \REG.mem_30_14 ;
    output \REG.mem_50_3 ;
    output \REG.mem_51_3 ;
    output \REG.mem_38_12 ;
    output \REG.mem_39_12 ;
    output \REG.mem_37_12 ;
    output \REG.mem_46_8 ;
    output \REG.mem_47_8 ;
    output \REG.mem_45_8 ;
    output \REG.mem_44_8 ;
    output \REG.mem_58_10 ;
    output \REG.mem_2_3 ;
    output \REG.mem_57_10 ;
    output \REG.mem_56_10 ;
    output \REG.mem_62_2 ;
    output \REG.mem_61_2 ;
    output \REG.mem_60_2 ;
    output \REG.mem_58_15 ;
    output \REG.mem_10_0 ;
    output \REG.mem_11_0 ;
    output \REG.mem_9_0 ;
    output \REG.mem_8_0 ;
    output \REG.mem_57_15 ;
    output \REG.mem_56_15 ;
    output \REG.mem_30_0 ;
    output \REG.mem_29_0 ;
    output \REG.mem_28_0 ;
    output \REG.mem_38_7 ;
    output \REG.mem_39_7 ;
    input FIFO_D13_c_13;
    output \REG.mem_37_7 ;
    output n58;
    input FIFO_D12_c_12;
    output \REG.mem_26_5 ;
    output \REG.mem_25_5 ;
    output \REG.mem_24_5 ;
    output n50;
    output \REG.mem_46_0 ;
    output \REG.mem_47_0 ;
    output \REG.mem_6_3 ;
    output \REG.mem_7_3 ;
    output \REG.mem_5_3 ;
    output \REG.mem_45_0 ;
    output \REG.mem_44_0 ;
    output \REG.mem_50_8 ;
    output \REG.mem_51_8 ;
    output n18;
    output \REG.mem_10_3 ;
    output \REG.mem_11_3 ;
    output \REG.mem_6_2 ;
    output \REG.mem_7_2 ;
    output \REG.mem_5_2 ;
    output \REG.mem_9_3 ;
    output \REG.mem_8_3 ;
    output \wr_addr_nxt_c[5] ;
    output \REG.mem_42_12 ;
    output \REG.mem_43_12 ;
    output \REG.mem_41_12 ;
    output \REG.mem_40_12 ;
    output \REG.mem_10_2 ;
    output \REG.mem_11_2 ;
    input n4169;
    output \REG.mem_2_15 ;
    output \REG.mem_9_2 ;
    output \REG.mem_8_2 ;
    input n4168;
    input n4167;
    output \REG.mem_2_13 ;
    input n4166;
    output \REG.mem_2_12 ;
    input n4165;
    output \REG.mem_2_11 ;
    input n4164;
    output \REG.mem_2_10 ;
    output \REG.mem_6_6 ;
    output \REG.mem_7_6 ;
    input n4163;
    output \REG.mem_2_9 ;
    output \REG.mem_5_6 ;
    output \REG.mem_30_3 ;
    output \REG.mem_29_3 ;
    output \REG.mem_28_3 ;
    output \REG.mem_22_13 ;
    output \REG.mem_23_13 ;
    output \REG.mem_21_13 ;
    output \REG.mem_54_3 ;
    output \REG.mem_55_3 ;
    output \REG.mem_53_3 ;
    output \REG.mem_42_10 ;
    output \REG.mem_43_10 ;
    output \REG.mem_41_10 ;
    output \REG.mem_40_10 ;
    output \REG.mem_56_4 ;
    output \REG.mem_57_4 ;
    output \REG.mem_6_15 ;
    output \REG.mem_7_15 ;
    output \REG.mem_58_4 ;
    output \REG.mem_26_15 ;
    output \REG.mem_5_15 ;
    output \REG.mem_25_15 ;
    output \REG.mem_24_15 ;
    output \REG.mem_58_3 ;
    output \REG.mem_57_3 ;
    output \REG.mem_56_3 ;
    output \REG.mem_62_3 ;
    output \REG.mem_62_4 ;
    output \REG.mem_60_4 ;
    output \REG.mem_61_4 ;
    output \REG.mem_61_3 ;
    output \REG.mem_60_3 ;
    output \rd_addr_r[6] ;
    output \rd_addr_nxt_c_6__N_176[5] ;
    output \REG.mem_22_8 ;
    output \REG.mem_23_8 ;
    output \rd_addr_nxt_c_6__N_176[3] ;
    output \REG.mem_21_8 ;
    output \REG.mem_54_8 ;
    output \REG.mem_55_8 ;
    input FIFO_D11_c_11;
    output \REG.mem_14_3 ;
    output \REG.mem_15_3 ;
    output \REG.mem_53_8 ;
    output \REG.mem_14_2 ;
    output \REG.mem_15_2 ;
    output \REG.mem_13_3 ;
    output \REG.mem_12_3 ;
    output \REG.mem_13_2 ;
    output \REG.mem_12_2 ;
    output \REG.mem_30_5 ;
    output \REG.mem_58_13 ;
    output \REG.mem_29_5 ;
    output \REG.mem_28_5 ;
    output \REG.mem_34_5 ;
    output \REG.mem_57_13 ;
    output \REG.mem_56_13 ;
    output \REG.mem_14_6 ;
    output \REG.mem_15_6 ;
    output \REG.mem_13_6 ;
    output \REG.mem_12_6 ;
    output \REG.mem_54_9 ;
    output \REG.mem_55_9 ;
    output \REG.mem_53_9 ;
    output \REG.mem_34_0 ;
    output \REG.mem_14_0 ;
    output \REG.mem_15_0 ;
    output \REG.mem_13_0 ;
    output \REG.mem_12_0 ;
    input FIFO_D10_c_10;
    output \REG.mem_42_14 ;
    output \REG.mem_43_14 ;
    output \REG.mem_41_14 ;
    output \REG.mem_40_14 ;
    input n4162;
    output \REG.mem_2_8 ;
    input n4161;
    output \REG.mem_2_7 ;
    input FIFO_D9_c_9;
    input n5327;
    input VCC_net;
    output \fifo_data_out[0] ;
    output \REG.mem_10_11 ;
    output \REG.mem_11_11 ;
    input FIFO_D8_c_8;
    input FIFO_D7_c_7;
    output \REG.mem_9_11 ;
    output \REG.mem_8_11 ;
    output \REG.mem_62_15 ;
    output \REG.mem_62_10 ;
    input n5305;
    output \fifo_data_out[15] ;
    output \REG.mem_46_12 ;
    output \REG.mem_47_12 ;
    input n5302;
    output \fifo_data_out[14] ;
    output \REG.mem_61_10 ;
    output \REG.mem_60_10 ;
    output \REG.mem_61_15 ;
    output \REG.mem_60_15 ;
    input n5299;
    output \fifo_data_out[13] ;
    input n5296;
    output \fifo_data_out[12] ;
    input n5293;
    output \fifo_data_out[11] ;
    input n5290;
    output \fifo_data_out[10] ;
    output \REG.mem_45_12 ;
    output \REG.mem_44_12 ;
    output \REG.mem_46_15 ;
    output \REG.mem_47_15 ;
    output \REG.mem_18_3 ;
    output \REG.mem_19_3 ;
    input n5255;
    output \fifo_data_out[9] ;
    input n5252;
    output \fifo_data_out[8] ;
    input n5249;
    output \fifo_data_out[7] ;
    output \REG.mem_45_15 ;
    output \REG.mem_44_15 ;
    input n4160;
    output \REG.mem_2_6 ;
    output \REG.mem_14_11 ;
    output \REG.mem_15_11 ;
    input n4159;
    output \REG.mem_2_5 ;
    input n5236;
    output \fifo_data_out[6] ;
    input n5233;
    output \fifo_data_out[5] ;
    output \REG.mem_13_11 ;
    output \REG.mem_12_11 ;
    input n5230;
    output \fifo_data_out[4] ;
    output \wr_grey_sync_r[5] ;
    output \wr_grey_sync_r[4] ;
    output \wr_grey_sync_r[3] ;
    input n5212;
    output \fifo_data_out[3] ;
    output \REG.mem_18_2 ;
    output \REG.mem_19_2 ;
    input n5208;
    input n5207;
    output \REG.mem_62_14 ;
    input n5206;
    output \REG.mem_62_13 ;
    input n5205;
    output \REG.mem_62_12 ;
    input n5204;
    output \REG.mem_62_11 ;
    input n5203;
    input n5202;
    output \REG.mem_62_9 ;
    input n5201;
    input n5200;
    output \wr_grey_sync_r[2] ;
    output \wr_grey_sync_r[1] ;
    input n5199;
    output \REG.mem_62_6 ;
    input n5198;
    input n5197;
    input n5196;
    input n5195;
    input n5194;
    output \REG.mem_62_1 ;
    input n5193;
    output \REG.mem_62_0 ;
    input n5192;
    input n5191;
    output \REG.mem_61_14 ;
    input n5190;
    output \REG.mem_61_13 ;
    input n5189;
    output \REG.mem_61_12 ;
    input n5188;
    output \REG.mem_61_11 ;
    input n5187;
    input n5186;
    output \REG.mem_61_9 ;
    input n5185;
    input n5184;
    input n5183;
    output \REG.mem_61_6 ;
    output \REG.mem_22_3 ;
    output \REG.mem_23_3 ;
    output \REG.mem_26_8 ;
    input n5182;
    output \REG.mem_21_3 ;
    input n5181;
    input n5180;
    input n5179;
    input n5178;
    output \REG.mem_61_1 ;
    input n5177;
    output \REG.mem_61_0 ;
    input n5176;
    input n5175;
    output \REG.mem_60_14 ;
    input n5174;
    output \REG.mem_60_13 ;
    input n5173;
    output \REG.mem_60_12 ;
    input n5172;
    output \REG.mem_60_11 ;
    input n5171;
    input n5170;
    output \REG.mem_60_9 ;
    input n5169;
    input n5168;
    input n5167;
    output \REG.mem_60_6 ;
    output \REG.mem_25_8 ;
    output \REG.mem_24_8 ;
    output \REG.mem_46_9 ;
    output \REG.mem_47_9 ;
    output \REG.mem_45_9 ;
    output \REG.mem_44_9 ;
    output \REG.mem_30_7 ;
    input n5166;
    input n5165;
    input n5164;
    input n5163;
    input n5162;
    output \REG.mem_60_1 ;
    input n5161;
    output \REG.mem_60_0 ;
    output \REG.mem_29_7 ;
    output \REG.mem_28_7 ;
    input n5144;
    input n5143;
    output \REG.mem_58_14 ;
    input n5142;
    input n5141;
    output \REG.mem_58_12 ;
    input n5140;
    input n5139;
    input n5138;
    output \REG.mem_58_9 ;
    input n5137;
    input n5136;
    input n5135;
    output \REG.mem_58_6 ;
    output \REG.mem_46_10 ;
    output \REG.mem_47_10 ;
    output \REG.mem_45_10 ;
    output \REG.mem_44_10 ;
    input n5134;
    output \REG.mem_58_5 ;
    output \REG.mem_30_9 ;
    input n5133;
    input n5132;
    input n5131;
    output \REG.mem_58_2 ;
    input n5130;
    output \REG.mem_58_1 ;
    input n5129;
    output \REG.mem_58_0 ;
    input n5128;
    input n5127;
    output \REG.mem_57_14 ;
    input n5126;
    input n5125;
    output \REG.mem_57_12 ;
    input n5124;
    input n5123;
    input n5122;
    output \REG.mem_57_9 ;
    input n5121;
    input n5120;
    input n5119;
    output \REG.mem_57_6 ;
    output \REG.mem_29_9 ;
    output \REG.mem_28_9 ;
    input n5118;
    output \REG.mem_57_5 ;
    input n5117;
    input n5116;
    input n5115;
    output \REG.mem_57_2 ;
    input n5114;
    output \REG.mem_57_1 ;
    input n5113;
    output \fifo_data_out[2] ;
    input n5110;
    output \REG.mem_57_0 ;
    input n5109;
    input n5108;
    output \REG.mem_56_14 ;
    input n5107;
    input n5106;
    output \REG.mem_56_12 ;
    input n5105;
    input n5104;
    input n5103;
    output \REG.mem_56_9 ;
    output \REG.mem_10_6 ;
    output \REG.mem_11_6 ;
    input n5102;
    output \REG.mem_9_6 ;
    output \REG.mem_8_6 ;
    input n5101;
    input n5100;
    output \REG.mem_56_6 ;
    input n5099;
    output \REG.mem_56_5 ;
    input n5098;
    input n5097;
    input n5096;
    output \REG.mem_56_2 ;
    input n5095;
    output \REG.mem_56_1 ;
    input n5094;
    output \fifo_data_out[1] ;
    input n5091;
    output \REG.mem_56_0 ;
    input n5090;
    output \REG.mem_55_15 ;
    input n5089;
    output \REG.mem_55_14 ;
    input n5088;
    output \REG.mem_55_13 ;
    input n5087;
    output \REG.mem_55_12 ;
    output \REG.mem_22_2 ;
    output \REG.mem_23_2 ;
    output \REG.mem_21_2 ;
    input n5086;
    output \REG.mem_55_11 ;
    input n5085;
    output \REG.mem_55_10 ;
    input n5084;
    input n5083;
    input n5082;
    output \REG.mem_55_7 ;
    input n5081;
    output \REG.mem_55_6 ;
    input n5080;
    output \REG.mem_55_5 ;
    input n5079;
    output \REG.mem_55_4 ;
    input n5078;
    input n5077;
    output \REG.mem_55_2 ;
    input n5076;
    output \REG.mem_55_1 ;
    input n5075;
    output \REG.mem_55_0 ;
    input n5074;
    output \REG.mem_54_15 ;
    input n5073;
    output \REG.mem_54_14 ;
    input n5072;
    output \REG.mem_54_13 ;
    output \num_words_in_buffer[6] ;
    output \num_words_in_buffer[5] ;
    output \num_words_in_buffer[4] ;
    input n5071;
    output \REG.mem_54_12 ;
    input n5070;
    output \REG.mem_54_11 ;
    input n5069;
    output \REG.mem_54_10 ;
    input n5068;
    input n5067;
    input n5066;
    output \REG.mem_54_7 ;
    input n5065;
    output \REG.mem_54_6 ;
    input n5064;
    output \REG.mem_54_5 ;
    input n5063;
    output \REG.mem_54_4 ;
    input n5062;
    input n5061;
    output \REG.mem_54_2 ;
    input n5060;
    output \REG.mem_54_1 ;
    input n5057;
    output \REG.mem_54_0 ;
    input n5056;
    output \REG.mem_53_15 ;
    input n5055;
    output \REG.mem_53_14 ;
    output \REG.mem_50_12 ;
    output \REG.mem_51_12 ;
    output \REG.mem_38_5 ;
    output \REG.mem_39_5 ;
    output \REG.mem_37_5 ;
    input n5054;
    output \REG.mem_53_13 ;
    input n5053;
    output \REG.mem_53_12 ;
    input n5052;
    output \REG.mem_53_11 ;
    input n5051;
    output \REG.mem_53_10 ;
    input n5050;
    input n5049;
    input n5048;
    output \REG.mem_53_7 ;
    input n5047;
    output \REG.mem_53_6 ;
    input n5046;
    output \REG.mem_53_5 ;
    input n5045;
    output \REG.mem_53_4 ;
    input n5044;
    input n5043;
    output \REG.mem_53_2 ;
    input n5042;
    output \REG.mem_53_1 ;
    input n5041;
    output \REG.mem_53_0 ;
    output \REG.mem_26_2 ;
    output \REG.mem_18_11 ;
    output \REG.mem_19_11 ;
    output \REG.mem_25_2 ;
    output \REG.mem_24_2 ;
    input n5024;
    output \REG.mem_51_15 ;
    input n5023;
    output \REG.mem_51_14 ;
    output n26;
    output \REG.mem_26_3 ;
    output \REG.mem_25_3 ;
    output \REG.mem_24_3 ;
    output \REG.mem_40_4 ;
    output \REG.mem_41_4 ;
    input n5022;
    output \REG.mem_51_13 ;
    input n5021;
    input n5020;
    output \REG.mem_51_11 ;
    input n5019;
    output \REG.mem_51_10 ;
    input n5018;
    output \REG.mem_51_9 ;
    input n5017;
    input n5016;
    output \REG.mem_51_7 ;
    input n5015;
    output \REG.mem_51_6 ;
    input n5014;
    output \REG.mem_51_5 ;
    input n5013;
    output \REG.mem_51_4 ;
    input n5012;
    input n5011;
    output \REG.mem_51_2 ;
    input n5010;
    output \REG.mem_51_1 ;
    input n5008;
    output \REG.mem_51_0 ;
    output \REG.mem_42_4 ;
    output \REG.mem_43_4 ;
    output \REG.mem_22_11 ;
    output \REG.mem_23_11 ;
    input n5007;
    output \REG.mem_50_15 ;
    input n5006;
    output \REG.mem_50_14 ;
    input n5005;
    output \REG.mem_50_13 ;
    input n5004;
    input n5003;
    output \REG.mem_50_11 ;
    input n5002;
    output \REG.mem_50_10 ;
    input n5001;
    output \REG.mem_50_9 ;
    input n5000;
    input n4999;
    output \REG.mem_50_7 ;
    input n4998;
    output \REG.mem_50_6 ;
    input n4997;
    output \REG.mem_50_5 ;
    input n4996;
    output \REG.mem_50_4 ;
    input n4995;
    input n4994;
    output \REG.mem_50_2 ;
    input n4993;
    output \REG.mem_50_1 ;
    input n4992;
    output \REG.mem_50_0 ;
    output \REG.mem_21_11 ;
    output \rd_addr_nxt_c_6__N_176[1] ;
    input n4158;
    output \REG.mem_2_4 ;
    output \REG.mem_30_15 ;
    output \REG.mem_29_15 ;
    output \REG.mem_28_15 ;
    output \REG.mem_30_8 ;
    output \REG.mem_29_8 ;
    output \REG.mem_28_8 ;
    output \REG.mem_46_4 ;
    output \REG.mem_47_4 ;
    input n4946;
    input n4945;
    output \REG.mem_47_14 ;
    input n4944;
    output \REG.mem_47_13 ;
    output \rd_grey_sync_r[5] ;
    output \rd_grey_sync_r[4] ;
    output \rd_grey_sync_r[3] ;
    output \rd_grey_sync_r[2] ;
    output \rd_grey_sync_r[1] ;
    input n4943;
    output \REG.mem_44_4 ;
    output \REG.mem_45_4 ;
    input n4942;
    output \REG.mem_47_11 ;
    input n4941;
    input n4940;
    input n4939;
    input n4938;
    output \REG.mem_47_7 ;
    input n4937;
    input n4936;
    output \REG.mem_47_5 ;
    input n4935;
    input n4934;
    output \REG.mem_47_3 ;
    input n4933;
    output \REG.mem_47_2 ;
    input n4932;
    output \REG.mem_47_1 ;
    input n4929;
    input n4928;
    input n4927;
    output \REG.mem_46_14 ;
    output \wr_addr_r[6] ;
    input n4926;
    output \REG.mem_46_13 ;
    input n4925;
    input n4924;
    output \REG.mem_46_11 ;
    input n4923;
    input n4922;
    input n4921;
    input n4920;
    output \REG.mem_46_7 ;
    input n4919;
    input n4918;
    output \REG.mem_46_5 ;
    input n4917;
    input n4916;
    output \REG.mem_46_3 ;
    input n4915;
    output \REG.mem_46_2 ;
    input n4914;
    output \REG.mem_46_1 ;
    input n4913;
    input n4912;
    input n4911;
    output \REG.mem_45_14 ;
    output n59;
    input n4910;
    output \REG.mem_45_13 ;
    input n4909;
    input n4908;
    output \REG.mem_45_11 ;
    input n4907;
    input n4906;
    input n4905;
    input n4904;
    output \REG.mem_45_7 ;
    input n4903;
    input n4902;
    output \REG.mem_45_5 ;
    input n4901;
    input n4900;
    output \REG.mem_45_3 ;
    input n4899;
    output \REG.mem_45_2 ;
    input n4898;
    output \REG.mem_45_1 ;
    input n4897;
    input n4896;
    output n27;
    input n4895;
    output \REG.mem_44_14 ;
    input n4894;
    output \REG.mem_44_13 ;
    input n4893;
    input n4892;
    output \REG.mem_44_11 ;
    input n4891;
    input n4890;
    input n4889;
    input n4888;
    output \REG.mem_44_7 ;
    input n4887;
    input n4886;
    output \REG.mem_44_5 ;
    input n4885;
    input n4884;
    output \REG.mem_44_3 ;
    input n4883;
    output \REG.mem_44_2 ;
    input n4882;
    output \REG.mem_44_1 ;
    input n4880;
    input n4879;
    input n4878;
    input n4877;
    output \REG.mem_43_13 ;
    input n4876;
    input n4875;
    output \REG.mem_43_11 ;
    input n4874;
    input n4873;
    input n4872;
    output \REG.mem_43_8 ;
    input n4871;
    output \REG.mem_43_7 ;
    input n4870;
    output \REG.mem_43_6 ;
    input n4869;
    output \REG.mem_43_5 ;
    input n4868;
    input n4867;
    output \REG.mem_43_3 ;
    input n4866;
    output \REG.mem_43_2 ;
    input n4865;
    output \REG.mem_43_1 ;
    input n4864;
    output \REG.mem_43_0 ;
    input n4863;
    output \REG.mem_30_2 ;
    input n4862;
    input n4861;
    output \REG.mem_42_13 ;
    input n4860;
    input n4859;
    output \REG.mem_42_11 ;
    input n4858;
    input n4857;
    input n4856;
    output \REG.mem_42_8 ;
    input n4855;
    output \REG.mem_42_7 ;
    input n4854;
    output \REG.mem_42_6 ;
    input n4853;
    output \REG.mem_42_5 ;
    input n4852;
    input n4851;
    output \REG.mem_42_3 ;
    input n4850;
    output \REG.mem_42_2 ;
    input n4849;
    output \REG.mem_42_1 ;
    input n4848;
    output \REG.mem_42_0 ;
    input n4847;
    output \REG.mem_29_2 ;
    output \REG.mem_28_2 ;
    output \REG.mem_26_11 ;
    output \REG.mem_6_7 ;
    output \REG.mem_7_7 ;
    output \REG.mem_5_7 ;
    input n4846;
    input n4845;
    output \REG.mem_41_13 ;
    input n4844;
    input n4843;
    output \REG.mem_41_11 ;
    input n4842;
    input n4841;
    input n4840;
    output \REG.mem_41_8 ;
    input n4839;
    output \REG.mem_41_7 ;
    input n4838;
    output \REG.mem_41_6 ;
    input n4837;
    output \REG.mem_41_5 ;
    input n4836;
    input n4835;
    output \REG.mem_41_3 ;
    input n4834;
    output \REG.mem_41_2 ;
    input n4833;
    output \REG.mem_41_1 ;
    input n4832;
    output \REG.mem_41_0 ;
    output \REG.mem_18_7 ;
    output \REG.mem_19_7 ;
    output \REG.mem_25_11 ;
    output \REG.mem_24_11 ;
    input n4157;
    input n4831;
    input n4830;
    input n4829;
    output \REG.mem_40_13 ;
    input n4828;
    input n4827;
    output \REG.mem_40_11 ;
    input n4826;
    input n4825;
    input n4824;
    output \REG.mem_40_8 ;
    input n4823;
    output \REG.mem_40_7 ;
    input n4822;
    output \REG.mem_40_6 ;
    input n4821;
    output \REG.mem_40_5 ;
    input n4820;
    input n4819;
    output \REG.mem_40_3 ;
    input n4818;
    output \REG.mem_40_2 ;
    input n4817;
    output \REG.mem_40_1 ;
    input n4814;
    output \REG.mem_40_0 ;
    input n4813;
    output \REG.mem_39_15 ;
    input n4812;
    output \REG.mem_39_14 ;
    output \REG.mem_22_7 ;
    output \REG.mem_23_7 ;
    input n4811;
    output \REG.mem_39_13 ;
    input n4810;
    input n4809;
    output \REG.mem_39_11 ;
    output \REG.mem_21_7 ;
    input n4808;
    output \REG.mem_30_11 ;
    input n4807;
    input n4806;
    output \REG.mem_39_8 ;
    input n4805;
    input n4804;
    output \REG.mem_39_6 ;
    input n4803;
    input n4802;
    output \REG.mem_39_4 ;
    input n4801;
    output \REG.mem_39_3 ;
    input n4800;
    output \REG.mem_39_2 ;
    input n4799;
    output \REG.mem_39_1 ;
    input n4798;
    output \REG.mem_39_0 ;
    input n4797;
    output \REG.mem_38_15 ;
    input n4796;
    output \REG.mem_38_14 ;
    input n4795;
    output \REG.mem_38_13 ;
    input n4794;
    input n4793;
    output \REG.mem_38_11 ;
    output \REG.mem_29_11 ;
    output \REG.mem_28_11 ;
    input n4792;
    output \REG.mem_34_2 ;
    input n4791;
    input n4790;
    output \REG.mem_38_8 ;
    input n4789;
    input n4788;
    output \REG.mem_38_6 ;
    input n4787;
    input n4786;
    output \REG.mem_38_4 ;
    input n4785;
    output \REG.mem_38_3 ;
    input n4784;
    output \REG.mem_38_2 ;
    input n4783;
    output \REG.mem_38_1 ;
    input n4782;
    output \REG.mem_38_0 ;
    input n4781;
    output \REG.mem_37_15 ;
    input n4780;
    output \REG.mem_37_14 ;
    input n4779;
    output \REG.mem_37_13 ;
    input n4778;
    input n4777;
    output \REG.mem_37_11 ;
    input n4776;
    input n4775;
    input n4774;
    output \REG.mem_37_8 ;
    input n4773;
    input n4772;
    output \REG.mem_37_6 ;
    input n4771;
    input n4770;
    output \REG.mem_37_4 ;
    input n4769;
    output \REG.mem_37_3 ;
    input n4768;
    output \REG.mem_37_2 ;
    input n4767;
    output \REG.mem_37_1 ;
    input n4766;
    output \REG.mem_37_0 ;
    input n4156;
    output \REG.mem_26_6 ;
    output \REG.mem_25_6 ;
    output \REG.mem_24_6 ;
    output \REG.mem_34_9 ;
    input n4733;
    output \REG.mem_34_15 ;
    input n4732;
    output \REG.mem_34_14 ;
    input n4731;
    output \REG.mem_34_13 ;
    input n4730;
    input n4729;
    output \REG.mem_34_11 ;
    input n4728;
    input n4727;
    input n4726;
    output \REG.mem_34_8 ;
    input n4725;
    input n4155;
    output \REG.mem_2_1 ;
    input n4154;
    output \REG.mem_24_4 ;
    output \REG.mem_25_4 ;
    output \REG.mem_26_4 ;
    input n4724;
    output \REG.mem_34_6 ;
    output \REG.mem_30_4 ;
    output \REG.mem_28_4 ;
    output \REG.mem_29_4 ;
    input n4723;
    input n4722;
    output \REG.mem_34_4 ;
    input n4721;
    output \REG.mem_34_3 ;
    input n4720;
    input n4719;
    output \REG.mem_34_1 ;
    input n4718;
    output \REG.mem_8_4 ;
    output \REG.mem_9_4 ;
    output \REG.mem_10_4 ;
    output \REG.mem_11_4 ;
    output \REG.mem_14_4 ;
    output \REG.mem_15_4 ;
    output \REG.mem_12_4 ;
    output \REG.mem_13_4 ;
    output \REG.mem_6_1 ;
    output \REG.mem_7_1 ;
    output \REG.mem_5_1 ;
    input n4677;
    output [6:0]rp_sync1_r;
    output \REG.mem_26_10 ;
    output \REG.mem_18_1 ;
    output \REG.mem_19_1 ;
    input n4676;
    input n4675;
    input n4674;
    input n4673;
    input n4672;
    output \REG.mem_25_10 ;
    output \REG.mem_24_10 ;
    output \REG.mem_22_1 ;
    output \REG.mem_23_1 ;
    output \REG.mem_21_1 ;
    output n46;
    output n14;
    input n4655;
    input n4654;
    input n4653;
    input n4652;
    input n4651;
    input n4650;
    input n4649;
    input n4648;
    input n4647;
    output \REG.mem_30_13 ;
    input n4646;
    output \REG.mem_30_12 ;
    input n4645;
    output n37;
    output n5;
    input n4644;
    input n4643;
    input n4642;
    input n4641;
    input n4640;
    output \REG.mem_30_6 ;
    input n4639;
    input n4638;
    input n4637;
    input n4636;
    input n4635;
    output \REG.mem_30_1 ;
    input n4634;
    input n4633;
    input n4631;
    input n4629;
    output \REG.mem_18_14 ;
    output \REG.mem_19_14 ;
    input n4627;
    output n51;
    input n4626;
    input n4625;
    output \REG.mem_29_13 ;
    output \REG.mem_22_14 ;
    output \REG.mem_23_14 ;
    output \REG.mem_21_14 ;
    input n4624;
    output \REG.mem_29_12 ;
    input n4623;
    input n4622;
    input n4621;
    input n4620;
    input n4619;
    input n4618;
    output \REG.mem_29_6 ;
    input n4617;
    input n4616;
    input n4615;
    input n4614;
    input n4613;
    output \REG.mem_29_1 ;
    input n4612;
    input n4611;
    input n4610;
    input n4609;
    output \REG.mem_28_13 ;
    output n19;
    input n4608;
    output \REG.mem_28_12 ;
    input n4607;
    output \REG.mem_18_12 ;
    output \REG.mem_19_12 ;
    output \REG.mem_22_12 ;
    output \REG.mem_23_12 ;
    input n4606;
    input n4605;
    input n4604;
    input n4603;
    input n4602;
    output \REG.mem_28_6 ;
    input n4601;
    input n4600;
    input n4599;
    input n4598;
    input n4597;
    output \REG.mem_28_1 ;
    input n4596;
    output \REG.mem_21_12 ;
    input n4579;
    input n4578;
    input n4577;
    output \REG.mem_26_13 ;
    input n4576;
    output \REG.mem_26_12 ;
    input n4575;
    input n4574;
    input n4573;
    input n4572;
    input n4571;
    output \REG.mem_26_7 ;
    input n4570;
    input n4569;
    input n4568;
    input n4567;
    output \REG.mem_6_13 ;
    output \REG.mem_7_13 ;
    input n4566;
    input n4565;
    output \REG.mem_26_1 ;
    input n4564;
    output \REG.mem_26_0 ;
    input n4563;
    output [6:0]wp_sync1_r;
    input n4562;
    input n4561;
    input n4560;
    input n4559;
    input n4558;
    input n4557;
    input n4556;
    output \REG.mem_25_13 ;
    input n4555;
    output \REG.mem_25_12 ;
    input n4554;
    input n4553;
    input n4552;
    input n4551;
    output \REG.mem_5_13 ;
    input n4550;
    output \REG.mem_25_7 ;
    input n4549;
    input n4548;
    input n4547;
    input n4546;
    input n4545;
    input n4544;
    output \REG.mem_25_1 ;
    input n4543;
    output \REG.mem_25_0 ;
    input n4542;
    input n4541;
    input n4540;
    input n4539;
    input n4538;
    input n4537;
    input n4536;
    input n4535;
    input n4534;
    output \REG.mem_18_0 ;
    output \REG.mem_19_0 ;
    output \REG.mem_22_0 ;
    output \REG.mem_23_0 ;
    output \REG.mem_21_0 ;
    input DEBUG_9_c;
    input n4533;
    output \REG.mem_24_13 ;
    input n4532;
    output \REG.mem_24_12 ;
    input n4531;
    input n4530;
    input n4529;
    input n4528;
    input n4527;
    output \REG.mem_24_7 ;
    input n4526;
    input n4525;
    input n4524;
    input n4523;
    input n4522;
    input n4521;
    output \REG.mem_24_1 ;
    input n4520;
    output \REG.mem_24_0 ;
    input n4519;
    output \REG.mem_23_15 ;
    input n4518;
    input n4517;
    input n4516;
    input n4515;
    input n4514;
    output \REG.mem_23_10 ;
    input n4513;
    output \REG.mem_23_9 ;
    input n4512;
    input n4511;
    input n4510;
    input n4509;
    input n4508;
    output \REG.mem_23_4 ;
    input n4507;
    input n4506;
    input n4505;
    input n4504;
    input n4503;
    output \REG.mem_22_15 ;
    input n4502;
    input n4501;
    input n4500;
    input n4499;
    input n4498;
    output \REG.mem_22_10 ;
    input n4497;
    output \REG.mem_22_9 ;
    input n4496;
    input n4495;
    input n4494;
    input n4493;
    input n4492;
    output \REG.mem_22_4 ;
    input n4491;
    input n4490;
    input n4489;
    input n4488;
    input n4487;
    output \REG.mem_21_15 ;
    input n4486;
    input n4485;
    input n4484;
    input n4483;
    input n4482;
    output \REG.mem_21_10 ;
    input n4481;
    output \REG.mem_21_9 ;
    input n4480;
    input n4479;
    input n4478;
    input n4477;
    input n4476;
    output \REG.mem_21_4 ;
    input n4475;
    input n4474;
    input n4473;
    output \REG.mem_6_12 ;
    output \REG.mem_7_12 ;
    input n4472;
    output \REG.out_raw[15] ;
    output \REG.out_raw[14] ;
    output \REG.out_raw[13] ;
    output \REG.mem_5_12 ;
    output \REG.out_raw[12] ;
    output \REG.out_raw[11] ;
    output \REG.out_raw[10] ;
    input n4455;
    output \REG.mem_19_15 ;
    input n4454;
    input n4453;
    input n4452;
    input n4451;
    input n4450;
    input n4449;
    output \REG.mem_19_9 ;
    input n4448;
    input n4447;
    input n4446;
    input n4445;
    input n4444;
    output \REG.mem_19_4 ;
    input n4443;
    input n4442;
    input n4441;
    input n4440;
    output \REG.out_raw[9] ;
    output \REG.out_raw[8] ;
    input n4439;
    output \REG.mem_18_15 ;
    output \REG.out_raw[7] ;
    output \REG.out_raw[6] ;
    output \REG.out_raw[5] ;
    output \REG.out_raw[4] ;
    output \REG.out_raw[3] ;
    input n4438;
    output \REG.mem_6_9 ;
    output \REG.mem_7_9 ;
    output n54;
    output \REG.mem_5_9 ;
    input n4437;
    input n4436;
    input n4435;
    input n4434;
    input n4433;
    output \REG.mem_18_9 ;
    input n4432;
    input n4431;
    input n4430;
    input n4429;
    input n4428;
    output \REG.mem_18_4 ;
    input n4427;
    input n4426;
    input n4425;
    input n4424;
    output \REG.out_raw[2] ;
    output n22;
    output n39;
    output \REG.mem_10_9 ;
    output \REG.mem_11_9 ;
    output \REG.mem_10_13 ;
    output \REG.mem_11_13 ;
    output n7;
    output n40;
    output \REG.mem_9_9 ;
    output \REG.mem_8_9 ;
    output \REG.mem_9_13 ;
    output \REG.mem_8_13 ;
    output n8;
    output \REG.mem_14_12 ;
    output \REG.mem_15_12 ;
    input n4391;
    output \REG.out_raw[1] ;
    input n4390;
    output \REG.mem_13_12 ;
    output \REG.mem_12_12 ;
    input n4389;
    output \REG.mem_15_13 ;
    input n4388;
    input n4387;
    input n4386;
    output \REG.mem_15_10 ;
    input n4385;
    output \REG.mem_15_9 ;
    input n4384;
    output \REG.mem_15_8 ;
    input n4383;
    output \REG.mem_15_7 ;
    input n4382;
    input n4381;
    output \REG.mem_15_5 ;
    input n4380;
    input n4379;
    input n4378;
    input n4377;
    output \REG.mem_15_1 ;
    input n4376;
    input n4375;
    input n4374;
    output \REG.mem_6_8 ;
    output \REG.mem_7_8 ;
    output \REG.mem_5_8 ;
    output \REG.mem_14_9 ;
    output \REG.mem_13_9 ;
    output \REG.mem_12_9 ;
    output \REG.mem_6_5 ;
    output \REG.mem_7_5 ;
    input n4373;
    output \REG.mem_14_13 ;
    input n4372;
    input n4371;
    input n4370;
    output \REG.mem_14_10 ;
    input n4369;
    input n4368;
    output \REG.mem_14_8 ;
    input n4367;
    output \REG.mem_14_7 ;
    output \REG.mem_5_5 ;
    input n4366;
    input n4365;
    output \REG.mem_14_5 ;
    input n4364;
    input n4363;
    input n4362;
    input n4361;
    output \REG.mem_14_1 ;
    input n4360;
    input n4359;
    input n4358;
    input n4357;
    output \REG.mem_13_13 ;
    input n4356;
    input n4355;
    input n4354;
    output \REG.mem_13_10 ;
    input n4353;
    input n4352;
    output \REG.mem_13_8 ;
    input n4351;
    output \REG.mem_13_7 ;
    input n4350;
    input n4349;
    output \REG.mem_13_5 ;
    input n4348;
    input n4347;
    input n4346;
    input n4345;
    output \REG.mem_13_1 ;
    input n4344;
    input n4343;
    input n4342;
    input n4341;
    output \REG.mem_12_13 ;
    input n4340;
    input n4339;
    input n4338;
    output \REG.mem_12_10 ;
    input n4337;
    input n4336;
    output \REG.mem_12_8 ;
    input n4335;
    output \REG.mem_12_7 ;
    input n4334;
    input n4333;
    output \REG.mem_12_5 ;
    input n4332;
    input n4331;
    input n4330;
    input n4329;
    output \REG.mem_12_1 ;
    input n4328;
    input n4327;
    input n4326;
    input n4325;
    input n4324;
    input n4323;
    output n60;
    input n4322;
    output n28;
    output n41;
    output n9;
    input n4321;
    input n4320;
    output \REG.mem_11_8 ;
    input n4319;
    output \REG.mem_11_7 ;
    input n4318;
    input n4317;
    output \REG.mem_11_5 ;
    input n4316;
    input n4315;
    input n4314;
    input n4313;
    output \REG.mem_11_1 ;
    input n4312;
    input n4311;
    output n42;
    input n4310;
    input n4309;
    input n4308;
    output n10;
    input n4307;
    input n4306;
    input n4305;
    input n4304;
    output \REG.mem_10_8 ;
    input n4303;
    output \REG.mem_10_7 ;
    input n4302;
    input n4301;
    output \REG.mem_10_5 ;
    input n4300;
    input n4299;
    input n4298;
    input n4297;
    output \REG.mem_10_1 ;
    input n4296;
    input n4130;
    output n57;
    output \REG.mem_9_5 ;
    output \REG.mem_8_5 ;
    input n4288;
    input n4287;
    input n4286;
    input n4285;
    input n4284;
    input n4283;
    input n4282;
    input n4281;
    input n4280;
    output \REG.mem_9_8 ;
    input n4279;
    output \REG.mem_9_7 ;
    input n4278;
    input n4277;
    input n4108;
    output n25;
    input n4276;
    output n43;
    output n11;
    output n44;
    output n12;
    input n4275;
    input n4274;
    input n4273;
    output \REG.mem_9_1 ;
    input n4272;
    input n4270;
    input n4268;
    input n4107;
    output \REG.mem_8_7 ;
    input n4265;
    input n4264;
    input n4263;
    input n4262;
    input n4261;
    output n52;
    input n4260;
    output \REG.mem_8_8 ;
    input n4259;
    input n4258;
    input n4257;
    input n4256;
    input n4255;
    input n4254;
    input n4253;
    input n4252;
    input n4251;
    output \REG.mem_8_1 ;
    input n4250;
    input n4249;
    input n4248;
    input n4247;
    input n4246;
    input n4245;
    output \REG.mem_7_11 ;
    input n4244;
    input n4243;
    input n4242;
    input n4241;
    input n4240;
    input n4239;
    input n4238;
    output \REG.mem_7_4 ;
    input n4237;
    input n4236;
    input n4235;
    input n4234;
    input n4233;
    input n4232;
    input n4231;
    input n4230;
    input n4229;
    output \REG.mem_6_11 ;
    input n4228;
    input n4227;
    input n4226;
    input n4225;
    input n4224;
    input n4223;
    input n4222;
    output \REG.mem_6_4 ;
    input n4221;
    input n4220;
    input n4219;
    input n4218;
    input n4217;
    input n4216;
    input n4215;
    input n4214;
    input n4213;
    output \REG.mem_5_11 ;
    input n4212;
    input n4211;
    input n4210;
    input n4209;
    input n4208;
    input n4207;
    input n4206;
    output \REG.mem_5_4 ;
    input n4205;
    input n4204;
    input n4203;
    input n4202;
    input n4103;
    output n20;
    output n53;
    input n4101;
    output n21;
    output n35;
    output n3;
    output n36;
    output n55;
    output n23;
    output n4;
    output n47;
    output n15;
    output n31;
    output n63;
    
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    wire DEBUG_6_c /* synthesis SET_AS_NETWORK=DEBUG_6_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    fifo_dc_32_lut_gen_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 lscc_fifo_dc_inst (.FIFO_D6_c_6(FIFO_D6_c_6), 
            .\REG.mem_42_15 (\REG.mem_42_15 ), .\REG.mem_43_15 (\REG.mem_43_15 ), 
            .FIFO_D5_c_5(FIFO_D5_c_5), .\REG.mem_29_14 (\REG.mem_29_14 ), 
            .\REG.mem_28_14 (\REG.mem_28_14 ), .FIFO_CLK_c(FIFO_CLK_c), 
            .\REG.mem_41_15 (\REG.mem_41_15 ), .\REG.mem_40_15 (\REG.mem_40_15 ), 
            .GND_net(GND_net), .\REG.mem_2_0 (\REG.mem_2_0 ), .\REG.mem_2_2 (\REG.mem_2_2 ), 
            .FIFO_D4_c_4(FIFO_D4_c_4), .\REG.mem_18_5 (\REG.mem_18_5 ), 
            .\REG.mem_19_5 (\REG.mem_19_5 ), .FIFO_D3_c_3(FIFO_D3_c_3), 
            .\REG.mem_62_5 (\REG.mem_62_5 ), .\REG.mem_61_5 (\REG.mem_61_5 ), 
            .\REG.mem_60_5 (\REG.mem_60_5 ), .FIFO_D2_c_2(FIFO_D2_c_2), 
            .t_rd_fifo_en_w(t_rd_fifo_en_w), .\REG.out_raw[0] (\REG.out_raw[0] ), 
            .DEBUG_6_c(DEBUG_6_c), .\REG.mem_30_10 (\REG.mem_30_10 ), .\REG.mem_29_10 (\REG.mem_29_10 ), 
            .\REG.mem_28_10 (\REG.mem_28_10 ), .\REG.mem_58_8 (\REG.mem_58_8 ), 
            .\REG.mem_57_8 (\REG.mem_57_8 ), .\REG.mem_56_8 (\REG.mem_56_8 ), 
            .FIFO_D1_c_1(FIFO_D1_c_1), .\REG.mem_2_14 (\REG.mem_2_14 ), 
            .FIFO_D0_c_0(FIFO_D0_c_0), .\REG.mem_14_15 (\REG.mem_14_15 ), 
            .\REG.mem_15_15 (\REG.mem_15_15 ), .\REG.mem_13_15 (\REG.mem_13_15 ), 
            .\REG.mem_12_15 (\REG.mem_12_15 ), .\REG.mem_10_15 (\REG.mem_10_15 ), 
            .\REG.mem_11_15 (\REG.mem_11_15 ), .n56(n56), .\REG.mem_62_8 (\REG.mem_62_8 ), 
            .\REG.mem_61_8 (\REG.mem_61_8 ), .\REG.mem_60_8 (\REG.mem_60_8 ), 
            .\REG.mem_46_6 (\REG.mem_46_6 ), .\REG.mem_47_6 (\REG.mem_47_6 ), 
            .n24(n24), .write_to_dc32_fifo(write_to_dc32_fifo), .reset_all(reset_all), 
            .\wr_addr_nxt_c[1] (\wr_addr_nxt_c[1] ), .\REG.mem_45_6 (\REG.mem_45_6 ), 
            .\REG.mem_44_6 (\REG.mem_44_6 ), .dc32_fifo_is_full(dc32_fifo_is_full), 
            .\REG.mem_34_10 (\REG.mem_34_10 ), .\REG.mem_18_8 (\REG.mem_18_8 ), 
            .\REG.mem_19_8 (\REG.mem_19_8 ), .\REG.mem_58_11 (\REG.mem_58_11 ), 
            .\rd_grey_sync_r[0] (\rd_grey_sync_r[0] ), .\REG.mem_57_11 (\REG.mem_57_11 ), 
            .\REG.mem_56_11 (\REG.mem_56_11 ), .\REG.mem_6_14 (\REG.mem_6_14 ), 
            .\REG.mem_7_14 (\REG.mem_7_14 ), .\REG.mem_5_14 (\REG.mem_5_14 ), 
            .\REG.mem_10_12 (\REG.mem_10_12 ), .\REG.mem_11_12 (\REG.mem_11_12 ), 
            .\REG.mem_9_12 (\REG.mem_9_12 ), .\REG.mem_8_12 (\REG.mem_8_12 ), 
            .\REG.mem_6_10 (\REG.mem_6_10 ), .\REG.mem_7_10 (\REG.mem_7_10 ), 
            .\REG.mem_26_9 (\REG.mem_26_9 ), .DEBUG_1_c(DEBUG_1_c), .\REG.mem_6_0 (\REG.mem_6_0 ), 
            .\REG.mem_7_0 (\REG.mem_7_0 ), .\REG.mem_5_0 (\REG.mem_5_0 ), 
            .\REG.mem_5_10 (\REG.mem_5_10 ), .\REG.mem_25_9 (\REG.mem_25_9 ), 
            .\REG.mem_24_9 (\REG.mem_24_9 ), .\REG.mem_56_7 (\REG.mem_56_7 ), 
            .\REG.mem_57_7 (\REG.mem_57_7 ), .\REG.mem_58_7 (\REG.mem_58_7 ), 
            .\num_words_in_buffer[3] (\num_words_in_buffer[3] ), .\wr_grey_sync_r[0] (\wr_grey_sync_r[0] ), 
            .\REG.mem_10_14 (\REG.mem_10_14 ), .\REG.mem_11_14 (\REG.mem_11_14 ), 
            .\REG.mem_9_14 (\REG.mem_9_14 ), .\REG.mem_8_14 (\REG.mem_8_14 ), 
            .\REG.mem_14_14 (\REG.mem_14_14 ), .\REG.mem_15_14 (\REG.mem_15_14 ), 
            .\REG.mem_13_14 (\REG.mem_13_14 ), .\REG.mem_12_14 (\REG.mem_12_14 ), 
            .\REG.mem_38_9 (\REG.mem_38_9 ), .\REG.mem_39_9 (\REG.mem_39_9 ), 
            .\REG.mem_37_9 (\REG.mem_37_9 ), .\REG.mem_34_7 (\REG.mem_34_7 ), 
            .\REG.mem_42_9 (\REG.mem_42_9 ), .\REG.mem_43_9 (\REG.mem_43_9 ), 
            .\REG.mem_10_10 (\REG.mem_10_10 ), .\REG.mem_11_10 (\REG.mem_11_10 ), 
            .\REG.mem_9_10 (\REG.mem_9_10 ), .\REG.mem_8_10 (\REG.mem_8_10 ), 
            .\REG.mem_41_9 (\REG.mem_41_9 ), .\REG.mem_40_9 (\REG.mem_40_9 ), 
            .\REG.mem_9_15 (\REG.mem_9_15 ), .\REG.mem_8_15 (\REG.mem_8_15 ), 
            .\REG.mem_18_6 (\REG.mem_18_6 ), .\REG.mem_19_6 (\REG.mem_19_6 ), 
            .\wr_addr_nxt_c[3] (\wr_addr_nxt_c[3] ), .FIFO_D15_c_15(FIFO_D15_c_15), 
            .\REG.mem_22_5 (\REG.mem_22_5 ), .\REG.mem_23_5 (\REG.mem_23_5 ), 
            .\REG.mem_21_5 (\REG.mem_21_5 ), .\REG.mem_38_10 (\REG.mem_38_10 ), 
            .\REG.mem_39_10 (\REG.mem_39_10 ), .\REG.mem_37_10 (\REG.mem_37_10 ), 
            .\REG.mem_18_10 (\REG.mem_18_10 ), .\REG.mem_19_10 (\REG.mem_19_10 ), 
            .FIFO_D14_c_14(FIFO_D14_c_14), .\REG.mem_34_12 (\REG.mem_34_12 ), 
            .\REG.mem_22_6 (\REG.mem_22_6 ), .\REG.mem_23_6 (\REG.mem_23_6 ), 
            .\REG.mem_26_14 (\REG.mem_26_14 ), .\REG.mem_25_14 (\REG.mem_25_14 ), 
            .\REG.mem_24_14 (\REG.mem_24_14 ), .\REG.mem_18_13 (\REG.mem_18_13 ), 
            .\REG.mem_19_13 (\REG.mem_19_13 ), .\REG.mem_62_7 (\REG.mem_62_7 ), 
            .\REG.mem_21_6 (\REG.mem_21_6 ), .\REG.mem_60_7 (\REG.mem_60_7 ), 
            .\REG.mem_61_7 (\REG.mem_61_7 ), .\REG.mem_30_14 (\REG.mem_30_14 ), 
            .\REG.mem_50_3 (\REG.mem_50_3 ), .\REG.mem_51_3 (\REG.mem_51_3 ), 
            .\REG.mem_38_12 (\REG.mem_38_12 ), .\REG.mem_39_12 (\REG.mem_39_12 ), 
            .\REG.mem_37_12 (\REG.mem_37_12 ), .\REG.mem_46_8 (\REG.mem_46_8 ), 
            .\REG.mem_47_8 (\REG.mem_47_8 ), .\REG.mem_45_8 (\REG.mem_45_8 ), 
            .\REG.mem_44_8 (\REG.mem_44_8 ), .\REG.mem_58_10 (\REG.mem_58_10 ), 
            .\REG.mem_2_3 (\REG.mem_2_3 ), .\REG.mem_57_10 (\REG.mem_57_10 ), 
            .\REG.mem_56_10 (\REG.mem_56_10 ), .\REG.mem_62_2 (\REG.mem_62_2 ), 
            .\REG.mem_61_2 (\REG.mem_61_2 ), .\REG.mem_60_2 (\REG.mem_60_2 ), 
            .\REG.mem_58_15 (\REG.mem_58_15 ), .\REG.mem_10_0 (\REG.mem_10_0 ), 
            .\REG.mem_11_0 (\REG.mem_11_0 ), .\REG.mem_9_0 (\REG.mem_9_0 ), 
            .\REG.mem_8_0 (\REG.mem_8_0 ), .\REG.mem_57_15 (\REG.mem_57_15 ), 
            .\REG.mem_56_15 (\REG.mem_56_15 ), .\REG.mem_30_0 (\REG.mem_30_0 ), 
            .\REG.mem_29_0 (\REG.mem_29_0 ), .\REG.mem_28_0 (\REG.mem_28_0 ), 
            .\REG.mem_38_7 (\REG.mem_38_7 ), .\REG.mem_39_7 (\REG.mem_39_7 ), 
            .FIFO_D13_c_13(FIFO_D13_c_13), .\REG.mem_37_7 (\REG.mem_37_7 ), 
            .n58(n58), .FIFO_D12_c_12(FIFO_D12_c_12), .\REG.mem_26_5 (\REG.mem_26_5 ), 
            .\REG.mem_25_5 (\REG.mem_25_5 ), .\REG.mem_24_5 (\REG.mem_24_5 ), 
            .n50(n50), .\REG.mem_46_0 (\REG.mem_46_0 ), .\REG.mem_47_0 (\REG.mem_47_0 ), 
            .\REG.mem_6_3 (\REG.mem_6_3 ), .\REG.mem_7_3 (\REG.mem_7_3 ), 
            .\REG.mem_5_3 (\REG.mem_5_3 ), .\REG.mem_45_0 (\REG.mem_45_0 ), 
            .\REG.mem_44_0 (\REG.mem_44_0 ), .\REG.mem_50_8 (\REG.mem_50_8 ), 
            .\REG.mem_51_8 (\REG.mem_51_8 ), .n18(n18), .\REG.mem_10_3 (\REG.mem_10_3 ), 
            .\REG.mem_11_3 (\REG.mem_11_3 ), .\REG.mem_6_2 (\REG.mem_6_2 ), 
            .\REG.mem_7_2 (\REG.mem_7_2 ), .\REG.mem_5_2 (\REG.mem_5_2 ), 
            .\REG.mem_9_3 (\REG.mem_9_3 ), .\REG.mem_8_3 (\REG.mem_8_3 ), 
            .\wr_addr_nxt_c[5] (\wr_addr_nxt_c[5] ), .\REG.mem_42_12 (\REG.mem_42_12 ), 
            .\REG.mem_43_12 (\REG.mem_43_12 ), .\REG.mem_41_12 (\REG.mem_41_12 ), 
            .\REG.mem_40_12 (\REG.mem_40_12 ), .\REG.mem_10_2 (\REG.mem_10_2 ), 
            .\REG.mem_11_2 (\REG.mem_11_2 ), .n4169(n4169), .\REG.mem_2_15 (\REG.mem_2_15 ), 
            .\REG.mem_9_2 (\REG.mem_9_2 ), .\REG.mem_8_2 (\REG.mem_8_2 ), 
            .n4168(n4168), .n4167(n4167), .\REG.mem_2_13 (\REG.mem_2_13 ), 
            .n4166(n4166), .\REG.mem_2_12 (\REG.mem_2_12 ), .n4165(n4165), 
            .\REG.mem_2_11 (\REG.mem_2_11 ), .n4164(n4164), .\REG.mem_2_10 (\REG.mem_2_10 ), 
            .\REG.mem_6_6 (\REG.mem_6_6 ), .\REG.mem_7_6 (\REG.mem_7_6 ), 
            .n4163(n4163), .\REG.mem_2_9 (\REG.mem_2_9 ), .\REG.mem_5_6 (\REG.mem_5_6 ), 
            .\REG.mem_30_3 (\REG.mem_30_3 ), .\REG.mem_29_3 (\REG.mem_29_3 ), 
            .\REG.mem_28_3 (\REG.mem_28_3 ), .\REG.mem_22_13 (\REG.mem_22_13 ), 
            .\REG.mem_23_13 (\REG.mem_23_13 ), .\REG.mem_21_13 (\REG.mem_21_13 ), 
            .\REG.mem_54_3 (\REG.mem_54_3 ), .\REG.mem_55_3 (\REG.mem_55_3 ), 
            .\REG.mem_53_3 (\REG.mem_53_3 ), .\REG.mem_42_10 (\REG.mem_42_10 ), 
            .\REG.mem_43_10 (\REG.mem_43_10 ), .\REG.mem_41_10 (\REG.mem_41_10 ), 
            .\REG.mem_40_10 (\REG.mem_40_10 ), .\REG.mem_56_4 (\REG.mem_56_4 ), 
            .\REG.mem_57_4 (\REG.mem_57_4 ), .\REG.mem_6_15 (\REG.mem_6_15 ), 
            .\REG.mem_7_15 (\REG.mem_7_15 ), .\REG.mem_58_4 (\REG.mem_58_4 ), 
            .\REG.mem_26_15 (\REG.mem_26_15 ), .\REG.mem_5_15 (\REG.mem_5_15 ), 
            .\REG.mem_25_15 (\REG.mem_25_15 ), .\REG.mem_24_15 (\REG.mem_24_15 ), 
            .\REG.mem_58_3 (\REG.mem_58_3 ), .\REG.mem_57_3 (\REG.mem_57_3 ), 
            .\REG.mem_56_3 (\REG.mem_56_3 ), .\REG.mem_62_3 (\REG.mem_62_3 ), 
            .\REG.mem_62_4 (\REG.mem_62_4 ), .\REG.mem_60_4 (\REG.mem_60_4 ), 
            .\REG.mem_61_4 (\REG.mem_61_4 ), .\REG.mem_61_3 (\REG.mem_61_3 ), 
            .\REG.mem_60_3 (\REG.mem_60_3 ), .\rd_addr_r[6] (\rd_addr_r[6] ), 
            .\rd_addr_nxt_c_6__N_176[5] (\rd_addr_nxt_c_6__N_176[5] ), .\REG.mem_22_8 (\REG.mem_22_8 ), 
            .\REG.mem_23_8 (\REG.mem_23_8 ), .\rd_addr_nxt_c_6__N_176[3] (\rd_addr_nxt_c_6__N_176[3] ), 
            .\REG.mem_21_8 (\REG.mem_21_8 ), .\REG.mem_54_8 (\REG.mem_54_8 ), 
            .\REG.mem_55_8 (\REG.mem_55_8 ), .FIFO_D11_c_11(FIFO_D11_c_11), 
            .\REG.mem_14_3 (\REG.mem_14_3 ), .\REG.mem_15_3 (\REG.mem_15_3 ), 
            .\REG.mem_53_8 (\REG.mem_53_8 ), .\REG.mem_14_2 (\REG.mem_14_2 ), 
            .\REG.mem_15_2 (\REG.mem_15_2 ), .\REG.mem_13_3 (\REG.mem_13_3 ), 
            .\REG.mem_12_3 (\REG.mem_12_3 ), .\REG.mem_13_2 (\REG.mem_13_2 ), 
            .\REG.mem_12_2 (\REG.mem_12_2 ), .\REG.mem_30_5 (\REG.mem_30_5 ), 
            .\REG.mem_58_13 (\REG.mem_58_13 ), .\REG.mem_29_5 (\REG.mem_29_5 ), 
            .\REG.mem_28_5 (\REG.mem_28_5 ), .\REG.mem_34_5 (\REG.mem_34_5 ), 
            .\REG.mem_57_13 (\REG.mem_57_13 ), .\REG.mem_56_13 (\REG.mem_56_13 ), 
            .\REG.mem_14_6 (\REG.mem_14_6 ), .\REG.mem_15_6 (\REG.mem_15_6 ), 
            .\REG.mem_13_6 (\REG.mem_13_6 ), .\REG.mem_12_6 (\REG.mem_12_6 ), 
            .\REG.mem_54_9 (\REG.mem_54_9 ), .\REG.mem_55_9 (\REG.mem_55_9 ), 
            .\REG.mem_53_9 (\REG.mem_53_9 ), .\REG.mem_34_0 (\REG.mem_34_0 ), 
            .\REG.mem_14_0 (\REG.mem_14_0 ), .\REG.mem_15_0 (\REG.mem_15_0 ), 
            .\REG.mem_13_0 (\REG.mem_13_0 ), .\REG.mem_12_0 (\REG.mem_12_0 ), 
            .FIFO_D10_c_10(FIFO_D10_c_10), .\REG.mem_42_14 (\REG.mem_42_14 ), 
            .\REG.mem_43_14 (\REG.mem_43_14 ), .\REG.mem_41_14 (\REG.mem_41_14 ), 
            .\REG.mem_40_14 (\REG.mem_40_14 ), .n4162(n4162), .\REG.mem_2_8 (\REG.mem_2_8 ), 
            .n4161(n4161), .\REG.mem_2_7 (\REG.mem_2_7 ), .FIFO_D9_c_9(FIFO_D9_c_9), 
            .n5327(n5327), .VCC_net(VCC_net), .\fifo_data_out[0] (\fifo_data_out[0] ), 
            .\REG.mem_10_11 (\REG.mem_10_11 ), .\REG.mem_11_11 (\REG.mem_11_11 ), 
            .FIFO_D8_c_8(FIFO_D8_c_8), .FIFO_D7_c_7(FIFO_D7_c_7), .\REG.mem_9_11 (\REG.mem_9_11 ), 
            .\REG.mem_8_11 (\REG.mem_8_11 ), .\REG.mem_62_15 (\REG.mem_62_15 ), 
            .\REG.mem_62_10 (\REG.mem_62_10 ), .n5305(n5305), .\fifo_data_out[15] (\fifo_data_out[15] ), 
            .\REG.mem_46_12 (\REG.mem_46_12 ), .\REG.mem_47_12 (\REG.mem_47_12 ), 
            .n5302(n5302), .\fifo_data_out[14] (\fifo_data_out[14] ), .\REG.mem_61_10 (\REG.mem_61_10 ), 
            .\REG.mem_60_10 (\REG.mem_60_10 ), .\REG.mem_61_15 (\REG.mem_61_15 ), 
            .\REG.mem_60_15 (\REG.mem_60_15 ), .n5299(n5299), .\fifo_data_out[13] (\fifo_data_out[13] ), 
            .n5296(n5296), .\fifo_data_out[12] (\fifo_data_out[12] ), .n5293(n5293), 
            .\fifo_data_out[11] (\fifo_data_out[11] ), .n5290(n5290), .\fifo_data_out[10] (\fifo_data_out[10] ), 
            .\REG.mem_45_12 (\REG.mem_45_12 ), .\REG.mem_44_12 (\REG.mem_44_12 ), 
            .\REG.mem_46_15 (\REG.mem_46_15 ), .\REG.mem_47_15 (\REG.mem_47_15 ), 
            .\REG.mem_18_3 (\REG.mem_18_3 ), .\REG.mem_19_3 (\REG.mem_19_3 ), 
            .n5255(n5255), .\fifo_data_out[9] (\fifo_data_out[9] ), .n5252(n5252), 
            .\fifo_data_out[8] (\fifo_data_out[8] ), .n5249(n5249), .\fifo_data_out[7] (\fifo_data_out[7] ), 
            .\REG.mem_45_15 (\REG.mem_45_15 ), .\REG.mem_44_15 (\REG.mem_44_15 ), 
            .n4160(n4160), .\REG.mem_2_6 (\REG.mem_2_6 ), .\REG.mem_14_11 (\REG.mem_14_11 ), 
            .\REG.mem_15_11 (\REG.mem_15_11 ), .n4159(n4159), .\REG.mem_2_5 (\REG.mem_2_5 ), 
            .n5236(n5236), .\fifo_data_out[6] (\fifo_data_out[6] ), .n5233(n5233), 
            .\fifo_data_out[5] (\fifo_data_out[5] ), .\REG.mem_13_11 (\REG.mem_13_11 ), 
            .\REG.mem_12_11 (\REG.mem_12_11 ), .n5230(n5230), .\fifo_data_out[4] (\fifo_data_out[4] ), 
            .\wr_grey_sync_r[5] (\wr_grey_sync_r[5] ), .\wr_grey_sync_r[4] (\wr_grey_sync_r[4] ), 
            .\wr_grey_sync_r[3] (\wr_grey_sync_r[3] ), .n5212(n5212), .\fifo_data_out[3] (\fifo_data_out[3] ), 
            .\REG.mem_18_2 (\REG.mem_18_2 ), .\REG.mem_19_2 (\REG.mem_19_2 ), 
            .n5208(n5208), .n5207(n5207), .\REG.mem_62_14 (\REG.mem_62_14 ), 
            .n5206(n5206), .\REG.mem_62_13 (\REG.mem_62_13 ), .n5205(n5205), 
            .\REG.mem_62_12 (\REG.mem_62_12 ), .n5204(n5204), .\REG.mem_62_11 (\REG.mem_62_11 ), 
            .n5203(n5203), .n5202(n5202), .\REG.mem_62_9 (\REG.mem_62_9 ), 
            .n5201(n5201), .n5200(n5200), .\wr_grey_sync_r[2] (\wr_grey_sync_r[2] ), 
            .\wr_grey_sync_r[1] (\wr_grey_sync_r[1] ), .n5199(n5199), .\REG.mem_62_6 (\REG.mem_62_6 ), 
            .n5198(n5198), .n5197(n5197), .n5196(n5196), .n5195(n5195), 
            .n5194(n5194), .\REG.mem_62_1 (\REG.mem_62_1 ), .n5193(n5193), 
            .\REG.mem_62_0 (\REG.mem_62_0 ), .n5192(n5192), .n5191(n5191), 
            .\REG.mem_61_14 (\REG.mem_61_14 ), .n5190(n5190), .\REG.mem_61_13 (\REG.mem_61_13 ), 
            .n5189(n5189), .\REG.mem_61_12 (\REG.mem_61_12 ), .n5188(n5188), 
            .\REG.mem_61_11 (\REG.mem_61_11 ), .n5187(n5187), .n5186(n5186), 
            .\REG.mem_61_9 (\REG.mem_61_9 ), .n5185(n5185), .n5184(n5184), 
            .n5183(n5183), .\REG.mem_61_6 (\REG.mem_61_6 ), .\REG.mem_22_3 (\REG.mem_22_3 ), 
            .\REG.mem_23_3 (\REG.mem_23_3 ), .\REG.mem_26_8 (\REG.mem_26_8 ), 
            .n5182(n5182), .\REG.mem_21_3 (\REG.mem_21_3 ), .n5181(n5181), 
            .n5180(n5180), .n5179(n5179), .n5178(n5178), .\REG.mem_61_1 (\REG.mem_61_1 ), 
            .n5177(n5177), .\REG.mem_61_0 (\REG.mem_61_0 ), .n5176(n5176), 
            .n5175(n5175), .\REG.mem_60_14 (\REG.mem_60_14 ), .n5174(n5174), 
            .\REG.mem_60_13 (\REG.mem_60_13 ), .n5173(n5173), .\REG.mem_60_12 (\REG.mem_60_12 ), 
            .n5172(n5172), .\REG.mem_60_11 (\REG.mem_60_11 ), .n5171(n5171), 
            .n5170(n5170), .\REG.mem_60_9 (\REG.mem_60_9 ), .n5169(n5169), 
            .n5168(n5168), .n5167(n5167), .\REG.mem_60_6 (\REG.mem_60_6 ), 
            .\REG.mem_25_8 (\REG.mem_25_8 ), .\REG.mem_24_8 (\REG.mem_24_8 ), 
            .\REG.mem_46_9 (\REG.mem_46_9 ), .\REG.mem_47_9 (\REG.mem_47_9 ), 
            .\REG.mem_45_9 (\REG.mem_45_9 ), .\REG.mem_44_9 (\REG.mem_44_9 ), 
            .\REG.mem_30_7 (\REG.mem_30_7 ), .n5166(n5166), .n5165(n5165), 
            .n5164(n5164), .n5163(n5163), .n5162(n5162), .\REG.mem_60_1 (\REG.mem_60_1 ), 
            .n5161(n5161), .\REG.mem_60_0 (\REG.mem_60_0 ), .\REG.mem_29_7 (\REG.mem_29_7 ), 
            .\REG.mem_28_7 (\REG.mem_28_7 ), .n5144(n5144), .n5143(n5143), 
            .\REG.mem_58_14 (\REG.mem_58_14 ), .n5142(n5142), .n5141(n5141), 
            .\REG.mem_58_12 (\REG.mem_58_12 ), .n5140(n5140), .n5139(n5139), 
            .n5138(n5138), .\REG.mem_58_9 (\REG.mem_58_9 ), .n5137(n5137), 
            .n5136(n5136), .n5135(n5135), .\REG.mem_58_6 (\REG.mem_58_6 ), 
            .\REG.mem_46_10 (\REG.mem_46_10 ), .\REG.mem_47_10 (\REG.mem_47_10 ), 
            .\REG.mem_45_10 (\REG.mem_45_10 ), .\REG.mem_44_10 (\REG.mem_44_10 ), 
            .n5134(n5134), .\REG.mem_58_5 (\REG.mem_58_5 ), .\REG.mem_30_9 (\REG.mem_30_9 ), 
            .n5133(n5133), .n5132(n5132), .n5131(n5131), .\REG.mem_58_2 (\REG.mem_58_2 ), 
            .n5130(n5130), .\REG.mem_58_1 (\REG.mem_58_1 ), .n5129(n5129), 
            .\REG.mem_58_0 (\REG.mem_58_0 ), .n5128(n5128), .n5127(n5127), 
            .\REG.mem_57_14 (\REG.mem_57_14 ), .n5126(n5126), .n5125(n5125), 
            .\REG.mem_57_12 (\REG.mem_57_12 ), .n5124(n5124), .n5123(n5123), 
            .n5122(n5122), .\REG.mem_57_9 (\REG.mem_57_9 ), .n5121(n5121), 
            .n5120(n5120), .n5119(n5119), .\REG.mem_57_6 (\REG.mem_57_6 ), 
            .\REG.mem_29_9 (\REG.mem_29_9 ), .\REG.mem_28_9 (\REG.mem_28_9 ), 
            .n5118(n5118), .\REG.mem_57_5 (\REG.mem_57_5 ), .n5117(n5117), 
            .n5116(n5116), .n5115(n5115), .\REG.mem_57_2 (\REG.mem_57_2 ), 
            .n5114(n5114), .\REG.mem_57_1 (\REG.mem_57_1 ), .n5113(n5113), 
            .\fifo_data_out[2] (\fifo_data_out[2] ), .n5110(n5110), .\REG.mem_57_0 (\REG.mem_57_0 ), 
            .n5109(n5109), .n5108(n5108), .\REG.mem_56_14 (\REG.mem_56_14 ), 
            .n5107(n5107), .n5106(n5106), .\REG.mem_56_12 (\REG.mem_56_12 ), 
            .n5105(n5105), .n5104(n5104), .n5103(n5103), .\REG.mem_56_9 (\REG.mem_56_9 ), 
            .\REG.mem_10_6 (\REG.mem_10_6 ), .\REG.mem_11_6 (\REG.mem_11_6 ), 
            .n5102(n5102), .\REG.mem_9_6 (\REG.mem_9_6 ), .\REG.mem_8_6 (\REG.mem_8_6 ), 
            .n5101(n5101), .n5100(n5100), .\REG.mem_56_6 (\REG.mem_56_6 ), 
            .n5099(n5099), .\REG.mem_56_5 (\REG.mem_56_5 ), .n5098(n5098), 
            .n5097(n5097), .n5096(n5096), .\REG.mem_56_2 (\REG.mem_56_2 ), 
            .n5095(n5095), .\REG.mem_56_1 (\REG.mem_56_1 ), .n5094(n5094), 
            .\fifo_data_out[1] (\fifo_data_out[1] ), .n5091(n5091), .\REG.mem_56_0 (\REG.mem_56_0 ), 
            .n5090(n5090), .\REG.mem_55_15 (\REG.mem_55_15 ), .n5089(n5089), 
            .\REG.mem_55_14 (\REG.mem_55_14 ), .n5088(n5088), .\REG.mem_55_13 (\REG.mem_55_13 ), 
            .n5087(n5087), .\REG.mem_55_12 (\REG.mem_55_12 ), .\REG.mem_22_2 (\REG.mem_22_2 ), 
            .\REG.mem_23_2 (\REG.mem_23_2 ), .\REG.mem_21_2 (\REG.mem_21_2 ), 
            .n5086(n5086), .\REG.mem_55_11 (\REG.mem_55_11 ), .n5085(n5085), 
            .\REG.mem_55_10 (\REG.mem_55_10 ), .n5084(n5084), .n5083(n5083), 
            .n5082(n5082), .\REG.mem_55_7 (\REG.mem_55_7 ), .n5081(n5081), 
            .\REG.mem_55_6 (\REG.mem_55_6 ), .n5080(n5080), .\REG.mem_55_5 (\REG.mem_55_5 ), 
            .n5079(n5079), .\REG.mem_55_4 (\REG.mem_55_4 ), .n5078(n5078), 
            .n5077(n5077), .\REG.mem_55_2 (\REG.mem_55_2 ), .n5076(n5076), 
            .\REG.mem_55_1 (\REG.mem_55_1 ), .n5075(n5075), .\REG.mem_55_0 (\REG.mem_55_0 ), 
            .n5074(n5074), .\REG.mem_54_15 (\REG.mem_54_15 ), .n5073(n5073), 
            .\REG.mem_54_14 (\REG.mem_54_14 ), .n5072(n5072), .\REG.mem_54_13 (\REG.mem_54_13 ), 
            .\num_words_in_buffer[6] (\num_words_in_buffer[6] ), .\num_words_in_buffer[5] (\num_words_in_buffer[5] ), 
            .\num_words_in_buffer[4] (\num_words_in_buffer[4] ), .n5071(n5071), 
            .\REG.mem_54_12 (\REG.mem_54_12 ), .n5070(n5070), .\REG.mem_54_11 (\REG.mem_54_11 ), 
            .n5069(n5069), .\REG.mem_54_10 (\REG.mem_54_10 ), .n5068(n5068), 
            .n5067(n5067), .n5066(n5066), .\REG.mem_54_7 (\REG.mem_54_7 ), 
            .n5065(n5065), .\REG.mem_54_6 (\REG.mem_54_6 ), .n5064(n5064), 
            .\REG.mem_54_5 (\REG.mem_54_5 ), .n5063(n5063), .\REG.mem_54_4 (\REG.mem_54_4 ), 
            .n5062(n5062), .n5061(n5061), .\REG.mem_54_2 (\REG.mem_54_2 ), 
            .n5060(n5060), .\REG.mem_54_1 (\REG.mem_54_1 ), .n5057(n5057), 
            .\REG.mem_54_0 (\REG.mem_54_0 ), .n5056(n5056), .\REG.mem_53_15 (\REG.mem_53_15 ), 
            .n5055(n5055), .\REG.mem_53_14 (\REG.mem_53_14 ), .\REG.mem_50_12 (\REG.mem_50_12 ), 
            .\REG.mem_51_12 (\REG.mem_51_12 ), .\REG.mem_38_5 (\REG.mem_38_5 ), 
            .\REG.mem_39_5 (\REG.mem_39_5 ), .\REG.mem_37_5 (\REG.mem_37_5 ), 
            .n5054(n5054), .\REG.mem_53_13 (\REG.mem_53_13 ), .n5053(n5053), 
            .\REG.mem_53_12 (\REG.mem_53_12 ), .n5052(n5052), .\REG.mem_53_11 (\REG.mem_53_11 ), 
            .n5051(n5051), .\REG.mem_53_10 (\REG.mem_53_10 ), .n5050(n5050), 
            .n5049(n5049), .n5048(n5048), .\REG.mem_53_7 (\REG.mem_53_7 ), 
            .n5047(n5047), .\REG.mem_53_6 (\REG.mem_53_6 ), .n5046(n5046), 
            .\REG.mem_53_5 (\REG.mem_53_5 ), .n5045(n5045), .\REG.mem_53_4 (\REG.mem_53_4 ), 
            .n5044(n5044), .n5043(n5043), .\REG.mem_53_2 (\REG.mem_53_2 ), 
            .n5042(n5042), .\REG.mem_53_1 (\REG.mem_53_1 ), .n5041(n5041), 
            .\REG.mem_53_0 (\REG.mem_53_0 ), .\REG.mem_26_2 (\REG.mem_26_2 ), 
            .\REG.mem_18_11 (\REG.mem_18_11 ), .\REG.mem_19_11 (\REG.mem_19_11 ), 
            .\REG.mem_25_2 (\REG.mem_25_2 ), .\REG.mem_24_2 (\REG.mem_24_2 ), 
            .n5024(n5024), .\REG.mem_51_15 (\REG.mem_51_15 ), .n5023(n5023), 
            .\REG.mem_51_14 (\REG.mem_51_14 ), .n26(n26), .\REG.mem_26_3 (\REG.mem_26_3 ), 
            .\REG.mem_25_3 (\REG.mem_25_3 ), .\REG.mem_24_3 (\REG.mem_24_3 ), 
            .\REG.mem_40_4 (\REG.mem_40_4 ), .\REG.mem_41_4 (\REG.mem_41_4 ), 
            .n5022(n5022), .\REG.mem_51_13 (\REG.mem_51_13 ), .n5021(n5021), 
            .n5020(n5020), .\REG.mem_51_11 (\REG.mem_51_11 ), .n5019(n5019), 
            .\REG.mem_51_10 (\REG.mem_51_10 ), .n5018(n5018), .\REG.mem_51_9 (\REG.mem_51_9 ), 
            .n5017(n5017), .n5016(n5016), .\REG.mem_51_7 (\REG.mem_51_7 ), 
            .n5015(n5015), .\REG.mem_51_6 (\REG.mem_51_6 ), .n5014(n5014), 
            .\REG.mem_51_5 (\REG.mem_51_5 ), .n5013(n5013), .\REG.mem_51_4 (\REG.mem_51_4 ), 
            .n5012(n5012), .n5011(n5011), .\REG.mem_51_2 (\REG.mem_51_2 ), 
            .n5010(n5010), .\REG.mem_51_1 (\REG.mem_51_1 ), .n5008(n5008), 
            .\REG.mem_51_0 (\REG.mem_51_0 ), .\REG.mem_42_4 (\REG.mem_42_4 ), 
            .\REG.mem_43_4 (\REG.mem_43_4 ), .\REG.mem_22_11 (\REG.mem_22_11 ), 
            .\REG.mem_23_11 (\REG.mem_23_11 ), .n5007(n5007), .\REG.mem_50_15 (\REG.mem_50_15 ), 
            .n5006(n5006), .\REG.mem_50_14 (\REG.mem_50_14 ), .n5005(n5005), 
            .\REG.mem_50_13 (\REG.mem_50_13 ), .n5004(n5004), .n5003(n5003), 
            .\REG.mem_50_11 (\REG.mem_50_11 ), .n5002(n5002), .\REG.mem_50_10 (\REG.mem_50_10 ), 
            .n5001(n5001), .\REG.mem_50_9 (\REG.mem_50_9 ), .n5000(n5000), 
            .n4999(n4999), .\REG.mem_50_7 (\REG.mem_50_7 ), .n4998(n4998), 
            .\REG.mem_50_6 (\REG.mem_50_6 ), .n4997(n4997), .\REG.mem_50_5 (\REG.mem_50_5 ), 
            .n4996(n4996), .\REG.mem_50_4 (\REG.mem_50_4 ), .n4995(n4995), 
            .n4994(n4994), .\REG.mem_50_2 (\REG.mem_50_2 ), .n4993(n4993), 
            .\REG.mem_50_1 (\REG.mem_50_1 ), .n4992(n4992), .\REG.mem_50_0 (\REG.mem_50_0 ), 
            .\REG.mem_21_11 (\REG.mem_21_11 ), .\rd_addr_nxt_c_6__N_176[1] (\rd_addr_nxt_c_6__N_176[1] ), 
            .n4158(n4158), .\REG.mem_2_4 (\REG.mem_2_4 ), .\REG.mem_30_15 (\REG.mem_30_15 ), 
            .\REG.mem_29_15 (\REG.mem_29_15 ), .\REG.mem_28_15 (\REG.mem_28_15 ), 
            .\REG.mem_30_8 (\REG.mem_30_8 ), .\REG.mem_29_8 (\REG.mem_29_8 ), 
            .\REG.mem_28_8 (\REG.mem_28_8 ), .\REG.mem_46_4 (\REG.mem_46_4 ), 
            .\REG.mem_47_4 (\REG.mem_47_4 ), .n4946(n4946), .n4945(n4945), 
            .\REG.mem_47_14 (\REG.mem_47_14 ), .n4944(n4944), .\REG.mem_47_13 (\REG.mem_47_13 ), 
            .\rd_grey_sync_r[5] (\rd_grey_sync_r[5] ), .\rd_grey_sync_r[4] (\rd_grey_sync_r[4] ), 
            .\rd_grey_sync_r[3] (\rd_grey_sync_r[3] ), .\rd_grey_sync_r[2] (\rd_grey_sync_r[2] ), 
            .\rd_grey_sync_r[1] (\rd_grey_sync_r[1] ), .n4943(n4943), .\REG.mem_44_4 (\REG.mem_44_4 ), 
            .\REG.mem_45_4 (\REG.mem_45_4 ), .n4942(n4942), .\REG.mem_47_11 (\REG.mem_47_11 ), 
            .n4941(n4941), .n4940(n4940), .n4939(n4939), .n4938(n4938), 
            .\REG.mem_47_7 (\REG.mem_47_7 ), .n4937(n4937), .n4936(n4936), 
            .\REG.mem_47_5 (\REG.mem_47_5 ), .n4935(n4935), .n4934(n4934), 
            .\REG.mem_47_3 (\REG.mem_47_3 ), .n4933(n4933), .\REG.mem_47_2 (\REG.mem_47_2 ), 
            .n4932(n4932), .\REG.mem_47_1 (\REG.mem_47_1 ), .n4929(n4929), 
            .n4928(n4928), .n4927(n4927), .\REG.mem_46_14 (\REG.mem_46_14 ), 
            .\wr_addr_r[6] (\wr_addr_r[6] ), .n4926(n4926), .\REG.mem_46_13 (\REG.mem_46_13 ), 
            .n4925(n4925), .n4924(n4924), .\REG.mem_46_11 (\REG.mem_46_11 ), 
            .n4923(n4923), .n4922(n4922), .n4921(n4921), .n4920(n4920), 
            .\REG.mem_46_7 (\REG.mem_46_7 ), .n4919(n4919), .n4918(n4918), 
            .\REG.mem_46_5 (\REG.mem_46_5 ), .n4917(n4917), .n4916(n4916), 
            .\REG.mem_46_3 (\REG.mem_46_3 ), .n4915(n4915), .\REG.mem_46_2 (\REG.mem_46_2 ), 
            .n4914(n4914), .\REG.mem_46_1 (\REG.mem_46_1 ), .n4913(n4913), 
            .n4912(n4912), .n4911(n4911), .\REG.mem_45_14 (\REG.mem_45_14 ), 
            .n59(n59), .n4910(n4910), .\REG.mem_45_13 (\REG.mem_45_13 ), 
            .n4909(n4909), .n4908(n4908), .\REG.mem_45_11 (\REG.mem_45_11 ), 
            .n4907(n4907), .n4906(n4906), .n4905(n4905), .n4904(n4904), 
            .\REG.mem_45_7 (\REG.mem_45_7 ), .n4903(n4903), .n4902(n4902), 
            .\REG.mem_45_5 (\REG.mem_45_5 ), .n4901(n4901), .n4900(n4900), 
            .\REG.mem_45_3 (\REG.mem_45_3 ), .n4899(n4899), .\REG.mem_45_2 (\REG.mem_45_2 ), 
            .n4898(n4898), .\REG.mem_45_1 (\REG.mem_45_1 ), .n4897(n4897), 
            .n4896(n4896), .n27(n27), .n4895(n4895), .\REG.mem_44_14 (\REG.mem_44_14 ), 
            .n4894(n4894), .\REG.mem_44_13 (\REG.mem_44_13 ), .n4893(n4893), 
            .n4892(n4892), .\REG.mem_44_11 (\REG.mem_44_11 ), .n4891(n4891), 
            .n4890(n4890), .n4889(n4889), .n4888(n4888), .\REG.mem_44_7 (\REG.mem_44_7 ), 
            .n4887(n4887), .n4886(n4886), .\REG.mem_44_5 (\REG.mem_44_5 ), 
            .n4885(n4885), .n4884(n4884), .\REG.mem_44_3 (\REG.mem_44_3 ), 
            .n4883(n4883), .\REG.mem_44_2 (\REG.mem_44_2 ), .n4882(n4882), 
            .\REG.mem_44_1 (\REG.mem_44_1 ), .n4880(n4880), .n4879(n4879), 
            .n4878(n4878), .n4877(n4877), .\REG.mem_43_13 (\REG.mem_43_13 ), 
            .n4876(n4876), .n4875(n4875), .\REG.mem_43_11 (\REG.mem_43_11 ), 
            .n4874(n4874), .n4873(n4873), .n4872(n4872), .\REG.mem_43_8 (\REG.mem_43_8 ), 
            .n4871(n4871), .\REG.mem_43_7 (\REG.mem_43_7 ), .n4870(n4870), 
            .\REG.mem_43_6 (\REG.mem_43_6 ), .n4869(n4869), .\REG.mem_43_5 (\REG.mem_43_5 ), 
            .n4868(n4868), .n4867(n4867), .\REG.mem_43_3 (\REG.mem_43_3 ), 
            .n4866(n4866), .\REG.mem_43_2 (\REG.mem_43_2 ), .n4865(n4865), 
            .\REG.mem_43_1 (\REG.mem_43_1 ), .n4864(n4864), .\REG.mem_43_0 (\REG.mem_43_0 ), 
            .n4863(n4863), .\REG.mem_30_2 (\REG.mem_30_2 ), .n4862(n4862), 
            .n4861(n4861), .\REG.mem_42_13 (\REG.mem_42_13 ), .n4860(n4860), 
            .n4859(n4859), .\REG.mem_42_11 (\REG.mem_42_11 ), .n4858(n4858), 
            .n4857(n4857), .n4856(n4856), .\REG.mem_42_8 (\REG.mem_42_8 ), 
            .n4855(n4855), .\REG.mem_42_7 (\REG.mem_42_7 ), .n4854(n4854), 
            .\REG.mem_42_6 (\REG.mem_42_6 ), .n4853(n4853), .\REG.mem_42_5 (\REG.mem_42_5 ), 
            .n4852(n4852), .n4851(n4851), .\REG.mem_42_3 (\REG.mem_42_3 ), 
            .n4850(n4850), .\REG.mem_42_2 (\REG.mem_42_2 ), .n4849(n4849), 
            .\REG.mem_42_1 (\REG.mem_42_1 ), .n4848(n4848), .\REG.mem_42_0 (\REG.mem_42_0 ), 
            .n4847(n4847), .\REG.mem_29_2 (\REG.mem_29_2 ), .\REG.mem_28_2 (\REG.mem_28_2 ), 
            .\REG.mem_26_11 (\REG.mem_26_11 ), .\REG.mem_6_7 (\REG.mem_6_7 ), 
            .\REG.mem_7_7 (\REG.mem_7_7 ), .\REG.mem_5_7 (\REG.mem_5_7 ), 
            .n4846(n4846), .n4845(n4845), .\REG.mem_41_13 (\REG.mem_41_13 ), 
            .n4844(n4844), .n4843(n4843), .\REG.mem_41_11 (\REG.mem_41_11 ), 
            .n4842(n4842), .n4841(n4841), .n4840(n4840), .\REG.mem_41_8 (\REG.mem_41_8 ), 
            .n4839(n4839), .\REG.mem_41_7 (\REG.mem_41_7 ), .n4838(n4838), 
            .\REG.mem_41_6 (\REG.mem_41_6 ), .n4837(n4837), .\REG.mem_41_5 (\REG.mem_41_5 ), 
            .n4836(n4836), .n4835(n4835), .\REG.mem_41_3 (\REG.mem_41_3 ), 
            .n4834(n4834), .\REG.mem_41_2 (\REG.mem_41_2 ), .n4833(n4833), 
            .\REG.mem_41_1 (\REG.mem_41_1 ), .n4832(n4832), .\REG.mem_41_0 (\REG.mem_41_0 ), 
            .\REG.mem_18_7 (\REG.mem_18_7 ), .\REG.mem_19_7 (\REG.mem_19_7 ), 
            .\REG.mem_25_11 (\REG.mem_25_11 ), .\REG.mem_24_11 (\REG.mem_24_11 ), 
            .n4157(n4157), .n4831(n4831), .n4830(n4830), .n4829(n4829), 
            .\REG.mem_40_13 (\REG.mem_40_13 ), .n4828(n4828), .n4827(n4827), 
            .\REG.mem_40_11 (\REG.mem_40_11 ), .n4826(n4826), .n4825(n4825), 
            .n4824(n4824), .\REG.mem_40_8 (\REG.mem_40_8 ), .n4823(n4823), 
            .\REG.mem_40_7 (\REG.mem_40_7 ), .n4822(n4822), .\REG.mem_40_6 (\REG.mem_40_6 ), 
            .n4821(n4821), .\REG.mem_40_5 (\REG.mem_40_5 ), .n4820(n4820), 
            .n4819(n4819), .\REG.mem_40_3 (\REG.mem_40_3 ), .n4818(n4818), 
            .\REG.mem_40_2 (\REG.mem_40_2 ), .n4817(n4817), .\REG.mem_40_1 (\REG.mem_40_1 ), 
            .n4814(n4814), .\REG.mem_40_0 (\REG.mem_40_0 ), .n4813(n4813), 
            .\REG.mem_39_15 (\REG.mem_39_15 ), .n4812(n4812), .\REG.mem_39_14 (\REG.mem_39_14 ), 
            .\REG.mem_22_7 (\REG.mem_22_7 ), .\REG.mem_23_7 (\REG.mem_23_7 ), 
            .n4811(n4811), .\REG.mem_39_13 (\REG.mem_39_13 ), .n4810(n4810), 
            .n4809(n4809), .\REG.mem_39_11 (\REG.mem_39_11 ), .\REG.mem_21_7 (\REG.mem_21_7 ), 
            .n4808(n4808), .\REG.mem_30_11 (\REG.mem_30_11 ), .n4807(n4807), 
            .n4806(n4806), .\REG.mem_39_8 (\REG.mem_39_8 ), .n4805(n4805), 
            .n4804(n4804), .\REG.mem_39_6 (\REG.mem_39_6 ), .n4803(n4803), 
            .n4802(n4802), .\REG.mem_39_4 (\REG.mem_39_4 ), .n4801(n4801), 
            .\REG.mem_39_3 (\REG.mem_39_3 ), .n4800(n4800), .\REG.mem_39_2 (\REG.mem_39_2 ), 
            .n4799(n4799), .\REG.mem_39_1 (\REG.mem_39_1 ), .n4798(n4798), 
            .\REG.mem_39_0 (\REG.mem_39_0 ), .n4797(n4797), .\REG.mem_38_15 (\REG.mem_38_15 ), 
            .n4796(n4796), .\REG.mem_38_14 (\REG.mem_38_14 ), .n4795(n4795), 
            .\REG.mem_38_13 (\REG.mem_38_13 ), .n4794(n4794), .n4793(n4793), 
            .\REG.mem_38_11 (\REG.mem_38_11 ), .\REG.mem_29_11 (\REG.mem_29_11 ), 
            .\REG.mem_28_11 (\REG.mem_28_11 ), .n4792(n4792), .\REG.mem_34_2 (\REG.mem_34_2 ), 
            .n4791(n4791), .n4790(n4790), .\REG.mem_38_8 (\REG.mem_38_8 ), 
            .n4789(n4789), .n4788(n4788), .\REG.mem_38_6 (\REG.mem_38_6 ), 
            .n4787(n4787), .n4786(n4786), .\REG.mem_38_4 (\REG.mem_38_4 ), 
            .n4785(n4785), .\REG.mem_38_3 (\REG.mem_38_3 ), .n4784(n4784), 
            .\REG.mem_38_2 (\REG.mem_38_2 ), .n4783(n4783), .\REG.mem_38_1 (\REG.mem_38_1 ), 
            .n4782(n4782), .\REG.mem_38_0 (\REG.mem_38_0 ), .n4781(n4781), 
            .\REG.mem_37_15 (\REG.mem_37_15 ), .n4780(n4780), .\REG.mem_37_14 (\REG.mem_37_14 ), 
            .n4779(n4779), .\REG.mem_37_13 (\REG.mem_37_13 ), .n4778(n4778), 
            .n4777(n4777), .\REG.mem_37_11 (\REG.mem_37_11 ), .n4776(n4776), 
            .n4775(n4775), .n4774(n4774), .\REG.mem_37_8 (\REG.mem_37_8 ), 
            .n4773(n4773), .n4772(n4772), .\REG.mem_37_6 (\REG.mem_37_6 ), 
            .n4771(n4771), .n4770(n4770), .\REG.mem_37_4 (\REG.mem_37_4 ), 
            .n4769(n4769), .\REG.mem_37_3 (\REG.mem_37_3 ), .n4768(n4768), 
            .\REG.mem_37_2 (\REG.mem_37_2 ), .n4767(n4767), .\REG.mem_37_1 (\REG.mem_37_1 ), 
            .n4766(n4766), .\REG.mem_37_0 (\REG.mem_37_0 ), .n4156(n4156), 
            .\REG.mem_26_6 (\REG.mem_26_6 ), .\REG.mem_25_6 (\REG.mem_25_6 ), 
            .\REG.mem_24_6 (\REG.mem_24_6 ), .\REG.mem_34_9 (\REG.mem_34_9 ), 
            .n4733(n4733), .\REG.mem_34_15 (\REG.mem_34_15 ), .n4732(n4732), 
            .\REG.mem_34_14 (\REG.mem_34_14 ), .n4731(n4731), .\REG.mem_34_13 (\REG.mem_34_13 ), 
            .n4730(n4730), .n4729(n4729), .\REG.mem_34_11 (\REG.mem_34_11 ), 
            .n4728(n4728), .n4727(n4727), .n4726(n4726), .\REG.mem_34_8 (\REG.mem_34_8 ), 
            .n4725(n4725), .n4155(n4155), .\REG.mem_2_1 (\REG.mem_2_1 ), 
            .n4154(n4154), .\REG.mem_24_4 (\REG.mem_24_4 ), .\REG.mem_25_4 (\REG.mem_25_4 ), 
            .\REG.mem_26_4 (\REG.mem_26_4 ), .n4724(n4724), .\REG.mem_34_6 (\REG.mem_34_6 ), 
            .\REG.mem_30_4 (\REG.mem_30_4 ), .\REG.mem_28_4 (\REG.mem_28_4 ), 
            .\REG.mem_29_4 (\REG.mem_29_4 ), .n4723(n4723), .n4722(n4722), 
            .\REG.mem_34_4 (\REG.mem_34_4 ), .n4721(n4721), .\REG.mem_34_3 (\REG.mem_34_3 ), 
            .n4720(n4720), .n4719(n4719), .\REG.mem_34_1 (\REG.mem_34_1 ), 
            .n4718(n4718), .\REG.mem_8_4 (\REG.mem_8_4 ), .\REG.mem_9_4 (\REG.mem_9_4 ), 
            .\REG.mem_10_4 (\REG.mem_10_4 ), .\REG.mem_11_4 (\REG.mem_11_4 ), 
            .\REG.mem_14_4 (\REG.mem_14_4 ), .\REG.mem_15_4 (\REG.mem_15_4 ), 
            .\REG.mem_12_4 (\REG.mem_12_4 ), .\REG.mem_13_4 (\REG.mem_13_4 ), 
            .\REG.mem_6_1 (\REG.mem_6_1 ), .\REG.mem_7_1 (\REG.mem_7_1 ), 
            .\REG.mem_5_1 (\REG.mem_5_1 ), .n4677(n4677), .rp_sync1_r({rp_sync1_r}), 
            .\REG.mem_26_10 (\REG.mem_26_10 ), .\REG.mem_18_1 (\REG.mem_18_1 ), 
            .\REG.mem_19_1 (\REG.mem_19_1 ), .n4676(n4676), .n4675(n4675), 
            .n4674(n4674), .n4673(n4673), .n4672(n4672), .\REG.mem_25_10 (\REG.mem_25_10 ), 
            .\REG.mem_24_10 (\REG.mem_24_10 ), .\REG.mem_22_1 (\REG.mem_22_1 ), 
            .\REG.mem_23_1 (\REG.mem_23_1 ), .\REG.mem_21_1 (\REG.mem_21_1 ), 
            .n46(n46), .n14(n14), .n4655(n4655), .n4654(n4654), .n4653(n4653), 
            .n4652(n4652), .n4651(n4651), .n4650(n4650), .n4649(n4649), 
            .n4648(n4648), .n4647(n4647), .\REG.mem_30_13 (\REG.mem_30_13 ), 
            .n4646(n4646), .\REG.mem_30_12 (\REG.mem_30_12 ), .n4645(n4645), 
            .n37(n37), .n5(n5), .n4644(n4644), .n4643(n4643), .n4642(n4642), 
            .n4641(n4641), .n4640(n4640), .\REG.mem_30_6 (\REG.mem_30_6 ), 
            .n4639(n4639), .n4638(n4638), .n4637(n4637), .n4636(n4636), 
            .n4635(n4635), .\REG.mem_30_1 (\REG.mem_30_1 ), .n4634(n4634), 
            .n4633(n4633), .n4631(n4631), .n4629(n4629), .\REG.mem_18_14 (\REG.mem_18_14 ), 
            .\REG.mem_19_14 (\REG.mem_19_14 ), .n4627(n4627), .n51(n51), 
            .n4626(n4626), .n4625(n4625), .\REG.mem_29_13 (\REG.mem_29_13 ), 
            .\REG.mem_22_14 (\REG.mem_22_14 ), .\REG.mem_23_14 (\REG.mem_23_14 ), 
            .\REG.mem_21_14 (\REG.mem_21_14 ), .n4624(n4624), .\REG.mem_29_12 (\REG.mem_29_12 ), 
            .n4623(n4623), .n4622(n4622), .n4621(n4621), .n4620(n4620), 
            .n4619(n4619), .n4618(n4618), .\REG.mem_29_6 (\REG.mem_29_6 ), 
            .n4617(n4617), .n4616(n4616), .n4615(n4615), .n4614(n4614), 
            .n4613(n4613), .\REG.mem_29_1 (\REG.mem_29_1 ), .n4612(n4612), 
            .n4611(n4611), .n4610(n4610), .n4609(n4609), .\REG.mem_28_13 (\REG.mem_28_13 ), 
            .n19(n19), .n4608(n4608), .\REG.mem_28_12 (\REG.mem_28_12 ), 
            .n4607(n4607), .\REG.mem_18_12 (\REG.mem_18_12 ), .\REG.mem_19_12 (\REG.mem_19_12 ), 
            .\REG.mem_22_12 (\REG.mem_22_12 ), .\REG.mem_23_12 (\REG.mem_23_12 ), 
            .n4606(n4606), .n4605(n4605), .n4604(n4604), .n4603(n4603), 
            .n4602(n4602), .\REG.mem_28_6 (\REG.mem_28_6 ), .n4601(n4601), 
            .n4600(n4600), .n4599(n4599), .n4598(n4598), .n4597(n4597), 
            .\REG.mem_28_1 (\REG.mem_28_1 ), .n4596(n4596), .\REG.mem_21_12 (\REG.mem_21_12 ), 
            .n4579(n4579), .n4578(n4578), .n4577(n4577), .\REG.mem_26_13 (\REG.mem_26_13 ), 
            .n4576(n4576), .\REG.mem_26_12 (\REG.mem_26_12 ), .n4575(n4575), 
            .n4574(n4574), .n4573(n4573), .n4572(n4572), .n4571(n4571), 
            .\REG.mem_26_7 (\REG.mem_26_7 ), .n4570(n4570), .n4569(n4569), 
            .n4568(n4568), .n4567(n4567), .\REG.mem_6_13 (\REG.mem_6_13 ), 
            .\REG.mem_7_13 (\REG.mem_7_13 ), .n4566(n4566), .n4565(n4565), 
            .\REG.mem_26_1 (\REG.mem_26_1 ), .n4564(n4564), .\REG.mem_26_0 (\REG.mem_26_0 ), 
            .n4563(n4563), .wp_sync1_r({wp_sync1_r}), .n4562(n4562), .n4561(n4561), 
            .n4560(n4560), .n4559(n4559), .n4558(n4558), .n4557(n4557), 
            .n4556(n4556), .\REG.mem_25_13 (\REG.mem_25_13 ), .n4555(n4555), 
            .\REG.mem_25_12 (\REG.mem_25_12 ), .n4554(n4554), .n4553(n4553), 
            .n4552(n4552), .n4551(n4551), .\REG.mem_5_13 (\REG.mem_5_13 ), 
            .n4550(n4550), .\REG.mem_25_7 (\REG.mem_25_7 ), .n4549(n4549), 
            .n4548(n4548), .n4547(n4547), .n4546(n4546), .n4545(n4545), 
            .n4544(n4544), .\REG.mem_25_1 (\REG.mem_25_1 ), .n4543(n4543), 
            .\REG.mem_25_0 (\REG.mem_25_0 ), .n4542(n4542), .n4541(n4541), 
            .n4540(n4540), .n4539(n4539), .n4538(n4538), .n4537(n4537), 
            .n4536(n4536), .n4535(n4535), .n4534(n4534), .\REG.mem_18_0 (\REG.mem_18_0 ), 
            .\REG.mem_19_0 (\REG.mem_19_0 ), .\REG.mem_22_0 (\REG.mem_22_0 ), 
            .\REG.mem_23_0 (\REG.mem_23_0 ), .\REG.mem_21_0 (\REG.mem_21_0 ), 
            .DEBUG_9_c(DEBUG_9_c), .n4533(n4533), .\REG.mem_24_13 (\REG.mem_24_13 ), 
            .n4532(n4532), .\REG.mem_24_12 (\REG.mem_24_12 ), .n4531(n4531), 
            .n4530(n4530), .n4529(n4529), .n4528(n4528), .n4527(n4527), 
            .\REG.mem_24_7 (\REG.mem_24_7 ), .n4526(n4526), .n4525(n4525), 
            .n4524(n4524), .n4523(n4523), .n4522(n4522), .n4521(n4521), 
            .\REG.mem_24_1 (\REG.mem_24_1 ), .n4520(n4520), .\REG.mem_24_0 (\REG.mem_24_0 ), 
            .n4519(n4519), .\REG.mem_23_15 (\REG.mem_23_15 ), .n4518(n4518), 
            .n4517(n4517), .n4516(n4516), .n4515(n4515), .n4514(n4514), 
            .\REG.mem_23_10 (\REG.mem_23_10 ), .n4513(n4513), .\REG.mem_23_9 (\REG.mem_23_9 ), 
            .n4512(n4512), .n4511(n4511), .n4510(n4510), .n4509(n4509), 
            .n4508(n4508), .\REG.mem_23_4 (\REG.mem_23_4 ), .n4507(n4507), 
            .n4506(n4506), .n4505(n4505), .n4504(n4504), .n4503(n4503), 
            .\REG.mem_22_15 (\REG.mem_22_15 ), .n4502(n4502), .n4501(n4501), 
            .n4500(n4500), .n4499(n4499), .n4498(n4498), .\REG.mem_22_10 (\REG.mem_22_10 ), 
            .n4497(n4497), .\REG.mem_22_9 (\REG.mem_22_9 ), .n4496(n4496), 
            .n4495(n4495), .n4494(n4494), .n4493(n4493), .n4492(n4492), 
            .\REG.mem_22_4 (\REG.mem_22_4 ), .n4491(n4491), .n4490(n4490), 
            .n4489(n4489), .n4488(n4488), .n4487(n4487), .\REG.mem_21_15 (\REG.mem_21_15 ), 
            .n4486(n4486), .n4485(n4485), .n4484(n4484), .n4483(n4483), 
            .n4482(n4482), .\REG.mem_21_10 (\REG.mem_21_10 ), .n4481(n4481), 
            .\REG.mem_21_9 (\REG.mem_21_9 ), .n4480(n4480), .n4479(n4479), 
            .n4478(n4478), .n4477(n4477), .n4476(n4476), .\REG.mem_21_4 (\REG.mem_21_4 ), 
            .n4475(n4475), .n4474(n4474), .n4473(n4473), .\REG.mem_6_12 (\REG.mem_6_12 ), 
            .\REG.mem_7_12 (\REG.mem_7_12 ), .n4472(n4472), .\REG.out_raw[15] (\REG.out_raw[15] ), 
            .\REG.out_raw[14] (\REG.out_raw[14] ), .\REG.out_raw[13] (\REG.out_raw[13] ), 
            .\REG.mem_5_12 (\REG.mem_5_12 ), .\REG.out_raw[12] (\REG.out_raw[12] ), 
            .\REG.out_raw[11] (\REG.out_raw[11] ), .\REG.out_raw[10] (\REG.out_raw[10] ), 
            .n4455(n4455), .\REG.mem_19_15 (\REG.mem_19_15 ), .n4454(n4454), 
            .n4453(n4453), .n4452(n4452), .n4451(n4451), .n4450(n4450), 
            .n4449(n4449), .\REG.mem_19_9 (\REG.mem_19_9 ), .n4448(n4448), 
            .n4447(n4447), .n4446(n4446), .n4445(n4445), .n4444(n4444), 
            .\REG.mem_19_4 (\REG.mem_19_4 ), .n4443(n4443), .n4442(n4442), 
            .n4441(n4441), .n4440(n4440), .\REG.out_raw[9] (\REG.out_raw[9] ), 
            .\REG.out_raw[8] (\REG.out_raw[8] ), .n4439(n4439), .\REG.mem_18_15 (\REG.mem_18_15 ), 
            .\REG.out_raw[7] (\REG.out_raw[7] ), .\REG.out_raw[6] (\REG.out_raw[6] ), 
            .\REG.out_raw[5] (\REG.out_raw[5] ), .\REG.out_raw[4] (\REG.out_raw[4] ), 
            .\REG.out_raw[3] (\REG.out_raw[3] ), .n4438(n4438), .\REG.mem_6_9 (\REG.mem_6_9 ), 
            .\REG.mem_7_9 (\REG.mem_7_9 ), .n54(n54), .\REG.mem_5_9 (\REG.mem_5_9 ), 
            .n4437(n4437), .n4436(n4436), .n4435(n4435), .n4434(n4434), 
            .n4433(n4433), .\REG.mem_18_9 (\REG.mem_18_9 ), .n4432(n4432), 
            .n4431(n4431), .n4430(n4430), .n4429(n4429), .n4428(n4428), 
            .\REG.mem_18_4 (\REG.mem_18_4 ), .n4427(n4427), .n4426(n4426), 
            .n4425(n4425), .n4424(n4424), .\REG.out_raw[2] (\REG.out_raw[2] ), 
            .n22(n22), .n39(n39), .\REG.mem_10_9 (\REG.mem_10_9 ), .\REG.mem_11_9 (\REG.mem_11_9 ), 
            .\REG.mem_10_13 (\REG.mem_10_13 ), .\REG.mem_11_13 (\REG.mem_11_13 ), 
            .n7(n7), .n40(n40), .\REG.mem_9_9 (\REG.mem_9_9 ), .\REG.mem_8_9 (\REG.mem_8_9 ), 
            .\REG.mem_9_13 (\REG.mem_9_13 ), .\REG.mem_8_13 (\REG.mem_8_13 ), 
            .n8(n8), .\REG.mem_14_12 (\REG.mem_14_12 ), .\REG.mem_15_12 (\REG.mem_15_12 ), 
            .n4391(n4391), .\REG.out_raw[1] (\REG.out_raw[1] ), .n4390(n4390), 
            .\REG.mem_13_12 (\REG.mem_13_12 ), .\REG.mem_12_12 (\REG.mem_12_12 ), 
            .n4389(n4389), .\REG.mem_15_13 (\REG.mem_15_13 ), .n4388(n4388), 
            .n4387(n4387), .n4386(n4386), .\REG.mem_15_10 (\REG.mem_15_10 ), 
            .n4385(n4385), .\REG.mem_15_9 (\REG.mem_15_9 ), .n4384(n4384), 
            .\REG.mem_15_8 (\REG.mem_15_8 ), .n4383(n4383), .\REG.mem_15_7 (\REG.mem_15_7 ), 
            .n4382(n4382), .n4381(n4381), .\REG.mem_15_5 (\REG.mem_15_5 ), 
            .n4380(n4380), .n4379(n4379), .n4378(n4378), .n4377(n4377), 
            .\REG.mem_15_1 (\REG.mem_15_1 ), .n4376(n4376), .n4375(n4375), 
            .n4374(n4374), .\REG.mem_6_8 (\REG.mem_6_8 ), .\REG.mem_7_8 (\REG.mem_7_8 ), 
            .\REG.mem_5_8 (\REG.mem_5_8 ), .\REG.mem_14_9 (\REG.mem_14_9 ), 
            .\REG.mem_13_9 (\REG.mem_13_9 ), .\REG.mem_12_9 (\REG.mem_12_9 ), 
            .\REG.mem_6_5 (\REG.mem_6_5 ), .\REG.mem_7_5 (\REG.mem_7_5 ), 
            .n4373(n4373), .\REG.mem_14_13 (\REG.mem_14_13 ), .n4372(n4372), 
            .n4371(n4371), .n4370(n4370), .\REG.mem_14_10 (\REG.mem_14_10 ), 
            .n4369(n4369), .n4368(n4368), .\REG.mem_14_8 (\REG.mem_14_8 ), 
            .n4367(n4367), .\REG.mem_14_7 (\REG.mem_14_7 ), .\REG.mem_5_5 (\REG.mem_5_5 ), 
            .n4366(n4366), .n4365(n4365), .\REG.mem_14_5 (\REG.mem_14_5 ), 
            .n4364(n4364), .n4363(n4363), .n4362(n4362), .n4361(n4361), 
            .\REG.mem_14_1 (\REG.mem_14_1 ), .n4360(n4360), .n4359(n4359), 
            .n4358(n4358), .n4357(n4357), .\REG.mem_13_13 (\REG.mem_13_13 ), 
            .n4356(n4356), .n4355(n4355), .n4354(n4354), .\REG.mem_13_10 (\REG.mem_13_10 ), 
            .n4353(n4353), .n4352(n4352), .\REG.mem_13_8 (\REG.mem_13_8 ), 
            .n4351(n4351), .\REG.mem_13_7 (\REG.mem_13_7 ), .n4350(n4350), 
            .n4349(n4349), .\REG.mem_13_5 (\REG.mem_13_5 ), .n4348(n4348), 
            .n4347(n4347), .n4346(n4346), .n4345(n4345), .\REG.mem_13_1 (\REG.mem_13_1 ), 
            .n4344(n4344), .n4343(n4343), .n4342(n4342), .n4341(n4341), 
            .\REG.mem_12_13 (\REG.mem_12_13 ), .n4340(n4340), .n4339(n4339), 
            .n4338(n4338), .\REG.mem_12_10 (\REG.mem_12_10 ), .n4337(n4337), 
            .n4336(n4336), .\REG.mem_12_8 (\REG.mem_12_8 ), .n4335(n4335), 
            .\REG.mem_12_7 (\REG.mem_12_7 ), .n4334(n4334), .n4333(n4333), 
            .\REG.mem_12_5 (\REG.mem_12_5 ), .n4332(n4332), .n4331(n4331), 
            .n4330(n4330), .n4329(n4329), .\REG.mem_12_1 (\REG.mem_12_1 ), 
            .n4328(n4328), .n4327(n4327), .n4326(n4326), .n4325(n4325), 
            .n4324(n4324), .n4323(n4323), .n60(n60), .n4322(n4322), 
            .n28(n28), .n41(n41), .n9(n9), .n4321(n4321), .n4320(n4320), 
            .\REG.mem_11_8 (\REG.mem_11_8 ), .n4319(n4319), .\REG.mem_11_7 (\REG.mem_11_7 ), 
            .n4318(n4318), .n4317(n4317), .\REG.mem_11_5 (\REG.mem_11_5 ), 
            .n4316(n4316), .n4315(n4315), .n4314(n4314), .n4313(n4313), 
            .\REG.mem_11_1 (\REG.mem_11_1 ), .n4312(n4312), .n4311(n4311), 
            .n42(n42), .n4310(n4310), .n4309(n4309), .n4308(n4308), 
            .n10(n10), .n4307(n4307), .n4306(n4306), .n4305(n4305), 
            .n4304(n4304), .\REG.mem_10_8 (\REG.mem_10_8 ), .n4303(n4303), 
            .\REG.mem_10_7 (\REG.mem_10_7 ), .n4302(n4302), .n4301(n4301), 
            .\REG.mem_10_5 (\REG.mem_10_5 ), .n4300(n4300), .n4299(n4299), 
            .n4298(n4298), .n4297(n4297), .\REG.mem_10_1 (\REG.mem_10_1 ), 
            .n4296(n4296), .n4130(n4130), .n57(n57), .\REG.mem_9_5 (\REG.mem_9_5 ), 
            .\REG.mem_8_5 (\REG.mem_8_5 ), .n4288(n4288), .n4287(n4287), 
            .n4286(n4286), .n4285(n4285), .n4284(n4284), .n4283(n4283), 
            .n4282(n4282), .n4281(n4281), .n4280(n4280), .\REG.mem_9_8 (\REG.mem_9_8 ), 
            .n4279(n4279), .\REG.mem_9_7 (\REG.mem_9_7 ), .n4278(n4278), 
            .n4277(n4277), .n4108(n4108), .n25(n25), .n4276(n4276), 
            .n43(n43), .n11(n11), .n44(n44), .n12(n12), .n4275(n4275), 
            .n4274(n4274), .n4273(n4273), .\REG.mem_9_1 (\REG.mem_9_1 ), 
            .n4272(n4272), .n4270(n4270), .n4268(n4268), .n4107(n4107), 
            .\REG.mem_8_7 (\REG.mem_8_7 ), .n4265(n4265), .n4264(n4264), 
            .n4263(n4263), .n4262(n4262), .n4261(n4261), .n52(n52), 
            .n4260(n4260), .\REG.mem_8_8 (\REG.mem_8_8 ), .n4259(n4259), 
            .n4258(n4258), .n4257(n4257), .n4256(n4256), .n4255(n4255), 
            .n4254(n4254), .n4253(n4253), .n4252(n4252), .n4251(n4251), 
            .\REG.mem_8_1 (\REG.mem_8_1 ), .n4250(n4250), .n4249(n4249), 
            .n4248(n4248), .n4247(n4247), .n4246(n4246), .n4245(n4245), 
            .\REG.mem_7_11 (\REG.mem_7_11 ), .n4244(n4244), .n4243(n4243), 
            .n4242(n4242), .n4241(n4241), .n4240(n4240), .n4239(n4239), 
            .n4238(n4238), .\REG.mem_7_4 (\REG.mem_7_4 ), .n4237(n4237), 
            .n4236(n4236), .n4235(n4235), .n4234(n4234), .n4233(n4233), 
            .n4232(n4232), .n4231(n4231), .n4230(n4230), .n4229(n4229), 
            .\REG.mem_6_11 (\REG.mem_6_11 ), .n4228(n4228), .n4227(n4227), 
            .n4226(n4226), .n4225(n4225), .n4224(n4224), .n4223(n4223), 
            .n4222(n4222), .\REG.mem_6_4 (\REG.mem_6_4 ), .n4221(n4221), 
            .n4220(n4220), .n4219(n4219), .n4218(n4218), .n4217(n4217), 
            .n4216(n4216), .n4215(n4215), .n4214(n4214), .n4213(n4213), 
            .\REG.mem_5_11 (\REG.mem_5_11 ), .n4212(n4212), .n4211(n4211), 
            .n4210(n4210), .n4209(n4209), .n4208(n4208), .n4207(n4207), 
            .n4206(n4206), .\REG.mem_5_4 (\REG.mem_5_4 ), .n4205(n4205), 
            .n4204(n4204), .n4203(n4203), .n4202(n4202), .n4103(n4103), 
            .n20(n20), .n53(n53), .n4101(n4101), .n21(n21), .n35(n35), 
            .n3(n3), .n36(n36), .n55(n55), .n23(n23), .n4(n4), .n47(n47), 
            .n15(n15), .n31(n31), .n63(n63)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_dc_32_lut_gen.v(51[33] 70[34])
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1
//

module fifo_dc_32_lut_gen_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 (FIFO_D6_c_6, 
            \REG.mem_42_15 , \REG.mem_43_15 , FIFO_D5_c_5, \REG.mem_29_14 , 
            \REG.mem_28_14 , FIFO_CLK_c, \REG.mem_41_15 , \REG.mem_40_15 , 
            GND_net, \REG.mem_2_0 , \REG.mem_2_2 , FIFO_D4_c_4, \REG.mem_18_5 , 
            \REG.mem_19_5 , FIFO_D3_c_3, \REG.mem_62_5 , \REG.mem_61_5 , 
            \REG.mem_60_5 , FIFO_D2_c_2, t_rd_fifo_en_w, \REG.out_raw[0] , 
            DEBUG_6_c, \REG.mem_30_10 , \REG.mem_29_10 , \REG.mem_28_10 , 
            \REG.mem_58_8 , \REG.mem_57_8 , \REG.mem_56_8 , FIFO_D1_c_1, 
            \REG.mem_2_14 , FIFO_D0_c_0, \REG.mem_14_15 , \REG.mem_15_15 , 
            \REG.mem_13_15 , \REG.mem_12_15 , \REG.mem_10_15 , \REG.mem_11_15 , 
            n56, \REG.mem_62_8 , \REG.mem_61_8 , \REG.mem_60_8 , \REG.mem_46_6 , 
            \REG.mem_47_6 , n24, write_to_dc32_fifo, reset_all, \wr_addr_nxt_c[1] , 
            \REG.mem_45_6 , \REG.mem_44_6 , dc32_fifo_is_full, \REG.mem_34_10 , 
            \REG.mem_18_8 , \REG.mem_19_8 , \REG.mem_58_11 , \rd_grey_sync_r[0] , 
            \REG.mem_57_11 , \REG.mem_56_11 , \REG.mem_6_14 , \REG.mem_7_14 , 
            \REG.mem_5_14 , \REG.mem_10_12 , \REG.mem_11_12 , \REG.mem_9_12 , 
            \REG.mem_8_12 , \REG.mem_6_10 , \REG.mem_7_10 , \REG.mem_26_9 , 
            DEBUG_1_c, \REG.mem_6_0 , \REG.mem_7_0 , \REG.mem_5_0 , 
            \REG.mem_5_10 , \REG.mem_25_9 , \REG.mem_24_9 , \REG.mem_56_7 , 
            \REG.mem_57_7 , \REG.mem_58_7 , \num_words_in_buffer[3] , 
            \wr_grey_sync_r[0] , \REG.mem_10_14 , \REG.mem_11_14 , \REG.mem_9_14 , 
            \REG.mem_8_14 , \REG.mem_14_14 , \REG.mem_15_14 , \REG.mem_13_14 , 
            \REG.mem_12_14 , \REG.mem_38_9 , \REG.mem_39_9 , \REG.mem_37_9 , 
            \REG.mem_34_7 , \REG.mem_42_9 , \REG.mem_43_9 , \REG.mem_10_10 , 
            \REG.mem_11_10 , \REG.mem_9_10 , \REG.mem_8_10 , \REG.mem_41_9 , 
            \REG.mem_40_9 , \REG.mem_9_15 , \REG.mem_8_15 , \REG.mem_18_6 , 
            \REG.mem_19_6 , \wr_addr_nxt_c[3] , FIFO_D15_c_15, \REG.mem_22_5 , 
            \REG.mem_23_5 , \REG.mem_21_5 , \REG.mem_38_10 , \REG.mem_39_10 , 
            \REG.mem_37_10 , \REG.mem_18_10 , \REG.mem_19_10 , FIFO_D14_c_14, 
            \REG.mem_34_12 , \REG.mem_22_6 , \REG.mem_23_6 , \REG.mem_26_14 , 
            \REG.mem_25_14 , \REG.mem_24_14 , \REG.mem_18_13 , \REG.mem_19_13 , 
            \REG.mem_62_7 , \REG.mem_21_6 , \REG.mem_60_7 , \REG.mem_61_7 , 
            \REG.mem_30_14 , \REG.mem_50_3 , \REG.mem_51_3 , \REG.mem_38_12 , 
            \REG.mem_39_12 , \REG.mem_37_12 , \REG.mem_46_8 , \REG.mem_47_8 , 
            \REG.mem_45_8 , \REG.mem_44_8 , \REG.mem_58_10 , \REG.mem_2_3 , 
            \REG.mem_57_10 , \REG.mem_56_10 , \REG.mem_62_2 , \REG.mem_61_2 , 
            \REG.mem_60_2 , \REG.mem_58_15 , \REG.mem_10_0 , \REG.mem_11_0 , 
            \REG.mem_9_0 , \REG.mem_8_0 , \REG.mem_57_15 , \REG.mem_56_15 , 
            \REG.mem_30_0 , \REG.mem_29_0 , \REG.mem_28_0 , \REG.mem_38_7 , 
            \REG.mem_39_7 , FIFO_D13_c_13, \REG.mem_37_7 , n58, FIFO_D12_c_12, 
            \REG.mem_26_5 , \REG.mem_25_5 , \REG.mem_24_5 , n50, \REG.mem_46_0 , 
            \REG.mem_47_0 , \REG.mem_6_3 , \REG.mem_7_3 , \REG.mem_5_3 , 
            \REG.mem_45_0 , \REG.mem_44_0 , \REG.mem_50_8 , \REG.mem_51_8 , 
            n18, \REG.mem_10_3 , \REG.mem_11_3 , \REG.mem_6_2 , \REG.mem_7_2 , 
            \REG.mem_5_2 , \REG.mem_9_3 , \REG.mem_8_3 , \wr_addr_nxt_c[5] , 
            \REG.mem_42_12 , \REG.mem_43_12 , \REG.mem_41_12 , \REG.mem_40_12 , 
            \REG.mem_10_2 , \REG.mem_11_2 , n4169, \REG.mem_2_15 , \REG.mem_9_2 , 
            \REG.mem_8_2 , n4168, n4167, \REG.mem_2_13 , n4166, \REG.mem_2_12 , 
            n4165, \REG.mem_2_11 , n4164, \REG.mem_2_10 , \REG.mem_6_6 , 
            \REG.mem_7_6 , n4163, \REG.mem_2_9 , \REG.mem_5_6 , \REG.mem_30_3 , 
            \REG.mem_29_3 , \REG.mem_28_3 , \REG.mem_22_13 , \REG.mem_23_13 , 
            \REG.mem_21_13 , \REG.mem_54_3 , \REG.mem_55_3 , \REG.mem_53_3 , 
            \REG.mem_42_10 , \REG.mem_43_10 , \REG.mem_41_10 , \REG.mem_40_10 , 
            \REG.mem_56_4 , \REG.mem_57_4 , \REG.mem_6_15 , \REG.mem_7_15 , 
            \REG.mem_58_4 , \REG.mem_26_15 , \REG.mem_5_15 , \REG.mem_25_15 , 
            \REG.mem_24_15 , \REG.mem_58_3 , \REG.mem_57_3 , \REG.mem_56_3 , 
            \REG.mem_62_3 , \REG.mem_62_4 , \REG.mem_60_4 , \REG.mem_61_4 , 
            \REG.mem_61_3 , \REG.mem_60_3 , \rd_addr_r[6] , \rd_addr_nxt_c_6__N_176[5] , 
            \REG.mem_22_8 , \REG.mem_23_8 , \rd_addr_nxt_c_6__N_176[3] , 
            \REG.mem_21_8 , \REG.mem_54_8 , \REG.mem_55_8 , FIFO_D11_c_11, 
            \REG.mem_14_3 , \REG.mem_15_3 , \REG.mem_53_8 , \REG.mem_14_2 , 
            \REG.mem_15_2 , \REG.mem_13_3 , \REG.mem_12_3 , \REG.mem_13_2 , 
            \REG.mem_12_2 , \REG.mem_30_5 , \REG.mem_58_13 , \REG.mem_29_5 , 
            \REG.mem_28_5 , \REG.mem_34_5 , \REG.mem_57_13 , \REG.mem_56_13 , 
            \REG.mem_14_6 , \REG.mem_15_6 , \REG.mem_13_6 , \REG.mem_12_6 , 
            \REG.mem_54_9 , \REG.mem_55_9 , \REG.mem_53_9 , \REG.mem_34_0 , 
            \REG.mem_14_0 , \REG.mem_15_0 , \REG.mem_13_0 , \REG.mem_12_0 , 
            FIFO_D10_c_10, \REG.mem_42_14 , \REG.mem_43_14 , \REG.mem_41_14 , 
            \REG.mem_40_14 , n4162, \REG.mem_2_8 , n4161, \REG.mem_2_7 , 
            FIFO_D9_c_9, n5327, VCC_net, \fifo_data_out[0] , \REG.mem_10_11 , 
            \REG.mem_11_11 , FIFO_D8_c_8, FIFO_D7_c_7, \REG.mem_9_11 , 
            \REG.mem_8_11 , \REG.mem_62_15 , \REG.mem_62_10 , n5305, 
            \fifo_data_out[15] , \REG.mem_46_12 , \REG.mem_47_12 , n5302, 
            \fifo_data_out[14] , \REG.mem_61_10 , \REG.mem_60_10 , \REG.mem_61_15 , 
            \REG.mem_60_15 , n5299, \fifo_data_out[13] , n5296, \fifo_data_out[12] , 
            n5293, \fifo_data_out[11] , n5290, \fifo_data_out[10] , 
            \REG.mem_45_12 , \REG.mem_44_12 , \REG.mem_46_15 , \REG.mem_47_15 , 
            \REG.mem_18_3 , \REG.mem_19_3 , n5255, \fifo_data_out[9] , 
            n5252, \fifo_data_out[8] , n5249, \fifo_data_out[7] , \REG.mem_45_15 , 
            \REG.mem_44_15 , n4160, \REG.mem_2_6 , \REG.mem_14_11 , 
            \REG.mem_15_11 , n4159, \REG.mem_2_5 , n5236, \fifo_data_out[6] , 
            n5233, \fifo_data_out[5] , \REG.mem_13_11 , \REG.mem_12_11 , 
            n5230, \fifo_data_out[4] , \wr_grey_sync_r[5] , \wr_grey_sync_r[4] , 
            \wr_grey_sync_r[3] , n5212, \fifo_data_out[3] , \REG.mem_18_2 , 
            \REG.mem_19_2 , n5208, n5207, \REG.mem_62_14 , n5206, 
            \REG.mem_62_13 , n5205, \REG.mem_62_12 , n5204, \REG.mem_62_11 , 
            n5203, n5202, \REG.mem_62_9 , n5201, n5200, \wr_grey_sync_r[2] , 
            \wr_grey_sync_r[1] , n5199, \REG.mem_62_6 , n5198, n5197, 
            n5196, n5195, n5194, \REG.mem_62_1 , n5193, \REG.mem_62_0 , 
            n5192, n5191, \REG.mem_61_14 , n5190, \REG.mem_61_13 , 
            n5189, \REG.mem_61_12 , n5188, \REG.mem_61_11 , n5187, 
            n5186, \REG.mem_61_9 , n5185, n5184, n5183, \REG.mem_61_6 , 
            \REG.mem_22_3 , \REG.mem_23_3 , \REG.mem_26_8 , n5182, \REG.mem_21_3 , 
            n5181, n5180, n5179, n5178, \REG.mem_61_1 , n5177, \REG.mem_61_0 , 
            n5176, n5175, \REG.mem_60_14 , n5174, \REG.mem_60_13 , 
            n5173, \REG.mem_60_12 , n5172, \REG.mem_60_11 , n5171, 
            n5170, \REG.mem_60_9 , n5169, n5168, n5167, \REG.mem_60_6 , 
            \REG.mem_25_8 , \REG.mem_24_8 , \REG.mem_46_9 , \REG.mem_47_9 , 
            \REG.mem_45_9 , \REG.mem_44_9 , \REG.mem_30_7 , n5166, n5165, 
            n5164, n5163, n5162, \REG.mem_60_1 , n5161, \REG.mem_60_0 , 
            \REG.mem_29_7 , \REG.mem_28_7 , n5144, n5143, \REG.mem_58_14 , 
            n5142, n5141, \REG.mem_58_12 , n5140, n5139, n5138, 
            \REG.mem_58_9 , n5137, n5136, n5135, \REG.mem_58_6 , \REG.mem_46_10 , 
            \REG.mem_47_10 , \REG.mem_45_10 , \REG.mem_44_10 , n5134, 
            \REG.mem_58_5 , \REG.mem_30_9 , n5133, n5132, n5131, \REG.mem_58_2 , 
            n5130, \REG.mem_58_1 , n5129, \REG.mem_58_0 , n5128, n5127, 
            \REG.mem_57_14 , n5126, n5125, \REG.mem_57_12 , n5124, 
            n5123, n5122, \REG.mem_57_9 , n5121, n5120, n5119, \REG.mem_57_6 , 
            \REG.mem_29_9 , \REG.mem_28_9 , n5118, \REG.mem_57_5 , n5117, 
            n5116, n5115, \REG.mem_57_2 , n5114, \REG.mem_57_1 , n5113, 
            \fifo_data_out[2] , n5110, \REG.mem_57_0 , n5109, n5108, 
            \REG.mem_56_14 , n5107, n5106, \REG.mem_56_12 , n5105, 
            n5104, n5103, \REG.mem_56_9 , \REG.mem_10_6 , \REG.mem_11_6 , 
            n5102, \REG.mem_9_6 , \REG.mem_8_6 , n5101, n5100, \REG.mem_56_6 , 
            n5099, \REG.mem_56_5 , n5098, n5097, n5096, \REG.mem_56_2 , 
            n5095, \REG.mem_56_1 , n5094, \fifo_data_out[1] , n5091, 
            \REG.mem_56_0 , n5090, \REG.mem_55_15 , n5089, \REG.mem_55_14 , 
            n5088, \REG.mem_55_13 , n5087, \REG.mem_55_12 , \REG.mem_22_2 , 
            \REG.mem_23_2 , \REG.mem_21_2 , n5086, \REG.mem_55_11 , 
            n5085, \REG.mem_55_10 , n5084, n5083, n5082, \REG.mem_55_7 , 
            n5081, \REG.mem_55_6 , n5080, \REG.mem_55_5 , n5079, \REG.mem_55_4 , 
            n5078, n5077, \REG.mem_55_2 , n5076, \REG.mem_55_1 , n5075, 
            \REG.mem_55_0 , n5074, \REG.mem_54_15 , n5073, \REG.mem_54_14 , 
            n5072, \REG.mem_54_13 , \num_words_in_buffer[6] , \num_words_in_buffer[5] , 
            \num_words_in_buffer[4] , n5071, \REG.mem_54_12 , n5070, 
            \REG.mem_54_11 , n5069, \REG.mem_54_10 , n5068, n5067, 
            n5066, \REG.mem_54_7 , n5065, \REG.mem_54_6 , n5064, \REG.mem_54_5 , 
            n5063, \REG.mem_54_4 , n5062, n5061, \REG.mem_54_2 , n5060, 
            \REG.mem_54_1 , n5057, \REG.mem_54_0 , n5056, \REG.mem_53_15 , 
            n5055, \REG.mem_53_14 , \REG.mem_50_12 , \REG.mem_51_12 , 
            \REG.mem_38_5 , \REG.mem_39_5 , \REG.mem_37_5 , n5054, \REG.mem_53_13 , 
            n5053, \REG.mem_53_12 , n5052, \REG.mem_53_11 , n5051, 
            \REG.mem_53_10 , n5050, n5049, n5048, \REG.mem_53_7 , 
            n5047, \REG.mem_53_6 , n5046, \REG.mem_53_5 , n5045, \REG.mem_53_4 , 
            n5044, n5043, \REG.mem_53_2 , n5042, \REG.mem_53_1 , n5041, 
            \REG.mem_53_0 , \REG.mem_26_2 , \REG.mem_18_11 , \REG.mem_19_11 , 
            \REG.mem_25_2 , \REG.mem_24_2 , n5024, \REG.mem_51_15 , 
            n5023, \REG.mem_51_14 , n26, \REG.mem_26_3 , \REG.mem_25_3 , 
            \REG.mem_24_3 , \REG.mem_40_4 , \REG.mem_41_4 , n5022, \REG.mem_51_13 , 
            n5021, n5020, \REG.mem_51_11 , n5019, \REG.mem_51_10 , 
            n5018, \REG.mem_51_9 , n5017, n5016, \REG.mem_51_7 , n5015, 
            \REG.mem_51_6 , n5014, \REG.mem_51_5 , n5013, \REG.mem_51_4 , 
            n5012, n5011, \REG.mem_51_2 , n5010, \REG.mem_51_1 , n5008, 
            \REG.mem_51_0 , \REG.mem_42_4 , \REG.mem_43_4 , \REG.mem_22_11 , 
            \REG.mem_23_11 , n5007, \REG.mem_50_15 , n5006, \REG.mem_50_14 , 
            n5005, \REG.mem_50_13 , n5004, n5003, \REG.mem_50_11 , 
            n5002, \REG.mem_50_10 , n5001, \REG.mem_50_9 , n5000, 
            n4999, \REG.mem_50_7 , n4998, \REG.mem_50_6 , n4997, \REG.mem_50_5 , 
            n4996, \REG.mem_50_4 , n4995, n4994, \REG.mem_50_2 , n4993, 
            \REG.mem_50_1 , n4992, \REG.mem_50_0 , \REG.mem_21_11 , 
            \rd_addr_nxt_c_6__N_176[1] , n4158, \REG.mem_2_4 , \REG.mem_30_15 , 
            \REG.mem_29_15 , \REG.mem_28_15 , \REG.mem_30_8 , \REG.mem_29_8 , 
            \REG.mem_28_8 , \REG.mem_46_4 , \REG.mem_47_4 , n4946, n4945, 
            \REG.mem_47_14 , n4944, \REG.mem_47_13 , \rd_grey_sync_r[5] , 
            \rd_grey_sync_r[4] , \rd_grey_sync_r[3] , \rd_grey_sync_r[2] , 
            \rd_grey_sync_r[1] , n4943, \REG.mem_44_4 , \REG.mem_45_4 , 
            n4942, \REG.mem_47_11 , n4941, n4940, n4939, n4938, 
            \REG.mem_47_7 , n4937, n4936, \REG.mem_47_5 , n4935, n4934, 
            \REG.mem_47_3 , n4933, \REG.mem_47_2 , n4932, \REG.mem_47_1 , 
            n4929, n4928, n4927, \REG.mem_46_14 , \wr_addr_r[6] , 
            n4926, \REG.mem_46_13 , n4925, n4924, \REG.mem_46_11 , 
            n4923, n4922, n4921, n4920, \REG.mem_46_7 , n4919, n4918, 
            \REG.mem_46_5 , n4917, n4916, \REG.mem_46_3 , n4915, \REG.mem_46_2 , 
            n4914, \REG.mem_46_1 , n4913, n4912, n4911, \REG.mem_45_14 , 
            n59, n4910, \REG.mem_45_13 , n4909, n4908, \REG.mem_45_11 , 
            n4907, n4906, n4905, n4904, \REG.mem_45_7 , n4903, n4902, 
            \REG.mem_45_5 , n4901, n4900, \REG.mem_45_3 , n4899, \REG.mem_45_2 , 
            n4898, \REG.mem_45_1 , n4897, n4896, n27, n4895, \REG.mem_44_14 , 
            n4894, \REG.mem_44_13 , n4893, n4892, \REG.mem_44_11 , 
            n4891, n4890, n4889, n4888, \REG.mem_44_7 , n4887, n4886, 
            \REG.mem_44_5 , n4885, n4884, \REG.mem_44_3 , n4883, \REG.mem_44_2 , 
            n4882, \REG.mem_44_1 , n4880, n4879, n4878, n4877, \REG.mem_43_13 , 
            n4876, n4875, \REG.mem_43_11 , n4874, n4873, n4872, 
            \REG.mem_43_8 , n4871, \REG.mem_43_7 , n4870, \REG.mem_43_6 , 
            n4869, \REG.mem_43_5 , n4868, n4867, \REG.mem_43_3 , n4866, 
            \REG.mem_43_2 , n4865, \REG.mem_43_1 , n4864, \REG.mem_43_0 , 
            n4863, \REG.mem_30_2 , n4862, n4861, \REG.mem_42_13 , 
            n4860, n4859, \REG.mem_42_11 , n4858, n4857, n4856, 
            \REG.mem_42_8 , n4855, \REG.mem_42_7 , n4854, \REG.mem_42_6 , 
            n4853, \REG.mem_42_5 , n4852, n4851, \REG.mem_42_3 , n4850, 
            \REG.mem_42_2 , n4849, \REG.mem_42_1 , n4848, \REG.mem_42_0 , 
            n4847, \REG.mem_29_2 , \REG.mem_28_2 , \REG.mem_26_11 , 
            \REG.mem_6_7 , \REG.mem_7_7 , \REG.mem_5_7 , n4846, n4845, 
            \REG.mem_41_13 , n4844, n4843, \REG.mem_41_11 , n4842, 
            n4841, n4840, \REG.mem_41_8 , n4839, \REG.mem_41_7 , n4838, 
            \REG.mem_41_6 , n4837, \REG.mem_41_5 , n4836, n4835, \REG.mem_41_3 , 
            n4834, \REG.mem_41_2 , n4833, \REG.mem_41_1 , n4832, \REG.mem_41_0 , 
            \REG.mem_18_7 , \REG.mem_19_7 , \REG.mem_25_11 , \REG.mem_24_11 , 
            n4157, n4831, n4830, n4829, \REG.mem_40_13 , n4828, 
            n4827, \REG.mem_40_11 , n4826, n4825, n4824, \REG.mem_40_8 , 
            n4823, \REG.mem_40_7 , n4822, \REG.mem_40_6 , n4821, \REG.mem_40_5 , 
            n4820, n4819, \REG.mem_40_3 , n4818, \REG.mem_40_2 , n4817, 
            \REG.mem_40_1 , n4814, \REG.mem_40_0 , n4813, \REG.mem_39_15 , 
            n4812, \REG.mem_39_14 , \REG.mem_22_7 , \REG.mem_23_7 , 
            n4811, \REG.mem_39_13 , n4810, n4809, \REG.mem_39_11 , 
            \REG.mem_21_7 , n4808, \REG.mem_30_11 , n4807, n4806, 
            \REG.mem_39_8 , n4805, n4804, \REG.mem_39_6 , n4803, n4802, 
            \REG.mem_39_4 , n4801, \REG.mem_39_3 , n4800, \REG.mem_39_2 , 
            n4799, \REG.mem_39_1 , n4798, \REG.mem_39_0 , n4797, \REG.mem_38_15 , 
            n4796, \REG.mem_38_14 , n4795, \REG.mem_38_13 , n4794, 
            n4793, \REG.mem_38_11 , \REG.mem_29_11 , \REG.mem_28_11 , 
            n4792, \REG.mem_34_2 , n4791, n4790, \REG.mem_38_8 , n4789, 
            n4788, \REG.mem_38_6 , n4787, n4786, \REG.mem_38_4 , n4785, 
            \REG.mem_38_3 , n4784, \REG.mem_38_2 , n4783, \REG.mem_38_1 , 
            n4782, \REG.mem_38_0 , n4781, \REG.mem_37_15 , n4780, 
            \REG.mem_37_14 , n4779, \REG.mem_37_13 , n4778, n4777, 
            \REG.mem_37_11 , n4776, n4775, n4774, \REG.mem_37_8 , 
            n4773, n4772, \REG.mem_37_6 , n4771, n4770, \REG.mem_37_4 , 
            n4769, \REG.mem_37_3 , n4768, \REG.mem_37_2 , n4767, \REG.mem_37_1 , 
            n4766, \REG.mem_37_0 , n4156, \REG.mem_26_6 , \REG.mem_25_6 , 
            \REG.mem_24_6 , \REG.mem_34_9 , n4733, \REG.mem_34_15 , 
            n4732, \REG.mem_34_14 , n4731, \REG.mem_34_13 , n4730, 
            n4729, \REG.mem_34_11 , n4728, n4727, n4726, \REG.mem_34_8 , 
            n4725, n4155, \REG.mem_2_1 , n4154, \REG.mem_24_4 , \REG.mem_25_4 , 
            \REG.mem_26_4 , n4724, \REG.mem_34_6 , \REG.mem_30_4 , \REG.mem_28_4 , 
            \REG.mem_29_4 , n4723, n4722, \REG.mem_34_4 , n4721, \REG.mem_34_3 , 
            n4720, n4719, \REG.mem_34_1 , n4718, \REG.mem_8_4 , \REG.mem_9_4 , 
            \REG.mem_10_4 , \REG.mem_11_4 , \REG.mem_14_4 , \REG.mem_15_4 , 
            \REG.mem_12_4 , \REG.mem_13_4 , \REG.mem_6_1 , \REG.mem_7_1 , 
            \REG.mem_5_1 , n4677, rp_sync1_r, \REG.mem_26_10 , \REG.mem_18_1 , 
            \REG.mem_19_1 , n4676, n4675, n4674, n4673, n4672, \REG.mem_25_10 , 
            \REG.mem_24_10 , \REG.mem_22_1 , \REG.mem_23_1 , \REG.mem_21_1 , 
            n46, n14, n4655, n4654, n4653, n4652, n4651, n4650, 
            n4649, n4648, n4647, \REG.mem_30_13 , n4646, \REG.mem_30_12 , 
            n4645, n37, n5, n4644, n4643, n4642, n4641, n4640, 
            \REG.mem_30_6 , n4639, n4638, n4637, n4636, n4635, \REG.mem_30_1 , 
            n4634, n4633, n4631, n4629, \REG.mem_18_14 , \REG.mem_19_14 , 
            n4627, n51, n4626, n4625, \REG.mem_29_13 , \REG.mem_22_14 , 
            \REG.mem_23_14 , \REG.mem_21_14 , n4624, \REG.mem_29_12 , 
            n4623, n4622, n4621, n4620, n4619, n4618, \REG.mem_29_6 , 
            n4617, n4616, n4615, n4614, n4613, \REG.mem_29_1 , n4612, 
            n4611, n4610, n4609, \REG.mem_28_13 , n19, n4608, \REG.mem_28_12 , 
            n4607, \REG.mem_18_12 , \REG.mem_19_12 , \REG.mem_22_12 , 
            \REG.mem_23_12 , n4606, n4605, n4604, n4603, n4602, 
            \REG.mem_28_6 , n4601, n4600, n4599, n4598, n4597, \REG.mem_28_1 , 
            n4596, \REG.mem_21_12 , n4579, n4578, n4577, \REG.mem_26_13 , 
            n4576, \REG.mem_26_12 , n4575, n4574, n4573, n4572, 
            n4571, \REG.mem_26_7 , n4570, n4569, n4568, n4567, \REG.mem_6_13 , 
            \REG.mem_7_13 , n4566, n4565, \REG.mem_26_1 , n4564, \REG.mem_26_0 , 
            n4563, wp_sync1_r, n4562, n4561, n4560, n4559, n4558, 
            n4557, n4556, \REG.mem_25_13 , n4555, \REG.mem_25_12 , 
            n4554, n4553, n4552, n4551, \REG.mem_5_13 , n4550, \REG.mem_25_7 , 
            n4549, n4548, n4547, n4546, n4545, n4544, \REG.mem_25_1 , 
            n4543, \REG.mem_25_0 , n4542, n4541, n4540, n4539, n4538, 
            n4537, n4536, n4535, n4534, \REG.mem_18_0 , \REG.mem_19_0 , 
            \REG.mem_22_0 , \REG.mem_23_0 , \REG.mem_21_0 , DEBUG_9_c, 
            n4533, \REG.mem_24_13 , n4532, \REG.mem_24_12 , n4531, 
            n4530, n4529, n4528, n4527, \REG.mem_24_7 , n4526, n4525, 
            n4524, n4523, n4522, n4521, \REG.mem_24_1 , n4520, \REG.mem_24_0 , 
            n4519, \REG.mem_23_15 , n4518, n4517, n4516, n4515, 
            n4514, \REG.mem_23_10 , n4513, \REG.mem_23_9 , n4512, 
            n4511, n4510, n4509, n4508, \REG.mem_23_4 , n4507, n4506, 
            n4505, n4504, n4503, \REG.mem_22_15 , n4502, n4501, 
            n4500, n4499, n4498, \REG.mem_22_10 , n4497, \REG.mem_22_9 , 
            n4496, n4495, n4494, n4493, n4492, \REG.mem_22_4 , n4491, 
            n4490, n4489, n4488, n4487, \REG.mem_21_15 , n4486, 
            n4485, n4484, n4483, n4482, \REG.mem_21_10 , n4481, 
            \REG.mem_21_9 , n4480, n4479, n4478, n4477, n4476, \REG.mem_21_4 , 
            n4475, n4474, n4473, \REG.mem_6_12 , \REG.mem_7_12 , n4472, 
            \REG.out_raw[15] , \REG.out_raw[14] , \REG.out_raw[13] , \REG.mem_5_12 , 
            \REG.out_raw[12] , \REG.out_raw[11] , \REG.out_raw[10] , n4455, 
            \REG.mem_19_15 , n4454, n4453, n4452, n4451, n4450, 
            n4449, \REG.mem_19_9 , n4448, n4447, n4446, n4445, n4444, 
            \REG.mem_19_4 , n4443, n4442, n4441, n4440, \REG.out_raw[9] , 
            \REG.out_raw[8] , n4439, \REG.mem_18_15 , \REG.out_raw[7] , 
            \REG.out_raw[6] , \REG.out_raw[5] , \REG.out_raw[4] , \REG.out_raw[3] , 
            n4438, \REG.mem_6_9 , \REG.mem_7_9 , n54, \REG.mem_5_9 , 
            n4437, n4436, n4435, n4434, n4433, \REG.mem_18_9 , n4432, 
            n4431, n4430, n4429, n4428, \REG.mem_18_4 , n4427, n4426, 
            n4425, n4424, \REG.out_raw[2] , n22, n39, \REG.mem_10_9 , 
            \REG.mem_11_9 , \REG.mem_10_13 , \REG.mem_11_13 , n7, n40, 
            \REG.mem_9_9 , \REG.mem_8_9 , \REG.mem_9_13 , \REG.mem_8_13 , 
            n8, \REG.mem_14_12 , \REG.mem_15_12 , n4391, \REG.out_raw[1] , 
            n4390, \REG.mem_13_12 , \REG.mem_12_12 , n4389, \REG.mem_15_13 , 
            n4388, n4387, n4386, \REG.mem_15_10 , n4385, \REG.mem_15_9 , 
            n4384, \REG.mem_15_8 , n4383, \REG.mem_15_7 , n4382, n4381, 
            \REG.mem_15_5 , n4380, n4379, n4378, n4377, \REG.mem_15_1 , 
            n4376, n4375, n4374, \REG.mem_6_8 , \REG.mem_7_8 , \REG.mem_5_8 , 
            \REG.mem_14_9 , \REG.mem_13_9 , \REG.mem_12_9 , \REG.mem_6_5 , 
            \REG.mem_7_5 , n4373, \REG.mem_14_13 , n4372, n4371, n4370, 
            \REG.mem_14_10 , n4369, n4368, \REG.mem_14_8 , n4367, 
            \REG.mem_14_7 , \REG.mem_5_5 , n4366, n4365, \REG.mem_14_5 , 
            n4364, n4363, n4362, n4361, \REG.mem_14_1 , n4360, n4359, 
            n4358, n4357, \REG.mem_13_13 , n4356, n4355, n4354, 
            \REG.mem_13_10 , n4353, n4352, \REG.mem_13_8 , n4351, 
            \REG.mem_13_7 , n4350, n4349, \REG.mem_13_5 , n4348, n4347, 
            n4346, n4345, \REG.mem_13_1 , n4344, n4343, n4342, n4341, 
            \REG.mem_12_13 , n4340, n4339, n4338, \REG.mem_12_10 , 
            n4337, n4336, \REG.mem_12_8 , n4335, \REG.mem_12_7 , n4334, 
            n4333, \REG.mem_12_5 , n4332, n4331, n4330, n4329, \REG.mem_12_1 , 
            n4328, n4327, n4326, n4325, n4324, n4323, n60, n4322, 
            n28, n41, n9, n4321, n4320, \REG.mem_11_8 , n4319, 
            \REG.mem_11_7 , n4318, n4317, \REG.mem_11_5 , n4316, n4315, 
            n4314, n4313, \REG.mem_11_1 , n4312, n4311, n42, n4310, 
            n4309, n4308, n10, n4307, n4306, n4305, n4304, \REG.mem_10_8 , 
            n4303, \REG.mem_10_7 , n4302, n4301, \REG.mem_10_5 , n4300, 
            n4299, n4298, n4297, \REG.mem_10_1 , n4296, n4130, n57, 
            \REG.mem_9_5 , \REG.mem_8_5 , n4288, n4287, n4286, n4285, 
            n4284, n4283, n4282, n4281, n4280, \REG.mem_9_8 , n4279, 
            \REG.mem_9_7 , n4278, n4277, n4108, n25, n4276, n43, 
            n11, n44, n12, n4275, n4274, n4273, \REG.mem_9_1 , 
            n4272, n4270, n4268, n4107, \REG.mem_8_7 , n4265, n4264, 
            n4263, n4262, n4261, n52, n4260, \REG.mem_8_8 , n4259, 
            n4258, n4257, n4256, n4255, n4254, n4253, n4252, n4251, 
            \REG.mem_8_1 , n4250, n4249, n4248, n4247, n4246, n4245, 
            \REG.mem_7_11 , n4244, n4243, n4242, n4241, n4240, n4239, 
            n4238, \REG.mem_7_4 , n4237, n4236, n4235, n4234, n4233, 
            n4232, n4231, n4230, n4229, \REG.mem_6_11 , n4228, n4227, 
            n4226, n4225, n4224, n4223, n4222, \REG.mem_6_4 , n4221, 
            n4220, n4219, n4218, n4217, n4216, n4215, n4214, n4213, 
            \REG.mem_5_11 , n4212, n4211, n4210, n4209, n4208, n4207, 
            n4206, \REG.mem_5_4 , n4205, n4204, n4203, n4202, n4103, 
            n20, n53, n4101, n21, n35, n3, n36, n55, n23, 
            n4, n47, n15, n31, n63) /* synthesis syn_module_defined=1 */ ;
    input FIFO_D6_c_6;
    output \REG.mem_42_15 ;
    output \REG.mem_43_15 ;
    input FIFO_D5_c_5;
    output \REG.mem_29_14 ;
    output \REG.mem_28_14 ;
    input FIFO_CLK_c;
    output \REG.mem_41_15 ;
    output \REG.mem_40_15 ;
    input GND_net;
    output \REG.mem_2_0 ;
    output \REG.mem_2_2 ;
    input FIFO_D4_c_4;
    output \REG.mem_18_5 ;
    output \REG.mem_19_5 ;
    input FIFO_D3_c_3;
    output \REG.mem_62_5 ;
    output \REG.mem_61_5 ;
    output \REG.mem_60_5 ;
    input FIFO_D2_c_2;
    output t_rd_fifo_en_w;
    output \REG.out_raw[0] ;
    input DEBUG_6_c;
    output \REG.mem_30_10 ;
    output \REG.mem_29_10 ;
    output \REG.mem_28_10 ;
    output \REG.mem_58_8 ;
    output \REG.mem_57_8 ;
    output \REG.mem_56_8 ;
    input FIFO_D1_c_1;
    output \REG.mem_2_14 ;
    input FIFO_D0_c_0;
    output \REG.mem_14_15 ;
    output \REG.mem_15_15 ;
    output \REG.mem_13_15 ;
    output \REG.mem_12_15 ;
    output \REG.mem_10_15 ;
    output \REG.mem_11_15 ;
    output n56;
    output \REG.mem_62_8 ;
    output \REG.mem_61_8 ;
    output \REG.mem_60_8 ;
    output \REG.mem_46_6 ;
    output \REG.mem_47_6 ;
    output n24;
    input write_to_dc32_fifo;
    input reset_all;
    output \wr_addr_nxt_c[1] ;
    output \REG.mem_45_6 ;
    output \REG.mem_44_6 ;
    output dc32_fifo_is_full;
    output \REG.mem_34_10 ;
    output \REG.mem_18_8 ;
    output \REG.mem_19_8 ;
    output \REG.mem_58_11 ;
    output \rd_grey_sync_r[0] ;
    output \REG.mem_57_11 ;
    output \REG.mem_56_11 ;
    output \REG.mem_6_14 ;
    output \REG.mem_7_14 ;
    output \REG.mem_5_14 ;
    output \REG.mem_10_12 ;
    output \REG.mem_11_12 ;
    output \REG.mem_9_12 ;
    output \REG.mem_8_12 ;
    output \REG.mem_6_10 ;
    output \REG.mem_7_10 ;
    output \REG.mem_26_9 ;
    output DEBUG_1_c;
    output \REG.mem_6_0 ;
    output \REG.mem_7_0 ;
    output \REG.mem_5_0 ;
    output \REG.mem_5_10 ;
    output \REG.mem_25_9 ;
    output \REG.mem_24_9 ;
    output \REG.mem_56_7 ;
    output \REG.mem_57_7 ;
    output \REG.mem_58_7 ;
    output \num_words_in_buffer[3] ;
    output \wr_grey_sync_r[0] ;
    output \REG.mem_10_14 ;
    output \REG.mem_11_14 ;
    output \REG.mem_9_14 ;
    output \REG.mem_8_14 ;
    output \REG.mem_14_14 ;
    output \REG.mem_15_14 ;
    output \REG.mem_13_14 ;
    output \REG.mem_12_14 ;
    output \REG.mem_38_9 ;
    output \REG.mem_39_9 ;
    output \REG.mem_37_9 ;
    output \REG.mem_34_7 ;
    output \REG.mem_42_9 ;
    output \REG.mem_43_9 ;
    output \REG.mem_10_10 ;
    output \REG.mem_11_10 ;
    output \REG.mem_9_10 ;
    output \REG.mem_8_10 ;
    output \REG.mem_41_9 ;
    output \REG.mem_40_9 ;
    output \REG.mem_9_15 ;
    output \REG.mem_8_15 ;
    output \REG.mem_18_6 ;
    output \REG.mem_19_6 ;
    output \wr_addr_nxt_c[3] ;
    input FIFO_D15_c_15;
    output \REG.mem_22_5 ;
    output \REG.mem_23_5 ;
    output \REG.mem_21_5 ;
    output \REG.mem_38_10 ;
    output \REG.mem_39_10 ;
    output \REG.mem_37_10 ;
    output \REG.mem_18_10 ;
    output \REG.mem_19_10 ;
    input FIFO_D14_c_14;
    output \REG.mem_34_12 ;
    output \REG.mem_22_6 ;
    output \REG.mem_23_6 ;
    output \REG.mem_26_14 ;
    output \REG.mem_25_14 ;
    output \REG.mem_24_14 ;
    output \REG.mem_18_13 ;
    output \REG.mem_19_13 ;
    output \REG.mem_62_7 ;
    output \REG.mem_21_6 ;
    output \REG.mem_60_7 ;
    output \REG.mem_61_7 ;
    output \REG.mem_30_14 ;
    output \REG.mem_50_3 ;
    output \REG.mem_51_3 ;
    output \REG.mem_38_12 ;
    output \REG.mem_39_12 ;
    output \REG.mem_37_12 ;
    output \REG.mem_46_8 ;
    output \REG.mem_47_8 ;
    output \REG.mem_45_8 ;
    output \REG.mem_44_8 ;
    output \REG.mem_58_10 ;
    output \REG.mem_2_3 ;
    output \REG.mem_57_10 ;
    output \REG.mem_56_10 ;
    output \REG.mem_62_2 ;
    output \REG.mem_61_2 ;
    output \REG.mem_60_2 ;
    output \REG.mem_58_15 ;
    output \REG.mem_10_0 ;
    output \REG.mem_11_0 ;
    output \REG.mem_9_0 ;
    output \REG.mem_8_0 ;
    output \REG.mem_57_15 ;
    output \REG.mem_56_15 ;
    output \REG.mem_30_0 ;
    output \REG.mem_29_0 ;
    output \REG.mem_28_0 ;
    output \REG.mem_38_7 ;
    output \REG.mem_39_7 ;
    input FIFO_D13_c_13;
    output \REG.mem_37_7 ;
    output n58;
    input FIFO_D12_c_12;
    output \REG.mem_26_5 ;
    output \REG.mem_25_5 ;
    output \REG.mem_24_5 ;
    output n50;
    output \REG.mem_46_0 ;
    output \REG.mem_47_0 ;
    output \REG.mem_6_3 ;
    output \REG.mem_7_3 ;
    output \REG.mem_5_3 ;
    output \REG.mem_45_0 ;
    output \REG.mem_44_0 ;
    output \REG.mem_50_8 ;
    output \REG.mem_51_8 ;
    output n18;
    output \REG.mem_10_3 ;
    output \REG.mem_11_3 ;
    output \REG.mem_6_2 ;
    output \REG.mem_7_2 ;
    output \REG.mem_5_2 ;
    output \REG.mem_9_3 ;
    output \REG.mem_8_3 ;
    output \wr_addr_nxt_c[5] ;
    output \REG.mem_42_12 ;
    output \REG.mem_43_12 ;
    output \REG.mem_41_12 ;
    output \REG.mem_40_12 ;
    output \REG.mem_10_2 ;
    output \REG.mem_11_2 ;
    input n4169;
    output \REG.mem_2_15 ;
    output \REG.mem_9_2 ;
    output \REG.mem_8_2 ;
    input n4168;
    input n4167;
    output \REG.mem_2_13 ;
    input n4166;
    output \REG.mem_2_12 ;
    input n4165;
    output \REG.mem_2_11 ;
    input n4164;
    output \REG.mem_2_10 ;
    output \REG.mem_6_6 ;
    output \REG.mem_7_6 ;
    input n4163;
    output \REG.mem_2_9 ;
    output \REG.mem_5_6 ;
    output \REG.mem_30_3 ;
    output \REG.mem_29_3 ;
    output \REG.mem_28_3 ;
    output \REG.mem_22_13 ;
    output \REG.mem_23_13 ;
    output \REG.mem_21_13 ;
    output \REG.mem_54_3 ;
    output \REG.mem_55_3 ;
    output \REG.mem_53_3 ;
    output \REG.mem_42_10 ;
    output \REG.mem_43_10 ;
    output \REG.mem_41_10 ;
    output \REG.mem_40_10 ;
    output \REG.mem_56_4 ;
    output \REG.mem_57_4 ;
    output \REG.mem_6_15 ;
    output \REG.mem_7_15 ;
    output \REG.mem_58_4 ;
    output \REG.mem_26_15 ;
    output \REG.mem_5_15 ;
    output \REG.mem_25_15 ;
    output \REG.mem_24_15 ;
    output \REG.mem_58_3 ;
    output \REG.mem_57_3 ;
    output \REG.mem_56_3 ;
    output \REG.mem_62_3 ;
    output \REG.mem_62_4 ;
    output \REG.mem_60_4 ;
    output \REG.mem_61_4 ;
    output \REG.mem_61_3 ;
    output \REG.mem_60_3 ;
    output \rd_addr_r[6] ;
    output \rd_addr_nxt_c_6__N_176[5] ;
    output \REG.mem_22_8 ;
    output \REG.mem_23_8 ;
    output \rd_addr_nxt_c_6__N_176[3] ;
    output \REG.mem_21_8 ;
    output \REG.mem_54_8 ;
    output \REG.mem_55_8 ;
    input FIFO_D11_c_11;
    output \REG.mem_14_3 ;
    output \REG.mem_15_3 ;
    output \REG.mem_53_8 ;
    output \REG.mem_14_2 ;
    output \REG.mem_15_2 ;
    output \REG.mem_13_3 ;
    output \REG.mem_12_3 ;
    output \REG.mem_13_2 ;
    output \REG.mem_12_2 ;
    output \REG.mem_30_5 ;
    output \REG.mem_58_13 ;
    output \REG.mem_29_5 ;
    output \REG.mem_28_5 ;
    output \REG.mem_34_5 ;
    output \REG.mem_57_13 ;
    output \REG.mem_56_13 ;
    output \REG.mem_14_6 ;
    output \REG.mem_15_6 ;
    output \REG.mem_13_6 ;
    output \REG.mem_12_6 ;
    output \REG.mem_54_9 ;
    output \REG.mem_55_9 ;
    output \REG.mem_53_9 ;
    output \REG.mem_34_0 ;
    output \REG.mem_14_0 ;
    output \REG.mem_15_0 ;
    output \REG.mem_13_0 ;
    output \REG.mem_12_0 ;
    input FIFO_D10_c_10;
    output \REG.mem_42_14 ;
    output \REG.mem_43_14 ;
    output \REG.mem_41_14 ;
    output \REG.mem_40_14 ;
    input n4162;
    output \REG.mem_2_8 ;
    input n4161;
    output \REG.mem_2_7 ;
    input FIFO_D9_c_9;
    input n5327;
    input VCC_net;
    output \fifo_data_out[0] ;
    output \REG.mem_10_11 ;
    output \REG.mem_11_11 ;
    input FIFO_D8_c_8;
    input FIFO_D7_c_7;
    output \REG.mem_9_11 ;
    output \REG.mem_8_11 ;
    output \REG.mem_62_15 ;
    output \REG.mem_62_10 ;
    input n5305;
    output \fifo_data_out[15] ;
    output \REG.mem_46_12 ;
    output \REG.mem_47_12 ;
    input n5302;
    output \fifo_data_out[14] ;
    output \REG.mem_61_10 ;
    output \REG.mem_60_10 ;
    output \REG.mem_61_15 ;
    output \REG.mem_60_15 ;
    input n5299;
    output \fifo_data_out[13] ;
    input n5296;
    output \fifo_data_out[12] ;
    input n5293;
    output \fifo_data_out[11] ;
    input n5290;
    output \fifo_data_out[10] ;
    output \REG.mem_45_12 ;
    output \REG.mem_44_12 ;
    output \REG.mem_46_15 ;
    output \REG.mem_47_15 ;
    output \REG.mem_18_3 ;
    output \REG.mem_19_3 ;
    input n5255;
    output \fifo_data_out[9] ;
    input n5252;
    output \fifo_data_out[8] ;
    input n5249;
    output \fifo_data_out[7] ;
    output \REG.mem_45_15 ;
    output \REG.mem_44_15 ;
    input n4160;
    output \REG.mem_2_6 ;
    output \REG.mem_14_11 ;
    output \REG.mem_15_11 ;
    input n4159;
    output \REG.mem_2_5 ;
    input n5236;
    output \fifo_data_out[6] ;
    input n5233;
    output \fifo_data_out[5] ;
    output \REG.mem_13_11 ;
    output \REG.mem_12_11 ;
    input n5230;
    output \fifo_data_out[4] ;
    output \wr_grey_sync_r[5] ;
    output \wr_grey_sync_r[4] ;
    output \wr_grey_sync_r[3] ;
    input n5212;
    output \fifo_data_out[3] ;
    output \REG.mem_18_2 ;
    output \REG.mem_19_2 ;
    input n5208;
    input n5207;
    output \REG.mem_62_14 ;
    input n5206;
    output \REG.mem_62_13 ;
    input n5205;
    output \REG.mem_62_12 ;
    input n5204;
    output \REG.mem_62_11 ;
    input n5203;
    input n5202;
    output \REG.mem_62_9 ;
    input n5201;
    input n5200;
    output \wr_grey_sync_r[2] ;
    output \wr_grey_sync_r[1] ;
    input n5199;
    output \REG.mem_62_6 ;
    input n5198;
    input n5197;
    input n5196;
    input n5195;
    input n5194;
    output \REG.mem_62_1 ;
    input n5193;
    output \REG.mem_62_0 ;
    input n5192;
    input n5191;
    output \REG.mem_61_14 ;
    input n5190;
    output \REG.mem_61_13 ;
    input n5189;
    output \REG.mem_61_12 ;
    input n5188;
    output \REG.mem_61_11 ;
    input n5187;
    input n5186;
    output \REG.mem_61_9 ;
    input n5185;
    input n5184;
    input n5183;
    output \REG.mem_61_6 ;
    output \REG.mem_22_3 ;
    output \REG.mem_23_3 ;
    output \REG.mem_26_8 ;
    input n5182;
    output \REG.mem_21_3 ;
    input n5181;
    input n5180;
    input n5179;
    input n5178;
    output \REG.mem_61_1 ;
    input n5177;
    output \REG.mem_61_0 ;
    input n5176;
    input n5175;
    output \REG.mem_60_14 ;
    input n5174;
    output \REG.mem_60_13 ;
    input n5173;
    output \REG.mem_60_12 ;
    input n5172;
    output \REG.mem_60_11 ;
    input n5171;
    input n5170;
    output \REG.mem_60_9 ;
    input n5169;
    input n5168;
    input n5167;
    output \REG.mem_60_6 ;
    output \REG.mem_25_8 ;
    output \REG.mem_24_8 ;
    output \REG.mem_46_9 ;
    output \REG.mem_47_9 ;
    output \REG.mem_45_9 ;
    output \REG.mem_44_9 ;
    output \REG.mem_30_7 ;
    input n5166;
    input n5165;
    input n5164;
    input n5163;
    input n5162;
    output \REG.mem_60_1 ;
    input n5161;
    output \REG.mem_60_0 ;
    output \REG.mem_29_7 ;
    output \REG.mem_28_7 ;
    input n5144;
    input n5143;
    output \REG.mem_58_14 ;
    input n5142;
    input n5141;
    output \REG.mem_58_12 ;
    input n5140;
    input n5139;
    input n5138;
    output \REG.mem_58_9 ;
    input n5137;
    input n5136;
    input n5135;
    output \REG.mem_58_6 ;
    output \REG.mem_46_10 ;
    output \REG.mem_47_10 ;
    output \REG.mem_45_10 ;
    output \REG.mem_44_10 ;
    input n5134;
    output \REG.mem_58_5 ;
    output \REG.mem_30_9 ;
    input n5133;
    input n5132;
    input n5131;
    output \REG.mem_58_2 ;
    input n5130;
    output \REG.mem_58_1 ;
    input n5129;
    output \REG.mem_58_0 ;
    input n5128;
    input n5127;
    output \REG.mem_57_14 ;
    input n5126;
    input n5125;
    output \REG.mem_57_12 ;
    input n5124;
    input n5123;
    input n5122;
    output \REG.mem_57_9 ;
    input n5121;
    input n5120;
    input n5119;
    output \REG.mem_57_6 ;
    output \REG.mem_29_9 ;
    output \REG.mem_28_9 ;
    input n5118;
    output \REG.mem_57_5 ;
    input n5117;
    input n5116;
    input n5115;
    output \REG.mem_57_2 ;
    input n5114;
    output \REG.mem_57_1 ;
    input n5113;
    output \fifo_data_out[2] ;
    input n5110;
    output \REG.mem_57_0 ;
    input n5109;
    input n5108;
    output \REG.mem_56_14 ;
    input n5107;
    input n5106;
    output \REG.mem_56_12 ;
    input n5105;
    input n5104;
    input n5103;
    output \REG.mem_56_9 ;
    output \REG.mem_10_6 ;
    output \REG.mem_11_6 ;
    input n5102;
    output \REG.mem_9_6 ;
    output \REG.mem_8_6 ;
    input n5101;
    input n5100;
    output \REG.mem_56_6 ;
    input n5099;
    output \REG.mem_56_5 ;
    input n5098;
    input n5097;
    input n5096;
    output \REG.mem_56_2 ;
    input n5095;
    output \REG.mem_56_1 ;
    input n5094;
    output \fifo_data_out[1] ;
    input n5091;
    output \REG.mem_56_0 ;
    input n5090;
    output \REG.mem_55_15 ;
    input n5089;
    output \REG.mem_55_14 ;
    input n5088;
    output \REG.mem_55_13 ;
    input n5087;
    output \REG.mem_55_12 ;
    output \REG.mem_22_2 ;
    output \REG.mem_23_2 ;
    output \REG.mem_21_2 ;
    input n5086;
    output \REG.mem_55_11 ;
    input n5085;
    output \REG.mem_55_10 ;
    input n5084;
    input n5083;
    input n5082;
    output \REG.mem_55_7 ;
    input n5081;
    output \REG.mem_55_6 ;
    input n5080;
    output \REG.mem_55_5 ;
    input n5079;
    output \REG.mem_55_4 ;
    input n5078;
    input n5077;
    output \REG.mem_55_2 ;
    input n5076;
    output \REG.mem_55_1 ;
    input n5075;
    output \REG.mem_55_0 ;
    input n5074;
    output \REG.mem_54_15 ;
    input n5073;
    output \REG.mem_54_14 ;
    input n5072;
    output \REG.mem_54_13 ;
    output \num_words_in_buffer[6] ;
    output \num_words_in_buffer[5] ;
    output \num_words_in_buffer[4] ;
    input n5071;
    output \REG.mem_54_12 ;
    input n5070;
    output \REG.mem_54_11 ;
    input n5069;
    output \REG.mem_54_10 ;
    input n5068;
    input n5067;
    input n5066;
    output \REG.mem_54_7 ;
    input n5065;
    output \REG.mem_54_6 ;
    input n5064;
    output \REG.mem_54_5 ;
    input n5063;
    output \REG.mem_54_4 ;
    input n5062;
    input n5061;
    output \REG.mem_54_2 ;
    input n5060;
    output \REG.mem_54_1 ;
    input n5057;
    output \REG.mem_54_0 ;
    input n5056;
    output \REG.mem_53_15 ;
    input n5055;
    output \REG.mem_53_14 ;
    output \REG.mem_50_12 ;
    output \REG.mem_51_12 ;
    output \REG.mem_38_5 ;
    output \REG.mem_39_5 ;
    output \REG.mem_37_5 ;
    input n5054;
    output \REG.mem_53_13 ;
    input n5053;
    output \REG.mem_53_12 ;
    input n5052;
    output \REG.mem_53_11 ;
    input n5051;
    output \REG.mem_53_10 ;
    input n5050;
    input n5049;
    input n5048;
    output \REG.mem_53_7 ;
    input n5047;
    output \REG.mem_53_6 ;
    input n5046;
    output \REG.mem_53_5 ;
    input n5045;
    output \REG.mem_53_4 ;
    input n5044;
    input n5043;
    output \REG.mem_53_2 ;
    input n5042;
    output \REG.mem_53_1 ;
    input n5041;
    output \REG.mem_53_0 ;
    output \REG.mem_26_2 ;
    output \REG.mem_18_11 ;
    output \REG.mem_19_11 ;
    output \REG.mem_25_2 ;
    output \REG.mem_24_2 ;
    input n5024;
    output \REG.mem_51_15 ;
    input n5023;
    output \REG.mem_51_14 ;
    output n26;
    output \REG.mem_26_3 ;
    output \REG.mem_25_3 ;
    output \REG.mem_24_3 ;
    output \REG.mem_40_4 ;
    output \REG.mem_41_4 ;
    input n5022;
    output \REG.mem_51_13 ;
    input n5021;
    input n5020;
    output \REG.mem_51_11 ;
    input n5019;
    output \REG.mem_51_10 ;
    input n5018;
    output \REG.mem_51_9 ;
    input n5017;
    input n5016;
    output \REG.mem_51_7 ;
    input n5015;
    output \REG.mem_51_6 ;
    input n5014;
    output \REG.mem_51_5 ;
    input n5013;
    output \REG.mem_51_4 ;
    input n5012;
    input n5011;
    output \REG.mem_51_2 ;
    input n5010;
    output \REG.mem_51_1 ;
    input n5008;
    output \REG.mem_51_0 ;
    output \REG.mem_42_4 ;
    output \REG.mem_43_4 ;
    output \REG.mem_22_11 ;
    output \REG.mem_23_11 ;
    input n5007;
    output \REG.mem_50_15 ;
    input n5006;
    output \REG.mem_50_14 ;
    input n5005;
    output \REG.mem_50_13 ;
    input n5004;
    input n5003;
    output \REG.mem_50_11 ;
    input n5002;
    output \REG.mem_50_10 ;
    input n5001;
    output \REG.mem_50_9 ;
    input n5000;
    input n4999;
    output \REG.mem_50_7 ;
    input n4998;
    output \REG.mem_50_6 ;
    input n4997;
    output \REG.mem_50_5 ;
    input n4996;
    output \REG.mem_50_4 ;
    input n4995;
    input n4994;
    output \REG.mem_50_2 ;
    input n4993;
    output \REG.mem_50_1 ;
    input n4992;
    output \REG.mem_50_0 ;
    output \REG.mem_21_11 ;
    output \rd_addr_nxt_c_6__N_176[1] ;
    input n4158;
    output \REG.mem_2_4 ;
    output \REG.mem_30_15 ;
    output \REG.mem_29_15 ;
    output \REG.mem_28_15 ;
    output \REG.mem_30_8 ;
    output \REG.mem_29_8 ;
    output \REG.mem_28_8 ;
    output \REG.mem_46_4 ;
    output \REG.mem_47_4 ;
    input n4946;
    input n4945;
    output \REG.mem_47_14 ;
    input n4944;
    output \REG.mem_47_13 ;
    output \rd_grey_sync_r[5] ;
    output \rd_grey_sync_r[4] ;
    output \rd_grey_sync_r[3] ;
    output \rd_grey_sync_r[2] ;
    output \rd_grey_sync_r[1] ;
    input n4943;
    output \REG.mem_44_4 ;
    output \REG.mem_45_4 ;
    input n4942;
    output \REG.mem_47_11 ;
    input n4941;
    input n4940;
    input n4939;
    input n4938;
    output \REG.mem_47_7 ;
    input n4937;
    input n4936;
    output \REG.mem_47_5 ;
    input n4935;
    input n4934;
    output \REG.mem_47_3 ;
    input n4933;
    output \REG.mem_47_2 ;
    input n4932;
    output \REG.mem_47_1 ;
    input n4929;
    input n4928;
    input n4927;
    output \REG.mem_46_14 ;
    output \wr_addr_r[6] ;
    input n4926;
    output \REG.mem_46_13 ;
    input n4925;
    input n4924;
    output \REG.mem_46_11 ;
    input n4923;
    input n4922;
    input n4921;
    input n4920;
    output \REG.mem_46_7 ;
    input n4919;
    input n4918;
    output \REG.mem_46_5 ;
    input n4917;
    input n4916;
    output \REG.mem_46_3 ;
    input n4915;
    output \REG.mem_46_2 ;
    input n4914;
    output \REG.mem_46_1 ;
    input n4913;
    input n4912;
    input n4911;
    output \REG.mem_45_14 ;
    output n59;
    input n4910;
    output \REG.mem_45_13 ;
    input n4909;
    input n4908;
    output \REG.mem_45_11 ;
    input n4907;
    input n4906;
    input n4905;
    input n4904;
    output \REG.mem_45_7 ;
    input n4903;
    input n4902;
    output \REG.mem_45_5 ;
    input n4901;
    input n4900;
    output \REG.mem_45_3 ;
    input n4899;
    output \REG.mem_45_2 ;
    input n4898;
    output \REG.mem_45_1 ;
    input n4897;
    input n4896;
    output n27;
    input n4895;
    output \REG.mem_44_14 ;
    input n4894;
    output \REG.mem_44_13 ;
    input n4893;
    input n4892;
    output \REG.mem_44_11 ;
    input n4891;
    input n4890;
    input n4889;
    input n4888;
    output \REG.mem_44_7 ;
    input n4887;
    input n4886;
    output \REG.mem_44_5 ;
    input n4885;
    input n4884;
    output \REG.mem_44_3 ;
    input n4883;
    output \REG.mem_44_2 ;
    input n4882;
    output \REG.mem_44_1 ;
    input n4880;
    input n4879;
    input n4878;
    input n4877;
    output \REG.mem_43_13 ;
    input n4876;
    input n4875;
    output \REG.mem_43_11 ;
    input n4874;
    input n4873;
    input n4872;
    output \REG.mem_43_8 ;
    input n4871;
    output \REG.mem_43_7 ;
    input n4870;
    output \REG.mem_43_6 ;
    input n4869;
    output \REG.mem_43_5 ;
    input n4868;
    input n4867;
    output \REG.mem_43_3 ;
    input n4866;
    output \REG.mem_43_2 ;
    input n4865;
    output \REG.mem_43_1 ;
    input n4864;
    output \REG.mem_43_0 ;
    input n4863;
    output \REG.mem_30_2 ;
    input n4862;
    input n4861;
    output \REG.mem_42_13 ;
    input n4860;
    input n4859;
    output \REG.mem_42_11 ;
    input n4858;
    input n4857;
    input n4856;
    output \REG.mem_42_8 ;
    input n4855;
    output \REG.mem_42_7 ;
    input n4854;
    output \REG.mem_42_6 ;
    input n4853;
    output \REG.mem_42_5 ;
    input n4852;
    input n4851;
    output \REG.mem_42_3 ;
    input n4850;
    output \REG.mem_42_2 ;
    input n4849;
    output \REG.mem_42_1 ;
    input n4848;
    output \REG.mem_42_0 ;
    input n4847;
    output \REG.mem_29_2 ;
    output \REG.mem_28_2 ;
    output \REG.mem_26_11 ;
    output \REG.mem_6_7 ;
    output \REG.mem_7_7 ;
    output \REG.mem_5_7 ;
    input n4846;
    input n4845;
    output \REG.mem_41_13 ;
    input n4844;
    input n4843;
    output \REG.mem_41_11 ;
    input n4842;
    input n4841;
    input n4840;
    output \REG.mem_41_8 ;
    input n4839;
    output \REG.mem_41_7 ;
    input n4838;
    output \REG.mem_41_6 ;
    input n4837;
    output \REG.mem_41_5 ;
    input n4836;
    input n4835;
    output \REG.mem_41_3 ;
    input n4834;
    output \REG.mem_41_2 ;
    input n4833;
    output \REG.mem_41_1 ;
    input n4832;
    output \REG.mem_41_0 ;
    output \REG.mem_18_7 ;
    output \REG.mem_19_7 ;
    output \REG.mem_25_11 ;
    output \REG.mem_24_11 ;
    input n4157;
    input n4831;
    input n4830;
    input n4829;
    output \REG.mem_40_13 ;
    input n4828;
    input n4827;
    output \REG.mem_40_11 ;
    input n4826;
    input n4825;
    input n4824;
    output \REG.mem_40_8 ;
    input n4823;
    output \REG.mem_40_7 ;
    input n4822;
    output \REG.mem_40_6 ;
    input n4821;
    output \REG.mem_40_5 ;
    input n4820;
    input n4819;
    output \REG.mem_40_3 ;
    input n4818;
    output \REG.mem_40_2 ;
    input n4817;
    output \REG.mem_40_1 ;
    input n4814;
    output \REG.mem_40_0 ;
    input n4813;
    output \REG.mem_39_15 ;
    input n4812;
    output \REG.mem_39_14 ;
    output \REG.mem_22_7 ;
    output \REG.mem_23_7 ;
    input n4811;
    output \REG.mem_39_13 ;
    input n4810;
    input n4809;
    output \REG.mem_39_11 ;
    output \REG.mem_21_7 ;
    input n4808;
    output \REG.mem_30_11 ;
    input n4807;
    input n4806;
    output \REG.mem_39_8 ;
    input n4805;
    input n4804;
    output \REG.mem_39_6 ;
    input n4803;
    input n4802;
    output \REG.mem_39_4 ;
    input n4801;
    output \REG.mem_39_3 ;
    input n4800;
    output \REG.mem_39_2 ;
    input n4799;
    output \REG.mem_39_1 ;
    input n4798;
    output \REG.mem_39_0 ;
    input n4797;
    output \REG.mem_38_15 ;
    input n4796;
    output \REG.mem_38_14 ;
    input n4795;
    output \REG.mem_38_13 ;
    input n4794;
    input n4793;
    output \REG.mem_38_11 ;
    output \REG.mem_29_11 ;
    output \REG.mem_28_11 ;
    input n4792;
    output \REG.mem_34_2 ;
    input n4791;
    input n4790;
    output \REG.mem_38_8 ;
    input n4789;
    input n4788;
    output \REG.mem_38_6 ;
    input n4787;
    input n4786;
    output \REG.mem_38_4 ;
    input n4785;
    output \REG.mem_38_3 ;
    input n4784;
    output \REG.mem_38_2 ;
    input n4783;
    output \REG.mem_38_1 ;
    input n4782;
    output \REG.mem_38_0 ;
    input n4781;
    output \REG.mem_37_15 ;
    input n4780;
    output \REG.mem_37_14 ;
    input n4779;
    output \REG.mem_37_13 ;
    input n4778;
    input n4777;
    output \REG.mem_37_11 ;
    input n4776;
    input n4775;
    input n4774;
    output \REG.mem_37_8 ;
    input n4773;
    input n4772;
    output \REG.mem_37_6 ;
    input n4771;
    input n4770;
    output \REG.mem_37_4 ;
    input n4769;
    output \REG.mem_37_3 ;
    input n4768;
    output \REG.mem_37_2 ;
    input n4767;
    output \REG.mem_37_1 ;
    input n4766;
    output \REG.mem_37_0 ;
    input n4156;
    output \REG.mem_26_6 ;
    output \REG.mem_25_6 ;
    output \REG.mem_24_6 ;
    output \REG.mem_34_9 ;
    input n4733;
    output \REG.mem_34_15 ;
    input n4732;
    output \REG.mem_34_14 ;
    input n4731;
    output \REG.mem_34_13 ;
    input n4730;
    input n4729;
    output \REG.mem_34_11 ;
    input n4728;
    input n4727;
    input n4726;
    output \REG.mem_34_8 ;
    input n4725;
    input n4155;
    output \REG.mem_2_1 ;
    input n4154;
    output \REG.mem_24_4 ;
    output \REG.mem_25_4 ;
    output \REG.mem_26_4 ;
    input n4724;
    output \REG.mem_34_6 ;
    output \REG.mem_30_4 ;
    output \REG.mem_28_4 ;
    output \REG.mem_29_4 ;
    input n4723;
    input n4722;
    output \REG.mem_34_4 ;
    input n4721;
    output \REG.mem_34_3 ;
    input n4720;
    input n4719;
    output \REG.mem_34_1 ;
    input n4718;
    output \REG.mem_8_4 ;
    output \REG.mem_9_4 ;
    output \REG.mem_10_4 ;
    output \REG.mem_11_4 ;
    output \REG.mem_14_4 ;
    output \REG.mem_15_4 ;
    output \REG.mem_12_4 ;
    output \REG.mem_13_4 ;
    output \REG.mem_6_1 ;
    output \REG.mem_7_1 ;
    output \REG.mem_5_1 ;
    input n4677;
    output [6:0]rp_sync1_r;
    output \REG.mem_26_10 ;
    output \REG.mem_18_1 ;
    output \REG.mem_19_1 ;
    input n4676;
    input n4675;
    input n4674;
    input n4673;
    input n4672;
    output \REG.mem_25_10 ;
    output \REG.mem_24_10 ;
    output \REG.mem_22_1 ;
    output \REG.mem_23_1 ;
    output \REG.mem_21_1 ;
    output n46;
    output n14;
    input n4655;
    input n4654;
    input n4653;
    input n4652;
    input n4651;
    input n4650;
    input n4649;
    input n4648;
    input n4647;
    output \REG.mem_30_13 ;
    input n4646;
    output \REG.mem_30_12 ;
    input n4645;
    output n37;
    output n5;
    input n4644;
    input n4643;
    input n4642;
    input n4641;
    input n4640;
    output \REG.mem_30_6 ;
    input n4639;
    input n4638;
    input n4637;
    input n4636;
    input n4635;
    output \REG.mem_30_1 ;
    input n4634;
    input n4633;
    input n4631;
    input n4629;
    output \REG.mem_18_14 ;
    output \REG.mem_19_14 ;
    input n4627;
    output n51;
    input n4626;
    input n4625;
    output \REG.mem_29_13 ;
    output \REG.mem_22_14 ;
    output \REG.mem_23_14 ;
    output \REG.mem_21_14 ;
    input n4624;
    output \REG.mem_29_12 ;
    input n4623;
    input n4622;
    input n4621;
    input n4620;
    input n4619;
    input n4618;
    output \REG.mem_29_6 ;
    input n4617;
    input n4616;
    input n4615;
    input n4614;
    input n4613;
    output \REG.mem_29_1 ;
    input n4612;
    input n4611;
    input n4610;
    input n4609;
    output \REG.mem_28_13 ;
    output n19;
    input n4608;
    output \REG.mem_28_12 ;
    input n4607;
    output \REG.mem_18_12 ;
    output \REG.mem_19_12 ;
    output \REG.mem_22_12 ;
    output \REG.mem_23_12 ;
    input n4606;
    input n4605;
    input n4604;
    input n4603;
    input n4602;
    output \REG.mem_28_6 ;
    input n4601;
    input n4600;
    input n4599;
    input n4598;
    input n4597;
    output \REG.mem_28_1 ;
    input n4596;
    output \REG.mem_21_12 ;
    input n4579;
    input n4578;
    input n4577;
    output \REG.mem_26_13 ;
    input n4576;
    output \REG.mem_26_12 ;
    input n4575;
    input n4574;
    input n4573;
    input n4572;
    input n4571;
    output \REG.mem_26_7 ;
    input n4570;
    input n4569;
    input n4568;
    input n4567;
    output \REG.mem_6_13 ;
    output \REG.mem_7_13 ;
    input n4566;
    input n4565;
    output \REG.mem_26_1 ;
    input n4564;
    output \REG.mem_26_0 ;
    input n4563;
    output [6:0]wp_sync1_r;
    input n4562;
    input n4561;
    input n4560;
    input n4559;
    input n4558;
    input n4557;
    input n4556;
    output \REG.mem_25_13 ;
    input n4555;
    output \REG.mem_25_12 ;
    input n4554;
    input n4553;
    input n4552;
    input n4551;
    output \REG.mem_5_13 ;
    input n4550;
    output \REG.mem_25_7 ;
    input n4549;
    input n4548;
    input n4547;
    input n4546;
    input n4545;
    input n4544;
    output \REG.mem_25_1 ;
    input n4543;
    output \REG.mem_25_0 ;
    input n4542;
    input n4541;
    input n4540;
    input n4539;
    input n4538;
    input n4537;
    input n4536;
    input n4535;
    input n4534;
    output \REG.mem_18_0 ;
    output \REG.mem_19_0 ;
    output \REG.mem_22_0 ;
    output \REG.mem_23_0 ;
    output \REG.mem_21_0 ;
    input DEBUG_9_c;
    input n4533;
    output \REG.mem_24_13 ;
    input n4532;
    output \REG.mem_24_12 ;
    input n4531;
    input n4530;
    input n4529;
    input n4528;
    input n4527;
    output \REG.mem_24_7 ;
    input n4526;
    input n4525;
    input n4524;
    input n4523;
    input n4522;
    input n4521;
    output \REG.mem_24_1 ;
    input n4520;
    output \REG.mem_24_0 ;
    input n4519;
    output \REG.mem_23_15 ;
    input n4518;
    input n4517;
    input n4516;
    input n4515;
    input n4514;
    output \REG.mem_23_10 ;
    input n4513;
    output \REG.mem_23_9 ;
    input n4512;
    input n4511;
    input n4510;
    input n4509;
    input n4508;
    output \REG.mem_23_4 ;
    input n4507;
    input n4506;
    input n4505;
    input n4504;
    input n4503;
    output \REG.mem_22_15 ;
    input n4502;
    input n4501;
    input n4500;
    input n4499;
    input n4498;
    output \REG.mem_22_10 ;
    input n4497;
    output \REG.mem_22_9 ;
    input n4496;
    input n4495;
    input n4494;
    input n4493;
    input n4492;
    output \REG.mem_22_4 ;
    input n4491;
    input n4490;
    input n4489;
    input n4488;
    input n4487;
    output \REG.mem_21_15 ;
    input n4486;
    input n4485;
    input n4484;
    input n4483;
    input n4482;
    output \REG.mem_21_10 ;
    input n4481;
    output \REG.mem_21_9 ;
    input n4480;
    input n4479;
    input n4478;
    input n4477;
    input n4476;
    output \REG.mem_21_4 ;
    input n4475;
    input n4474;
    input n4473;
    output \REG.mem_6_12 ;
    output \REG.mem_7_12 ;
    input n4472;
    output \REG.out_raw[15] ;
    output \REG.out_raw[14] ;
    output \REG.out_raw[13] ;
    output \REG.mem_5_12 ;
    output \REG.out_raw[12] ;
    output \REG.out_raw[11] ;
    output \REG.out_raw[10] ;
    input n4455;
    output \REG.mem_19_15 ;
    input n4454;
    input n4453;
    input n4452;
    input n4451;
    input n4450;
    input n4449;
    output \REG.mem_19_9 ;
    input n4448;
    input n4447;
    input n4446;
    input n4445;
    input n4444;
    output \REG.mem_19_4 ;
    input n4443;
    input n4442;
    input n4441;
    input n4440;
    output \REG.out_raw[9] ;
    output \REG.out_raw[8] ;
    input n4439;
    output \REG.mem_18_15 ;
    output \REG.out_raw[7] ;
    output \REG.out_raw[6] ;
    output \REG.out_raw[5] ;
    output \REG.out_raw[4] ;
    output \REG.out_raw[3] ;
    input n4438;
    output \REG.mem_6_9 ;
    output \REG.mem_7_9 ;
    output n54;
    output \REG.mem_5_9 ;
    input n4437;
    input n4436;
    input n4435;
    input n4434;
    input n4433;
    output \REG.mem_18_9 ;
    input n4432;
    input n4431;
    input n4430;
    input n4429;
    input n4428;
    output \REG.mem_18_4 ;
    input n4427;
    input n4426;
    input n4425;
    input n4424;
    output \REG.out_raw[2] ;
    output n22;
    output n39;
    output \REG.mem_10_9 ;
    output \REG.mem_11_9 ;
    output \REG.mem_10_13 ;
    output \REG.mem_11_13 ;
    output n7;
    output n40;
    output \REG.mem_9_9 ;
    output \REG.mem_8_9 ;
    output \REG.mem_9_13 ;
    output \REG.mem_8_13 ;
    output n8;
    output \REG.mem_14_12 ;
    output \REG.mem_15_12 ;
    input n4391;
    output \REG.out_raw[1] ;
    input n4390;
    output \REG.mem_13_12 ;
    output \REG.mem_12_12 ;
    input n4389;
    output \REG.mem_15_13 ;
    input n4388;
    input n4387;
    input n4386;
    output \REG.mem_15_10 ;
    input n4385;
    output \REG.mem_15_9 ;
    input n4384;
    output \REG.mem_15_8 ;
    input n4383;
    output \REG.mem_15_7 ;
    input n4382;
    input n4381;
    output \REG.mem_15_5 ;
    input n4380;
    input n4379;
    input n4378;
    input n4377;
    output \REG.mem_15_1 ;
    input n4376;
    input n4375;
    input n4374;
    output \REG.mem_6_8 ;
    output \REG.mem_7_8 ;
    output \REG.mem_5_8 ;
    output \REG.mem_14_9 ;
    output \REG.mem_13_9 ;
    output \REG.mem_12_9 ;
    output \REG.mem_6_5 ;
    output \REG.mem_7_5 ;
    input n4373;
    output \REG.mem_14_13 ;
    input n4372;
    input n4371;
    input n4370;
    output \REG.mem_14_10 ;
    input n4369;
    input n4368;
    output \REG.mem_14_8 ;
    input n4367;
    output \REG.mem_14_7 ;
    output \REG.mem_5_5 ;
    input n4366;
    input n4365;
    output \REG.mem_14_5 ;
    input n4364;
    input n4363;
    input n4362;
    input n4361;
    output \REG.mem_14_1 ;
    input n4360;
    input n4359;
    input n4358;
    input n4357;
    output \REG.mem_13_13 ;
    input n4356;
    input n4355;
    input n4354;
    output \REG.mem_13_10 ;
    input n4353;
    input n4352;
    output \REG.mem_13_8 ;
    input n4351;
    output \REG.mem_13_7 ;
    input n4350;
    input n4349;
    output \REG.mem_13_5 ;
    input n4348;
    input n4347;
    input n4346;
    input n4345;
    output \REG.mem_13_1 ;
    input n4344;
    input n4343;
    input n4342;
    input n4341;
    output \REG.mem_12_13 ;
    input n4340;
    input n4339;
    input n4338;
    output \REG.mem_12_10 ;
    input n4337;
    input n4336;
    output \REG.mem_12_8 ;
    input n4335;
    output \REG.mem_12_7 ;
    input n4334;
    input n4333;
    output \REG.mem_12_5 ;
    input n4332;
    input n4331;
    input n4330;
    input n4329;
    output \REG.mem_12_1 ;
    input n4328;
    input n4327;
    input n4326;
    input n4325;
    input n4324;
    input n4323;
    output n60;
    input n4322;
    output n28;
    output n41;
    output n9;
    input n4321;
    input n4320;
    output \REG.mem_11_8 ;
    input n4319;
    output \REG.mem_11_7 ;
    input n4318;
    input n4317;
    output \REG.mem_11_5 ;
    input n4316;
    input n4315;
    input n4314;
    input n4313;
    output \REG.mem_11_1 ;
    input n4312;
    input n4311;
    output n42;
    input n4310;
    input n4309;
    input n4308;
    output n10;
    input n4307;
    input n4306;
    input n4305;
    input n4304;
    output \REG.mem_10_8 ;
    input n4303;
    output \REG.mem_10_7 ;
    input n4302;
    input n4301;
    output \REG.mem_10_5 ;
    input n4300;
    input n4299;
    input n4298;
    input n4297;
    output \REG.mem_10_1 ;
    input n4296;
    input n4130;
    output n57;
    output \REG.mem_9_5 ;
    output \REG.mem_8_5 ;
    input n4288;
    input n4287;
    input n4286;
    input n4285;
    input n4284;
    input n4283;
    input n4282;
    input n4281;
    input n4280;
    output \REG.mem_9_8 ;
    input n4279;
    output \REG.mem_9_7 ;
    input n4278;
    input n4277;
    input n4108;
    output n25;
    input n4276;
    output n43;
    output n11;
    output n44;
    output n12;
    input n4275;
    input n4274;
    input n4273;
    output \REG.mem_9_1 ;
    input n4272;
    input n4270;
    input n4268;
    input n4107;
    output \REG.mem_8_7 ;
    input n4265;
    input n4264;
    input n4263;
    input n4262;
    input n4261;
    output n52;
    input n4260;
    output \REG.mem_8_8 ;
    input n4259;
    input n4258;
    input n4257;
    input n4256;
    input n4255;
    input n4254;
    input n4253;
    input n4252;
    input n4251;
    output \REG.mem_8_1 ;
    input n4250;
    input n4249;
    input n4248;
    input n4247;
    input n4246;
    input n4245;
    output \REG.mem_7_11 ;
    input n4244;
    input n4243;
    input n4242;
    input n4241;
    input n4240;
    input n4239;
    input n4238;
    output \REG.mem_7_4 ;
    input n4237;
    input n4236;
    input n4235;
    input n4234;
    input n4233;
    input n4232;
    input n4231;
    input n4230;
    input n4229;
    output \REG.mem_6_11 ;
    input n4228;
    input n4227;
    input n4226;
    input n4225;
    input n4224;
    input n4223;
    input n4222;
    output \REG.mem_6_4 ;
    input n4221;
    input n4220;
    input n4219;
    input n4218;
    input n4217;
    input n4216;
    input n4215;
    input n4214;
    input n4213;
    output \REG.mem_5_11 ;
    input n4212;
    input n4211;
    input n4210;
    input n4209;
    input n4208;
    input n4207;
    input n4206;
    output \REG.mem_5_4 ;
    input n4205;
    input n4204;
    input n4203;
    input n4202;
    input n4103;
    output n20;
    output n53;
    input n4101;
    output n21;
    output n35;
    output n3;
    output n36;
    output n55;
    output n23;
    output n4;
    output n47;
    output n15;
    output n31;
    output n63;
    
    wire FIFO_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=FIFO_CLK_c */ ;   // src/top.v(84[12:20])
    wire DEBUG_6_c /* synthesis SET_AS_NETWORK=DEBUG_6_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n37_c;
    wire [6:0]wr_addr_r;   // src/fifo_dc_32_lut_gen.v(194[29:38])
    
    wire \REG.mem_48_6 , n4958;
    wire [6:0]rd_addr_r;   // src/fifo_dc_32_lut_gen.v(215[29:38])
    
    wire n11568, \REG.mem_48_5 , n4957, n12222, n12225, n10929, 
        n10863, n11022, n10971, n11019, n11025, n4179, \REG.mem_3_9 , 
        n11571, n9_c, n33, \REG.mem_3_0 , n10818, n11073, n10947, 
        n12216, \REG.mem_3_2 , n11562, \REG.mem_48_4 , n4956, n11016, 
        \REG.mem_48_3 , n4955, \REG.mem_1_0 , \REG.mem_0_0 , n10821, 
        n10905, n10719, n12396, \REG.mem_1_2 , \REG.mem_0_2 , n10088, 
        n11001, n11253;
    wire [31:0]\REG.out_raw_31__N_237 ;
    
    wire \REG.mem_63_5 , n12390, n9842, \REG.mem_48_2 , n4954, n11175, 
        n11277, n10346, \REG.mem_17_5 , \REG.mem_16_5 , n10275, n10276, 
        n11010, n10267, n10266, n11013, n10182, n10183, n11004, 
        n4178, \REG.mem_3_8 , \REG.mem_31_10 , n12384, n9845, \REG.mem_59_8 , 
        n12378, n10274, n10138, n10137, n11007, n10833, n10797, 
        n12372, n9770, n10998, n9722, n9629, n10887, n10911, \REG.mem_48_1 , 
        n4953, n4177, \REG.mem_3_7 , \REG.mem_3_14 , n12366, \REG.mem_48_0 , 
        n4952, \REG.mem_1_14 , \REG.mem_0_14 , n10286, n10428, n10429, 
        n10992, n12360, n12363, n10812, n23_c, \REG.mem_63_8 , n12354, 
        n10426, n10425, n10995, n10289, n9512, n9515, n12210, 
        n10001, n10073, n11556, n10365, n10366, n10986, n9506, 
        n10827, n10357, n10356, n10989, n9935, n9890, n10520, 
        n12348;
    wire [6:0]wr_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(198[30:42])
    
    wire n4271;
    wire [6:0]wr_grey_w;   // src/fifo_dc_32_lut_gen.v(201[38:47])
    
    wire n12351, full_nxt_c_N_303, \REG.mem_35_10 , n12342, \REG.mem_33_10 , 
        \REG.mem_32_10 , n9866, n11550, n4176, \REG.mem_3_6 , \REG.mem_59_11 , 
        n12336;
    wire [6:0]rd_grey_w;   // src/fifo_dc_32_lut_gen.v(222[38:47])
    
    wire n12339, n12330, \REG.mem_4_14 , n10298, \REG.mem_17_8 , \REG.mem_16_8 , 
        n11553, n10980, n10983, n11544, \REG.mem_27_9 , n12324, 
        empty_nxt_c_N_306, n12198, \REG.mem_4_0 , n12201, \REG.mem_4_10 , 
        n10523, n9491, n9903, \REG.mem_59_7 , n9904;
    wire [6:0]rd_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(231[30:44])
    
    wire n4175, \REG.mem_3_5 , n12318, n4174, \REG.mem_3_4 , n10301, 
        n12312, n10307, n11517, n10051, n11538, n12306, \REG.mem_36_9 , 
        n9887, n10039, n11499, n11541, n12_c, n31_c, \REG.mem_35_7 , 
        n10974, n12192, n12300, n9494, n9932, \REG.mem_33_7 , \REG.mem_32_7 , 
        n10977, n10815, n12294, \REG.mem_17_6 , \REG.mem_16_6 , n10881, 
        n10803, n12186, n11793, n11769, n12288, n11805, n11829, 
        n10313, n4173, \REG.mem_3_3 , n9852, n9853, n12282, n9850, 
        n9849, n9895, n9894, n12276, n9880, n9879, n12279, n67, 
        \REG.mem_31_15 , n4671, n11655, n11589, n12270, n11781, 
        n11823, n10322, n10968, \REG.mem_20_5 , n11127, n11061, 
        n12264, n9867, n9868, n11532, n10893, n10953, n9638, n11139, 
        n11229, n9626, n9847, n9846, n11535, n12258, \REG.mem_36_10 , 
        n9911, n12252, n10323, n10324, n10962, \REG.mem_17_10 , 
        \REG.mem_16_10 , \REG.mem_31_14 , n4670, \REG.mem_35_12 , n12246, 
        n4172, \REG.mem_33_12 , \REG.mem_32_12 , n9914, n12180, \REG.mem_27_14 , 
        n12240, n10008, n10009, n11526, n12243, n10309, n10308, 
        n10965, n11367, n11307, n12234, n11427, n10334, n10956, 
        n10302, n10303, n12228, n10294, n10293, n9520, \REG.mem_63_7 , 
        n9919, n10006, n10005, n11529, \REG.mem_20_6 , n9918, n9972, 
        n9973, n11520, n9970, n9969, n11523, \REG.mem_17_13 , \REG.mem_16_13 , 
        n10959, n10950, n9942, n9943, n11514, n12174, \REG.mem_36_12 , 
        n9938, n9940, n9939, \REG.mem_49_3 , n12168, n10944, n10731, 
        n10785, \REG.mem_59_10 , n11508, n12081, n11931, n9544, 
        n12162, n10094, \REG.mem_1_3 , \REG.mem_0_3 , n9527, \REG.mem_63_2 , 
        n10938, n10217, \REG.mem_59_15 , n10932, n12156, n12159, 
        n10935, \REG.mem_31_0 , n11502, n11505, n10806, \REG.mem_31_13 , 
        n4669, \REG.mem_36_7 , n10809, n36_c, \REG.mem_31_12 , n4668, 
        \REG.mem_27_5 , n10926, n9915, n9916, n11496, n35_c, n10920, 
        n12144, \REG.mem_4_3 , n9533, n9907, n9906, n10923, n10914, 
        n12138, n9660, n9661, n11490, n9658, n9657, n9739, n9947, 
        n9968, n11484, n10097, n11433, n9964, n11478, n9949, n11415, 
        n11481, n9882, n9883, n11472, n9871, n9870, n11475, n11466, 
        \REG.mem_4_2 , n10100, \REG.mem_49_8 , \REG.mem_48_8 , n10917, 
        n4171, \REG.mem_3_1 , n9687, n9688, n11460, n9685, n9684, 
        n9742, n9536, n10103, n10112, n10908;
    wire [6:0]n1;
    
    wire n12132, n4170, n11454, n9956, n9980, n10902, n12120, 
        \REG.mem_4_6 , n9539, \REG.mem_31_3 , n11448, n9569, n10896, 
        \REG.mem_20_13 , n10899, n10013, n10037, n11442, n10004, 
        n9983, n10106, n10890, \REG.mem_52_3 , n12108, n10136, n10148, 
        n10884, n10133, n10124, n9729, n11436, \REG.mem_59_4 , n9730, 
        \REG.mem_27_15 , n12102, \REG.mem_4_15 , n11439, n12105, \REG.mem_59_3 , 
        n10878, n9690, n9691, n11430, n10317, n10318, n10872, 
        n10282, n10281, n10875, \REG.mem_63_3 , n10800, \REG.mem_63_4 , 
        n9733, n9732;
    wire [6:0]rd_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(219[30:42])
    
    wire rd_fifo_en_w, n4628, n9655, n9654, n12009, n12090, n4630, 
        n11424, n11733, n11757, n10373, \REG.mem_20_8 , n10866, 
        \REG.mem_31_11 , n4667, n12084, \REG.mem_52_8 , n10869, n11418, 
        n9548, n10202, n10794, \REG.mem_31_5 , n10860, \REG.mem_59_13 , 
        n12078, n9564, n9565, n11412, \REG.mem_35_5 , n10854, \REG.mem_33_5 , 
        \REG.mem_32_5 , n9812, n10848, n9529, n9528, n10851, n12072, 
        n11406, n10382, \REG.mem_52_9 , n11409, \REG.mem_35_0 , n11400, 
        n12066, n10199, n10190, \REG.mem_33_0 , \REG.mem_32_0 , n11403, 
        n12069, n4666, n12060, n9708, n9709, n11394, n12063, n9706, 
        n9705, n9751, n46_c, n4201, n4200, \REG.mem_4_13 , n4199, 
        \REG.mem_4_12 , n4198, \REG.mem_4_11 , n4197, n4196, \REG.mem_4_9 , 
        n4195, \REG.mem_31_9 , n4665, n12054, \REG.mem_4_8 , n4194, 
        \REG.mem_4_7 , n4193, n12057, n4192, \REG.mem_63_15 , n10842, 
        \REG.mem_4_5 , n4191, \REG.mem_63_10 , n11388, n12048, n10118, 
        n10845, n9518, n9563, n10836, n11382, n12042, n10502, 
        \REG.mem_4_4 , n4190, \REG.mem_17_3 , \REG.mem_16_3 , n9551, 
        n11385, n10172, n10181, n10830, n10169, n10154, n11376, 
        n12036, n4189, n4188, n10824, \REG.mem_4_1 , n4187, n11955, 
        n11901, n9562, n11091, n10773, n9517, n12039, n9754, n5227, 
        n5226, \REG.mem_63_14 , n5225, \REG.mem_63_13 , n5224, \REG.mem_63_12 , 
        n5223, \REG.mem_63_11 , n4186, n5222, n5221, \REG.mem_63_9 , 
        n5220, n5219, n5218, \REG.mem_63_6 , n5217, n5216, n11055, 
        n12030, n5215, n5214, n5213, \REG.mem_63_1 , n5209, \REG.mem_63_0 , 
        n11370, n12033, n38, n4140, \REG.mem_17_2 , \REG.mem_16_2 , 
        \REG.mem_0_15 , n4112, n4113, \REG.mem_0_13 , n4114, n12024, 
        \REG.mem_0_12 , n4119, \REG.mem_0_11 , n4120, \REG.mem_27_8 , 
        n11364, \REG.mem_0_10 , n4124, \REG.mem_20_3 , n9557, \REG.mem_0_9 , 
        n4125, \REG.mem_0_8 , n4126, n12018, n9977, \REG.mem_31_7 , 
        n11358, \REG.mem_0_7 , n4131, n5160, n5159, \REG.mem_59_14 , 
        n5158, n5157, \REG.mem_59_12 , n5156, n5155, n5154, \REG.mem_59_9 , 
        n5153, n5152, n5151, \REG.mem_59_6 , n11361, \REG.mem_0_6 , 
        n4132, \REG.mem_0_5 , n4133, \REG.mem_0_4 , n4134, n5150, 
        \REG.mem_59_5 , n4136, n5149, n5148, n5147, \REG.mem_59_2 , 
        n5146, \REG.mem_59_1 , n5145, \REG.mem_59_0 , n11352, n12012, 
        n4138, n10076, n10061, n12006, \REG.mem_0_1 , n4139, n11325, 
        n9874, n11346, \REG.mem_16_15 , n4407, n10752, \REG.mem_49_0 , 
        n10755, \REG.mem_16_14 , n4406, n4405, \REG.mem_16_12 , n4404, 
        n9862, n9861, n11349, n12000, \REG.mem_16_11 , n4403, n4402, 
        n9677, \REG.mem_16_9 , n4401, n8728, n4400, n11340, \REG.mem_20_2 , 
        \REG.mem_16_7 , n4399, n4398, n4397, \REG.mem_16_4 , n4396, 
        n4395, n4394, \REG.mem_16_1 , n4393, \REG.mem_16_0 , n4392, 
        \REG.mem_3_15 , n11994, n8729, n8727, n39_c, \REG.mem_17_15 , 
        n4423, \REG.mem_1_15 , n11997, \REG.mem_17_14 , n4422, n8726, 
        n11988, n10788, \REG.mem_49_12 , \REG.mem_48_12 , n4421, \REG.mem_36_5 , 
        n9824, n11247, n11334, n5040, \REG.mem_52_15 , n5039, \REG.mem_52_14 , 
        n11241, n11337, n9858, n9859, n11982, \REG.mem_17_12 , n4420, 
        n9838, n9837, n9985, \REG.mem_27_2 , n11328, \REG.mem_17_11 , 
        n4419, n4418, \REG.mem_17_9 , n4417, n11976, n10397, n5038, 
        \REG.mem_52_13 , n5037, \REG.mem_52_12 , n5036, \REG.mem_52_11 , 
        n5035, \REG.mem_52_10 , n5034, n5033, n5032, \REG.mem_52_7 , 
        n5031, \REG.mem_52_6 , n5030, \REG.mem_52_5 , n5029, \REG.mem_52_4 , 
        n5028, n5027, \REG.mem_52_2 , n5026, \REG.mem_52_1 , n5025, 
        \REG.mem_52_0 , \REG.mem_27_3 , n11970, n9702, n9703, n11322, 
        n9560, n10782, n9682, n9681, n4416, n11964;
    wire [6:0]wp_sync2_r;   // src/fifo_dc_32_lut_gen.v(221[37:47])
    
    wire n8742, \REG.mem_17_7 , n4415;
    wire [6:0]wp_sync_w;   // src/fifo_dc_32_lut_gen.v(224[30:39])
    
    wire n8741, n8725, n4414, n4413, n8740, n11316, n8724, n4990, 
        \REG.mem_49_15 , n4989, \REG.mem_49_14 , n4988, \REG.mem_49_13 , 
        n4987, n4986, \REG.mem_49_11 , n4985, \REG.mem_49_10 , n4984, 
        \REG.mem_49_9 , n4983, n4982, \REG.mem_49_7 , n4981, \REG.mem_49_6 , 
        n4980, \REG.mem_49_5 , n4979, \REG.mem_49_4 , n4978, n4977, 
        \REG.mem_49_2 , n4976, \REG.mem_49_1 , \REG.mem_1_5 , n11319, 
        \REG.mem_20_11 , n10400, n4632, \REG.mem_17_4 , n4412, n4975, 
        \REG.mem_3_13 , n11310, \REG.mem_1_13 , n11313, n4411, n4410, 
        \REG.mem_17_1 , n4409, \REG.mem_17_0 , n4408, n45, \REG.mem_20_15 , 
        n4471, \REG.mem_20_14 , n4470, n4968, \REG.mem_48_15 , n4966, 
        \REG.mem_48_14 , n4965, \REG.mem_48_13 , n4964, n4963, \REG.mem_48_11 , 
        n4962, \REG.mem_48_10 , n4961, \REG.mem_48_9 , n4960, n4959, 
        \REG.mem_48_7 , n11958, n11961, n4469, \REG.mem_20_12 , n4468, 
        \REG.mem_31_8 , n11304, n11952, n4467, \REG.mem_20_10 , n4466, 
        n8739, n8738, n8723, \REG.mem_20_9 , n4465, n8737, n8722, 
        n4664, n34, n4663, n8721, n4464, \REG.mem_20_7 , n4463, 
        n4462, n11946, \REG.mem_1_7 , n8720, \REG.mem_31_2 , n11298, 
        n8719, n4461, n9997, \REG.mem_31_6 , n4662, \REG.mem_20_4 , 
        n4460, \REG.mem_27_11 , n11940, n11292, n11295, n10406, 
        n4459, n4458, \REG.mem_20_1 , n4457, \REG.mem_20_0 , n4456, 
        n59_adj_1060, n4595, n8718, n4594, \REG.mem_27_13 , n4593, 
        n11934, n10409, \REG.mem_27_12 , n4592, n4591, \REG.mem_27_10 , 
        n4590, n4589, n11928, \REG.mem_35_2 , n11286, n4588, \REG.mem_33_2 , 
        \REG.mem_32_2 , \REG.mem_27_7 , n4587, \REG.mem_27_6 , n4586, 
        n4585, \REG.mem_27_4 , n4584, n4765, \REG.mem_36_15 , n4764, 
        \REG.mem_36_14 , n4763, \REG.mem_36_13 , n4762, n4761, \REG.mem_36_11 , 
        n4760, n4759, n4583, n4661, n4582, \REG.mem_27_1 , n4581, 
        n11922, \REG.mem_27_0 , n4580, n4758, \REG.mem_36_8 , n4757, 
        n44_c, n4756, \REG.mem_36_6 , n4755, n4754, \REG.mem_36_4 , 
        n4753, \REG.mem_36_3 , n4752, \REG.mem_36_2 , n4751, \REG.mem_36_1 , 
        n4750, \REG.mem_36_0 , n4749, \REG.mem_35_15 , n4748, \REG.mem_35_14 , 
        n4747, \REG.mem_35_13 , n4746, n4745, \REG.mem_35_11 , n4744, 
        n4743, \REG.mem_35_9 , n4742, \REG.mem_35_8 , n4741, n11280, 
        n4740, \REG.mem_35_6 , n4739, n4738, \REG.mem_35_4 , n4737, 
        \REG.mem_35_3 , n4736, n4735, \REG.mem_35_1 , n4734, n4153, 
        \REG.mem_33_9 , \REG.mem_32_9 , n11283, n4152, n4151, n4150, 
        \REG.mem_1_12 , n11916, \REG.mem_31_4 , n4717, \REG.mem_33_15 , 
        n4716, \REG.mem_33_14 , n4715, \REG.mem_33_13 , n4714, n4713, 
        \REG.mem_33_11 , n4712, n4711, n4710, \REG.mem_33_8 , n4709, 
        n4708, \REG.mem_33_6 , n11919, n11274, n11685, n10761, n11595, 
        n11910, \REG.mem_32_8 , n4707, n4706, \REG.mem_33_4 , n4705, 
        \REG.mem_33_3 , n4704, n4703, \REG.mem_33_1 , n4702, n4700, 
        \REG.mem_32_15 , n4698, \REG.mem_32_14 , n4697, \REG.mem_32_13 , 
        n4696, n4695, \REG.mem_32_11 , n4694, n4693, n4149, \REG.mem_1_11 , 
        n4185, n4148, \REG.mem_1_10 , n11268, n4184, n4692, n11271, 
        \REG.mem_1_1 , n4183, n4691, n4690, \REG.mem_32_6 , n4689, 
        n4688, \REG.mem_32_4 , n4687, \REG.mem_32_3 , n4686, n4685, 
        \REG.mem_32_1 , n4684, n10776, \REG.mem_3_12 , n4182, \REG.mem_3_11 , 
        n4181, n11262, n11904, \REG.mem_3_10 , n4180, n4660, n20_c, 
        n4659, n4658, n4657, \REG.mem_31_1 , n4656;
    wire [6:0]rp_sync2_r;   // src/fifo_dc_32_lut_gen.v(200[37:47])
    
    wire n29, n10779, n11898, n10_c, n11_c, n11892, n11223, n11256, 
        n11217, n11259, n11109, n11250, n11886, n9984, n11889, 
        n10511, n9921, n9922, n11880, n11181, n11133, n9892, n9891, 
        n9717, n9718, n11244, n10725, n9715, n9714, n11874, n11877, 
        n11868, n10022, n9696, n9697, n11238, n11862, n11865, 
        n9694, n9693, n11856, n11232, n10025, n11235, n11226, 
        n3571, n11838, n11841, n9386, n9382, n3560, n10_adj_1064, 
        n8_adj_1065, n12_adj_1066, n9378, n9478, n8847, n9669, n9670, 
        n11220, n9667, n9666, n11826, \REG.mem_1_9 , n9648, n9649, 
        n11214, n11820, n9646, n9645, \REG.mem_1_8 , n11814, n11208, 
        n10454, n11808, n4147, n11211, n4146, n11802, n11202, 
        n9927, n9928, n11796, n9925, n9924, n11196, n25_c, n11790, 
        n10722, n11190, n11193, n11784, n10463, n9827, n10746, 
        n10740, n40_adj_1070, n10716, n10743, n10734, n10737, n3567, 
        n10046, n11178, n3563, n3550, n10728, n11778, n3597, n9366, 
        n9412, n9432, n9_adj_1071, n11772, n3584, n3586, n11766, 
        n11172, n11760, n11166, n11763, n9396, n9380, n10527, 
        n9390, n9480, n11169, n9505, n11754, n9632, n9653, n11748, 
        n10512, n10513, n11160, n11079, n9542, n9514, n11742, 
        n32, n21_c, n10507, n10506, n11163, n10472, n9511, n10770, 
        n11154, n9960, n9961, n11736, n10482, n10483, n11148, 
        n9952, n9951, n10477, n10476, n11151, n11730, n11142, 
        \genblk16.rd_prev_r , n11145, n11115, n11724, n11136, n10481, 
        n4118, n4117, n10710, n9993, n9994, n11718, n9988, n9987, 
        n10054, n11130, n11712, n10487, n11706, n11709, n11700, 
        n11703, n11124, n11694, n10493, n11679, n11118, n10422, 
        n10423, n11688, n11121, n11112, n4269, n10351, n10350, 
        n11691, n11682, n4266, n11676, n11106, n11607, n11670, 
        n11100, n11673, n11094, n11097, n10749, n11664, n11625, 
        n10392, n10393, n11088, n10375, n10374, n9507, n9508, 
        n11082, n11658, n4106, \REG.mem_1_4 , n4104, n10764, n4105, 
        n11619, n4075, \REG.mem_1_6 , n4102, n10713, n11652, n4070, 
        n10432, n10431, n11085, n4074, n4092, n10029, n10030, 
        n11646, n10018, n10017, n10066, n11076, n11640, n11583, 
        n11634, n11070, n11628, n11622, n10758, n11616, n11610, 
        n11058, n10338, n10339, n11052, n9900, n9901, n11604, 
        n9877, n9876, n11598, n10327, n10326, n10335, n10336, 
        n11046, n10315, n10314, n11049, n11040, n11592, n11043, 
        n11586, n11034, n11580, n11574, n11577, n11028, n26_adj_1085, 
        n9631, n9652, n9541;
    
    SB_LUT4 i3869_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_48_6 ), .O(n4958));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3869_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9890 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_15 ), 
            .I2(\REG.mem_43_15 ), .I3(rd_addr_r[1]), .O(n11568));
    defparam rd_addr_r_0__bdd_4_lut_9890.LUT_INIT = 16'he4aa;
    SB_LUT4 i3868_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_48_5 ), .O(n4957));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3868_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12222_bdd_4_lut (.I0(n12222), .I1(\REG.mem_29_14 ), .I2(\REG.mem_28_14 ), 
            .I3(rd_addr_r[1]), .O(n12225));
    defparam n12222_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9470 (.I0(rd_addr_r[2]), .I1(n10929), 
            .I2(n10863), .I3(rd_addr_r[3]), .O(n11022));
    defparam rd_addr_r_2__bdd_4_lut_9470.LUT_INIT = 16'he4aa;
    SB_LUT4 n11022_bdd_4_lut (.I0(n11022), .I1(n10971), .I2(n11019), .I3(rd_addr_r[3]), 
            .O(n11025));
    defparam n11022_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i353_354 (.Q(\REG.mem_3_9 ), .C(FIFO_CLK_c), .D(n4179));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11568_bdd_4_lut (.I0(n11568), .I1(\REG.mem_41_15 ), .I2(\REG.mem_40_15 ), 
            .I3(rd_addr_r[1]), .O(n11571));
    defparam n11568_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i33_2_lut_3_lut (.I0(n9_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n33));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i33_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9278 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_0 ), 
            .I2(\REG.mem_3_0 ), .I3(rd_addr_r[1]), .O(n10818));
    defparam rd_addr_r_0__bdd_4_lut_9278.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10434 (.I0(rd_addr_r[2]), .I1(n11073), 
            .I2(n10947), .I3(rd_addr_r[3]), .O(n12216));
    defparam rd_addr_r_2__bdd_4_lut_10434.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9880 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_2 ), 
            .I2(\REG.mem_3_2 ), .I3(rd_addr_r[1]), .O(n11562));
    defparam rd_addr_r_0__bdd_4_lut_9880.LUT_INIT = 16'he4aa;
    SB_LUT4 i3867_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_48_4 ), .O(n4956));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3867_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9431 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_5 ), 
            .I2(\REG.mem_19_5 ), .I3(rd_addr_r[1]), .O(n11016));
    defparam rd_addr_r_0__bdd_4_lut_9431.LUT_INIT = 16'he4aa;
    SB_LUT4 i3866_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_48_3 ), .O(n4955));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3866_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n10818_bdd_4_lut (.I0(n10818), .I1(\REG.mem_1_0 ), .I2(\REG.mem_0_0 ), 
            .I3(rd_addr_r[1]), .O(n10821));
    defparam n10818_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_4__bdd_4_lut (.I0(rd_addr_r[4]), .I1(n10905), .I2(n10719), 
            .I3(rd_addr_r[5]), .O(n12396));
    defparam rd_addr_r_4__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n11562_bdd_4_lut (.I0(n11562), .I1(\REG.mem_1_2 ), .I2(\REG.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(n10088));
    defparam n11562_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12396_bdd_4_lut (.I0(n12396), .I1(n11001), .I2(n11253), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_237 [10]));
    defparam n12396_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\REG.mem_62_5 ), 
            .I2(\REG.mem_63_5 ), .I3(rd_addr_r[1]), .O(n12390));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n12390_bdd_4_lut (.I0(n12390), .I1(\REG.mem_61_5 ), .I2(\REG.mem_60_5 ), 
            .I3(rd_addr_r[1]), .O(n9842));
    defparam n12390_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3865_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_48_2 ), .O(n4954));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3865_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12216_bdd_4_lut (.I0(n12216), .I1(n11175), .I2(n11277), .I3(rd_addr_r[3]), 
            .O(n10346));
    defparam n12216_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11016_bdd_4_lut (.I0(n11016), .I1(\REG.mem_17_5 ), .I2(\REG.mem_16_5 ), 
            .I3(rd_addr_r[1]), .O(n11019));
    defparam n11016_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9446 (.I0(rd_addr_r[1]), .I1(n10275), 
            .I2(n10276), .I3(rd_addr_r[2]), .O(n11010));
    defparam rd_addr_r_1__bdd_4_lut_9446.LUT_INIT = 16'he4aa;
    SB_DFFE \REG.out_raw__i1  (.Q(\REG.out_raw[0] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [0]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_LUT4 n11010_bdd_4_lut (.I0(n11010), .I1(n10267), .I2(n10266), .I3(rd_addr_r[2]), 
            .O(n11013));
    defparam n11010_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9416 (.I0(rd_addr_r[1]), .I1(n10182), 
            .I2(n10183), .I3(rd_addr_r[2]), .O(n11004));
    defparam rd_addr_r_1__bdd_4_lut_9416.LUT_INIT = 16'he4aa;
    SB_DFF i350_351 (.Q(\REG.mem_3_8 ), .C(FIFO_CLK_c), .D(n4178));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10564 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_10 ), 
            .I2(\REG.mem_31_10 ), .I3(rd_addr_r[1]), .O(n12384));
    defparam rd_addr_r_0__bdd_4_lut_10564.LUT_INIT = 16'he4aa;
    SB_LUT4 n12384_bdd_4_lut (.I0(n12384), .I1(\REG.mem_29_10 ), .I2(\REG.mem_28_10 ), 
            .I3(rd_addr_r[1]), .O(n9845));
    defparam n12384_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10559 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_8 ), 
            .I2(\REG.mem_59_8 ), .I3(rd_addr_r[1]), .O(n12378));
    defparam rd_addr_r_0__bdd_4_lut_10559.LUT_INIT = 16'he4aa;
    SB_LUT4 n12378_bdd_4_lut (.I0(n12378), .I1(\REG.mem_57_8 ), .I2(\REG.mem_56_8 ), 
            .I3(rd_addr_r[1]), .O(n10274));
    defparam n12378_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11004_bdd_4_lut (.I0(n11004), .I1(n10138), .I2(n10137), .I3(rd_addr_r[2]), 
            .O(n11007));
    defparam n11004_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10569 (.I0(rd_addr_r[4]), .I1(n10833), 
            .I2(n10797), .I3(rd_addr_r[5]), .O(n12372));
    defparam rd_addr_r_4__bdd_4_lut_10569.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9426 (.I0(rd_addr_r[2]), .I1(n9770), 
            .I2(n9845), .I3(rd_addr_r[3]), .O(n10998));
    defparam rd_addr_r_2__bdd_4_lut_9426.LUT_INIT = 16'he4aa;
    SB_LUT4 n10998_bdd_4_lut (.I0(n10998), .I1(n9722), .I2(n9629), .I3(rd_addr_r[3]), 
            .O(n11001));
    defparam n10998_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12372_bdd_4_lut (.I0(n12372), .I1(n10887), .I2(n10911), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_237 [2]));
    defparam n12372_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3864_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_48_1 ), .O(n4953));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3864_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i347_348 (.Q(\REG.mem_3_7 ), .C(FIFO_CLK_c), .D(n4177));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10554 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_14 ), 
            .I2(\REG.mem_3_14 ), .I3(rd_addr_r[1]), .O(n12366));
    defparam rd_addr_r_0__bdd_4_lut_10554.LUT_INIT = 16'he4aa;
    SB_LUT4 i3863_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_48_0 ), .O(n4952));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3863_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12366_bdd_4_lut (.I0(n12366), .I1(\REG.mem_1_14 ), .I2(\REG.mem_0_14 ), 
            .I3(rd_addr_r[1]), .O(n10286));
    defparam n12366_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9411 (.I0(rd_addr_r[1]), .I1(n10428), 
            .I2(n10429), .I3(rd_addr_r[2]), .O(n10992));
    defparam rd_addr_r_1__bdd_4_lut_9411.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10544 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_15 ), 
            .I2(\REG.mem_15_15 ), .I3(rd_addr_r[1]), .O(n12360));
    defparam rd_addr_r_0__bdd_4_lut_10544.LUT_INIT = 16'he4aa;
    SB_LUT4 n12360_bdd_4_lut (.I0(n12360), .I1(\REG.mem_13_15 ), .I2(\REG.mem_12_15 ), 
            .I3(rd_addr_r[1]), .O(n12363));
    defparam n12360_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9259 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_15 ), 
            .I2(\REG.mem_11_15 ), .I3(rd_addr_r[1]), .O(n10812));
    defparam rd_addr_r_0__bdd_4_lut_9259.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i88_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n56));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i88_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10539 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_8 ), 
            .I2(\REG.mem_63_8 ), .I3(rd_addr_r[1]), .O(n12354));
    defparam rd_addr_r_0__bdd_4_lut_10539.LUT_INIT = 16'he4aa;
    SB_LUT4 n10992_bdd_4_lut (.I0(n10992), .I1(n10426), .I2(n10425), .I3(rd_addr_r[2]), 
            .O(n10995));
    defparam n10992_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12354_bdd_4_lut (.I0(n12354), .I1(\REG.mem_61_8 ), .I2(\REG.mem_60_8 ), 
            .I3(rd_addr_r[1]), .O(n10289));
    defparam n12354_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10549 (.I0(rd_addr_r[4]), .I1(n9512), 
            .I2(n9515), .I3(rd_addr_r[5]), .O(n12210));
    defparam rd_addr_r_4__bdd_4_lut_10549.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9925 (.I0(rd_addr_r[2]), .I1(n10001), 
            .I2(n10073), .I3(rd_addr_r[3]), .O(n11556));
    defparam rd_addr_r_2__bdd_4_lut_9925.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9401 (.I0(rd_addr_r[1]), .I1(n10365), 
            .I2(n10366), .I3(rd_addr_r[2]), .O(n10986));
    defparam rd_addr_r_1__bdd_4_lut_9401.LUT_INIT = 16'he4aa;
    SB_LUT4 n12210_bdd_4_lut (.I0(n12210), .I1(n9506), .I2(n10827), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_237 [14]));
    defparam n12210_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10986_bdd_4_lut (.I0(n10986), .I1(n10357), .I2(n10356), .I3(rd_addr_r[2]), 
            .O(n10989));
    defparam n10986_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11556_bdd_4_lut (.I0(n11556), .I1(n9935), .I2(n9890), .I3(rd_addr_r[3]), 
            .O(n10520));
    defparam n11556_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10534 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_6 ), 
            .I2(\REG.mem_47_6 ), .I3(rd_addr_r[1]), .O(n12348));
    defparam rd_addr_r_0__bdd_4_lut_10534.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i87_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n24));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i87_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i3182_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(write_to_dc32_fifo), .I3(reset_all), .O(n4271));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam i3182_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 wr_addr_nxt_c_6__I_0_128_i2_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(write_to_dc32_fifo), .I3(\wr_addr_nxt_c[1] ), .O(wr_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam wr_addr_nxt_c_6__I_0_128_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n12348_bdd_4_lut (.I0(n12348), .I1(\REG.mem_45_6 ), .I2(\REG.mem_44_6 ), 
            .I3(rd_addr_r[1]), .O(n12351));
    defparam n12348_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR full_ext_r_100 (.Q(dc32_fifo_is_full), .C(FIFO_CLK_c), .D(full_nxt_c_N_303), 
            .R(reset_all));   // src/fifo_dc_32_lut_gen.v(308[21] 324[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10529 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_10 ), 
            .I2(\REG.mem_35_10 ), .I3(rd_addr_r[1]), .O(n12342));
    defparam rd_addr_r_0__bdd_4_lut_10529.LUT_INIT = 16'he4aa;
    SB_LUT4 n12342_bdd_4_lut (.I0(n12342), .I1(\REG.mem_33_10 ), .I2(\REG.mem_32_10 ), 
            .I3(rd_addr_r[1]), .O(n9866));
    defparam n12342_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9875 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_8 ), 
            .I2(\REG.mem_19_8 ), .I3(rd_addr_r[1]), .O(n11550));
    defparam rd_addr_r_0__bdd_4_lut_9875.LUT_INIT = 16'he4aa;
    SB_DFF i344_345 (.Q(\REG.mem_3_6 ), .C(FIFO_CLK_c), .D(n4176));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10524 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_11 ), 
            .I2(\REG.mem_59_11 ), .I3(rd_addr_r[1]), .O(n12336));
    defparam rd_addr_r_0__bdd_4_lut_10524.LUT_INIT = 16'he4aa;
    SB_DFFSR rd_grey_sync_r__i0 (.Q(\rd_grey_sync_r[0] ), .C(DEBUG_6_c), 
            .D(rd_grey_w[0]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(506[21] 516[24])
    SB_LUT4 n12336_bdd_4_lut (.I0(n12336), .I1(\REG.mem_57_11 ), .I2(\REG.mem_56_11 ), 
            .I3(rd_addr_r[1]), .O(n12339));
    defparam n12336_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10519 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_14 ), 
            .I2(\REG.mem_7_14 ), .I3(rd_addr_r[1]), .O(n12330));
    defparam rd_addr_r_0__bdd_4_lut_10519.LUT_INIT = 16'he4aa;
    SB_LUT4 n12330_bdd_4_lut (.I0(n12330), .I1(\REG.mem_5_14 ), .I2(\REG.mem_4_14 ), 
            .I3(rd_addr_r[1]), .O(n10298));
    defparam n12330_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11550_bdd_4_lut (.I0(n11550), .I1(\REG.mem_17_8 ), .I2(\REG.mem_16_8 ), 
            .I3(rd_addr_r[1]), .O(n11553));
    defparam n11550_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9421 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_12 ), 
            .I2(\REG.mem_11_12 ), .I3(rd_addr_r[1]), .O(n10980));
    defparam rd_addr_r_0__bdd_4_lut_9421.LUT_INIT = 16'he4aa;
    SB_LUT4 n10980_bdd_4_lut (.I0(n10980), .I1(\REG.mem_9_12 ), .I2(\REG.mem_8_12 ), 
            .I3(rd_addr_r[1]), .O(n10983));
    defparam n10980_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9865 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_10 ), 
            .I2(\REG.mem_7_10 ), .I3(rd_addr_r[1]), .O(n11544));
    defparam rd_addr_r_0__bdd_4_lut_9865.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10514 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_9 ), 
            .I2(\REG.mem_27_9 ), .I3(rd_addr_r[1]), .O(n12324));
    defparam rd_addr_r_0__bdd_4_lut_10514.LUT_INIT = 16'he4aa;
    SB_DFFSS empty_ext_r_105 (.Q(DEBUG_1_c), .C(DEBUG_6_c), .D(empty_nxt_c_N_306), 
            .S(reset_all));   // src/fifo_dc_32_lut_gen.v(558[21] 574[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10424 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_0 ), 
            .I2(\REG.mem_7_0 ), .I3(rd_addr_r[1]), .O(n12198));
    defparam rd_addr_r_0__bdd_4_lut_10424.LUT_INIT = 16'he4aa;
    SB_LUT4 n12198_bdd_4_lut (.I0(n12198), .I1(\REG.mem_5_0 ), .I2(\REG.mem_4_0 ), 
            .I3(rd_addr_r[1]), .O(n12201));
    defparam n12198_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11544_bdd_4_lut (.I0(n11544), .I1(\REG.mem_5_10 ), .I2(\REG.mem_4_10 ), 
            .I3(rd_addr_r[1]), .O(n10523));
    defparam n11544_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12324_bdd_4_lut (.I0(n12324), .I1(\REG.mem_25_9 ), .I2(\REG.mem_24_9 ), 
            .I3(rd_addr_r[1]), .O(n9491));
    defparam n12324_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8361_3_lut (.I0(\REG.mem_56_7 ), .I1(\REG.mem_57_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9903));
    defparam i8361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8362_3_lut (.I0(\REG.mem_58_7 ), .I1(\REG.mem_59_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9904));
    defparam i8362_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR \en_rd_cnt.rd_counter_r__i1  (.Q(\num_words_in_buffer[3] ), .C(DEBUG_6_c), 
            .D(rd_sig_diff0_w[3]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(704[29] 714[32])
    SB_DFFSR wr_grey_sync_r__i0 (.Q(\wr_grey_sync_r[0] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[0]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(255[21] 265[24])
    SB_DFF i341_342 (.Q(\REG.mem_3_5 ), .C(FIFO_CLK_c), .D(n4175));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10509 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_14 ), 
            .I2(\REG.mem_11_14 ), .I3(rd_addr_r[1]), .O(n12318));
    defparam rd_addr_r_0__bdd_4_lut_10509.LUT_INIT = 16'he4aa;
    SB_DFF i338_339 (.Q(\REG.mem_3_4 ), .C(FIFO_CLK_c), .D(n4174));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n12318_bdd_4_lut (.I0(n12318), .I1(\REG.mem_9_14 ), .I2(\REG.mem_8_14 ), 
            .I3(rd_addr_r[1]), .O(n10301));
    defparam n12318_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10504 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_14 ), 
            .I2(\REG.mem_15_14 ), .I3(rd_addr_r[1]), .O(n12312));
    defparam rd_addr_r_0__bdd_4_lut_10504.LUT_INIT = 16'he4aa;
    SB_LUT4 n12312_bdd_4_lut (.I0(n12312), .I1(\REG.mem_13_14 ), .I2(\REG.mem_12_14 ), 
            .I3(rd_addr_r[1]), .O(n10307));
    defparam n12312_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_9885 (.I0(rd_addr_r[3]), .I1(n11517), 
            .I2(n10051), .I3(rd_addr_r[4]), .O(n11538));
    defparam rd_addr_r_3__bdd_4_lut_9885.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10499 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_9 ), 
            .I2(\REG.mem_39_9 ), .I3(rd_addr_r[1]), .O(n12306));
    defparam rd_addr_r_0__bdd_4_lut_10499.LUT_INIT = 16'he4aa;
    SB_LUT4 n12306_bdd_4_lut (.I0(n12306), .I1(\REG.mem_37_9 ), .I2(\REG.mem_36_9 ), 
            .I3(rd_addr_r[1]), .O(n9887));
    defparam n12306_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11538_bdd_4_lut (.I0(n11538), .I1(n10039), .I2(n11499), .I3(rd_addr_r[4]), 
            .O(n11541));
    defparam n11538_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i31_2_lut_3_lut (.I0(n12_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n31_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i31_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9391 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_7 ), 
            .I2(\REG.mem_35_7 ), .I3(rd_addr_r[1]), .O(n10974));
    defparam rd_addr_r_0__bdd_4_lut_9391.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10404 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_9 ), 
            .I2(\REG.mem_43_9 ), .I3(rd_addr_r[1]), .O(n12192));
    defparam rd_addr_r_0__bdd_4_lut_10404.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10494 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_10 ), 
            .I2(\REG.mem_11_10 ), .I3(rd_addr_r[1]), .O(n12300));
    defparam rd_addr_r_0__bdd_4_lut_10494.LUT_INIT = 16'he4aa;
    SB_LUT4 n12300_bdd_4_lut (.I0(n12300), .I1(\REG.mem_9_10 ), .I2(\REG.mem_8_10 ), 
            .I3(rd_addr_r[1]), .O(n9494));
    defparam n12300_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12192_bdd_4_lut (.I0(n12192), .I1(\REG.mem_41_9 ), .I2(\REG.mem_40_9 ), 
            .I3(rd_addr_r[1]), .O(n9932));
    defparam n12192_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10974_bdd_4_lut (.I0(n10974), .I1(\REG.mem_33_7 ), .I2(\REG.mem_32_7 ), 
            .I3(rd_addr_r[1]), .O(n10977));
    defparam n10974_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10812_bdd_4_lut (.I0(n10812), .I1(\REG.mem_9_15 ), .I2(\REG.mem_8_15 ), 
            .I3(rd_addr_r[1]), .O(n10815));
    defparam n10812_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10489 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_6 ), 
            .I2(\REG.mem_19_6 ), .I3(rd_addr_r[1]), .O(n12294));
    defparam rd_addr_r_0__bdd_4_lut_10489.LUT_INIT = 16'he4aa;
    SB_LUT4 n12294_bdd_4_lut (.I0(n12294), .I1(\REG.mem_17_6 ), .I2(\REG.mem_16_6 ), 
            .I3(rd_addr_r[1]), .O(n9890));
    defparam n12294_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10419 (.I0(rd_addr_r[2]), .I1(n10881), 
            .I2(n10803), .I3(rd_addr_r[3]), .O(n12186));
    defparam rd_addr_r_2__bdd_4_lut_10419.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut (.I0(rd_addr_r[2]), .I1(n11793), .I2(n11769), 
            .I3(rd_addr_r[3]), .O(n12288));
    defparam rd_addr_r_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n12288_bdd_4_lut (.I0(n12288), .I1(n11805), .I2(n11829), .I3(rd_addr_r[3]), 
            .O(n10313));
    defparam n12288_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i335_336 (.Q(\REG.mem_3_3 ), .C(FIFO_CLK_c), .D(n4173));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut (.I0(rd_addr_r[1]), .I1(n9852), .I2(n9853), 
            .I3(rd_addr_r[2]), .O(n12282));
    defparam rd_addr_r_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n12282_bdd_4_lut (.I0(n12282), .I1(n9850), .I2(n9849), .I3(rd_addr_r[2]), 
            .O(n9895));
    defparam n12282_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_nxt_c_6__I_0_128_i3_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(write_to_dc32_fifo), .I3(\wr_addr_nxt_c[3] ), .O(wr_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam wr_addr_nxt_c_6__I_0_128_i3_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_r_3__bdd_4_lut (.I0(rd_addr_r[3]), .I1(n9894), .I2(n9895), 
            .I3(rd_addr_r[4]), .O(n12276));
    defparam rd_addr_r_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n12276_bdd_4_lut (.I0(n12276), .I1(n9880), .I2(n9879), .I3(rd_addr_r[4]), 
            .O(n12279));
    defparam n12276_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3582_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_31_15 ), .O(n4671));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3582_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10479 (.I0(rd_addr_r[2]), .I1(n11655), 
            .I2(n11589), .I3(rd_addr_r[3]), .O(n12270));
    defparam rd_addr_r_2__bdd_4_lut_10479.LUT_INIT = 16'he4aa;
    SB_LUT4 n12270_bdd_4_lut (.I0(n12270), .I1(n11781), .I2(n11823), .I3(rd_addr_r[3]), 
            .O(n10322));
    defparam n12270_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9386 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_5 ), 
            .I2(\REG.mem_23_5 ), .I3(rd_addr_r[1]), .O(n10968));
    defparam rd_addr_r_0__bdd_4_lut_9386.LUT_INIT = 16'he4aa;
    SB_LUT4 n10968_bdd_4_lut (.I0(n10968), .I1(\REG.mem_21_5 ), .I2(\REG.mem_20_5 ), 
            .I3(rd_addr_r[1]), .O(n10971));
    defparam n10968_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10464 (.I0(rd_addr_r[2]), .I1(n11127), 
            .I2(n11061), .I3(rd_addr_r[3]), .O(n12264));
    defparam rd_addr_r_2__bdd_4_lut_10464.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9910 (.I0(rd_addr_r[1]), .I1(n9867), 
            .I2(n9868), .I3(rd_addr_r[2]), .O(n11532));
    defparam rd_addr_r_1__bdd_4_lut_9910.LUT_INIT = 16'he4aa;
    SB_LUT4 n12186_bdd_4_lut (.I0(n12186), .I1(n10893), .I2(n10953), .I3(rd_addr_r[3]), 
            .O(n9638));
    defparam n12186_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12264_bdd_4_lut (.I0(n12264), .I1(n11139), .I2(n11229), .I3(rd_addr_r[3]), 
            .O(n9626));
    defparam n12264_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11532_bdd_4_lut (.I0(n11532), .I1(n9847), .I2(n9846), .I3(rd_addr_r[2]), 
            .O(n11535));
    defparam n11532_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10484 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_10 ), 
            .I2(\REG.mem_39_10 ), .I3(rd_addr_r[1]), .O(n12258));
    defparam rd_addr_r_0__bdd_4_lut_10484.LUT_INIT = 16'he4aa;
    SB_LUT4 n12258_bdd_4_lut (.I0(n12258), .I1(\REG.mem_37_10 ), .I2(\REG.mem_36_10 ), 
            .I3(rd_addr_r[1]), .O(n9911));
    defparam n12258_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10454 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_10 ), 
            .I2(\REG.mem_19_10 ), .I3(rd_addr_r[1]), .O(n12252));
    defparam rd_addr_r_0__bdd_4_lut_10454.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9396 (.I0(rd_addr_r[1]), .I1(n10323), 
            .I2(n10324), .I3(rd_addr_r[2]), .O(n10962));
    defparam rd_addr_r_1__bdd_4_lut_9396.LUT_INIT = 16'he4aa;
    SB_LUT4 n12252_bdd_4_lut (.I0(n12252), .I1(\REG.mem_17_10 ), .I2(\REG.mem_16_10 ), 
            .I3(rd_addr_r[1]), .O(n9629));
    defparam n12252_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3581_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_31_14 ), .O(n4670));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3581_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10449 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_12 ), 
            .I2(\REG.mem_35_12 ), .I3(rd_addr_r[1]), .O(n12246));
    defparam rd_addr_r_0__bdd_4_lut_10449.LUT_INIT = 16'he4aa;
    SB_DFF i332_333 (.Q(\REG.mem_3_2 ), .C(FIFO_CLK_c), .D(n4172));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n12246_bdd_4_lut (.I0(n12246), .I1(\REG.mem_33_12 ), .I2(\REG.mem_32_12 ), 
            .I3(rd_addr_r[1]), .O(n9914));
    defparam n12246_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10399 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_6 ), 
            .I2(\REG.mem_23_6 ), .I3(rd_addr_r[1]), .O(n12180));
    defparam rd_addr_r_0__bdd_4_lut_10399.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10444 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_14 ), 
            .I2(\REG.mem_27_14 ), .I3(rd_addr_r[1]), .O(n12240));
    defparam rd_addr_r_0__bdd_4_lut_10444.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9850 (.I0(rd_addr_r[1]), .I1(n10008), 
            .I2(n10009), .I3(rd_addr_r[2]), .O(n11526));
    defparam rd_addr_r_1__bdd_4_lut_9850.LUT_INIT = 16'he4aa;
    SB_LUT4 n12240_bdd_4_lut (.I0(n12240), .I1(\REG.mem_25_14 ), .I2(\REG.mem_24_14 ), 
            .I3(rd_addr_r[1]), .O(n12243));
    defparam n12240_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10962_bdd_4_lut (.I0(n10962), .I1(n10309), .I2(n10308), .I3(rd_addr_r[2]), 
            .O(n10965));
    defparam n10962_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10459 (.I0(rd_addr_r[2]), .I1(n11367), 
            .I2(n11307), .I3(rd_addr_r[3]), .O(n12234));
    defparam rd_addr_r_2__bdd_4_lut_10459.LUT_INIT = 16'he4aa;
    SB_LUT4 n12234_bdd_4_lut (.I0(n12234), .I1(n11427), .I2(n11553), .I3(rd_addr_r[3]), 
            .O(n10334));
    defparam n12234_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9381 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_13 ), 
            .I2(\REG.mem_19_13 ), .I3(rd_addr_r[1]), .O(n10956));
    defparam rd_addr_r_0__bdd_4_lut_9381.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10474 (.I0(rd_addr_r[1]), .I1(n10302), 
            .I2(n10303), .I3(rd_addr_r[2]), .O(n12228));
    defparam rd_addr_r_1__bdd_4_lut_10474.LUT_INIT = 16'he4aa;
    SB_LUT4 n12228_bdd_4_lut (.I0(n12228), .I1(n10294), .I2(n10293), .I3(rd_addr_r[2]), 
            .O(n9520));
    defparam n12228_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8377_3_lut (.I0(\REG.mem_62_7 ), .I1(\REG.mem_63_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9919));
    defparam i8377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11526_bdd_4_lut (.I0(n11526), .I1(n10006), .I2(n10005), .I3(rd_addr_r[2]), 
            .O(n11529));
    defparam n11526_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12180_bdd_4_lut (.I0(n12180), .I1(\REG.mem_21_6 ), .I2(\REG.mem_20_6 ), 
            .I3(rd_addr_r[1]), .O(n9935));
    defparam n12180_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8376_3_lut (.I0(\REG.mem_60_7 ), .I1(\REG.mem_61_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9918));
    defparam i8376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9845 (.I0(rd_addr_r[1]), .I1(n9972), 
            .I2(n9973), .I3(rd_addr_r[2]), .O(n11520));
    defparam rd_addr_r_1__bdd_4_lut_9845.LUT_INIT = 16'he4aa;
    SB_LUT4 n11520_bdd_4_lut (.I0(n11520), .I1(n9970), .I2(n9969), .I3(rd_addr_r[2]), 
            .O(n11523));
    defparam n11520_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10956_bdd_4_lut (.I0(n10956), .I1(\REG.mem_17_13 ), .I2(\REG.mem_16_13 ), 
            .I3(rd_addr_r[1]), .O(n10959));
    defparam n10956_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_r_6__I_0_114_i4_3_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(write_to_dc32_fifo), .I3(GND_net), .O(\wr_addr_nxt_c[3] ));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam wr_addr_r_6__I_0_114_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10439 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_14 ), 
            .I2(\REG.mem_31_14 ), .I3(rd_addr_r[1]), .O(n12222));
    defparam rd_addr_r_0__bdd_4_lut_10439.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9372 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_3 ), 
            .I2(\REG.mem_51_3 ), .I3(rd_addr_r[1]), .O(n10950));
    defparam rd_addr_r_0__bdd_4_lut_9372.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9840 (.I0(rd_addr_r[1]), .I1(n9942), 
            .I2(n9943), .I3(rd_addr_r[2]), .O(n11514));
    defparam rd_addr_r_1__bdd_4_lut_9840.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10389 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_12 ), 
            .I2(\REG.mem_39_12 ), .I3(rd_addr_r[1]), .O(n12174));
    defparam rd_addr_r_0__bdd_4_lut_10389.LUT_INIT = 16'he4aa;
    SB_LUT4 n12174_bdd_4_lut (.I0(n12174), .I1(\REG.mem_37_12 ), .I2(\REG.mem_36_12 ), 
            .I3(rd_addr_r[1]), .O(n9938));
    defparam n12174_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11514_bdd_4_lut (.I0(n11514), .I1(n9940), .I2(n9939), .I3(rd_addr_r[2]), 
            .O(n11517));
    defparam n11514_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10950_bdd_4_lut (.I0(n10950), .I1(\REG.mem_49_3 ), .I2(\REG.mem_48_3 ), 
            .I3(rd_addr_r[1]), .O(n10953));
    defparam n10950_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10414 (.I0(rd_addr_r[4]), .I1(n9626), 
            .I2(n9638), .I3(rd_addr_r[5]), .O(n12168));
    defparam rd_addr_r_4__bdd_4_lut_10414.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9367 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_8 ), 
            .I2(\REG.mem_47_8 ), .I3(rd_addr_r[1]), .O(n10944));
    defparam rd_addr_r_0__bdd_4_lut_9367.LUT_INIT = 16'he4aa;
    SB_LUT4 n12168_bdd_4_lut (.I0(n12168), .I1(n10731), .I2(n10785), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_237 [3]));
    defparam n12168_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10944_bdd_4_lut (.I0(n10944), .I1(\REG.mem_45_8 ), .I2(\REG.mem_44_8 ), 
            .I3(rd_addr_r[1]), .O(n10947));
    defparam n10944_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9860 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_10 ), 
            .I2(\REG.mem_59_10 ), .I3(rd_addr_r[1]), .O(n11508));
    defparam rd_addr_r_0__bdd_4_lut_9860.LUT_INIT = 16'he4aa;
    SB_LUT4 i8002_3_lut (.I0(n12081), .I1(n11931), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9544));
    defparam i8002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10384 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_3 ), 
            .I2(\REG.mem_3_3 ), .I3(rd_addr_r[1]), .O(n12162));
    defparam rd_addr_r_0__bdd_4_lut_10384.LUT_INIT = 16'he4aa;
    SB_LUT4 n11508_bdd_4_lut (.I0(n11508), .I1(\REG.mem_57_10 ), .I2(\REG.mem_56_10 ), 
            .I3(rd_addr_r[1]), .O(n10094));
    defparam n11508_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12162_bdd_4_lut (.I0(n12162), .I1(\REG.mem_1_3 ), .I2(\REG.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(n9527));
    defparam n12162_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9362 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_2 ), 
            .I2(\REG.mem_63_2 ), .I3(rd_addr_r[1]), .O(n10938));
    defparam rd_addr_r_0__bdd_4_lut_9362.LUT_INIT = 16'he4aa;
    SB_LUT4 n10938_bdd_4_lut (.I0(n10938), .I1(\REG.mem_61_2 ), .I2(\REG.mem_60_2 ), 
            .I3(rd_addr_r[1]), .O(n10217));
    defparam n10938_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9357 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_15 ), 
            .I2(\REG.mem_59_15 ), .I3(rd_addr_r[1]), .O(n10932));
    defparam rd_addr_r_0__bdd_4_lut_9357.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10374 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_0 ), 
            .I2(\REG.mem_11_0 ), .I3(rd_addr_r[1]), .O(n12156));
    defparam rd_addr_r_0__bdd_4_lut_10374.LUT_INIT = 16'he4aa;
    SB_LUT4 n12156_bdd_4_lut (.I0(n12156), .I1(\REG.mem_9_0 ), .I2(\REG.mem_8_0 ), 
            .I3(rd_addr_r[1]), .O(n12159));
    defparam n12156_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10932_bdd_4_lut (.I0(n10932), .I1(\REG.mem_57_15 ), .I2(\REG.mem_56_15 ), 
            .I3(rd_addr_r[1]), .O(n10935));
    defparam n10932_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9830 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_0 ), 
            .I2(\REG.mem_31_0 ), .I3(rd_addr_r[1]), .O(n11502));
    defparam rd_addr_r_0__bdd_4_lut_9830.LUT_INIT = 16'he4aa;
    SB_LUT4 n11502_bdd_4_lut (.I0(n11502), .I1(\REG.mem_29_0 ), .I2(\REG.mem_28_0 ), 
            .I3(rd_addr_r[1]), .O(n11505));
    defparam n11502_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9254 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_7 ), 
            .I2(\REG.mem_39_7 ), .I3(rd_addr_r[1]), .O(n10806));
    defparam rd_addr_r_0__bdd_4_lut_9254.LUT_INIT = 16'he4aa;
    SB_LUT4 i3580_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_31_13 ), .O(n4669));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3580_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n10806_bdd_4_lut (.I0(n10806), .I1(\REG.mem_37_7 ), .I2(\REG.mem_36_7 ), 
            .I3(rd_addr_r[1]), .O(n10809));
    defparam n10806_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i84_2_lut_3_lut (.I0(n36_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n58));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i84_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i3579_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_31_12 ), .O(n4668));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3579_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9352 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_5 ), 
            .I2(\REG.mem_27_5 ), .I3(rd_addr_r[1]), .O(n10926));
    defparam rd_addr_r_0__bdd_4_lut_9352.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9835 (.I0(rd_addr_r[1]), .I1(n9915), 
            .I2(n9916), .I3(rd_addr_r[2]), .O(n11496));
    defparam rd_addr_r_1__bdd_4_lut_9835.LUT_INIT = 16'he4aa;
    SB_LUT4 n10926_bdd_4_lut (.I0(n10926), .I1(\REG.mem_25_5 ), .I2(\REG.mem_24_5 ), 
            .I3(rd_addr_r[1]), .O(n10929));
    defparam n10926_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i100_2_lut_3_lut (.I0(n35_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n50));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i100_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9347 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_0 ), 
            .I2(\REG.mem_47_0 ), .I3(rd_addr_r[1]), .O(n10920));
    defparam rd_addr_r_0__bdd_4_lut_9347.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10369 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_3 ), 
            .I2(\REG.mem_7_3 ), .I3(rd_addr_r[1]), .O(n12144));
    defparam rd_addr_r_0__bdd_4_lut_10369.LUT_INIT = 16'he4aa;
    SB_LUT4 n12144_bdd_4_lut (.I0(n12144), .I1(\REG.mem_5_3 ), .I2(\REG.mem_4_3 ), 
            .I3(rd_addr_r[1]), .O(n9533));
    defparam n12144_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11496_bdd_4_lut (.I0(n11496), .I1(n9907), .I2(n9906), .I3(rd_addr_r[2]), 
            .O(n11499));
    defparam n11496_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10920_bdd_4_lut (.I0(n10920), .I1(\REG.mem_45_0 ), .I2(\REG.mem_44_0 ), 
            .I3(rd_addr_r[1]), .O(n10923));
    defparam n10920_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9342 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_8 ), 
            .I2(\REG.mem_51_8 ), .I3(rd_addr_r[1]), .O(n10914));
    defparam rd_addr_r_0__bdd_4_lut_9342.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i99_2_lut_3_lut (.I0(n35_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n18));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i99_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10359 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_3 ), 
            .I2(\REG.mem_11_3 ), .I3(rd_addr_r[1]), .O(n12138));
    defparam rd_addr_r_0__bdd_4_lut_10359.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9820 (.I0(rd_addr_r[1]), .I1(n9660), 
            .I2(n9661), .I3(rd_addr_r[2]), .O(n11490));
    defparam rd_addr_r_1__bdd_4_lut_9820.LUT_INIT = 16'he4aa;
    SB_LUT4 n11490_bdd_4_lut (.I0(n11490), .I1(n9658), .I2(n9657), .I3(rd_addr_r[2]), 
            .O(n9739));
    defparam n11490_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9870 (.I0(rd_addr_r[2]), .I1(n9947), 
            .I2(n9968), .I3(rd_addr_r[3]), .O(n11484));
    defparam rd_addr_r_2__bdd_4_lut_9870.LUT_INIT = 16'he4aa;
    SB_LUT4 n11484_bdd_4_lut (.I0(n11484), .I1(n9938), .I2(n9914), .I3(rd_addr_r[3]), 
            .O(n10097));
    defparam n11484_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_9855 (.I0(rd_addr_r[3]), .I1(n11433), 
            .I2(n9964), .I3(rd_addr_r[4]), .O(n11478));
    defparam rd_addr_r_3__bdd_4_lut_9855.LUT_INIT = 16'he4aa;
    SB_LUT4 n11478_bdd_4_lut (.I0(n11478), .I1(n9949), .I2(n11415), .I3(rd_addr_r[4]), 
            .O(n11481));
    defparam n11478_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9815 (.I0(rd_addr_r[1]), .I1(n9882), 
            .I2(n9883), .I3(rd_addr_r[2]), .O(n11472));
    defparam rd_addr_r_1__bdd_4_lut_9815.LUT_INIT = 16'he4aa;
    SB_LUT4 n11472_bdd_4_lut (.I0(n11472), .I1(n9871), .I2(n9870), .I3(rd_addr_r[2]), 
            .O(n11475));
    defparam n11472_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9825 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_2 ), 
            .I2(\REG.mem_7_2 ), .I3(rd_addr_r[1]), .O(n11466));
    defparam rd_addr_r_0__bdd_4_lut_9825.LUT_INIT = 16'he4aa;
    SB_LUT4 n11466_bdd_4_lut (.I0(n11466), .I1(\REG.mem_5_2 ), .I2(\REG.mem_4_2 ), 
            .I3(rd_addr_r[1]), .O(n10100));
    defparam n11466_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10914_bdd_4_lut (.I0(n10914), .I1(\REG.mem_49_8 ), .I2(\REG.mem_48_8 ), 
            .I3(rd_addr_r[1]), .O(n10917));
    defparam n10914_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i329_330 (.Q(\REG.mem_3_1 ), .C(FIFO_CLK_c), .D(n4171));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9800 (.I0(rd_addr_r[1]), .I1(n9687), 
            .I2(n9688), .I3(rd_addr_r[2]), .O(n11460));
    defparam rd_addr_r_1__bdd_4_lut_9800.LUT_INIT = 16'he4aa;
    SB_LUT4 n11460_bdd_4_lut (.I0(n11460), .I1(n9685), .I2(n9684), .I3(rd_addr_r[2]), 
            .O(n9742));
    defparam n11460_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12138_bdd_4_lut (.I0(n12138), .I1(\REG.mem_9_3 ), .I2(\REG.mem_8_3 ), 
            .I3(rd_addr_r[1]), .O(n9536));
    defparam n12138_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9406 (.I0(rd_addr_r[2]), .I1(n10103), 
            .I2(n10112), .I3(rd_addr_r[3]), .O(n10908));
    defparam rd_addr_r_2__bdd_4_lut_9406.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_r_6__I_0_114_i6_3_lut (.I0(wr_addr_r[5]), .I1(wr_addr_p1_w[5]), 
            .I2(write_to_dc32_fifo), .I3(GND_net), .O(\wr_addr_nxt_c[5] ));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam wr_addr_r_6__I_0_114_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n10908_bdd_4_lut (.I0(n10908), .I1(n10100), .I2(n10088), .I3(rd_addr_r[3]), 
            .O(n10911));
    defparam n10908_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_6__I_0_127_inv_0_i1_1_lut (.I0(rd_addr_r[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // src/fifo_dc_32_lut_gen.v(231[47:78])
    defparam wp_sync2_r_6__I_0_127_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10354 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_12 ), 
            .I2(\REG.mem_43_12 ), .I3(rd_addr_r[1]), .O(n12132));
    defparam rd_addr_r_0__bdd_4_lut_10354.LUT_INIT = 16'he4aa;
    SB_LUT4 n12132_bdd_4_lut (.I0(n12132), .I1(\REG.mem_41_12 ), .I2(\REG.mem_40_12 ), 
            .I3(rd_addr_r[1]), .O(n9947));
    defparam n12132_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i326_327 (.Q(\REG.mem_3_0 ), .C(FIFO_CLK_c), .D(n4170));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9795 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_2 ), 
            .I2(\REG.mem_11_2 ), .I3(rd_addr_r[1]), .O(n11454));
    defparam rd_addr_r_0__bdd_4_lut_9795.LUT_INIT = 16'he4aa;
    SB_DFF i275_276 (.Q(\REG.mem_2_15 ), .C(FIFO_CLK_c), .D(n4169));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11454_bdd_4_lut (.I0(n11454), .I1(\REG.mem_9_2 ), .I2(\REG.mem_8_2 ), 
            .I3(rd_addr_r[1]), .O(n10103));
    defparam n11454_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i272_273 (.Q(\REG.mem_2_14 ), .C(FIFO_CLK_c), .D(n4168));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i269_270 (.Q(\REG.mem_2_13 ), .C(FIFO_CLK_c), .D(n4167));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i266_267 (.Q(\REG.mem_2_12 ), .C(FIFO_CLK_c), .D(n4166));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i263_264 (.Q(\REG.mem_2_11 ), .C(FIFO_CLK_c), .D(n4165));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i260_261 (.Q(\REG.mem_2_10 ), .C(FIFO_CLK_c), .D(n4164));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9332 (.I0(rd_addr_r[2]), .I1(n9956), 
            .I2(n9980), .I3(rd_addr_r[3]), .O(n10902));
    defparam rd_addr_r_2__bdd_4_lut_9332.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10349 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_6 ), 
            .I2(\REG.mem_7_6 ), .I3(rd_addr_r[1]), .O(n12120));
    defparam rd_addr_r_0__bdd_4_lut_10349.LUT_INIT = 16'he4aa;
    SB_DFF i257_258 (.Q(\REG.mem_2_9 ), .C(FIFO_CLK_c), .D(n4163));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n10902_bdd_4_lut (.I0(n10902), .I1(n9911), .I2(n9866), .I3(rd_addr_r[3]), 
            .O(n10905));
    defparam n10902_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12120_bdd_4_lut (.I0(n12120), .I1(\REG.mem_5_6 ), .I2(\REG.mem_4_6 ), 
            .I3(rd_addr_r[1]), .O(n9539));
    defparam n12120_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9785 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_3 ), 
            .I2(\REG.mem_31_3 ), .I3(rd_addr_r[1]), .O(n11448));
    defparam rd_addr_r_0__bdd_4_lut_9785.LUT_INIT = 16'he4aa;
    SB_LUT4 n11448_bdd_4_lut (.I0(n11448), .I1(\REG.mem_29_3 ), .I2(\REG.mem_28_3 ), 
            .I3(rd_addr_r[1]), .O(n9569));
    defparam n11448_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9337 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_13 ), 
            .I2(\REG.mem_23_13 ), .I3(rd_addr_r[1]), .O(n10896));
    defparam rd_addr_r_0__bdd_4_lut_9337.LUT_INIT = 16'he4aa;
    SB_LUT4 n10896_bdd_4_lut (.I0(n10896), .I1(\REG.mem_21_13 ), .I2(\REG.mem_20_13 ), 
            .I3(rd_addr_r[1]), .O(n10899));
    defparam n10896_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9810 (.I0(rd_addr_r[2]), .I1(n10013), 
            .I2(n10037), .I3(rd_addr_r[3]), .O(n11442));
    defparam rd_addr_r_2__bdd_4_lut_9810.LUT_INIT = 16'he4aa;
    SB_LUT4 n11442_bdd_4_lut (.I0(n11442), .I1(n10004), .I2(n9983), .I3(rd_addr_r[3]), 
            .O(n10106));
    defparam n11442_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9322 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_3 ), 
            .I2(\REG.mem_55_3 ), .I3(rd_addr_r[1]), .O(n10890));
    defparam rd_addr_r_0__bdd_4_lut_9322.LUT_INIT = 16'he4aa;
    SB_LUT4 n10890_bdd_4_lut (.I0(n10890), .I1(\REG.mem_53_3 ), .I2(\REG.mem_52_3 ), 
            .I3(rd_addr_r[1]), .O(n10893));
    defparam n10890_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10339 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_10 ), 
            .I2(\REG.mem_43_10 ), .I3(rd_addr_r[1]), .O(n12108));
    defparam rd_addr_r_0__bdd_4_lut_10339.LUT_INIT = 16'he4aa;
    SB_LUT4 wp_sync2_r_6__I_0_127_inv_0_i2_1_lut (.I0(rd_addr_r[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // src/fifo_dc_32_lut_gen.v(231[47:78])
    defparam wp_sync2_r_6__I_0_127_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9327 (.I0(rd_addr_r[2]), .I1(n10136), 
            .I2(n10148), .I3(rd_addr_r[3]), .O(n10884));
    defparam rd_addr_r_2__bdd_4_lut_9327.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i67_2_lut (.I0(n35_c), .I1(wr_addr_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n67));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n10884_bdd_4_lut (.I0(n10884), .I1(n10133), .I2(n10124), .I3(rd_addr_r[3]), 
            .O(n10887));
    defparam n10884_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12108_bdd_4_lut (.I0(n12108), .I1(\REG.mem_41_10 ), .I2(\REG.mem_40_10 ), 
            .I3(rd_addr_r[1]), .O(n9956));
    defparam n12108_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_6__I_0_127_inv_0_i3_1_lut (.I0(rd_addr_r[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // src/fifo_dc_32_lut_gen.v(231[47:78])
    defparam wp_sync2_r_6__I_0_127_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8187_3_lut (.I0(\REG.mem_56_4 ), .I1(\REG.mem_57_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9729));
    defparam i8187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9780 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_15 ), 
            .I2(\REG.mem_7_15 ), .I3(rd_addr_r[1]), .O(n11436));
    defparam rd_addr_r_0__bdd_4_lut_9780.LUT_INIT = 16'he4aa;
    SB_LUT4 i8188_3_lut (.I0(\REG.mem_58_4 ), .I1(\REG.mem_59_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9730));
    defparam i8188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10329 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_15 ), 
            .I2(\REG.mem_27_15 ), .I3(rd_addr_r[1]), .O(n12102));
    defparam rd_addr_r_0__bdd_4_lut_10329.LUT_INIT = 16'he4aa;
    SB_LUT4 n11436_bdd_4_lut (.I0(n11436), .I1(\REG.mem_5_15 ), .I2(\REG.mem_4_15 ), 
            .I3(rd_addr_r[1]), .O(n11439));
    defparam n11436_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12102_bdd_4_lut (.I0(n12102), .I1(\REG.mem_25_15 ), .I2(\REG.mem_24_15 ), 
            .I3(rd_addr_r[1]), .O(n12105));
    defparam n12102_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9317 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_3 ), 
            .I2(\REG.mem_59_3 ), .I3(rd_addr_r[1]), .O(n10878));
    defparam rd_addr_r_0__bdd_4_lut_9317.LUT_INIT = 16'he4aa;
    SB_LUT4 n10878_bdd_4_lut (.I0(n10878), .I1(\REG.mem_57_3 ), .I2(\REG.mem_56_3 ), 
            .I3(rd_addr_r[1]), .O(n10881));
    defparam n10878_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9790 (.I0(rd_addr_r[1]), .I1(n9690), 
            .I2(n9691), .I3(rd_addr_r[2]), .O(n11430));
    defparam rd_addr_r_1__bdd_4_lut_9790.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_9475 (.I0(rd_addr_r[3]), .I1(n10317), 
            .I2(n10318), .I3(rd_addr_r[4]), .O(n10872));
    defparam rd_addr_r_3__bdd_4_lut_9475.LUT_INIT = 16'he4aa;
    SB_LUT4 n10872_bdd_4_lut (.I0(n10872), .I1(n10282), .I2(n10281), .I3(rd_addr_r[4]), 
            .O(n10875));
    defparam n10872_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9249 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_3 ), 
            .I2(\REG.mem_63_3 ), .I3(rd_addr_r[1]), .O(n10800));
    defparam rd_addr_r_0__bdd_4_lut_9249.LUT_INIT = 16'he4aa;
    SB_LUT4 i8191_3_lut (.I0(\REG.mem_62_4 ), .I1(\REG.mem_63_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9733));
    defparam i8191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8190_3_lut (.I0(\REG.mem_60_4 ), .I1(\REG.mem_61_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9732));
    defparam i8190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n10800_bdd_4_lut (.I0(n10800), .I1(\REG.mem_61_3 ), .I2(\REG.mem_60_3 ), 
            .I3(rd_addr_r[1]), .O(n10803));
    defparam n10800_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3539_2_lut_4_lut (.I0(\rd_addr_r[6] ), .I1(rd_addr_p1_w[6]), 
            .I2(rd_fifo_en_w), .I3(reset_all), .O(n4628));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam i3539_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 n11430_bdd_4_lut (.I0(n11430), .I1(n9655), .I2(n9654), .I3(rd_addr_r[2]), 
            .O(n11433));
    defparam n11430_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_nxt_c_6__I_0_130_i6_2_lut_4_lut (.I0(\rd_addr_r[6] ), 
            .I1(rd_addr_p1_w[6]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_176[5] ), 
            .O(rd_grey_w[5]));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam rd_addr_nxt_c_6__I_0_130_i6_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10394 (.I0(rd_addr_r[2]), .I1(n9491), 
            .I2(n12009), .I3(rd_addr_r[3]), .O(n12090));
    defparam rd_addr_r_2__bdd_4_lut_10394.LUT_INIT = 16'he4aa;
    SB_LUT4 i3541_2_lut_4_lut (.I0(rd_addr_r[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(reset_all), .O(n4630));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam i3541_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9770 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_8 ), 
            .I2(\REG.mem_23_8 ), .I3(rd_addr_r[1]), .O(n11424));
    defparam rd_addr_r_0__bdd_4_lut_9770.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_6__I_0_130_i4_2_lut_4_lut (.I0(rd_addr_r[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_176[3] ), .O(rd_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam rd_addr_nxt_c_6__I_0_130_i4_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n12090_bdd_4_lut (.I0(n12090), .I1(n11733), .I2(n11757), .I3(rd_addr_r[3]), 
            .O(n10373));
    defparam n12090_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11424_bdd_4_lut (.I0(n11424), .I1(\REG.mem_21_8 ), .I2(\REG.mem_20_8 ), 
            .I3(rd_addr_r[1]), .O(n11427));
    defparam n11424_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9307 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_8 ), 
            .I2(\REG.mem_55_8 ), .I3(rd_addr_r[1]), .O(n10866));
    defparam rd_addr_r_0__bdd_4_lut_9307.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_6__I_0_130_i5_2_lut_4_lut (.I0(rd_addr_r[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_176[5] ), .O(rd_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam rd_addr_nxt_c_6__I_0_130_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i3578_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_31_11 ), .O(n4667));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3578_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10324 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_3 ), 
            .I2(\REG.mem_15_3 ), .I3(rd_addr_r[1]), .O(n12084));
    defparam rd_addr_r_0__bdd_4_lut_10324.LUT_INIT = 16'he4aa;
    SB_LUT4 n10866_bdd_4_lut (.I0(n10866), .I1(\REG.mem_53_8 ), .I2(\REG.mem_52_8 ), 
            .I3(rd_addr_r[1]), .O(n10869));
    defparam n10866_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9760 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_2 ), 
            .I2(\REG.mem_15_2 ), .I3(rd_addr_r[1]), .O(n11418));
    defparam rd_addr_r_0__bdd_4_lut_9760.LUT_INIT = 16'he4aa;
    SB_LUT4 n12084_bdd_4_lut (.I0(n12084), .I1(\REG.mem_13_3 ), .I2(\REG.mem_12_3 ), 
            .I3(rd_addr_r[1]), .O(n9548));
    defparam n12084_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9264 (.I0(rd_addr_r[2]), .I1(n10202), 
            .I2(n10217), .I3(rd_addr_r[3]), .O(n10794));
    defparam rd_addr_r_2__bdd_4_lut_9264.LUT_INIT = 16'he4aa;
    SB_LUT4 n11418_bdd_4_lut (.I0(n11418), .I1(\REG.mem_13_2 ), .I2(\REG.mem_12_2 ), 
            .I3(rd_addr_r[1]), .O(n10112));
    defparam n11418_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9298 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_5 ), 
            .I2(\REG.mem_31_5 ), .I3(rd_addr_r[1]), .O(n10860));
    defparam rd_addr_r_0__bdd_4_lut_9298.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10309 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_13 ), 
            .I2(\REG.mem_59_13 ), .I3(rd_addr_r[1]), .O(n12078));
    defparam rd_addr_r_0__bdd_4_lut_10309.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9765 (.I0(rd_addr_r[1]), .I1(n9564), 
            .I2(n9565), .I3(rd_addr_r[2]), .O(n11412));
    defparam rd_addr_r_1__bdd_4_lut_9765.LUT_INIT = 16'he4aa;
    SB_LUT4 n10860_bdd_4_lut (.I0(n10860), .I1(\REG.mem_29_5 ), .I2(\REG.mem_28_5 ), 
            .I3(rd_addr_r[1]), .O(n10863));
    defparam n10860_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9293 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_5 ), 
            .I2(\REG.mem_35_5 ), .I3(rd_addr_r[1]), .O(n10854));
    defparam rd_addr_r_0__bdd_4_lut_9293.LUT_INIT = 16'he4aa;
    SB_LUT4 n10854_bdd_4_lut (.I0(n10854), .I1(\REG.mem_33_5 ), .I2(\REG.mem_32_5 ), 
            .I3(rd_addr_r[1]), .O(n9812));
    defparam n10854_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12078_bdd_4_lut (.I0(n12078), .I1(\REG.mem_57_13 ), .I2(\REG.mem_56_13 ), 
            .I3(rd_addr_r[1]), .O(n12081));
    defparam n12078_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9288 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_6 ), 
            .I2(\REG.mem_15_6 ), .I3(rd_addr_r[1]), .O(n10848));
    defparam rd_addr_r_0__bdd_4_lut_9288.LUT_INIT = 16'he4aa;
    SB_LUT4 n11412_bdd_4_lut (.I0(n11412), .I1(n9529), .I2(n9528), .I3(rd_addr_r[2]), 
            .O(n11415));
    defparam n11412_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10848_bdd_4_lut (.I0(n10848), .I1(\REG.mem_13_6 ), .I2(\REG.mem_12_6 ), 
            .I3(rd_addr_r[1]), .O(n10851));
    defparam n10848_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10314 (.I0(rd_addr_r[2]), .I1(n10274), 
            .I2(n10289), .I3(rd_addr_r[3]), .O(n12072));
    defparam rd_addr_r_2__bdd_4_lut_10314.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9755 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_9 ), 
            .I2(\REG.mem_55_9 ), .I3(rd_addr_r[1]), .O(n11406));
    defparam rd_addr_r_0__bdd_4_lut_9755.LUT_INIT = 16'he4aa;
    SB_LUT4 n12072_bdd_4_lut (.I0(n12072), .I1(n10869), .I2(n10917), .I3(rd_addr_r[3]), 
            .O(n10382));
    defparam n12072_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11406_bdd_4_lut (.I0(n11406), .I1(\REG.mem_53_9 ), .I2(\REG.mem_52_9 ), 
            .I3(rd_addr_r[1]), .O(n11409));
    defparam n11406_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9745 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_0 ), 
            .I2(\REG.mem_35_0 ), .I3(rd_addr_r[1]), .O(n11400));
    defparam rd_addr_r_0__bdd_4_lut_9745.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10304 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_0 ), 
            .I2(\REG.mem_15_0 ), .I3(rd_addr_r[1]), .O(n12066));
    defparam rd_addr_r_0__bdd_4_lut_10304.LUT_INIT = 16'he4aa;
    SB_LUT4 n10794_bdd_4_lut (.I0(n10794), .I1(n10199), .I2(n10190), .I3(rd_addr_r[3]), 
            .O(n10797));
    defparam n10794_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11400_bdd_4_lut (.I0(n11400), .I1(\REG.mem_33_0 ), .I2(\REG.mem_32_0 ), 
            .I3(rd_addr_r[1]), .O(n11403));
    defparam n11400_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12066_bdd_4_lut (.I0(n12066), .I1(\REG.mem_13_0 ), .I2(\REG.mem_12_0 ), 
            .I3(rd_addr_r[1]), .O(n12069));
    defparam n12066_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3577_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_31_10 ), .O(n4666));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3577_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10294 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_14 ), 
            .I2(\REG.mem_43_14 ), .I3(rd_addr_r[1]), .O(n12060));
    defparam rd_addr_r_0__bdd_4_lut_10294.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9750 (.I0(rd_addr_r[1]), .I1(n9708), 
            .I2(n9709), .I3(rd_addr_r[2]), .O(n11394));
    defparam rd_addr_r_1__bdd_4_lut_9750.LUT_INIT = 16'he4aa;
    SB_LUT4 n12060_bdd_4_lut (.I0(n12060), .I1(\REG.mem_41_14 ), .I2(\REG.mem_40_14 ), 
            .I3(rd_addr_r[1]), .O(n12063));
    defparam n12060_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11394_bdd_4_lut (.I0(n11394), .I1(n9706), .I2(n9705), .I3(rd_addr_r[2]), 
            .O(n9751));
    defparam n11394_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3112_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_4_15 ), .O(n4201));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3112_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3111_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_4_14 ), .O(n4200));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3111_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3110_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_4_13 ), .O(n4199));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3110_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3109_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_4_12 ), .O(n4198));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3109_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i254_255 (.Q(\REG.mem_2_8 ), .C(FIFO_CLK_c), .D(n4162));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i251_252 (.Q(\REG.mem_2_7 ), .C(FIFO_CLK_c), .D(n4161));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3108_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_4_11 ), .O(n4197));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3108_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3107_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_4_10 ), .O(n4196));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3107_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3106_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_4_9 ), .O(n4195));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3106_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_buffer__i0  (.Q(\fifo_data_out[0] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5327));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_LUT4 i3576_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_31_9 ), .O(n4665));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3576_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10289 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_11 ), 
            .I2(\REG.mem_11_11 ), .I3(rd_addr_r[1]), .O(n12054));
    defparam rd_addr_r_0__bdd_4_lut_10289.LUT_INIT = 16'he4aa;
    SB_LUT4 i3105_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_4_8 ), .O(n4194));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3105_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3104_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_4_7 ), .O(n4193));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3104_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n12054_bdd_4_lut (.I0(n12054), .I1(\REG.mem_9_11 ), .I2(\REG.mem_8_11 ), 
            .I3(rd_addr_r[1]), .O(n12057));
    defparam n12054_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3103_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_4_6 ), .O(n4192));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3103_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9283 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_15 ), 
            .I2(\REG.mem_63_15 ), .I3(rd_addr_r[1]), .O(n10842));
    defparam rd_addr_r_0__bdd_4_lut_9283.LUT_INIT = 16'he4aa;
    SB_LUT4 i3102_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_4_5 ), .O(n4191));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3102_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9740 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_10 ), 
            .I2(\REG.mem_63_10 ), .I3(rd_addr_r[1]), .O(n11388));
    defparam rd_addr_r_0__bdd_4_lut_9740.LUT_INIT = 16'he4aa;
    SB_DFFE \REG.out_buffer__i15  (.Q(\fifo_data_out[15] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5305));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10284 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_12 ), 
            .I2(\REG.mem_47_12 ), .I3(rd_addr_r[1]), .O(n12048));
    defparam rd_addr_r_0__bdd_4_lut_10284.LUT_INIT = 16'he4aa;
    SB_DFFE \REG.out_buffer__i14  (.Q(\fifo_data_out[14] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5302));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_LUT4 n11388_bdd_4_lut (.I0(n11388), .I1(\REG.mem_61_10 ), .I2(\REG.mem_60_10 ), 
            .I3(rd_addr_r[1]), .O(n10118));
    defparam n11388_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10842_bdd_4_lut (.I0(n10842), .I1(\REG.mem_61_15 ), .I2(\REG.mem_60_15 ), 
            .I3(rd_addr_r[1]), .O(n10845));
    defparam n10842_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \REG.out_buffer__i13  (.Q(\fifo_data_out[13] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5299));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_LUT4 wp_sync2_r_6__I_0_127_inv_0_i4_1_lut (.I0(rd_addr_r[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // src/fifo_dc_32_lut_gen.v(231[47:78])
    defparam wp_sync2_r_6__I_0_127_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE \REG.out_buffer__i12  (.Q(\fifo_data_out[12] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5296));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_DFFE \REG.out_buffer__i11  (.Q(\fifo_data_out[11] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5293));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_LUT4 rd_addr_r_4__bdd_4_lut_9700 (.I0(rd_addr_r[4]), .I1(n9518), 
            .I2(n9563), .I3(rd_addr_r[5]), .O(n10836));
    defparam rd_addr_r_4__bdd_4_lut_9700.LUT_INIT = 16'he4aa;
    SB_DFFE \REG.out_buffer__i10  (.Q(\fifo_data_out[10] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5290));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_LUT4 rd_addr_r_6__I_0_i4_3_lut (.I0(rd_addr_r[3]), .I1(rd_addr_p1_w[3]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_176[3] ));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam rd_addr_r_6__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12048_bdd_4_lut (.I0(n12048), .I1(\REG.mem_45_12 ), .I2(\REG.mem_44_12 ), 
            .I3(rd_addr_r[1]), .O(n9968));
    defparam n12048_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9730 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_15 ), 
            .I2(\REG.mem_47_15 ), .I3(rd_addr_r[1]), .O(n11382));
    defparam rd_addr_r_0__bdd_4_lut_9730.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10279 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_3 ), 
            .I2(\REG.mem_19_3 ), .I3(rd_addr_r[1]), .O(n12042));
    defparam rd_addr_r_0__bdd_4_lut_10279.LUT_INIT = 16'he4aa;
    SB_LUT4 n10836_bdd_4_lut (.I0(n10836), .I1(n10520), .I2(n10502), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_237 [6]));
    defparam n10836_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3101_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_4_4 ), .O(n4190));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3101_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_buffer__i9  (.Q(\fifo_data_out[9] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5255));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_DFFE \REG.out_buffer__i8  (.Q(\fifo_data_out[8] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5252));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_LUT4 n12042_bdd_4_lut (.I0(n12042), .I1(\REG.mem_17_3 ), .I2(\REG.mem_16_3 ), 
            .I3(rd_addr_r[1]), .O(n9551));
    defparam n12042_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \REG.out_buffer__i7  (.Q(\fifo_data_out[7] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5249));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_LUT4 n11382_bdd_4_lut (.I0(n11382), .I1(\REG.mem_45_15 ), .I2(\REG.mem_44_15 ), 
            .I3(rd_addr_r[1]), .O(n11385));
    defparam n11382_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i248_249 (.Q(\REG.mem_2_6 ), .C(FIFO_CLK_c), .D(n4160));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_6__I_0_i6_3_lut (.I0(rd_addr_r[5]), .I1(rd_addr_p1_w[5]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_176[5] ));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam rd_addr_r_6__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9312 (.I0(rd_addr_r[2]), .I1(n10172), 
            .I2(n10181), .I3(rd_addr_r[3]), .O(n10830));
    defparam rd_addr_r_2__bdd_4_lut_9312.LUT_INIT = 16'he4aa;
    SB_LUT4 n10830_bdd_4_lut (.I0(n10830), .I1(n10169), .I2(n10154), .I3(rd_addr_r[3]), 
            .O(n10833));
    defparam n10830_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9735 (.I0(rd_addr_r[1]), .I1(n9732), 
            .I2(n9733), .I3(rd_addr_r[2]), .O(n11376));
    defparam rd_addr_r_1__bdd_4_lut_9735.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10274 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_11 ), 
            .I2(\REG.mem_15_11 ), .I3(rd_addr_r[1]), .O(n12036));
    defparam rd_addr_r_0__bdd_4_lut_10274.LUT_INIT = 16'he4aa;
    SB_DFF i245_246 (.Q(\REG.mem_2_5 ), .C(FIFO_CLK_c), .D(n4159));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3100_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_4_3 ), .O(n4189));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3100_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3099_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_4_2 ), .O(n4188));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3099_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9269 (.I0(rd_addr_r[2]), .I1(n10301), 
            .I2(n10307), .I3(rd_addr_r[3]), .O(n10824));
    defparam rd_addr_r_2__bdd_4_lut_9269.LUT_INIT = 16'he4aa;
    SB_LUT4 i3098_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_4_1 ), .O(n4187));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3098_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8020_3_lut (.I0(n11955), .I1(n11901), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9562));
    defparam i8020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8021_3_lut (.I0(n11091), .I1(n9562), .I2(rd_addr_r[3]), .I3(GND_net), 
            .O(n9563));
    defparam i8021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7975_3_lut (.I0(n10773), .I1(n12351), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9517));
    defparam i7975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7976_3_lut (.I0(n11007), .I1(n9517), .I2(rd_addr_r[3]), .I3(GND_net), 
            .O(n9518));
    defparam i7976_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE \REG.out_buffer__i6  (.Q(\fifo_data_out[6] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5236));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_DFFE \REG.out_buffer__i5  (.Q(\fifo_data_out[5] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5233));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_LUT4 n12036_bdd_4_lut (.I0(n12036), .I1(\REG.mem_13_11 ), .I2(\REG.mem_12_11 ), 
            .I3(rd_addr_r[1]), .O(n12039));
    defparam n12036_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \REG.out_buffer__i4  (.Q(\fifo_data_out[4] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5230));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_LUT4 n11376_bdd_4_lut (.I0(n11376), .I1(n9730), .I2(n9729), .I3(rd_addr_r[2]), 
            .O(n9754));
    defparam n11376_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i6131_6132 (.Q(\REG.mem_63_15 ), .C(FIFO_CLK_c), .D(n5227));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6128_6129 (.Q(\REG.mem_63_14 ), .C(FIFO_CLK_c), .D(n5226));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6125_6126 (.Q(\REG.mem_63_13 ), .C(FIFO_CLK_c), .D(n5225));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6122_6123 (.Q(\REG.mem_63_12 ), .C(FIFO_CLK_c), .D(n5224));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6119_6120 (.Q(\REG.mem_63_11 ), .C(FIFO_CLK_c), .D(n5223));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3097_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_4_0 ), .O(n4186));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3097_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFSR wr_grey_sync_r__i5 (.Q(\wr_grey_sync_r[5] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[5]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(255[21] 265[24])
    SB_DFF i6116_6117 (.Q(\REG.mem_63_10 ), .C(FIFO_CLK_c), .D(n5222));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6113_6114 (.Q(\REG.mem_63_9 ), .C(FIFO_CLK_c), .D(n5221));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6110_6111 (.Q(\REG.mem_63_8 ), .C(FIFO_CLK_c), .D(n5220));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6107_6108 (.Q(\REG.mem_63_7 ), .C(FIFO_CLK_c), .D(n5219));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6104_6105 (.Q(\REG.mem_63_6 ), .C(FIFO_CLK_c), .D(n5218));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6101_6102 (.Q(\REG.mem_63_5 ), .C(FIFO_CLK_c), .D(n5217));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6098_6099 (.Q(\REG.mem_63_4 ), .C(FIFO_CLK_c), .D(n5216));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFFSR wr_grey_sync_r__i4 (.Q(\wr_grey_sync_r[4] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[4]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(255[21] 265[24])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10469 (.I0(rd_addr_r[3]), .I1(n11055), 
            .I2(n9544), .I3(rd_addr_r[4]), .O(n12030));
    defparam rd_addr_r_3__bdd_4_lut_10469.LUT_INIT = 16'he4aa;
    SB_DFFSR wr_grey_sync_r__i3 (.Q(\wr_grey_sync_r[3] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[3]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(255[21] 265[24])
    SB_DFF i6095_6096 (.Q(\REG.mem_63_3 ), .C(FIFO_CLK_c), .D(n5215));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6092_6093 (.Q(\REG.mem_63_2 ), .C(FIFO_CLK_c), .D(n5214));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6089_6090 (.Q(\REG.mem_63_1 ), .C(FIFO_CLK_c), .D(n5213));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFFE \REG.out_buffer__i3  (.Q(\fifo_data_out[3] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5212));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_DFF i6086_6087 (.Q(\REG.mem_63_0 ), .C(FIFO_CLK_c), .D(n5209));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9725 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_2 ), 
            .I2(\REG.mem_19_2 ), .I3(rd_addr_r[1]), .O(n11370));
    defparam rd_addr_r_0__bdd_4_lut_9725.LUT_INIT = 16'he4aa;
    SB_DFF i6035_6036 (.Q(\REG.mem_62_15 ), .C(FIFO_CLK_c), .D(n5208));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6032_6033 (.Q(\REG.mem_62_14 ), .C(FIFO_CLK_c), .D(n5207));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6029_6030 (.Q(\REG.mem_62_13 ), .C(FIFO_CLK_c), .D(n5206));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6026_6027 (.Q(\REG.mem_62_12 ), .C(FIFO_CLK_c), .D(n5205));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6023_6024 (.Q(\REG.mem_62_11 ), .C(FIFO_CLK_c), .D(n5204));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6020_6021 (.Q(\REG.mem_62_10 ), .C(FIFO_CLK_c), .D(n5203));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6017_6018 (.Q(\REG.mem_62_9 ), .C(FIFO_CLK_c), .D(n5202));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6014_6015 (.Q(\REG.mem_62_8 ), .C(FIFO_CLK_c), .D(n5201));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6011_6012 (.Q(\REG.mem_62_7 ), .C(FIFO_CLK_c), .D(n5200));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFFSR wr_grey_sync_r__i2 (.Q(\wr_grey_sync_r[2] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[2]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(255[21] 265[24])
    SB_DFFSR wr_grey_sync_r__i1 (.Q(\wr_grey_sync_r[1] ), .C(FIFO_CLK_c), 
            .D(wr_grey_w[1]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(255[21] 265[24])
    SB_DFF i6008_6009 (.Q(\REG.mem_62_6 ), .C(FIFO_CLK_c), .D(n5199));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n12030_bdd_4_lut (.I0(n12030), .I1(n9520), .I2(n11013), .I3(rd_addr_r[4]), 
            .O(n12033));
    defparam n12030_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10824_bdd_4_lut (.I0(n10824), .I1(n10298), .I2(n10286), .I3(rd_addr_r[3]), 
            .O(n10827));
    defparam n10824_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3051_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_0_0 ), .O(n4140));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3051_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11370_bdd_4_lut (.I0(n11370), .I1(\REG.mem_17_2 ), .I2(\REG.mem_16_2 ), 
            .I3(rd_addr_r[1]), .O(n10124));
    defparam n11370_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3023_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_0_15 ), .O(n4112));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3023_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3024_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_0_14 ), .O(n4113));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3024_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i6005_6006 (.Q(\REG.mem_62_5 ), .C(FIFO_CLK_c), .D(n5198));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i6002_6003 (.Q(\REG.mem_62_4 ), .C(FIFO_CLK_c), .D(n5197));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5999_6000 (.Q(\REG.mem_62_3 ), .C(FIFO_CLK_c), .D(n5196));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5996_5997 (.Q(\REG.mem_62_2 ), .C(FIFO_CLK_c), .D(n5195));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5993_5994 (.Q(\REG.mem_62_1 ), .C(FIFO_CLK_c), .D(n5194));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5990_5991 (.Q(\REG.mem_62_0 ), .C(FIFO_CLK_c), .D(n5193));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5939_5940 (.Q(\REG.mem_61_15 ), .C(FIFO_CLK_c), .D(n5192));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5936_5937 (.Q(\REG.mem_61_14 ), .C(FIFO_CLK_c), .D(n5191));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5933_5934 (.Q(\REG.mem_61_13 ), .C(FIFO_CLK_c), .D(n5190));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5930_5931 (.Q(\REG.mem_61_12 ), .C(FIFO_CLK_c), .D(n5189));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5927_5928 (.Q(\REG.mem_61_11 ), .C(FIFO_CLK_c), .D(n5188));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5924_5925 (.Q(\REG.mem_61_10 ), .C(FIFO_CLK_c), .D(n5187));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5921_5922 (.Q(\REG.mem_61_9 ), .C(FIFO_CLK_c), .D(n5186));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5918_5919 (.Q(\REG.mem_61_8 ), .C(FIFO_CLK_c), .D(n5185));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5915_5916 (.Q(\REG.mem_61_7 ), .C(FIFO_CLK_c), .D(n5184));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5912_5913 (.Q(\REG.mem_61_6 ), .C(FIFO_CLK_c), .D(n5183));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3025_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_0_13 ), .O(n4114));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3025_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10269 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_3 ), 
            .I2(\REG.mem_23_3 ), .I3(rd_addr_r[1]), .O(n12024));
    defparam rd_addr_r_0__bdd_4_lut_10269.LUT_INIT = 16'he4aa;
    SB_LUT4 i3030_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_0_12 ), .O(n4119));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3030_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3031_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_0_11 ), .O(n4120));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3031_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9715 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_8 ), 
            .I2(\REG.mem_27_8 ), .I3(rd_addr_r[1]), .O(n11364));
    defparam rd_addr_r_0__bdd_4_lut_9715.LUT_INIT = 16'he4aa;
    SB_LUT4 i3035_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_0_10 ), .O(n4124));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3035_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5909_5910 (.Q(\REG.mem_61_5 ), .C(FIFO_CLK_c), .D(n5182));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n12024_bdd_4_lut (.I0(n12024), .I1(\REG.mem_21_3 ), .I2(\REG.mem_20_3 ), 
            .I3(rd_addr_r[1]), .O(n9557));
    defparam n12024_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5906_5907 (.Q(\REG.mem_61_4 ), .C(FIFO_CLK_c), .D(n5181));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5903_5904 (.Q(\REG.mem_61_3 ), .C(FIFO_CLK_c), .D(n5180));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5900_5901 (.Q(\REG.mem_61_2 ), .C(FIFO_CLK_c), .D(n5179));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5897_5898 (.Q(\REG.mem_61_1 ), .C(FIFO_CLK_c), .D(n5178));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5894_5895 (.Q(\REG.mem_61_0 ), .C(FIFO_CLK_c), .D(n5177));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5843_5844 (.Q(\REG.mem_60_15 ), .C(FIFO_CLK_c), .D(n5176));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5840_5841 (.Q(\REG.mem_60_14 ), .C(FIFO_CLK_c), .D(n5175));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5837_5838 (.Q(\REG.mem_60_13 ), .C(FIFO_CLK_c), .D(n5174));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5834_5835 (.Q(\REG.mem_60_12 ), .C(FIFO_CLK_c), .D(n5173));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5831_5832 (.Q(\REG.mem_60_11 ), .C(FIFO_CLK_c), .D(n5172));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5828_5829 (.Q(\REG.mem_60_10 ), .C(FIFO_CLK_c), .D(n5171));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5825_5826 (.Q(\REG.mem_60_9 ), .C(FIFO_CLK_c), .D(n5170));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5822_5823 (.Q(\REG.mem_60_8 ), .C(FIFO_CLK_c), .D(n5169));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5819_5820 (.Q(\REG.mem_60_7 ), .C(FIFO_CLK_c), .D(n5168));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5816_5817 (.Q(\REG.mem_60_6 ), .C(FIFO_CLK_c), .D(n5167));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3036_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_0_9 ), .O(n4125));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3036_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11364_bdd_4_lut (.I0(n11364), .I1(\REG.mem_25_8 ), .I2(\REG.mem_24_8 ), 
            .I3(rd_addr_r[1]), .O(n11367));
    defparam n11364_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3037_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_0_8 ), .O(n4126));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3037_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10259 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_9 ), 
            .I2(\REG.mem_47_9 ), .I3(rd_addr_r[1]), .O(n12018));
    defparam rd_addr_r_0__bdd_4_lut_10259.LUT_INIT = 16'he4aa;
    SB_LUT4 n12018_bdd_4_lut (.I0(n12018), .I1(\REG.mem_45_9 ), .I2(\REG.mem_44_9 ), 
            .I3(rd_addr_r[1]), .O(n9977));
    defparam n12018_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9710 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_7 ), 
            .I2(\REG.mem_31_7 ), .I3(rd_addr_r[1]), .O(n11358));
    defparam rd_addr_r_0__bdd_4_lut_9710.LUT_INIT = 16'he4aa;
    SB_DFF i5813_5814 (.Q(\REG.mem_60_5 ), .C(FIFO_CLK_c), .D(n5166));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3042_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_0_7 ), .O(n4131));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3042_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5810_5811 (.Q(\REG.mem_60_4 ), .C(FIFO_CLK_c), .D(n5165));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5807_5808 (.Q(\REG.mem_60_3 ), .C(FIFO_CLK_c), .D(n5164));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5804_5805 (.Q(\REG.mem_60_2 ), .C(FIFO_CLK_c), .D(n5163));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5801_5802 (.Q(\REG.mem_60_1 ), .C(FIFO_CLK_c), .D(n5162));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5798_5799 (.Q(\REG.mem_60_0 ), .C(FIFO_CLK_c), .D(n5161));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5747_5748 (.Q(\REG.mem_59_15 ), .C(FIFO_CLK_c), .D(n5160));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5744_5745 (.Q(\REG.mem_59_14 ), .C(FIFO_CLK_c), .D(n5159));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5741_5742 (.Q(\REG.mem_59_13 ), .C(FIFO_CLK_c), .D(n5158));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5738_5739 (.Q(\REG.mem_59_12 ), .C(FIFO_CLK_c), .D(n5157));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5735_5736 (.Q(\REG.mem_59_11 ), .C(FIFO_CLK_c), .D(n5156));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5732_5733 (.Q(\REG.mem_59_10 ), .C(FIFO_CLK_c), .D(n5155));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5729_5730 (.Q(\REG.mem_59_9 ), .C(FIFO_CLK_c), .D(n5154));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5726_5727 (.Q(\REG.mem_59_8 ), .C(FIFO_CLK_c), .D(n5153));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5723_5724 (.Q(\REG.mem_59_7 ), .C(FIFO_CLK_c), .D(n5152));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5720_5721 (.Q(\REG.mem_59_6 ), .C(FIFO_CLK_c), .D(n5151));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11358_bdd_4_lut (.I0(n11358), .I1(\REG.mem_29_7 ), .I2(\REG.mem_28_7 ), 
            .I3(rd_addr_r[1]), .O(n11361));
    defparam n11358_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3043_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_0_6 ), .O(n4132));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3043_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3044_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_0_5 ), .O(n4133));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3044_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3045_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_0_4 ), .O(n4134));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3045_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5717_5718 (.Q(\REG.mem_59_5 ), .C(FIFO_CLK_c), .D(n5150));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3047_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_0_3 ), .O(n4136));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3047_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5714_5715 (.Q(\REG.mem_59_4 ), .C(FIFO_CLK_c), .D(n5149));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5711_5712 (.Q(\REG.mem_59_3 ), .C(FIFO_CLK_c), .D(n5148));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5708_5709 (.Q(\REG.mem_59_2 ), .C(FIFO_CLK_c), .D(n5147));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5705_5706 (.Q(\REG.mem_59_1 ), .C(FIFO_CLK_c), .D(n5146));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5702_5703 (.Q(\REG.mem_59_0 ), .C(FIFO_CLK_c), .D(n5145));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5651_5652 (.Q(\REG.mem_58_15 ), .C(FIFO_CLK_c), .D(n5144));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5648_5649 (.Q(\REG.mem_58_14 ), .C(FIFO_CLK_c), .D(n5143));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5645_5646 (.Q(\REG.mem_58_13 ), .C(FIFO_CLK_c), .D(n5142));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5642_5643 (.Q(\REG.mem_58_12 ), .C(FIFO_CLK_c), .D(n5141));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5639_5640 (.Q(\REG.mem_58_11 ), .C(FIFO_CLK_c), .D(n5140));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5636_5637 (.Q(\REG.mem_58_10 ), .C(FIFO_CLK_c), .D(n5139));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5633_5634 (.Q(\REG.mem_58_9 ), .C(FIFO_CLK_c), .D(n5138));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5630_5631 (.Q(\REG.mem_58_8 ), .C(FIFO_CLK_c), .D(n5137));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5627_5628 (.Q(\REG.mem_58_7 ), .C(FIFO_CLK_c), .D(n5136));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5624_5625 (.Q(\REG.mem_58_6 ), .C(FIFO_CLK_c), .D(n5135));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_4__bdd_4_lut_9935 (.I0(rd_addr_r[4]), .I1(n10097), 
            .I2(n10106), .I3(rd_addr_r[5]), .O(n11352));
    defparam rd_addr_r_4__bdd_4_lut_9935.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10254 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_10 ), 
            .I2(\REG.mem_47_10 ), .I3(rd_addr_r[1]), .O(n12012));
    defparam rd_addr_r_0__bdd_4_lut_10254.LUT_INIT = 16'he4aa;
    SB_LUT4 n12012_bdd_4_lut (.I0(n12012), .I1(\REG.mem_45_10 ), .I2(\REG.mem_44_10 ), 
            .I3(rd_addr_r[1]), .O(n9980));
    defparam n12012_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3049_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_0_2 ), .O(n4138));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3049_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11352_bdd_4_lut (.I0(n11352), .I1(n10076), .I2(n10061), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_237 [12]));
    defparam n11352_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5621_5622 (.Q(\REG.mem_58_5 ), .C(FIFO_CLK_c), .D(n5134));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10249 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_9 ), 
            .I2(\REG.mem_31_9 ), .I3(rd_addr_r[1]), .O(n12006));
    defparam rd_addr_r_0__bdd_4_lut_10249.LUT_INIT = 16'he4aa;
    SB_DFF i5618_5619 (.Q(\REG.mem_58_4 ), .C(FIFO_CLK_c), .D(n5133));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5615_5616 (.Q(\REG.mem_58_3 ), .C(FIFO_CLK_c), .D(n5132));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5612_5613 (.Q(\REG.mem_58_2 ), .C(FIFO_CLK_c), .D(n5131));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5609_5610 (.Q(\REG.mem_58_1 ), .C(FIFO_CLK_c), .D(n5130));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5606_5607 (.Q(\REG.mem_58_0 ), .C(FIFO_CLK_c), .D(n5129));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5555_5556 (.Q(\REG.mem_57_15 ), .C(FIFO_CLK_c), .D(n5128));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5552_5553 (.Q(\REG.mem_57_14 ), .C(FIFO_CLK_c), .D(n5127));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5549_5550 (.Q(\REG.mem_57_13 ), .C(FIFO_CLK_c), .D(n5126));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5546_5547 (.Q(\REG.mem_57_12 ), .C(FIFO_CLK_c), .D(n5125));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5543_5544 (.Q(\REG.mem_57_11 ), .C(FIFO_CLK_c), .D(n5124));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5540_5541 (.Q(\REG.mem_57_10 ), .C(FIFO_CLK_c), .D(n5123));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5537_5538 (.Q(\REG.mem_57_9 ), .C(FIFO_CLK_c), .D(n5122));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5534_5535 (.Q(\REG.mem_57_8 ), .C(FIFO_CLK_c), .D(n5121));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5531_5532 (.Q(\REG.mem_57_7 ), .C(FIFO_CLK_c), .D(n5120));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5528_5529 (.Q(\REG.mem_57_6 ), .C(FIFO_CLK_c), .D(n5119));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3050_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_0_1 ), .O(n4139));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3050_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_9805 (.I0(rd_addr_r[3]), .I1(n11325), 
            .I2(n9874), .I3(rd_addr_r[4]), .O(n11346));
    defparam rd_addr_r_3__bdd_4_lut_9805.LUT_INIT = 16'he4aa;
    SB_LUT4 n12006_bdd_4_lut (.I0(n12006), .I1(\REG.mem_29_9 ), .I2(\REG.mem_28_9 ), 
            .I3(rd_addr_r[1]), .O(n12009));
    defparam n12006_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3318_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_16_15 ), .O(n4407));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3318_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n10752_bdd_4_lut (.I0(n10752), .I1(\REG.mem_49_0 ), .I2(\REG.mem_48_0 ), 
            .I3(rd_addr_r[1]), .O(n10755));
    defparam n10752_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5525_5526 (.Q(\REG.mem_57_5 ), .C(FIFO_CLK_c), .D(n5118));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3317_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_16_14 ), .O(n4406));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3317_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5522_5523 (.Q(\REG.mem_57_4 ), .C(FIFO_CLK_c), .D(n5117));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5519_5520 (.Q(\REG.mem_57_3 ), .C(FIFO_CLK_c), .D(n5116));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5516_5517 (.Q(\REG.mem_57_2 ), .C(FIFO_CLK_c), .D(n5115));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5513_5514 (.Q(\REG.mem_57_1 ), .C(FIFO_CLK_c), .D(n5114));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFFE \REG.out_buffer__i2  (.Q(\fifo_data_out[2] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5113));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_DFF i5510_5511 (.Q(\REG.mem_57_0 ), .C(FIFO_CLK_c), .D(n5110));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3316_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_16_13 ), .O(n4405));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3316_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5459_5460 (.Q(\REG.mem_56_15 ), .C(FIFO_CLK_c), .D(n5109));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5456_5457 (.Q(\REG.mem_56_14 ), .C(FIFO_CLK_c), .D(n5108));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5453_5454 (.Q(\REG.mem_56_13 ), .C(FIFO_CLK_c), .D(n5107));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5450_5451 (.Q(\REG.mem_56_12 ), .C(FIFO_CLK_c), .D(n5106));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5447_5448 (.Q(\REG.mem_56_11 ), .C(FIFO_CLK_c), .D(n5105));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5444_5445 (.Q(\REG.mem_56_10 ), .C(FIFO_CLK_c), .D(n5104));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5441_5442 (.Q(\REG.mem_56_9 ), .C(FIFO_CLK_c), .D(n5103));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3315_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_16_12 ), .O(n4404));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3315_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11346_bdd_4_lut (.I0(n11346), .I1(n9862), .I2(n9861), .I3(rd_addr_r[4]), 
            .O(n11349));
    defparam n11346_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10244 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_6 ), 
            .I2(\REG.mem_11_6 ), .I3(rd_addr_r[1]), .O(n12000));
    defparam rd_addr_r_0__bdd_4_lut_10244.LUT_INIT = 16'he4aa;
    SB_LUT4 i3314_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_16_11 ), .O(n4403));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3314_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3313_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_16_10 ), .O(n4402));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3313_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5438_5439 (.Q(\REG.mem_56_8 ), .C(FIFO_CLK_c), .D(n5102));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n12000_bdd_4_lut (.I0(n12000), .I1(\REG.mem_9_6 ), .I2(\REG.mem_8_6 ), 
            .I3(rd_addr_r[1]), .O(n9677));
    defparam n12000_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5435_5436 (.Q(\REG.mem_56_7 ), .C(FIFO_CLK_c), .D(n5101));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5432_5433 (.Q(\REG.mem_56_6 ), .C(FIFO_CLK_c), .D(n5100));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5429_5430 (.Q(\REG.mem_56_5 ), .C(FIFO_CLK_c), .D(n5099));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5426_5427 (.Q(\REG.mem_56_4 ), .C(FIFO_CLK_c), .D(n5098));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5423_5424 (.Q(\REG.mem_56_3 ), .C(FIFO_CLK_c), .D(n5097));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5420_5421 (.Q(\REG.mem_56_2 ), .C(FIFO_CLK_c), .D(n5096));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5417_5418 (.Q(\REG.mem_56_1 ), .C(FIFO_CLK_c), .D(n5095));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFFE \REG.out_buffer__i1  (.Q(\fifo_data_out[1] ), .C(DEBUG_6_c), 
            .E(VCC_net), .D(n5094));   // src/fifo_dc_32_lut_gen.v(920[41] 931[44])
    SB_DFF i5414_5415 (.Q(\REG.mem_56_0 ), .C(FIFO_CLK_c), .D(n5091));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3312_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_16_9 ), .O(n4401));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3312_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5363_5364 (.Q(\REG.mem_55_15 ), .C(FIFO_CLK_c), .D(n5090));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5360_5361 (.Q(\REG.mem_55_14 ), .C(FIFO_CLK_c), .D(n5089));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5357_5358 (.Q(\REG.mem_55_13 ), .C(FIFO_CLK_c), .D(n5088));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5354_5355 (.Q(\REG.mem_55_12 ), .C(FIFO_CLK_c), .D(n5087));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_6__I_0_129_7_lut (.I0(GND_net), .I1(rd_addr_r[5]), 
            .I2(GND_net), .I3(n8728), .O(rd_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_129_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3311_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_16_8 ), .O(n4400));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3311_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9705 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_2 ), 
            .I2(\REG.mem_23_2 ), .I3(rd_addr_r[1]), .O(n11340));
    defparam rd_addr_r_0__bdd_4_lut_9705.LUT_INIT = 16'he4aa;
    SB_LUT4 n11340_bdd_4_lut (.I0(n11340), .I1(\REG.mem_21_2 ), .I2(\REG.mem_20_2 ), 
            .I3(rd_addr_r[1]), .O(n10133));
    defparam n11340_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5351_5352 (.Q(\REG.mem_55_11 ), .C(FIFO_CLK_c), .D(n5086));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5348_5349 (.Q(\REG.mem_55_10 ), .C(FIFO_CLK_c), .D(n5085));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5345_5346 (.Q(\REG.mem_55_9 ), .C(FIFO_CLK_c), .D(n5084));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5342_5343 (.Q(\REG.mem_55_8 ), .C(FIFO_CLK_c), .D(n5083));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5339_5340 (.Q(\REG.mem_55_7 ), .C(FIFO_CLK_c), .D(n5082));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5336_5337 (.Q(\REG.mem_55_6 ), .C(FIFO_CLK_c), .D(n5081));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5333_5334 (.Q(\REG.mem_55_5 ), .C(FIFO_CLK_c), .D(n5080));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5330_5331 (.Q(\REG.mem_55_4 ), .C(FIFO_CLK_c), .D(n5079));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5327_5328 (.Q(\REG.mem_55_3 ), .C(FIFO_CLK_c), .D(n5078));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5324_5325 (.Q(\REG.mem_55_2 ), .C(FIFO_CLK_c), .D(n5077));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5321_5322 (.Q(\REG.mem_55_1 ), .C(FIFO_CLK_c), .D(n5076));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5318_5319 (.Q(\REG.mem_55_0 ), .C(FIFO_CLK_c), .D(n5075));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5267_5268 (.Q(\REG.mem_54_15 ), .C(FIFO_CLK_c), .D(n5074));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5264_5265 (.Q(\REG.mem_54_14 ), .C(FIFO_CLK_c), .D(n5073));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5261_5262 (.Q(\REG.mem_54_13 ), .C(FIFO_CLK_c), .D(n5072));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFFSR \en_rd_cnt.rd_counter_r__i4  (.Q(\num_words_in_buffer[6] ), .C(DEBUG_6_c), 
            .D(rd_sig_diff0_w[6]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(704[29] 714[32])
    SB_LUT4 i3310_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_16_7 ), .O(n4399));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3310_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3309_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_16_6 ), .O(n4398));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3309_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3308_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_16_5 ), .O(n4397));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3308_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3307_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_16_4 ), .O(n4396));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3307_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3306_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_16_3 ), .O(n4395));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3306_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3305_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_16_2 ), .O(n4394));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3305_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFSR \en_rd_cnt.rd_counter_r__i3  (.Q(\num_words_in_buffer[5] ), .C(DEBUG_6_c), 
            .D(rd_sig_diff0_w[5]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(704[29] 714[32])
    SB_DFFSR \en_rd_cnt.rd_counter_r__i2  (.Q(\num_words_in_buffer[4] ), .C(DEBUG_6_c), 
            .D(rd_sig_diff0_w[4]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(704[29] 714[32])
    SB_DFF i5258_5259 (.Q(\REG.mem_54_12 ), .C(FIFO_CLK_c), .D(n5071));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3304_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_16_1 ), .O(n4393));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3304_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3303_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_16_0 ), .O(n4392));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3303_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10239 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_15 ), 
            .I2(\REG.mem_3_15 ), .I3(rd_addr_r[1]), .O(n11994));
    defparam rd_addr_r_0__bdd_4_lut_10239.LUT_INIT = 16'he4aa;
    SB_CARRY rd_addr_r_6__I_0_129_7 (.CI(n8728), .I0(rd_addr_r[5]), .I1(GND_net), 
            .CO(n8729));
    SB_LUT4 rd_addr_r_6__I_0_129_6_lut (.I0(GND_net), .I1(rd_addr_r[4]), 
            .I2(GND_net), .I3(n8727), .O(rd_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_129_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3334_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_17_15 ), .O(n4423));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3334_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5255_5256 (.Q(\REG.mem_54_11 ), .C(FIFO_CLK_c), .D(n5070));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5252_5253 (.Q(\REG.mem_54_10 ), .C(FIFO_CLK_c), .D(n5069));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5249_5250 (.Q(\REG.mem_54_9 ), .C(FIFO_CLK_c), .D(n5068));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5246_5247 (.Q(\REG.mem_54_8 ), .C(FIFO_CLK_c), .D(n5067));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5243_5244 (.Q(\REG.mem_54_7 ), .C(FIFO_CLK_c), .D(n5066));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5240_5241 (.Q(\REG.mem_54_6 ), .C(FIFO_CLK_c), .D(n5065));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5237_5238 (.Q(\REG.mem_54_5 ), .C(FIFO_CLK_c), .D(n5064));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5234_5235 (.Q(\REG.mem_54_4 ), .C(FIFO_CLK_c), .D(n5063));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5231_5232 (.Q(\REG.mem_54_3 ), .C(FIFO_CLK_c), .D(n5062));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5228_5229 (.Q(\REG.mem_54_2 ), .C(FIFO_CLK_c), .D(n5061));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5225_5226 (.Q(\REG.mem_54_1 ), .C(FIFO_CLK_c), .D(n5060));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5222_5223 (.Q(\REG.mem_54_0 ), .C(FIFO_CLK_c), .D(n5057));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5171_5172 (.Q(\REG.mem_53_15 ), .C(FIFO_CLK_c), .D(n5056));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5168_5169 (.Q(\REG.mem_53_14 ), .C(FIFO_CLK_c), .D(n5055));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11994_bdd_4_lut (.I0(n11994), .I1(\REG.mem_1_15 ), .I2(\REG.mem_0_15 ), 
            .I3(rd_addr_r[1]), .O(n11997));
    defparam n11994_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY rd_addr_r_6__I_0_129_6 (.CI(n8727), .I0(rd_addr_r[4]), .I1(GND_net), 
            .CO(n8728));
    SB_LUT4 i3333_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_17_14 ), .O(n4422));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3333_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_6__I_0_129_5_lut (.I0(GND_net), .I1(rd_addr_r[3]), 
            .I2(GND_net), .I3(n8726), .O(rd_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_129_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10234 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_12 ), 
            .I2(\REG.mem_51_12 ), .I3(rd_addr_r[1]), .O(n11988));
    defparam rd_addr_r_0__bdd_4_lut_10234.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9244 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_5 ), 
            .I2(\REG.mem_39_5 ), .I3(rd_addr_r[1]), .O(n10788));
    defparam rd_addr_r_0__bdd_4_lut_9244.LUT_INIT = 16'he4aa;
    SB_LUT4 n11988_bdd_4_lut (.I0(n11988), .I1(\REG.mem_49_12 ), .I2(\REG.mem_48_12 ), 
            .I3(rd_addr_r[1]), .O(n9983));
    defparam n11988_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3332_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_17_13 ), .O(n4421));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3332_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n10788_bdd_4_lut (.I0(n10788), .I1(\REG.mem_37_5 ), .I2(\REG.mem_36_5 ), 
            .I3(rd_addr_r[1]), .O(n9824));
    defparam n10788_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_9695 (.I0(rd_addr_r[3]), .I1(n11247), 
            .I2(n9754), .I3(rd_addr_r[4]), .O(n11334));
    defparam rd_addr_r_3__bdd_4_lut_9695.LUT_INIT = 16'he4aa;
    SB_DFF i5165_5166 (.Q(\REG.mem_53_13 ), .C(FIFO_CLK_c), .D(n5054));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5162_5163 (.Q(\REG.mem_53_12 ), .C(FIFO_CLK_c), .D(n5053));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5159_5160 (.Q(\REG.mem_53_11 ), .C(FIFO_CLK_c), .D(n5052));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5156_5157 (.Q(\REG.mem_53_10 ), .C(FIFO_CLK_c), .D(n5051));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5153_5154 (.Q(\REG.mem_53_9 ), .C(FIFO_CLK_c), .D(n5050));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5150_5151 (.Q(\REG.mem_53_8 ), .C(FIFO_CLK_c), .D(n5049));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5147_5148 (.Q(\REG.mem_53_7 ), .C(FIFO_CLK_c), .D(n5048));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5144_5145 (.Q(\REG.mem_53_6 ), .C(FIFO_CLK_c), .D(n5047));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5141_5142 (.Q(\REG.mem_53_5 ), .C(FIFO_CLK_c), .D(n5046));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5138_5139 (.Q(\REG.mem_53_4 ), .C(FIFO_CLK_c), .D(n5045));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5135_5136 (.Q(\REG.mem_53_3 ), .C(FIFO_CLK_c), .D(n5044));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5132_5133 (.Q(\REG.mem_53_2 ), .C(FIFO_CLK_c), .D(n5043));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5129_5130 (.Q(\REG.mem_53_1 ), .C(FIFO_CLK_c), .D(n5042));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5126_5127 (.Q(\REG.mem_53_0 ), .C(FIFO_CLK_c), .D(n5041));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5075_5076 (.Q(\REG.mem_52_15 ), .C(FIFO_CLK_c), .D(n5040));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5072_5073 (.Q(\REG.mem_52_14 ), .C(FIFO_CLK_c), .D(n5039));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11334_bdd_4_lut (.I0(n11334), .I1(n9751), .I2(n11241), .I3(rd_addr_r[4]), 
            .O(n11337));
    defparam n11334_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10429 (.I0(rd_addr_r[1]), .I1(n9858), 
            .I2(n9859), .I3(rd_addr_r[2]), .O(n11982));
    defparam rd_addr_r_1__bdd_4_lut_10429.LUT_INIT = 16'he4aa;
    SB_LUT4 i3331_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_17_12 ), .O(n4420));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3331_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11982_bdd_4_lut (.I0(n11982), .I1(n9838), .I2(n9837), .I3(rd_addr_r[2]), 
            .O(n9985));
    defparam n11982_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9690 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_2 ), 
            .I2(\REG.mem_27_2 ), .I3(rd_addr_r[1]), .O(n11328));
    defparam rd_addr_r_0__bdd_4_lut_9690.LUT_INIT = 16'he4aa;
    SB_LUT4 i3330_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_17_11 ), .O(n4419));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3330_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3329_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_17_10 ), .O(n4418));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3329_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3328_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_17_9 ), .O(n4417));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3328_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10229 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_11 ), 
            .I2(\REG.mem_19_11 ), .I3(rd_addr_r[1]), .O(n11976));
    defparam rd_addr_r_0__bdd_4_lut_10229.LUT_INIT = 16'he4aa;
    SB_LUT4 n11328_bdd_4_lut (.I0(n11328), .I1(\REG.mem_25_2 ), .I2(\REG.mem_24_2 ), 
            .I3(rd_addr_r[1]), .O(n10136));
    defparam n11328_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11976_bdd_4_lut (.I0(n11976), .I1(\REG.mem_17_11 ), .I2(\REG.mem_16_11 ), 
            .I3(rd_addr_r[1]), .O(n10397));
    defparam n11976_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5069_5070 (.Q(\REG.mem_52_13 ), .C(FIFO_CLK_c), .D(n5038));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5066_5067 (.Q(\REG.mem_52_12 ), .C(FIFO_CLK_c), .D(n5037));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5063_5064 (.Q(\REG.mem_52_11 ), .C(FIFO_CLK_c), .D(n5036));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5060_5061 (.Q(\REG.mem_52_10 ), .C(FIFO_CLK_c), .D(n5035));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5057_5058 (.Q(\REG.mem_52_9 ), .C(FIFO_CLK_c), .D(n5034));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5054_5055 (.Q(\REG.mem_52_8 ), .C(FIFO_CLK_c), .D(n5033));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5051_5052 (.Q(\REG.mem_52_7 ), .C(FIFO_CLK_c), .D(n5032));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5048_5049 (.Q(\REG.mem_52_6 ), .C(FIFO_CLK_c), .D(n5031));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5045_5046 (.Q(\REG.mem_52_5 ), .C(FIFO_CLK_c), .D(n5030));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5042_5043 (.Q(\REG.mem_52_4 ), .C(FIFO_CLK_c), .D(n5029));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5039_5040 (.Q(\REG.mem_52_3 ), .C(FIFO_CLK_c), .D(n5028));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5036_5037 (.Q(\REG.mem_52_2 ), .C(FIFO_CLK_c), .D(n5027));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5033_5034 (.Q(\REG.mem_52_1 ), .C(FIFO_CLK_c), .D(n5026));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i5030_5031 (.Q(\REG.mem_52_0 ), .C(FIFO_CLK_c), .D(n5025));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4979_4980 (.Q(\REG.mem_51_15 ), .C(FIFO_CLK_c), .D(n5024));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4976_4977 (.Q(\REG.mem_51_14 ), .C(FIFO_CLK_c), .D(n5023));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i83_2_lut_3_lut (.I0(n36_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n26));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i83_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10219 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_3 ), 
            .I2(\REG.mem_27_3 ), .I3(rd_addr_r[1]), .O(n11970));
    defparam rd_addr_r_0__bdd_4_lut_10219.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9720 (.I0(rd_addr_r[1]), .I1(n9702), 
            .I2(n9703), .I3(rd_addr_r[2]), .O(n11322));
    defparam rd_addr_r_1__bdd_4_lut_9720.LUT_INIT = 16'he4aa;
    SB_LUT4 n11970_bdd_4_lut (.I0(n11970), .I1(\REG.mem_25_3 ), .I2(\REG.mem_24_3 ), 
            .I3(rd_addr_r[1]), .O(n9560));
    defparam n11970_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9239 (.I0(rd_addr_r[2]), .I1(n9536), 
            .I2(n9548), .I3(rd_addr_r[3]), .O(n10782));
    defparam rd_addr_r_2__bdd_4_lut_9239.LUT_INIT = 16'he4aa;
    SB_LUT4 n11322_bdd_4_lut (.I0(n11322), .I1(n9682), .I2(n9681), .I3(rd_addr_r[2]), 
            .O(n11325));
    defparam n11322_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8163_3_lut (.I0(\REG.mem_40_4 ), .I1(\REG.mem_41_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9705));
    defparam i8163_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i4973_4974 (.Q(\REG.mem_51_13 ), .C(FIFO_CLK_c), .D(n5022));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4970_4971 (.Q(\REG.mem_51_12 ), .C(FIFO_CLK_c), .D(n5021));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4967_4968 (.Q(\REG.mem_51_11 ), .C(FIFO_CLK_c), .D(n5020));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4964_4965 (.Q(\REG.mem_51_10 ), .C(FIFO_CLK_c), .D(n5019));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4961_4962 (.Q(\REG.mem_51_9 ), .C(FIFO_CLK_c), .D(n5018));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4958_4959 (.Q(\REG.mem_51_8 ), .C(FIFO_CLK_c), .D(n5017));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4955_4956 (.Q(\REG.mem_51_7 ), .C(FIFO_CLK_c), .D(n5016));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4952_4953 (.Q(\REG.mem_51_6 ), .C(FIFO_CLK_c), .D(n5015));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4949_4950 (.Q(\REG.mem_51_5 ), .C(FIFO_CLK_c), .D(n5014));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4946_4947 (.Q(\REG.mem_51_4 ), .C(FIFO_CLK_c), .D(n5013));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4943_4944 (.Q(\REG.mem_51_3 ), .C(FIFO_CLK_c), .D(n5012));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4940_4941 (.Q(\REG.mem_51_2 ), .C(FIFO_CLK_c), .D(n5011));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4937_4938 (.Q(\REG.mem_51_1 ), .C(FIFO_CLK_c), .D(n5010));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4934_4935 (.Q(\REG.mem_51_0 ), .C(FIFO_CLK_c), .D(n5008));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8164_3_lut (.I0(\REG.mem_42_4 ), .I1(\REG.mem_43_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9706));
    defparam i8164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3327_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_17_8 ), .O(n4416));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3327_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10214 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_11 ), 
            .I2(\REG.mem_23_11 ), .I3(rd_addr_r[1]), .O(n11964));
    defparam rd_addr_r_0__bdd_4_lut_10214.LUT_INIT = 16'he4aa;
    SB_DFF i4883_4884 (.Q(\REG.mem_50_15 ), .C(FIFO_CLK_c), .D(n5007));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 wp_sync2_r_6__I_0_127_add_2_8_lut (.I0(GND_net), .I1(wp_sync2_r[6]), 
            .I2(n1[6]), .I3(n8742), .O(rd_sig_diff0_w[6])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_127_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3326_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_17_7 ), .O(n4415));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3326_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wp_sync2_r_6__I_0_127_add_2_7_lut (.I0(GND_net), .I1(wp_sync_w[5]), 
            .I2(n1[5]), .I3(n8741), .O(rd_sig_diff0_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_127_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF i4880_4881 (.Q(\REG.mem_50_14 ), .C(FIFO_CLK_c), .D(n5006));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_CARRY rd_addr_r_6__I_0_129_5 (.CI(n8726), .I0(rd_addr_r[3]), .I1(GND_net), 
            .CO(n8727));
    SB_DFF i4877_4878 (.Q(\REG.mem_50_13 ), .C(FIFO_CLK_c), .D(n5005));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4874_4875 (.Q(\REG.mem_50_12 ), .C(FIFO_CLK_c), .D(n5004));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4871_4872 (.Q(\REG.mem_50_11 ), .C(FIFO_CLK_c), .D(n5003));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4868_4869 (.Q(\REG.mem_50_10 ), .C(FIFO_CLK_c), .D(n5002));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4865_4866 (.Q(\REG.mem_50_9 ), .C(FIFO_CLK_c), .D(n5001));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4862_4863 (.Q(\REG.mem_50_8 ), .C(FIFO_CLK_c), .D(n5000));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4859_4860 (.Q(\REG.mem_50_7 ), .C(FIFO_CLK_c), .D(n4999));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4856_4857 (.Q(\REG.mem_50_6 ), .C(FIFO_CLK_c), .D(n4998));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4853_4854 (.Q(\REG.mem_50_5 ), .C(FIFO_CLK_c), .D(n4997));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4850_4851 (.Q(\REG.mem_50_4 ), .C(FIFO_CLK_c), .D(n4996));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4847_4848 (.Q(\REG.mem_50_3 ), .C(FIFO_CLK_c), .D(n4995));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4844_4845 (.Q(\REG.mem_50_2 ), .C(FIFO_CLK_c), .D(n4994));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4841_4842 (.Q(\REG.mem_50_1 ), .C(FIFO_CLK_c), .D(n4993));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4838_4839 (.Q(\REG.mem_50_0 ), .C(FIFO_CLK_c), .D(n4992));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_6__I_0_129_4_lut (.I0(GND_net), .I1(rd_addr_r[2]), 
            .I2(GND_net), .I3(n8725), .O(rd_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_129_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3325_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_17_6 ), .O(n4414));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3325_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY wp_sync2_r_6__I_0_127_add_2_7 (.CI(n8741), .I0(wp_sync_w[5]), 
            .I1(n1[5]), .CO(n8742));
    SB_LUT4 i3324_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_17_5 ), .O(n4413));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3324_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wp_sync2_r_6__I_0_127_add_2_6_lut (.I0(GND_net), .I1(wp_sync_w[4]), 
            .I2(n1[4]), .I3(n8740), .O(rd_sig_diff0_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_127_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rd_addr_r_6__I_0_129_4 (.CI(n8725), .I0(rd_addr_r[2]), .I1(GND_net), 
            .CO(n8726));
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9680 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_5 ), 
            .I2(\REG.mem_3_5 ), .I3(rd_addr_r[1]), .O(n11316));
    defparam rd_addr_r_0__bdd_4_lut_9680.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_6__I_0_129_3_lut (.I0(GND_net), .I1(rd_addr_r[1]), 
            .I2(GND_net), .I3(n8724), .O(rd_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_129_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF i4787_4788 (.Q(\REG.mem_49_15 ), .C(FIFO_CLK_c), .D(n4990));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4784_4785 (.Q(\REG.mem_49_14 ), .C(FIFO_CLK_c), .D(n4989));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4781_4782 (.Q(\REG.mem_49_13 ), .C(FIFO_CLK_c), .D(n4988));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4778_4779 (.Q(\REG.mem_49_12 ), .C(FIFO_CLK_c), .D(n4987));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4775_4776 (.Q(\REG.mem_49_11 ), .C(FIFO_CLK_c), .D(n4986));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4772_4773 (.Q(\REG.mem_49_10 ), .C(FIFO_CLK_c), .D(n4985));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4769_4770 (.Q(\REG.mem_49_9 ), .C(FIFO_CLK_c), .D(n4984));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4766_4767 (.Q(\REG.mem_49_8 ), .C(FIFO_CLK_c), .D(n4983));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4763_4764 (.Q(\REG.mem_49_7 ), .C(FIFO_CLK_c), .D(n4982));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4760_4761 (.Q(\REG.mem_49_6 ), .C(FIFO_CLK_c), .D(n4981));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4757_4758 (.Q(\REG.mem_49_5 ), .C(FIFO_CLK_c), .D(n4980));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4754_4755 (.Q(\REG.mem_49_4 ), .C(FIFO_CLK_c), .D(n4979));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4751_4752 (.Q(\REG.mem_49_3 ), .C(FIFO_CLK_c), .D(n4978));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4748_4749 (.Q(\REG.mem_49_2 ), .C(FIFO_CLK_c), .D(n4977));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4745_4746 (.Q(\REG.mem_49_1 ), .C(FIFO_CLK_c), .D(n4976));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11316_bdd_4_lut (.I0(n11316), .I1(\REG.mem_1_5 ), .I2(\REG.mem_0_5 ), 
            .I3(rd_addr_r[1]), .O(n11319));
    defparam n11316_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11964_bdd_4_lut (.I0(n11964), .I1(\REG.mem_21_11 ), .I2(\REG.mem_20_11 ), 
            .I3(rd_addr_r[1]), .O(n10400));
    defparam n11964_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3543_2_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(reset_all), .O(n4632));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam i3543_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i3323_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_17_4 ), .O(n4412));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3323_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_nxt_c_6__I_0_130_i2_2_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_176[1] ), .O(rd_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam rd_addr_nxt_c_6__I_0_130_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_DFF i242_243 (.Q(\REG.mem_2_4 ), .C(FIFO_CLK_c), .D(n4158));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4742_4743 (.Q(\REG.mem_49_0 ), .C(FIFO_CLK_c), .D(n4975));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9670 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_13 ), 
            .I2(\REG.mem_3_13 ), .I3(rd_addr_r[1]), .O(n11310));
    defparam rd_addr_r_0__bdd_4_lut_9670.LUT_INIT = 16'he4aa;
    SB_LUT4 n11310_bdd_4_lut (.I0(n11310), .I1(\REG.mem_1_13 ), .I2(\REG.mem_0_13 ), 
            .I3(rd_addr_r[1]), .O(n11313));
    defparam n11310_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3322_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_17_3 ), .O(n4411));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3322_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3321_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_17_2 ), .O(n4410));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3321_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3320_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_17_1 ), .O(n4409));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3320_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3319_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_17_0 ), .O(n4408));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3319_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3382_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_20_15 ), .O(n4471));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3382_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_nxt_c_6__I_0_130_i3_2_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_176[3] ), .O(rd_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam rd_addr_nxt_c_6__I_0_130_i3_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i3381_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_20_14 ), .O(n4470));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3381_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4691_4692 (.Q(\REG.mem_48_15 ), .C(FIFO_CLK_c), .D(n4968));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4688_4689 (.Q(\REG.mem_48_14 ), .C(FIFO_CLK_c), .D(n4966));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4685_4686 (.Q(\REG.mem_48_13 ), .C(FIFO_CLK_c), .D(n4965));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4682_4683 (.Q(\REG.mem_48_12 ), .C(FIFO_CLK_c), .D(n4964));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4679_4680 (.Q(\REG.mem_48_11 ), .C(FIFO_CLK_c), .D(n4963));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4676_4677 (.Q(\REG.mem_48_10 ), .C(FIFO_CLK_c), .D(n4962));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4673_4674 (.Q(\REG.mem_48_9 ), .C(FIFO_CLK_c), .D(n4961));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4670_4671 (.Q(\REG.mem_48_8 ), .C(FIFO_CLK_c), .D(n4960));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4667_4668 (.Q(\REG.mem_48_7 ), .C(FIFO_CLK_c), .D(n4959));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10209 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_15 ), 
            .I2(\REG.mem_31_15 ), .I3(rd_addr_r[1]), .O(n11958));
    defparam rd_addr_r_0__bdd_4_lut_10209.LUT_INIT = 16'he4aa;
    SB_LUT4 n11958_bdd_4_lut (.I0(n11958), .I1(\REG.mem_29_15 ), .I2(\REG.mem_28_15 ), 
            .I3(rd_addr_r[1]), .O(n11961));
    defparam n11958_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3380_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_20_13 ), .O(n4469));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3380_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3379_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_20_12 ), .O(n4468));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3379_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9665 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_8 ), 
            .I2(\REG.mem_31_8 ), .I3(rd_addr_r[1]), .O(n11304));
    defparam rd_addr_r_0__bdd_4_lut_9665.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10204 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_6 ), 
            .I2(\REG.mem_59_6 ), .I3(rd_addr_r[1]), .O(n11952));
    defparam rd_addr_r_0__bdd_4_lut_10204.LUT_INIT = 16'he4aa;
    SB_LUT4 i3378_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_20_11 ), .O(n4467));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3378_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11304_bdd_4_lut (.I0(n11304), .I1(\REG.mem_29_8 ), .I2(\REG.mem_28_8 ), 
            .I3(rd_addr_r[1]), .O(n11307));
    defparam n11304_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3377_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_20_10 ), .O(n4466));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3377_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8167_3_lut (.I0(\REG.mem_46_4 ), .I1(\REG.mem_47_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9709));
    defparam i8167_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i4664_4665 (.Q(\REG.mem_48_6 ), .C(FIFO_CLK_c), .D(n4958));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4661_4662 (.Q(\REG.mem_48_5 ), .C(FIFO_CLK_c), .D(n4957));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4658_4659 (.Q(\REG.mem_48_4 ), .C(FIFO_CLK_c), .D(n4956));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4655_4656 (.Q(\REG.mem_48_3 ), .C(FIFO_CLK_c), .D(n4955));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4652_4653 (.Q(\REG.mem_48_2 ), .C(FIFO_CLK_c), .D(n4954));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4649_4650 (.Q(\REG.mem_48_1 ), .C(FIFO_CLK_c), .D(n4953));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4646_4647 (.Q(\REG.mem_48_0 ), .C(FIFO_CLK_c), .D(n4952));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4595_4596 (.Q(\REG.mem_47_15 ), .C(FIFO_CLK_c), .D(n4946));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4592_4593 (.Q(\REG.mem_47_14 ), .C(FIFO_CLK_c), .D(n4945));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4589_4590 (.Q(\REG.mem_47_13 ), .C(FIFO_CLK_c), .D(n4944));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFFSR rd_grey_sync_r__i5 (.Q(\rd_grey_sync_r[5] ), .C(DEBUG_6_c), 
            .D(rd_grey_w[5]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(506[21] 516[24])
    SB_DFFSR rd_grey_sync_r__i4 (.Q(\rd_grey_sync_r[4] ), .C(DEBUG_6_c), 
            .D(rd_grey_w[4]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(506[21] 516[24])
    SB_DFFSR rd_grey_sync_r__i3 (.Q(\rd_grey_sync_r[3] ), .C(DEBUG_6_c), 
            .D(rd_grey_w[3]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(506[21] 516[24])
    SB_DFFSR rd_grey_sync_r__i2 (.Q(\rd_grey_sync_r[2] ), .C(DEBUG_6_c), 
            .D(rd_grey_w[2]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(506[21] 516[24])
    SB_DFFSR rd_grey_sync_r__i1 (.Q(\rd_grey_sync_r[1] ), .C(DEBUG_6_c), 
            .D(rd_grey_w[1]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(506[21] 516[24])
    SB_DFF i4586_4587 (.Q(\REG.mem_47_12 ), .C(FIFO_CLK_c), .D(n4943));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_CARRY rd_addr_r_6__I_0_129_3 (.CI(n8724), .I0(rd_addr_r[1]), .I1(GND_net), 
            .CO(n8725));
    SB_LUT4 i8166_3_lut (.I0(\REG.mem_44_4 ), .I1(\REG.mem_45_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9708));
    defparam i8166_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY wp_sync2_r_6__I_0_127_add_2_6 (.CI(n8740), .I0(wp_sync_w[4]), 
            .I1(n1[4]), .CO(n8741));
    SB_LUT4 wp_sync2_r_6__I_0_127_add_2_5_lut (.I0(GND_net), .I1(wp_sync_w[3]), 
            .I2(n1[3]), .I3(n8739), .O(rd_sig_diff0_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_127_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_6__I_0_129_2_lut (.I0(GND_net), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(VCC_net), .O(rd_addr_p1_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_129_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wp_sync2_r_6__I_0_127_add_2_5 (.CI(n8739), .I0(wp_sync_w[3]), 
            .I1(n1[3]), .CO(n8740));
    SB_DFF i4583_4584 (.Q(\REG.mem_47_11 ), .C(FIFO_CLK_c), .D(n4942));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4580_4581 (.Q(\REG.mem_47_10 ), .C(FIFO_CLK_c), .D(n4941));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4577_4578 (.Q(\REG.mem_47_9 ), .C(FIFO_CLK_c), .D(n4940));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4574_4575 (.Q(\REG.mem_47_8 ), .C(FIFO_CLK_c), .D(n4939));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4571_4572 (.Q(\REG.mem_47_7 ), .C(FIFO_CLK_c), .D(n4938));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4568_4569 (.Q(\REG.mem_47_6 ), .C(FIFO_CLK_c), .D(n4937));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4565_4566 (.Q(\REG.mem_47_5 ), .C(FIFO_CLK_c), .D(n4936));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4562_4563 (.Q(\REG.mem_47_4 ), .C(FIFO_CLK_c), .D(n4935));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4559_4560 (.Q(\REG.mem_47_3 ), .C(FIFO_CLK_c), .D(n4934));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4556_4557 (.Q(\REG.mem_47_2 ), .C(FIFO_CLK_c), .D(n4933));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4553_4554 (.Q(\REG.mem_47_1 ), .C(FIFO_CLK_c), .D(n4932));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4550_4551 (.Q(\REG.mem_47_0 ), .C(FIFO_CLK_c), .D(n4929));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4499_4500 (.Q(\REG.mem_46_15 ), .C(FIFO_CLK_c), .D(n4928));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_CARRY wp_sync2_r_6__I_0_127_add_2_4 (.CI(n8738), .I0(wp_sync_w[2]), 
            .I1(n1[2]), .CO(n8739));
    SB_DFF i4496_4497 (.Q(\REG.mem_46_14 ), .C(FIFO_CLK_c), .D(n4927));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_CARRY rd_addr_r_6__I_0_129_2 (.CI(VCC_net), .I0(rd_addr_r[0]), .I1(GND_net), 
            .CO(n8724));
    SB_LUT4 wr_addr_r_6__I_0_8_lut (.I0(GND_net), .I1(\wr_addr_r[6] ), .I2(GND_net), 
            .I3(n8723), .O(wr_addr_p1_w[6])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3376_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_20_9 ), .O(n4465));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3376_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY wp_sync2_r_6__I_0_127_add_2_3 (.CI(n8737), .I0(wp_sync_w[1]), 
            .I1(n1[1]), .CO(n8738));
    SB_DFF i4493_4494 (.Q(\REG.mem_46_13 ), .C(FIFO_CLK_c), .D(n4926));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4490_4491 (.Q(\REG.mem_46_12 ), .C(FIFO_CLK_c), .D(n4925));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4487_4488 (.Q(\REG.mem_46_11 ), .C(FIFO_CLK_c), .D(n4924));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4484_4485 (.Q(\REG.mem_46_10 ), .C(FIFO_CLK_c), .D(n4923));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4481_4482 (.Q(\REG.mem_46_9 ), .C(FIFO_CLK_c), .D(n4922));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4478_4479 (.Q(\REG.mem_46_8 ), .C(FIFO_CLK_c), .D(n4921));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4475_4476 (.Q(\REG.mem_46_7 ), .C(FIFO_CLK_c), .D(n4920));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4472_4473 (.Q(\REG.mem_46_6 ), .C(FIFO_CLK_c), .D(n4919));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4469_4470 (.Q(\REG.mem_46_5 ), .C(FIFO_CLK_c), .D(n4918));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4466_4467 (.Q(\REG.mem_46_4 ), .C(FIFO_CLK_c), .D(n4917));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4463_4464 (.Q(\REG.mem_46_3 ), .C(FIFO_CLK_c), .D(n4916));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4460_4461 (.Q(\REG.mem_46_2 ), .C(FIFO_CLK_c), .D(n4915));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4457_4458 (.Q(\REG.mem_46_1 ), .C(FIFO_CLK_c), .D(n4914));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4454_4455 (.Q(\REG.mem_46_0 ), .C(FIFO_CLK_c), .D(n4913));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4403_4404 (.Q(\REG.mem_45_15 ), .C(FIFO_CLK_c), .D(n4912));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4400_4401 (.Q(\REG.mem_45_14 ), .C(FIFO_CLK_c), .D(n4911));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 wr_addr_r_6__I_0_7_lut (.I0(GND_net), .I1(wr_addr_r[5]), .I2(GND_net), 
            .I3(n8722), .O(wr_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3575_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_31_8 ), .O(n4664));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3575_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY wp_sync2_r_6__I_0_127_add_2_2 (.CI(VCC_net), .I0(wp_sync_w[0]), 
            .I1(n1[0]), .CO(n8737));
    SB_LUT4 EnabledDecoder_2_i82_2_lut_3_lut (.I0(n34), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n59));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i82_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_DFF i4397_4398 (.Q(\REG.mem_45_13 ), .C(FIFO_CLK_c), .D(n4910));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_CARRY wr_addr_r_6__I_0_7 (.CI(n8722), .I0(wr_addr_r[5]), .I1(GND_net), 
            .CO(n8723));
    SB_DFF i4394_4395 (.Q(\REG.mem_45_12 ), .C(FIFO_CLK_c), .D(n4909));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4391_4392 (.Q(\REG.mem_45_11 ), .C(FIFO_CLK_c), .D(n4908));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4388_4389 (.Q(\REG.mem_45_10 ), .C(FIFO_CLK_c), .D(n4907));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4385_4386 (.Q(\REG.mem_45_9 ), .C(FIFO_CLK_c), .D(n4906));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4382_4383 (.Q(\REG.mem_45_8 ), .C(FIFO_CLK_c), .D(n4905));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4379_4380 (.Q(\REG.mem_45_7 ), .C(FIFO_CLK_c), .D(n4904));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4376_4377 (.Q(\REG.mem_45_6 ), .C(FIFO_CLK_c), .D(n4903));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4373_4374 (.Q(\REG.mem_45_5 ), .C(FIFO_CLK_c), .D(n4902));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4370_4371 (.Q(\REG.mem_45_4 ), .C(FIFO_CLK_c), .D(n4901));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4367_4368 (.Q(\REG.mem_45_3 ), .C(FIFO_CLK_c), .D(n4900));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4364_4365 (.Q(\REG.mem_45_2 ), .C(FIFO_CLK_c), .D(n4899));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4361_4362 (.Q(\REG.mem_45_1 ), .C(FIFO_CLK_c), .D(n4898));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4358_4359 (.Q(\REG.mem_45_0 ), .C(FIFO_CLK_c), .D(n4897));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4307_4308 (.Q(\REG.mem_44_15 ), .C(FIFO_CLK_c), .D(n4896));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i81_2_lut_3_lut (.I0(n34), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n27));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i81_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i3574_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_31_7 ), .O(n4663));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3574_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_r_6__I_0_6_lut (.I0(GND_net), .I1(wr_addr_r[4]), .I2(GND_net), 
            .I3(n8721), .O(wr_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_6 (.CI(n8721), .I0(wr_addr_r[4]), .I1(GND_net), 
            .CO(n8722));
    SB_DFF i4304_4305 (.Q(\REG.mem_44_14 ), .C(FIFO_CLK_c), .D(n4895));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4301_4302 (.Q(\REG.mem_44_13 ), .C(FIFO_CLK_c), .D(n4894));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4298_4299 (.Q(\REG.mem_44_12 ), .C(FIFO_CLK_c), .D(n4893));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4295_4296 (.Q(\REG.mem_44_11 ), .C(FIFO_CLK_c), .D(n4892));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4292_4293 (.Q(\REG.mem_44_10 ), .C(FIFO_CLK_c), .D(n4891));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4289_4290 (.Q(\REG.mem_44_9 ), .C(FIFO_CLK_c), .D(n4890));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4286_4287 (.Q(\REG.mem_44_8 ), .C(FIFO_CLK_c), .D(n4889));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4283_4284 (.Q(\REG.mem_44_7 ), .C(FIFO_CLK_c), .D(n4888));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4280_4281 (.Q(\REG.mem_44_6 ), .C(FIFO_CLK_c), .D(n4887));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4277_4278 (.Q(\REG.mem_44_5 ), .C(FIFO_CLK_c), .D(n4886));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4274_4275 (.Q(\REG.mem_44_4 ), .C(FIFO_CLK_c), .D(n4885));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4271_4272 (.Q(\REG.mem_44_3 ), .C(FIFO_CLK_c), .D(n4884));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4268_4269 (.Q(\REG.mem_44_2 ), .C(FIFO_CLK_c), .D(n4883));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4265_4266 (.Q(\REG.mem_44_1 ), .C(FIFO_CLK_c), .D(n4882));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4262_4263 (.Q(\REG.mem_44_0 ), .C(FIFO_CLK_c), .D(n4880));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4211_4212 (.Q(\REG.mem_43_15 ), .C(FIFO_CLK_c), .D(n4879));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3375_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_20_8 ), .O(n4464));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3375_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3374_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_20_7 ), .O(n4463));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3374_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11952_bdd_4_lut (.I0(n11952), .I1(\REG.mem_57_6 ), .I2(\REG.mem_56_6 ), 
            .I3(rd_addr_r[1]), .O(n11955));
    defparam n11952_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3373_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_20_6 ), .O(n4462));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3373_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10224 (.I0(rd_addr_r[1]), .I1(n9918), 
            .I2(n9919), .I3(rd_addr_r[2]), .O(n11946));
    defparam rd_addr_r_1__bdd_4_lut_10224.LUT_INIT = 16'he4aa;
    SB_DFF i4208_4209 (.Q(\REG.mem_43_14 ), .C(FIFO_CLK_c), .D(n4878));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4205_4206 (.Q(\REG.mem_43_13 ), .C(FIFO_CLK_c), .D(n4877));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4202_4203 (.Q(\REG.mem_43_12 ), .C(FIFO_CLK_c), .D(n4876));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4199_4200 (.Q(\REG.mem_43_11 ), .C(FIFO_CLK_c), .D(n4875));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4196_4197 (.Q(\REG.mem_43_10 ), .C(FIFO_CLK_c), .D(n4874));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4193_4194 (.Q(\REG.mem_43_9 ), .C(FIFO_CLK_c), .D(n4873));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4190_4191 (.Q(\REG.mem_43_8 ), .C(FIFO_CLK_c), .D(n4872));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4187_4188 (.Q(\REG.mem_43_7 ), .C(FIFO_CLK_c), .D(n4871));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4184_4185 (.Q(\REG.mem_43_6 ), .C(FIFO_CLK_c), .D(n4870));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4181_4182 (.Q(\REG.mem_43_5 ), .C(FIFO_CLK_c), .D(n4869));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4178_4179 (.Q(\REG.mem_43_4 ), .C(FIFO_CLK_c), .D(n4868));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4175_4176 (.Q(\REG.mem_43_3 ), .C(FIFO_CLK_c), .D(n4867));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4172_4173 (.Q(\REG.mem_43_2 ), .C(FIFO_CLK_c), .D(n4866));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4169_4170 (.Q(\REG.mem_43_1 ), .C(FIFO_CLK_c), .D(n4865));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4166_4167 (.Q(\REG.mem_43_0 ), .C(FIFO_CLK_c), .D(n4864));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4115_4116 (.Q(\REG.mem_42_15 ), .C(FIFO_CLK_c), .D(n4863));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i7986_3_lut (.I0(\REG.mem_0_7 ), .I1(\REG.mem_1_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9528));
    defparam i7986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_5_lut (.I0(GND_net), .I1(wr_addr_r[3]), .I2(GND_net), 
            .I3(n8720), .O(wr_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_5 (.CI(n8720), .I0(wr_addr_r[3]), .I1(GND_net), 
            .CO(n8721));
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9660 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_2 ), 
            .I2(\REG.mem_31_2 ), .I3(rd_addr_r[1]), .O(n11298));
    defparam rd_addr_r_0__bdd_4_lut_9660.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_r_6__I_0_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), .I2(GND_net), 
            .I3(n8719), .O(wr_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7987_3_lut (.I0(\REG.mem_2_7 ), .I1(\REG.mem_3_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9529));
    defparam i7987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n10782_bdd_4_lut (.I0(n10782), .I1(n9533), .I2(n9527), .I3(rd_addr_r[3]), 
            .O(n10785));
    defparam n10782_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY wr_addr_r_6__I_0_4 (.CI(n8719), .I0(wr_addr_r[2]), .I1(GND_net), 
            .CO(n8720));
    SB_DFF i4112_4113 (.Q(\REG.mem_42_14 ), .C(FIFO_CLK_c), .D(n4862));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4109_4110 (.Q(\REG.mem_42_13 ), .C(FIFO_CLK_c), .D(n4861));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4106_4107 (.Q(\REG.mem_42_12 ), .C(FIFO_CLK_c), .D(n4860));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4103_4104 (.Q(\REG.mem_42_11 ), .C(FIFO_CLK_c), .D(n4859));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4100_4101 (.Q(\REG.mem_42_10 ), .C(FIFO_CLK_c), .D(n4858));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4097_4098 (.Q(\REG.mem_42_9 ), .C(FIFO_CLK_c), .D(n4857));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4094_4095 (.Q(\REG.mem_42_8 ), .C(FIFO_CLK_c), .D(n4856));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4091_4092 (.Q(\REG.mem_42_7 ), .C(FIFO_CLK_c), .D(n4855));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4088_4089 (.Q(\REG.mem_42_6 ), .C(FIFO_CLK_c), .D(n4854));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4085_4086 (.Q(\REG.mem_42_5 ), .C(FIFO_CLK_c), .D(n4853));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4082_4083 (.Q(\REG.mem_42_4 ), .C(FIFO_CLK_c), .D(n4852));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4079_4080 (.Q(\REG.mem_42_3 ), .C(FIFO_CLK_c), .D(n4851));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4076_4077 (.Q(\REG.mem_42_2 ), .C(FIFO_CLK_c), .D(n4850));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4073_4074 (.Q(\REG.mem_42_1 ), .C(FIFO_CLK_c), .D(n4849));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4070_4071 (.Q(\REG.mem_42_0 ), .C(FIFO_CLK_c), .D(n4848));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4019_4020 (.Q(\REG.mem_41_15 ), .C(FIFO_CLK_c), .D(n4847));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3372_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_20_5 ), .O(n4461));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3372_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11946_bdd_4_lut (.I0(n11946), .I1(n9904), .I2(n9903), .I3(rd_addr_r[2]), 
            .O(n9997));
    defparam n11946_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11298_bdd_4_lut (.I0(n11298), .I1(\REG.mem_29_2 ), .I2(\REG.mem_28_2 ), 
            .I3(rd_addr_r[1]), .O(n10148));
    defparam n11298_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3573_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_31_6 ), .O(n4662));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3573_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wp_sync2_r_6__I_0_127_inv_0_i5_1_lut (.I0(rd_addr_r[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // src/fifo_dc_32_lut_gen.v(231[47:78])
    defparam wp_sync2_r_6__I_0_127_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3371_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_20_4 ), .O(n4460));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3371_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10199 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_11 ), 
            .I2(\REG.mem_27_11 ), .I3(rd_addr_r[1]), .O(n11940));
    defparam rd_addr_r_0__bdd_4_lut_10199.LUT_INIT = 16'he4aa;
    SB_LUT4 i8023_3_lut (.I0(\REG.mem_6_7 ), .I1(\REG.mem_7_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9565));
    defparam i8023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9655 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_15 ), 
            .I2(\REG.mem_51_15 ), .I3(rd_addr_r[1]), .O(n11292));
    defparam rd_addr_r_0__bdd_4_lut_9655.LUT_INIT = 16'he4aa;
    SB_LUT4 i8022_3_lut (.I0(\REG.mem_4_7 ), .I1(\REG.mem_5_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9564));
    defparam i8022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11292_bdd_4_lut (.I0(n11292), .I1(\REG.mem_49_15 ), .I2(\REG.mem_48_15 ), 
            .I3(rd_addr_r[1]), .O(n11295));
    defparam n11292_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4016_4017 (.Q(\REG.mem_41_14 ), .C(FIFO_CLK_c), .D(n4846));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4013_4014 (.Q(\REG.mem_41_13 ), .C(FIFO_CLK_c), .D(n4845));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4010_4011 (.Q(\REG.mem_41_12 ), .C(FIFO_CLK_c), .D(n4844));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4007_4008 (.Q(\REG.mem_41_11 ), .C(FIFO_CLK_c), .D(n4843));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4004_4005 (.Q(\REG.mem_41_10 ), .C(FIFO_CLK_c), .D(n4842));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i4001_4002 (.Q(\REG.mem_41_9 ), .C(FIFO_CLK_c), .D(n4841));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3998_3999 (.Q(\REG.mem_41_8 ), .C(FIFO_CLK_c), .D(n4840));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3995_3996 (.Q(\REG.mem_41_7 ), .C(FIFO_CLK_c), .D(n4839));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3992_3993 (.Q(\REG.mem_41_6 ), .C(FIFO_CLK_c), .D(n4838));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3989_3990 (.Q(\REG.mem_41_5 ), .C(FIFO_CLK_c), .D(n4837));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3986_3987 (.Q(\REG.mem_41_4 ), .C(FIFO_CLK_c), .D(n4836));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3983_3984 (.Q(\REG.mem_41_3 ), .C(FIFO_CLK_c), .D(n4835));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3980_3981 (.Q(\REG.mem_41_2 ), .C(FIFO_CLK_c), .D(n4834));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3977_3978 (.Q(\REG.mem_41_1 ), .C(FIFO_CLK_c), .D(n4833));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3974_3975 (.Q(\REG.mem_41_0 ), .C(FIFO_CLK_c), .D(n4832));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8112_3_lut (.I0(\REG.mem_16_7 ), .I1(\REG.mem_17_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9654));
    defparam i8112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8113_3_lut (.I0(\REG.mem_18_7 ), .I1(\REG.mem_19_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9655));
    defparam i8113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11940_bdd_4_lut (.I0(n11940), .I1(\REG.mem_25_11 ), .I2(\REG.mem_24_11 ), 
            .I3(rd_addr_r[1]), .O(n10406));
    defparam n11940_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3370_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_20_3 ), .O(n4459));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3370_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8739_3_lut (.I0(n11997), .I1(n11439), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10281));
    defparam i8739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8740_3_lut (.I0(n10815), .I1(n12363), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10282));
    defparam i8740_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i239_240 (.Q(\REG.mem_2_3 ), .C(FIFO_CLK_c), .D(n4157));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3369_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_20_2 ), .O(n4458));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3369_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3923_3924 (.Q(\REG.mem_40_15 ), .C(FIFO_CLK_c), .D(n4831));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3368_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_20_1 ), .O(n4457));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3368_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3920_3921 (.Q(\REG.mem_40_14 ), .C(FIFO_CLK_c), .D(n4830));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3367_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_20_0 ), .O(n4456));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3367_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3917_3918 (.Q(\REG.mem_40_13 ), .C(FIFO_CLK_c), .D(n4829));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3914_3915 (.Q(\REG.mem_40_12 ), .C(FIFO_CLK_c), .D(n4828));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3911_3912 (.Q(\REG.mem_40_11 ), .C(FIFO_CLK_c), .D(n4827));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3908_3909 (.Q(\REG.mem_40_10 ), .C(FIFO_CLK_c), .D(n4826));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3905_3906 (.Q(\REG.mem_40_9 ), .C(FIFO_CLK_c), .D(n4825));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3902_3903 (.Q(\REG.mem_40_8 ), .C(FIFO_CLK_c), .D(n4824));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3899_3900 (.Q(\REG.mem_40_7 ), .C(FIFO_CLK_c), .D(n4823));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3896_3897 (.Q(\REG.mem_40_6 ), .C(FIFO_CLK_c), .D(n4822));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3893_3894 (.Q(\REG.mem_40_5 ), .C(FIFO_CLK_c), .D(n4821));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3890_3891 (.Q(\REG.mem_40_4 ), .C(FIFO_CLK_c), .D(n4820));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3887_3888 (.Q(\REG.mem_40_3 ), .C(FIFO_CLK_c), .D(n4819));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3884_3885 (.Q(\REG.mem_40_2 ), .C(FIFO_CLK_c), .D(n4818));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3881_3882 (.Q(\REG.mem_40_1 ), .C(FIFO_CLK_c), .D(n4817));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3878_3879 (.Q(\REG.mem_40_0 ), .C(FIFO_CLK_c), .D(n4814));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3827_3828 (.Q(\REG.mem_39_15 ), .C(FIFO_CLK_c), .D(n4813));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8776_3_lut (.I0(n12105), .I1(n11961), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10318));
    defparam i8776_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3824_3825 (.Q(\REG.mem_39_14 ), .C(FIFO_CLK_c), .D(n4812));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8149_3_lut (.I0(\REG.mem_22_7 ), .I1(\REG.mem_23_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9691));
    defparam i8149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3506_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_27_15 ), .O(n4595));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3506_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_r_6__I_0_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), .I2(GND_net), 
            .I3(n8718), .O(wr_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF i3821_3822 (.Q(\REG.mem_39_13 ), .C(FIFO_CLK_c), .D(n4811));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_CARRY wr_addr_r_6__I_0_3 (.CI(n8718), .I0(wr_addr_r[1]), .I1(GND_net), 
            .CO(n8719));
    SB_DFF i3818_3819 (.Q(\REG.mem_39_12 ), .C(FIFO_CLK_c), .D(n4810));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3505_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_27_14 ), .O(n4594));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3505_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3815_3816 (.Q(\REG.mem_39_11 ), .C(FIFO_CLK_c), .D(n4809));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8148_3_lut (.I0(\REG.mem_20_7 ), .I1(\REG.mem_21_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9690));
    defparam i8148_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3812_3813 (.Q(\REG.mem_39_10 ), .C(FIFO_CLK_c), .D(n4808));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3504_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_27_13 ), .O(n4593));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3504_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10189 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_11 ), 
            .I2(\REG.mem_31_11 ), .I3(rd_addr_r[1]), .O(n11934));
    defparam rd_addr_r_0__bdd_4_lut_10189.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_r_6__I_0_2_lut (.I0(GND_net), .I1(wr_addr_r[0]), .I2(GND_net), 
            .I3(VCC_net), .O(wr_addr_p1_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF i3809_3810 (.Q(\REG.mem_39_9 ), .C(FIFO_CLK_c), .D(n4807));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3806_3807 (.Q(\REG.mem_39_8 ), .C(FIFO_CLK_c), .D(n4806));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3803_3804 (.Q(\REG.mem_39_7 ), .C(FIFO_CLK_c), .D(n4805));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3800_3801 (.Q(\REG.mem_39_6 ), .C(FIFO_CLK_c), .D(n4804));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3797_3798 (.Q(\REG.mem_39_5 ), .C(FIFO_CLK_c), .D(n4803));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3794_3795 (.Q(\REG.mem_39_4 ), .C(FIFO_CLK_c), .D(n4802));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3791_3792 (.Q(\REG.mem_39_3 ), .C(FIFO_CLK_c), .D(n4801));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3788_3789 (.Q(\REG.mem_39_2 ), .C(FIFO_CLK_c), .D(n4800));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3785_3786 (.Q(\REG.mem_39_1 ), .C(FIFO_CLK_c), .D(n4799));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3782_3783 (.Q(\REG.mem_39_0 ), .C(FIFO_CLK_c), .D(n4798));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3731_3732 (.Q(\REG.mem_38_15 ), .C(FIFO_CLK_c), .D(n4797));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3728_3729 (.Q(\REG.mem_38_14 ), .C(FIFO_CLK_c), .D(n4796));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3725_3726 (.Q(\REG.mem_38_13 ), .C(FIFO_CLK_c), .D(n4795));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3722_3723 (.Q(\REG.mem_38_12 ), .C(FIFO_CLK_c), .D(n4794));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3719_3720 (.Q(\REG.mem_38_11 ), .C(FIFO_CLK_c), .D(n4793));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11934_bdd_4_lut (.I0(n11934), .I1(\REG.mem_29_11 ), .I2(\REG.mem_28_11 ), 
            .I3(rd_addr_r[1]), .O(n10409));
    defparam n11934_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3503_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_27_12 ), .O(n4592));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3503_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3716_3717 (.Q(\REG.mem_38_10 ), .C(FIFO_CLK_c), .D(n4792));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3502_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_27_11 ), .O(n4591));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3502_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3501_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_27_10 ), .O(n4590));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3501_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3500_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_27_9 ), .O(n4589));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3500_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10184 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_13 ), 
            .I2(\REG.mem_63_13 ), .I3(rd_addr_r[1]), .O(n11928));
    defparam rd_addr_r_0__bdd_4_lut_10184.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9650 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_2 ), 
            .I2(\REG.mem_35_2 ), .I3(rd_addr_r[1]), .O(n11286));
    defparam rd_addr_r_0__bdd_4_lut_9650.LUT_INIT = 16'he4aa;
    SB_LUT4 i3499_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_27_8 ), .O(n4588));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3499_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11928_bdd_4_lut (.I0(n11928), .I1(\REG.mem_61_13 ), .I2(\REG.mem_60_13 ), 
            .I3(rd_addr_r[1]), .O(n11931));
    defparam n11928_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11286_bdd_4_lut (.I0(n11286), .I1(\REG.mem_33_2 ), .I2(\REG.mem_32_2 ), 
            .I3(rd_addr_r[1]), .O(n10154));
    defparam n11286_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3498_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_27_7 ), .O(n4587));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3498_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3713_3714 (.Q(\REG.mem_38_9 ), .C(FIFO_CLK_c), .D(n4791));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3710_3711 (.Q(\REG.mem_38_8 ), .C(FIFO_CLK_c), .D(n4790));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3707_3708 (.Q(\REG.mem_38_7 ), .C(FIFO_CLK_c), .D(n4789));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3704_3705 (.Q(\REG.mem_38_6 ), .C(FIFO_CLK_c), .D(n4788));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3701_3702 (.Q(\REG.mem_38_5 ), .C(FIFO_CLK_c), .D(n4787));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3698_3699 (.Q(\REG.mem_38_4 ), .C(FIFO_CLK_c), .D(n4786));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3695_3696 (.Q(\REG.mem_38_3 ), .C(FIFO_CLK_c), .D(n4785));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3692_3693 (.Q(\REG.mem_38_2 ), .C(FIFO_CLK_c), .D(n4784));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3689_3690 (.Q(\REG.mem_38_1 ), .C(FIFO_CLK_c), .D(n4783));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3686_3687 (.Q(\REG.mem_38_0 ), .C(FIFO_CLK_c), .D(n4782));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3635_3636 (.Q(\REG.mem_37_15 ), .C(FIFO_CLK_c), .D(n4781));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3632_3633 (.Q(\REG.mem_37_14 ), .C(FIFO_CLK_c), .D(n4780));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3629_3630 (.Q(\REG.mem_37_13 ), .C(FIFO_CLK_c), .D(n4779));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3626_3627 (.Q(\REG.mem_37_12 ), .C(FIFO_CLK_c), .D(n4778));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3623_3624 (.Q(\REG.mem_37_11 ), .C(FIFO_CLK_c), .D(n4777));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3620_3621 (.Q(\REG.mem_37_10 ), .C(FIFO_CLK_c), .D(n4776));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3497_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_27_6 ), .O(n4586));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3497_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3496_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_27_5 ), .O(n4585));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3496_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3617_3618 (.Q(\REG.mem_37_9 ), .C(FIFO_CLK_c), .D(n4775));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3614_3615 (.Q(\REG.mem_37_8 ), .C(FIFO_CLK_c), .D(n4774));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3495_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_27_4 ), .O(n4584));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3495_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY wr_addr_r_6__I_0_2 (.CI(VCC_net), .I0(wr_addr_r[0]), .I1(GND_net), 
            .CO(n8718));
    SB_DFF i3611_3612 (.Q(\REG.mem_37_7 ), .C(FIFO_CLK_c), .D(n4773));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3608_3609 (.Q(\REG.mem_37_6 ), .C(FIFO_CLK_c), .D(n4772));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3605_3606 (.Q(\REG.mem_37_5 ), .C(FIFO_CLK_c), .D(n4771));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3602_3603 (.Q(\REG.mem_37_4 ), .C(FIFO_CLK_c), .D(n4770));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3599_3600 (.Q(\REG.mem_37_3 ), .C(FIFO_CLK_c), .D(n4769));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3596_3597 (.Q(\REG.mem_37_2 ), .C(FIFO_CLK_c), .D(n4768));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3593_3594 (.Q(\REG.mem_37_1 ), .C(FIFO_CLK_c), .D(n4767));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3590_3591 (.Q(\REG.mem_37_0 ), .C(FIFO_CLK_c), .D(n4766));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3539_3540 (.Q(\REG.mem_36_15 ), .C(FIFO_CLK_c), .D(n4765));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3536_3537 (.Q(\REG.mem_36_14 ), .C(FIFO_CLK_c), .D(n4764));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3533_3534 (.Q(\REG.mem_36_13 ), .C(FIFO_CLK_c), .D(n4763));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3530_3531 (.Q(\REG.mem_36_12 ), .C(FIFO_CLK_c), .D(n4762));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3527_3528 (.Q(\REG.mem_36_11 ), .C(FIFO_CLK_c), .D(n4761));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3524_3525 (.Q(\REG.mem_36_10 ), .C(FIFO_CLK_c), .D(n4760));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3521_3522 (.Q(\REG.mem_36_9 ), .C(FIFO_CLK_c), .D(n4759));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i236_237 (.Q(\REG.mem_2_2 ), .C(FIFO_CLK_c), .D(n4156));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3494_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_27_3 ), .O(n4583));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3494_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3572_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_31_5 ), .O(n4661));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3572_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3493_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_27_2 ), .O(n4582));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3493_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3492_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_27_1 ), .O(n4581));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3492_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10179 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_6 ), 
            .I2(\REG.mem_27_6 ), .I3(rd_addr_r[1]), .O(n11922));
    defparam rd_addr_r_0__bdd_4_lut_10179.LUT_INIT = 16'he4aa;
    SB_LUT4 i3491_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_27_0 ), .O(n4580));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3491_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3518_3519 (.Q(\REG.mem_36_8 ), .C(FIFO_CLK_c), .D(n4758));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3515_3516 (.Q(\REG.mem_36_7 ), .C(FIFO_CLK_c), .D(n4757));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3090_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_3_9 ), .O(n4179));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3090_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3512_3513 (.Q(\REG.mem_36_6 ), .C(FIFO_CLK_c), .D(n4756));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3509_3510 (.Q(\REG.mem_36_5 ), .C(FIFO_CLK_c), .D(n4755));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3506_3507 (.Q(\REG.mem_36_4 ), .C(FIFO_CLK_c), .D(n4754));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3503_3504 (.Q(\REG.mem_36_3 ), .C(FIFO_CLK_c), .D(n4753));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3500_3501 (.Q(\REG.mem_36_2 ), .C(FIFO_CLK_c), .D(n4752));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3497_3498 (.Q(\REG.mem_36_1 ), .C(FIFO_CLK_c), .D(n4751));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3494_3495 (.Q(\REG.mem_36_0 ), .C(FIFO_CLK_c), .D(n4750));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3443_3444 (.Q(\REG.mem_35_15 ), .C(FIFO_CLK_c), .D(n4749));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3440_3441 (.Q(\REG.mem_35_14 ), .C(FIFO_CLK_c), .D(n4748));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3437_3438 (.Q(\REG.mem_35_13 ), .C(FIFO_CLK_c), .D(n4747));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3434_3435 (.Q(\REG.mem_35_12 ), .C(FIFO_CLK_c), .D(n4746));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3431_3432 (.Q(\REG.mem_35_11 ), .C(FIFO_CLK_c), .D(n4745));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3428_3429 (.Q(\REG.mem_35_10 ), .C(FIFO_CLK_c), .D(n4744));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3425_3426 (.Q(\REG.mem_35_9 ), .C(FIFO_CLK_c), .D(n4743));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3422_3423 (.Q(\REG.mem_35_8 ), .C(FIFO_CLK_c), .D(n4742));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3089_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_3_8 ), .O(n4178));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3089_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3088_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_3_7 ), .O(n4177));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3088_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3087_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_3_6 ), .O(n4176));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3087_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3086_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_3_5 ), .O(n4175));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3086_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3419_3420 (.Q(\REG.mem_35_7 ), .C(FIFO_CLK_c), .D(n4741));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11922_bdd_4_lut (.I0(n11922), .I1(\REG.mem_25_6 ), .I2(\REG.mem_24_6 ), 
            .I3(rd_addr_r[1]), .O(n10001));
    defparam n11922_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9645 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_9 ), 
            .I2(\REG.mem_35_9 ), .I3(rd_addr_r[1]), .O(n11280));
    defparam rd_addr_r_0__bdd_4_lut_9645.LUT_INIT = 16'he4aa;
    SB_LUT4 i3085_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_3_4 ), .O(n4174));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3085_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3416_3417 (.Q(\REG.mem_35_6 ), .C(FIFO_CLK_c), .D(n4740));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3413_3414 (.Q(\REG.mem_35_5 ), .C(FIFO_CLK_c), .D(n4739));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3410_3411 (.Q(\REG.mem_35_4 ), .C(FIFO_CLK_c), .D(n4738));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3407_3408 (.Q(\REG.mem_35_3 ), .C(FIFO_CLK_c), .D(n4737));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3404_3405 (.Q(\REG.mem_35_2 ), .C(FIFO_CLK_c), .D(n4736));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3401_3402 (.Q(\REG.mem_35_1 ), .C(FIFO_CLK_c), .D(n4735));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3398_3399 (.Q(\REG.mem_35_0 ), .C(FIFO_CLK_c), .D(n4734));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3347_3348 (.Q(\REG.mem_34_15 ), .C(FIFO_CLK_c), .D(n4733));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3344_3345 (.Q(\REG.mem_34_14 ), .C(FIFO_CLK_c), .D(n4732));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3341_3342 (.Q(\REG.mem_34_13 ), .C(FIFO_CLK_c), .D(n4731));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3338_3339 (.Q(\REG.mem_34_12 ), .C(FIFO_CLK_c), .D(n4730));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3335_3336 (.Q(\REG.mem_34_11 ), .C(FIFO_CLK_c), .D(n4729));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3332_3333 (.Q(\REG.mem_34_10 ), .C(FIFO_CLK_c), .D(n4728));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3329_3330 (.Q(\REG.mem_34_9 ), .C(FIFO_CLK_c), .D(n4727));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3326_3327 (.Q(\REG.mem_34_8 ), .C(FIFO_CLK_c), .D(n4726));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3323_3324 (.Q(\REG.mem_34_7 ), .C(FIFO_CLK_c), .D(n4725));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i233_234 (.Q(\REG.mem_2_1 ), .C(FIFO_CLK_c), .D(n4155));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i230_231 (.Q(\REG.mem_2_0 ), .C(FIFO_CLK_c), .D(n4154));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3084_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_3_3 ), .O(n4173));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3084_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i179_180 (.Q(\REG.mem_1_15 ), .C(FIFO_CLK_c), .D(n4153));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11280_bdd_4_lut (.I0(n11280), .I1(\REG.mem_33_9 ), .I2(\REG.mem_32_9 ), 
            .I3(rd_addr_r[1]), .O(n11283));
    defparam n11280_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i176_177 (.Q(\REG.mem_1_14 ), .C(FIFO_CLK_c), .D(n4152));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i173_174 (.Q(\REG.mem_1_13 ), .C(FIFO_CLK_c), .D(n4151));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i170_171 (.Q(\REG.mem_1_12 ), .C(FIFO_CLK_c), .D(n4150));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8142_3_lut (.I0(\REG.mem_24_4 ), .I1(\REG.mem_25_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9684));
    defparam i8142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10174 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_14 ), 
            .I2(\REG.mem_47_14 ), .I3(rd_addr_r[1]), .O(n11916));
    defparam rd_addr_r_0__bdd_4_lut_10174.LUT_INIT = 16'he4aa;
    SB_LUT4 i8143_3_lut (.I0(\REG.mem_26_4 ), .I1(\REG.mem_27_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9685));
    defparam i8143_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3320_3321 (.Q(\REG.mem_34_6 ), .C(FIFO_CLK_c), .D(n4724));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8146_3_lut (.I0(\REG.mem_30_4 ), .I1(\REG.mem_31_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9688));
    defparam i8146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8145_3_lut (.I0(\REG.mem_28_4 ), .I1(\REG.mem_29_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9687));
    defparam i8145_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3317_3318 (.Q(\REG.mem_34_5 ), .C(FIFO_CLK_c), .D(n4723));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3314_3315 (.Q(\REG.mem_34_4 ), .C(FIFO_CLK_c), .D(n4722));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3311_3312 (.Q(\REG.mem_34_3 ), .C(FIFO_CLK_c), .D(n4721));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3308_3309 (.Q(\REG.mem_34_2 ), .C(FIFO_CLK_c), .D(n4720));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3305_3306 (.Q(\REG.mem_34_1 ), .C(FIFO_CLK_c), .D(n4719));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3302_3303 (.Q(\REG.mem_34_0 ), .C(FIFO_CLK_c), .D(n4718));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3251_3252 (.Q(\REG.mem_33_15 ), .C(FIFO_CLK_c), .D(n4717));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3248_3249 (.Q(\REG.mem_33_14 ), .C(FIFO_CLK_c), .D(n4716));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3245_3246 (.Q(\REG.mem_33_13 ), .C(FIFO_CLK_c), .D(n4715));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3242_3243 (.Q(\REG.mem_33_12 ), .C(FIFO_CLK_c), .D(n4714));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3239_3240 (.Q(\REG.mem_33_11 ), .C(FIFO_CLK_c), .D(n4713));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3236_3237 (.Q(\REG.mem_33_10 ), .C(FIFO_CLK_c), .D(n4712));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3233_3234 (.Q(\REG.mem_33_9 ), .C(FIFO_CLK_c), .D(n4711));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3230_3231 (.Q(\REG.mem_33_8 ), .C(FIFO_CLK_c), .D(n4710));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3227_3228 (.Q(\REG.mem_33_7 ), .C(FIFO_CLK_c), .D(n4709));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3224_3225 (.Q(\REG.mem_33_6 ), .C(FIFO_CLK_c), .D(n4708));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3083_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_3_2 ), .O(n4172));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3083_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8328_3_lut (.I0(\REG.mem_48_7 ), .I1(\REG.mem_49_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9870));
    defparam i8328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3082_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_3_1 ), .O(n4171));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3082_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8329_3_lut (.I0(\REG.mem_50_7 ), .I1(\REG.mem_51_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9871));
    defparam i8329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8341_3_lut (.I0(\REG.mem_54_7 ), .I1(\REG.mem_55_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9883));
    defparam i8341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3081_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_3_0 ), .O(n4170));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3081_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8340_3_lut (.I0(\REG.mem_52_7 ), .I1(\REG.mem_53_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9882));
    defparam i8340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11916_bdd_4_lut (.I0(n11916), .I1(\REG.mem_45_14 ), .I2(\REG.mem_44_14 ), 
            .I3(rd_addr_r[1]), .O(n11919));
    defparam n11916_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9640 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_8 ), 
            .I2(\REG.mem_35_8 ), .I3(rd_addr_r[1]), .O(n11274));
    defparam rd_addr_r_0__bdd_4_lut_9640.LUT_INIT = 16'he4aa;
    SB_LUT4 i8407_3_lut (.I0(n11685), .I1(n10761), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9949));
    defparam i8407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8422_3_lut (.I0(n11595), .I1(n11361), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9964));
    defparam i8422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_6__I_0_127_inv_0_i6_1_lut (.I0(rd_addr_r[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // src/fifo_dc_32_lut_gen.v(231[47:78])
    defparam wp_sync2_r_6__I_0_127_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10169 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_12 ), 
            .I2(\REG.mem_55_12 ), .I3(rd_addr_r[1]), .O(n11910));
    defparam rd_addr_r_0__bdd_4_lut_10169.LUT_INIT = 16'he4aa;
    SB_LUT4 i8115_3_lut (.I0(\REG.mem_8_4 ), .I1(\REG.mem_9_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9657));
    defparam i8115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11274_bdd_4_lut (.I0(n11274), .I1(\REG.mem_33_8 ), .I2(\REG.mem_32_8 ), 
            .I3(rd_addr_r[1]), .O(n11277));
    defparam n11274_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11910_bdd_4_lut (.I0(n11910), .I1(\REG.mem_53_12 ), .I2(\REG.mem_52_12 ), 
            .I3(rd_addr_r[1]), .O(n10004));
    defparam n11910_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_6__I_0_121_i1_2_lut (.I0(wp_sync2_r[5]), .I1(wp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(wp_sync_w[5]));   // src/fifo_dc_32_lut_gen.v(537[38:77])
    defparam wp_sync2_r_6__I_0_121_i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8116_3_lut (.I0(\REG.mem_10_4 ), .I1(\REG.mem_11_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9658));
    defparam i8116_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3221_3222 (.Q(\REG.mem_33_5 ), .C(FIFO_CLK_c), .D(n4707));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8119_3_lut (.I0(\REG.mem_14_4 ), .I1(\REG.mem_15_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9661));
    defparam i8119_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3218_3219 (.Q(\REG.mem_33_4 ), .C(FIFO_CLK_c), .D(n4706));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3215_3216 (.Q(\REG.mem_33_3 ), .C(FIFO_CLK_c), .D(n4705));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3212_3213 (.Q(\REG.mem_33_2 ), .C(FIFO_CLK_c), .D(n4704));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3209_3210 (.Q(\REG.mem_33_1 ), .C(FIFO_CLK_c), .D(n4703));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3206_3207 (.Q(\REG.mem_33_0 ), .C(FIFO_CLK_c), .D(n4702));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3155_3156 (.Q(\REG.mem_32_15 ), .C(FIFO_CLK_c), .D(n4700));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3152_3153 (.Q(\REG.mem_32_14 ), .C(FIFO_CLK_c), .D(n4698));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3149_3150 (.Q(\REG.mem_32_13 ), .C(FIFO_CLK_c), .D(n4697));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3146_3147 (.Q(\REG.mem_32_12 ), .C(FIFO_CLK_c), .D(n4696));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3143_3144 (.Q(\REG.mem_32_11 ), .C(FIFO_CLK_c), .D(n4695));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3140_3141 (.Q(\REG.mem_32_10 ), .C(FIFO_CLK_c), .D(n4694));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3137_3138 (.Q(\REG.mem_32_9 ), .C(FIFO_CLK_c), .D(n4693));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i167_168 (.Q(\REG.mem_1_11 ), .C(FIFO_CLK_c), .D(n4149));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 wp_sync2_r_6__I_0_127_inv_0_i7_1_lut (.I0(\rd_addr_r[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // src/fifo_dc_32_lut_gen.v(231[47:78])
    defparam wp_sync2_r_6__I_0_127_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3096_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_3_15 ), .O(n4185));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3096_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i164_165 (.Q(\REG.mem_1_10 ), .C(FIFO_CLK_c), .D(n4148));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9635 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_9 ), 
            .I2(\REG.mem_59_9 ), .I3(rd_addr_r[1]), .O(n11268));
    defparam rd_addr_r_0__bdd_4_lut_9635.LUT_INIT = 16'he4aa;
    SB_LUT4 i3095_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_3_14 ), .O(n4184));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3095_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8118_3_lut (.I0(\REG.mem_12_4 ), .I1(\REG.mem_13_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9660));
    defparam i8118_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3134_3135 (.Q(\REG.mem_32_8 ), .C(FIFO_CLK_c), .D(n4692));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11268_bdd_4_lut (.I0(n11268), .I1(\REG.mem_57_9 ), .I2(\REG.mem_56_9 ), 
            .I3(rd_addr_r[1]), .O(n11271));
    defparam n11268_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8364_3_lut (.I0(\REG.mem_0_1 ), .I1(\REG.mem_1_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9906));
    defparam i8364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8365_3_lut (.I0(\REG.mem_2_1 ), .I1(\REG.mem_3_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9907));
    defparam i8365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8374_3_lut (.I0(\REG.mem_6_1 ), .I1(\REG.mem_7_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9916));
    defparam i8374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3094_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_3_13 ), .O(n4183));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3094_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8373_3_lut (.I0(\REG.mem_4_1 ), .I1(\REG.mem_5_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9915));
    defparam i8373_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3131_3132 (.Q(\REG.mem_32_7 ), .C(FIFO_CLK_c), .D(n4691));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8397_3_lut (.I0(\REG.mem_16_1 ), .I1(\REG.mem_17_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9939));
    defparam i8397_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3128_3129 (.Q(\REG.mem_32_6 ), .C(FIFO_CLK_c), .D(n4690));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3125_3126 (.Q(\REG.mem_32_5 ), .C(FIFO_CLK_c), .D(n4689));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3122_3123 (.Q(\REG.mem_32_4 ), .C(FIFO_CLK_c), .D(n4688));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3119_3120 (.Q(\REG.mem_32_3 ), .C(FIFO_CLK_c), .D(n4687));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3116_3117 (.Q(\REG.mem_32_2 ), .C(FIFO_CLK_c), .D(n4686));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3113_3114 (.Q(\REG.mem_32_1 ), .C(FIFO_CLK_c), .D(n4685));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3110_3111 (.Q(\REG.mem_32_0 ), .C(FIFO_CLK_c), .D(n4684));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF rp_sync1_r__i1 (.Q(rp_sync1_r[1]), .C(FIFO_CLK_c), .D(n4677));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9234 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_9 ), 
            .I2(\REG.mem_63_9 ), .I3(rd_addr_r[1]), .O(n10776));
    defparam rd_addr_r_0__bdd_4_lut_9234.LUT_INIT = 16'he4aa;
    SB_LUT4 i3093_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_3_12 ), .O(n4182));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3093_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3092_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_3_11 ), .O(n4181));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3092_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_6__I_0_129_8_lut (.I0(GND_net), .I1(\rd_addr_r[6] ), 
            .I2(GND_net), .I3(n8729), .O(rd_addr_p1_w[6])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_129_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9630 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_10 ), 
            .I2(\REG.mem_27_10 ), .I3(rd_addr_r[1]), .O(n11262));
    defparam rd_addr_r_0__bdd_4_lut_9630.LUT_INIT = 16'he4aa;
    SB_LUT4 i8398_3_lut (.I0(\REG.mem_18_1 ), .I1(\REG.mem_19_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9940));
    defparam i8398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10379 (.I0(rd_addr_r[4]), .I1(n10346), 
            .I2(n10382), .I3(rd_addr_r[5]), .O(n11904));
    defparam rd_addr_r_4__bdd_4_lut_10379.LUT_INIT = 16'he4aa;
    SB_LUT4 i3091_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_3_10 ), .O(n4180));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3091_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF rp_sync1_r__i2 (.Q(rp_sync1_r[2]), .C(FIFO_CLK_c), .D(n4676));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_DFF rp_sync1_r__i3 (.Q(rp_sync1_r[3]), .C(FIFO_CLK_c), .D(n4675));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_DFF rp_sync1_r__i4 (.Q(rp_sync1_r[4]), .C(FIFO_CLK_c), .D(n4674));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_DFF rp_sync1_r__i5 (.Q(rp_sync1_r[5]), .C(FIFO_CLK_c), .D(n4673));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_DFF rp_sync1_r__i6 (.Q(rp_sync1_r[6]), .C(FIFO_CLK_c), .D(n4672));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_DFF i3059_3060 (.Q(\REG.mem_31_15 ), .C(FIFO_CLK_c), .D(n4671));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3056_3057 (.Q(\REG.mem_31_14 ), .C(FIFO_CLK_c), .D(n4670));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3053_3054 (.Q(\REG.mem_31_13 ), .C(FIFO_CLK_c), .D(n4669));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3050_3051 (.Q(\REG.mem_31_12 ), .C(FIFO_CLK_c), .D(n4668));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3047_3048 (.Q(\REG.mem_31_11 ), .C(FIFO_CLK_c), .D(n4667));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3044_3045 (.Q(\REG.mem_31_10 ), .C(FIFO_CLK_c), .D(n4666));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3041_3042 (.Q(\REG.mem_31_9 ), .C(FIFO_CLK_c), .D(n4665));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3038_3039 (.Q(\REG.mem_31_8 ), .C(FIFO_CLK_c), .D(n4664));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3035_3036 (.Q(\REG.mem_31_7 ), .C(FIFO_CLK_c), .D(n4663));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3032_3033 (.Q(\REG.mem_31_6 ), .C(FIFO_CLK_c), .D(n4662));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3029_3030 (.Q(\REG.mem_31_5 ), .C(FIFO_CLK_c), .D(n4661));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11262_bdd_4_lut (.I0(n11262), .I1(\REG.mem_25_10 ), .I2(\REG.mem_24_10 ), 
            .I3(rd_addr_r[1]), .O(n9770));
    defparam n11262_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8401_3_lut (.I0(\REG.mem_22_1 ), .I1(\REG.mem_23_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9943));
    defparam i8401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3571_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_31_4 ), .O(n4660));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3571_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11904_bdd_4_lut (.I0(n11904), .I1(n10334), .I2(n10322), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_237 [8]));
    defparam n11904_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8400_3_lut (.I0(\REG.mem_20_1 ), .I1(\REG.mem_21_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9942));
    defparam i8400_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3026_3027 (.Q(\REG.mem_31_4 ), .C(FIFO_CLK_c), .D(n4660));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i108_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n46));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i108_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i8427_3_lut (.I0(\REG.mem_32_1 ), .I1(\REG.mem_33_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9969));
    defparam i8427_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3023_3024 (.Q(\REG.mem_31_3 ), .C(FIFO_CLK_c), .D(n4659));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i107_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n14));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i107_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_DFF i3020_3021 (.Q(\REG.mem_31_2 ), .C(FIFO_CLK_c), .D(n4658));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3017_3018 (.Q(\REG.mem_31_1 ), .C(FIFO_CLK_c), .D(n4657));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i3014_3015 (.Q(\REG.mem_31_0 ), .C(FIFO_CLK_c), .D(n4656));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF rp_sync2_r__i1 (.Q(rp_sync2_r[1]), .C(FIFO_CLK_c), .D(n4655));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_DFF rp_sync2_r__i2 (.Q(rp_sync2_r[2]), .C(FIFO_CLK_c), .D(n4654));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_DFF rp_sync2_r__i3 (.Q(rp_sync2_r[3]), .C(FIFO_CLK_c), .D(n4653));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_DFF rp_sync2_r__i4 (.Q(rp_sync2_r[4]), .C(FIFO_CLK_c), .D(n4652));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_DFF rp_sync2_r__i5 (.Q(rp_sync2_r[5]), .C(FIFO_CLK_c), .D(n4651));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_DFF rp_sync2_r__i6 (.Q(rp_sync2_r[6]), .C(FIFO_CLK_c), .D(n4650));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_DFF i2963_2964 (.Q(\REG.mem_30_15 ), .C(FIFO_CLK_c), .D(n4649));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2960_2961 (.Q(\REG.mem_30_14 ), .C(FIFO_CLK_c), .D(n4648));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2957_2958 (.Q(\REG.mem_30_13 ), .C(FIFO_CLK_c), .D(n4647));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2954_2955 (.Q(\REG.mem_30_12 ), .C(FIFO_CLK_c), .D(n4646));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2951_2952 (.Q(\REG.mem_30_11 ), .C(FIFO_CLK_c), .D(n4645));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i126_2_lut_3_lut (.I0(n29), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n37));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i126_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i8428_3_lut (.I0(\REG.mem_34_1 ), .I1(\REG.mem_35_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9970));
    defparam i8428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i125_2_lut_3_lut (.I0(n29), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n5));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i125_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n10776_bdd_4_lut (.I0(n10776), .I1(\REG.mem_61_9 ), .I2(\REG.mem_60_9 ), 
            .I3(rd_addr_r[1]), .O(n10779));
    defparam n10776_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8431_3_lut (.I0(\REG.mem_38_1 ), .I1(\REG.mem_39_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9973));
    defparam i8431_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2948_2949 (.Q(\REG.mem_30_10 ), .C(FIFO_CLK_c), .D(n4644));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10164 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_6 ), 
            .I2(\REG.mem_63_6 ), .I3(rd_addr_r[1]), .O(n11898));
    defparam rd_addr_r_0__bdd_4_lut_10164.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i29_2_lut_3_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n29));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i29_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i46_2_lut_3_lut_4_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n46_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i46_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i45_2_lut_3_lut_4_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n45));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i45_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i8430_3_lut (.I0(\REG.mem_36_1 ), .I1(\REG.mem_37_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9972));
    defparam i8430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8463_3_lut (.I0(\REG.mem_48_1 ), .I1(\REG.mem_49_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10005));
    defparam i8463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8464_3_lut (.I0(\REG.mem_50_1 ), .I1(\REG.mem_51_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10006));
    defparam i8464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8751_3_lut (.I0(\REG.mem_40_13 ), .I1(\REG.mem_41_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10293));
    defparam i8751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8752_3_lut (.I0(\REG.mem_42_13 ), .I1(\REG.mem_43_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10294));
    defparam i8752_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2945_2946 (.Q(\REG.mem_30_9 ), .C(FIFO_CLK_c), .D(n4643));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2942_2943 (.Q(\REG.mem_30_8 ), .C(FIFO_CLK_c), .D(n4642));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2939_2940 (.Q(\REG.mem_30_7 ), .C(FIFO_CLK_c), .D(n4641));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2936_2937 (.Q(\REG.mem_30_6 ), .C(FIFO_CLK_c), .D(n4640));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2933_2934 (.Q(\REG.mem_30_5 ), .C(FIFO_CLK_c), .D(n4639));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2930_2931 (.Q(\REG.mem_30_4 ), .C(FIFO_CLK_c), .D(n4638));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2927_2928 (.Q(\REG.mem_30_3 ), .C(FIFO_CLK_c), .D(n4637));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2924_2925 (.Q(\REG.mem_30_2 ), .C(FIFO_CLK_c), .D(n4636));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2921_2922 (.Q(\REG.mem_30_1 ), .C(FIFO_CLK_c), .D(n4635));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2918_2919 (.Q(\REG.mem_30_0 ), .C(FIFO_CLK_c), .D(n4634));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(DEBUG_6_c), .D(n4633));   // src/fifo_dc_32_lut_gen.v(558[21] 574[24])
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r[2]), .C(DEBUG_6_c), .D(n4632));   // src/fifo_dc_32_lut_gen.v(558[21] 574[24])
    SB_DFF rd_addr_r__i3 (.Q(rd_addr_r[3]), .C(DEBUG_6_c), .D(n4631));   // src/fifo_dc_32_lut_gen.v(558[21] 574[24])
    SB_DFF rd_addr_r__i4 (.Q(rd_addr_r[4]), .C(DEBUG_6_c), .D(n4630));   // src/fifo_dc_32_lut_gen.v(558[21] 574[24])
    SB_DFF rd_addr_r__i5 (.Q(rd_addr_r[5]), .C(DEBUG_6_c), .D(n4629));   // src/fifo_dc_32_lut_gen.v(558[21] 574[24])
    SB_DFF rd_addr_r__i6 (.Q(\rd_addr_r[6] ), .C(DEBUG_6_c), .D(n4628));   // src/fifo_dc_32_lut_gen.v(558[21] 574[24])
    SB_LUT4 EnabledDecoder_2_i12_2_lut_3_lut (.I0(write_to_dc32_fifo), .I1(wr_addr_r[0]), 
            .I2(wr_addr_r[1]), .I3(GND_net), .O(n12_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i12_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i8761_3_lut (.I0(\REG.mem_46_13 ), .I1(\REG.mem_47_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10303));
    defparam i8761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i11_2_lut_3_lut (.I0(write_to_dc32_fifo), .I1(wr_addr_r[0]), 
            .I2(wr_addr_r[1]), .I3(GND_net), .O(n11_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i11_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i8760_3_lut (.I0(\REG.mem_44_13 ), .I1(\REG.mem_45_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10302));
    defparam i8760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8766_3_lut (.I0(\REG.mem_16_14 ), .I1(\REG.mem_17_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10308));
    defparam i8766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8767_3_lut (.I0(\REG.mem_18_14 ), .I1(\REG.mem_19_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10309));
    defparam i8767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8467_3_lut (.I0(\REG.mem_54_1 ), .I1(\REG.mem_55_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10009));
    defparam i8467_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2867_2868 (.Q(\REG.mem_29_15 ), .C(FIFO_CLK_c), .D(n4627));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11898_bdd_4_lut (.I0(n11898), .I1(\REG.mem_61_6 ), .I2(\REG.mem_60_6 ), 
            .I3(rd_addr_r[1]), .O(n11901));
    defparam n11898_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i98_2_lut_3_lut (.I0(n33), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n51));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i98_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_DFF i2864_2865 (.Q(\REG.mem_29_14 ), .C(FIFO_CLK_c), .D(n4626));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8466_3_lut (.I0(\REG.mem_52_1 ), .I1(\REG.mem_53_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10008));
    defparam i8466_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2861_2862 (.Q(\REG.mem_29_13 ), .C(FIFO_CLK_c), .D(n4625));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8782_3_lut (.I0(\REG.mem_22_14 ), .I1(\REG.mem_23_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10324));
    defparam i8782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8781_3_lut (.I0(\REG.mem_20_14 ), .I1(\REG.mem_21_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10323));
    defparam i8781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10154 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_12 ), 
            .I2(\REG.mem_59_12 ), .I3(rd_addr_r[1]), .O(n11892));
    defparam rd_addr_r_0__bdd_4_lut_10154.LUT_INIT = 16'he4aa;
    SB_DFF i2858_2859 (.Q(\REG.mem_29_12 ), .C(FIFO_CLK_c), .D(n4624));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2855_2856 (.Q(\REG.mem_29_11 ), .C(FIFO_CLK_c), .D(n4623));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2852_2853 (.Q(\REG.mem_29_10 ), .C(FIFO_CLK_c), .D(n4622));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2849_2850 (.Q(\REG.mem_29_9 ), .C(FIFO_CLK_c), .D(n4621));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2846_2847 (.Q(\REG.mem_29_8 ), .C(FIFO_CLK_c), .D(n4620));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2843_2844 (.Q(\REG.mem_29_7 ), .C(FIFO_CLK_c), .D(n4619));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2840_2841 (.Q(\REG.mem_29_6 ), .C(FIFO_CLK_c), .D(n4618));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2837_2838 (.Q(\REG.mem_29_5 ), .C(FIFO_CLK_c), .D(n4617));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2834_2835 (.Q(\REG.mem_29_4 ), .C(FIFO_CLK_c), .D(n4616));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2831_2832 (.Q(\REG.mem_29_3 ), .C(FIFO_CLK_c), .D(n4615));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2828_2829 (.Q(\REG.mem_29_2 ), .C(FIFO_CLK_c), .D(n4614));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2825_2826 (.Q(\REG.mem_29_1 ), .C(FIFO_CLK_c), .D(n4613));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2822_2823 (.Q(\REG.mem_29_0 ), .C(FIFO_CLK_c), .D(n4612));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2771_2772 (.Q(\REG.mem_28_15 ), .C(FIFO_CLK_c), .D(n4611));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2768_2769 (.Q(\REG.mem_28_14 ), .C(FIFO_CLK_c), .D(n4610));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2765_2766 (.Q(\REG.mem_28_13 ), .C(FIFO_CLK_c), .D(n4609));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_9685 (.I0(rd_addr_r[3]), .I1(n11223), 
            .I2(n9742), .I3(rd_addr_r[4]), .O(n11256));
    defparam rd_addr_r_3__bdd_4_lut_9685.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i97_2_lut_3_lut (.I0(n33), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n19));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i97_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i2762_2763 (.Q(\REG.mem_28_12 ), .C(FIFO_CLK_c), .D(n4608));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11892_bdd_4_lut (.I0(n11892), .I1(\REG.mem_57_12 ), .I2(\REG.mem_56_12 ), 
            .I3(rd_addr_r[1]), .O(n10013));
    defparam n11892_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11256_bdd_4_lut (.I0(n11256), .I1(n9739), .I2(n11217), .I3(rd_addr_r[4]), 
            .O(n11259));
    defparam n11256_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8304_3_lut (.I0(\REG.mem_16_12 ), .I1(\REG.mem_17_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9846));
    defparam i8304_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2759_2760 (.Q(\REG.mem_28_11 ), .C(FIFO_CLK_c), .D(n4607));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i4071_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_59_15 ), .O(n5160));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4071_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9775 (.I0(rd_addr_r[2]), .I1(n9494), 
            .I2(n11109), .I3(rd_addr_r[3]), .O(n11250));
    defparam rd_addr_r_2__bdd_4_lut_9775.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10264 (.I0(rd_addr_r[3]), .I1(n11475), 
            .I2(n9997), .I3(rd_addr_r[4]), .O(n11886));
    defparam rd_addr_r_3__bdd_4_lut_10264.LUT_INIT = 16'he4aa;
    SB_LUT4 n11886_bdd_4_lut (.I0(n11886), .I1(n9985), .I2(n9984), .I3(rd_addr_r[4]), 
            .O(n11889));
    defparam n11886_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8305_3_lut (.I0(\REG.mem_18_12 ), .I1(\REG.mem_19_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9847));
    defparam i8305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4070_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_59_14 ), .O(n5159));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4070_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8326_3_lut (.I0(\REG.mem_22_12 ), .I1(\REG.mem_23_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9868));
    defparam i8326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4069_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_59_13 ), .O(n5158));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4069_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11250_bdd_4_lut (.I0(n11250), .I1(n10523), .I2(n10511), .I3(rd_addr_r[3]), 
            .O(n11253));
    defparam n11250_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2756_2757 (.Q(\REG.mem_28_10 ), .C(FIFO_CLK_c), .D(n4606));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10194 (.I0(rd_addr_r[1]), .I1(n9921), 
            .I2(n9922), .I3(rd_addr_r[2]), .O(n11880));
    defparam rd_addr_r_1__bdd_4_lut_10194.LUT_INIT = 16'he4aa;
    SB_DFF i2753_2754 (.Q(\REG.mem_28_9 ), .C(FIFO_CLK_c), .D(n4605));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2750_2751 (.Q(\REG.mem_28_8 ), .C(FIFO_CLK_c), .D(n4604));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2747_2748 (.Q(\REG.mem_28_7 ), .C(FIFO_CLK_c), .D(n4603));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2744_2745 (.Q(\REG.mem_28_6 ), .C(FIFO_CLK_c), .D(n4602));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2741_2742 (.Q(\REG.mem_28_5 ), .C(FIFO_CLK_c), .D(n4601));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2738_2739 (.Q(\REG.mem_28_4 ), .C(FIFO_CLK_c), .D(n4600));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2735_2736 (.Q(\REG.mem_28_3 ), .C(FIFO_CLK_c), .D(n4599));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2732_2733 (.Q(\REG.mem_28_2 ), .C(FIFO_CLK_c), .D(n4598));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2729_2730 (.Q(\REG.mem_28_1 ), .C(FIFO_CLK_c), .D(n4597));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2726_2727 (.Q(\REG.mem_28_0 ), .C(FIFO_CLK_c), .D(n4596));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2675_2676 (.Q(\REG.mem_27_15 ), .C(FIFO_CLK_c), .D(n4595));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2672_2673 (.Q(\REG.mem_27_14 ), .C(FIFO_CLK_c), .D(n4594));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2669_2670 (.Q(\REG.mem_27_13 ), .C(FIFO_CLK_c), .D(n4593));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2666_2667 (.Q(\REG.mem_27_12 ), .C(FIFO_CLK_c), .D(n4592));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2663_2664 (.Q(\REG.mem_27_11 ), .C(FIFO_CLK_c), .D(n4591));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8325_3_lut (.I0(\REG.mem_20_12 ), .I1(\REG.mem_21_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9867));
    defparam i8325_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2660_2661 (.Q(\REG.mem_27_10 ), .C(FIFO_CLK_c), .D(n4590));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8337_3_lut (.I0(n11403), .I1(n11181), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9879));
    defparam i8337_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2657_2658 (.Q(\REG.mem_27_9 ), .C(FIFO_CLK_c), .D(n4589));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2654_2655 (.Q(\REG.mem_27_8 ), .C(FIFO_CLK_c), .D(n4588));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2651_2652 (.Q(\REG.mem_27_7 ), .C(FIFO_CLK_c), .D(n4587));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8338_3_lut (.I0(n11133), .I1(n10923), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9880));
    defparam i8338_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2648_2649 (.Q(\REG.mem_27_6 ), .C(FIFO_CLK_c), .D(n4586));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11880_bdd_4_lut (.I0(n11880), .I1(n9892), .I2(n9891), .I3(rd_addr_r[2]), 
            .O(n10317));
    defparam n11880_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9675 (.I0(rd_addr_r[1]), .I1(n9717), 
            .I2(n9718), .I3(rd_addr_r[2]), .O(n11244));
    defparam rd_addr_r_1__bdd_4_lut_9675.LUT_INIT = 16'he4aa;
    SB_LUT4 i4068_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_59_12 ), .O(n5157));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4068_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2645_2646 (.Q(\REG.mem_27_5 ), .C(FIFO_CLK_c), .D(n4585));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8352_3_lut (.I0(n10755), .I1(n10725), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9894));
    defparam i8352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8307_3_lut (.I0(\REG.mem_56_0 ), .I1(\REG.mem_57_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9849));
    defparam i8307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8308_3_lut (.I0(\REG.mem_58_0 ), .I1(\REG.mem_59_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9850));
    defparam i8308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8311_3_lut (.I0(\REG.mem_62_0 ), .I1(\REG.mem_63_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9853));
    defparam i8311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8310_3_lut (.I0(\REG.mem_60_0 ), .I1(\REG.mem_61_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9852));
    defparam i8310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4067_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_59_11 ), .O(n5156));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4067_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11244_bdd_4_lut (.I0(n11244), .I1(n9715), .I2(n9714), .I3(rd_addr_r[2]), 
            .O(n11247));
    defparam n11244_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2642_2643 (.Q(\REG.mem_27_4 ), .C(FIFO_CLK_c), .D(n4584));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10149 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_14 ), 
            .I2(\REG.mem_59_14 ), .I3(rd_addr_r[1]), .O(n11874));
    defparam rd_addr_r_0__bdd_4_lut_10149.LUT_INIT = 16'he4aa;
    SB_DFF i2639_2640 (.Q(\REG.mem_27_3 ), .C(FIFO_CLK_c), .D(n4583));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2636_2637 (.Q(\REG.mem_27_2 ), .C(FIFO_CLK_c), .D(n4582));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2633_2634 (.Q(\REG.mem_27_1 ), .C(FIFO_CLK_c), .D(n4581));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2630_2631 (.Q(\REG.mem_27_0 ), .C(FIFO_CLK_c), .D(n4580));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2579_2580 (.Q(\REG.mem_26_15 ), .C(FIFO_CLK_c), .D(n4579));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2576_2577 (.Q(\REG.mem_26_14 ), .C(FIFO_CLK_c), .D(n4578));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2573_2574 (.Q(\REG.mem_26_13 ), .C(FIFO_CLK_c), .D(n4577));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2570_2571 (.Q(\REG.mem_26_12 ), .C(FIFO_CLK_c), .D(n4576));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2567_2568 (.Q(\REG.mem_26_11 ), .C(FIFO_CLK_c), .D(n4575));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2564_2565 (.Q(\REG.mem_26_10 ), .C(FIFO_CLK_c), .D(n4574));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2561_2562 (.Q(\REG.mem_26_9 ), .C(FIFO_CLK_c), .D(n4573));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2558_2559 (.Q(\REG.mem_26_8 ), .C(FIFO_CLK_c), .D(n4572));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2555_2556 (.Q(\REG.mem_26_7 ), .C(FIFO_CLK_c), .D(n4571));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2552_2553 (.Q(\REG.mem_26_6 ), .C(FIFO_CLK_c), .D(n4570));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2549_2550 (.Q(\REG.mem_26_5 ), .C(FIFO_CLK_c), .D(n4569));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11874_bdd_4_lut (.I0(n11874), .I1(\REG.mem_57_14 ), .I2(\REG.mem_56_14 ), 
            .I3(rd_addr_r[1]), .O(n11877));
    defparam n11874_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4066_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_59_10 ), .O(n5155));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4066_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10134 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_9 ), 
            .I2(\REG.mem_51_9 ), .I3(rd_addr_r[1]), .O(n11868));
    defparam rd_addr_r_0__bdd_4_lut_10134.LUT_INIT = 16'he4aa;
    SB_LUT4 i4065_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_59_9 ), .O(n5154));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4065_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11868_bdd_4_lut (.I0(n11868), .I1(\REG.mem_49_9 ), .I2(\REG.mem_48_9 ), 
            .I3(rd_addr_r[1]), .O(n10022));
    defparam n11868_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9610 (.I0(rd_addr_r[1]), .I1(n9696), 
            .I2(n9697), .I3(rd_addr_r[2]), .O(n11238));
    defparam rd_addr_r_1__bdd_4_lut_9610.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_r_6__I_0_114_i2_3_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(write_to_dc32_fifo), .I3(GND_net), .O(\wr_addr_nxt_c[1] ));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam wr_addr_r_6__I_0_114_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10129 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_14 ), 
            .I2(\REG.mem_63_14 ), .I3(rd_addr_r[1]), .O(n11862));
    defparam rd_addr_r_0__bdd_4_lut_10129.LUT_INIT = 16'he4aa;
    SB_LUT4 n11862_bdd_4_lut (.I0(n11862), .I1(\REG.mem_61_14 ), .I2(\REG.mem_60_14 ), 
            .I3(rd_addr_r[1]), .O(n11865));
    defparam n11862_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11238_bdd_4_lut (.I0(n11238), .I1(n9694), .I2(n9693), .I3(rd_addr_r[2]), 
            .O(n11241));
    defparam n11238_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2546_2547 (.Q(\REG.mem_26_4 ), .C(FIFO_CLK_c), .D(n4568));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10124 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_10 ), 
            .I2(\REG.mem_51_10 ), .I3(rd_addr_r[1]), .O(n11856));
    defparam rd_addr_r_0__bdd_4_lut_10124.LUT_INIT = 16'he4aa;
    SB_DFF i2543_2544 (.Q(\REG.mem_26_3 ), .C(FIFO_CLK_c), .D(n4567));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9625 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_13 ), 
            .I2(\REG.mem_7_13 ), .I3(rd_addr_r[1]), .O(n11232));
    defparam rd_addr_r_0__bdd_4_lut_9625.LUT_INIT = 16'he4aa;
    SB_DFF i2540_2541 (.Q(\REG.mem_26_2 ), .C(FIFO_CLK_c), .D(n4566));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2537_2538 (.Q(\REG.mem_26_1 ), .C(FIFO_CLK_c), .D(n4565));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2534_2535 (.Q(\REG.mem_26_0 ), .C(FIFO_CLK_c), .D(n4564));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF wp_sync1_r__i1 (.Q(wp_sync1_r[1]), .C(DEBUG_6_c), .D(n4563));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_DFF wp_sync1_r__i2 (.Q(wp_sync1_r[2]), .C(DEBUG_6_c), .D(n4562));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_DFF wp_sync1_r__i3 (.Q(wp_sync1_r[3]), .C(DEBUG_6_c), .D(n4561));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_DFF wp_sync1_r__i4 (.Q(wp_sync1_r[4]), .C(DEBUG_6_c), .D(n4560));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_DFF i2483_2484 (.Q(\REG.mem_25_15 ), .C(FIFO_CLK_c), .D(n4559));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF wp_sync1_r__i5 (.Q(wp_sync1_r[5]), .C(DEBUG_6_c), .D(n4558));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_DFF i2480_2481 (.Q(\REG.mem_25_14 ), .C(FIFO_CLK_c), .D(n4557));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2477_2478 (.Q(\REG.mem_25_13 ), .C(FIFO_CLK_c), .D(n4556));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2474_2475 (.Q(\REG.mem_25_12 ), .C(FIFO_CLK_c), .D(n4555));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2471_2472 (.Q(\REG.mem_25_11 ), .C(FIFO_CLK_c), .D(n4554));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2468_2469 (.Q(\REG.mem_25_10 ), .C(FIFO_CLK_c), .D(n4553));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2465_2466 (.Q(\REG.mem_25_9 ), .C(FIFO_CLK_c), .D(n4552));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11856_bdd_4_lut (.I0(n11856), .I1(\REG.mem_49_10 ), .I2(\REG.mem_48_10 ), 
            .I3(rd_addr_r[1]), .O(n10025));
    defparam n11856_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2462_2463 (.Q(\REG.mem_25_8 ), .C(FIFO_CLK_c), .D(n4551));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11232_bdd_4_lut (.I0(n11232), .I1(\REG.mem_5_13 ), .I2(\REG.mem_4_13 ), 
            .I3(rd_addr_r[1]), .O(n11235));
    defparam n11232_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut (.I0(wp_sync2_r[1]), .I1(wp_sync_w[2]), .I2(GND_net), 
            .I3(GND_net), .O(wp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(537[38:77])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9600 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_3 ), 
            .I2(\REG.mem_35_3 ), .I3(rd_addr_r[1]), .O(n11226));
    defparam rd_addr_r_0__bdd_4_lut_9600.LUT_INIT = 16'he4aa;
    SB_LUT4 n11226_bdd_4_lut (.I0(n11226), .I1(\REG.mem_33_3 ), .I2(\REG.mem_32_3 ), 
            .I3(rd_addr_r[1]), .O(n11229));
    defparam n11226_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_27 (.I0(wp_sync2_r[6]), .I1(wp_sync2_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n3571));   // src/fifo_dc_32_lut_gen.v(537[38:77])
    defparam i1_2_lut_adj_27.LUT_INIT = 16'h6666;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10119 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_15 ), 
            .I2(\REG.mem_35_15 ), .I3(rd_addr_r[1]), .O(n11838));
    defparam rd_addr_r_0__bdd_4_lut_10119.LUT_INIT = 16'he4aa;
    SB_LUT4 n11838_bdd_4_lut (.I0(n11838), .I1(\REG.mem_33_15 ), .I2(\REG.mem_32_15 ), 
            .I3(rd_addr_r[1]), .O(n11841));
    defparam n11838_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2459_2460 (.Q(\REG.mem_25_7 ), .C(FIFO_CLK_c), .D(n4550));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i7846_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_r[4]), .I2(wp_sync_w[0]), 
            .I3(wp_sync_w[4]), .O(n9386));
    defparam i7846_4_lut.LUT_INIT = 16'h7bde;
    SB_DFF i2456_2457 (.Q(\REG.mem_25_6 ), .C(FIFO_CLK_c), .D(n4549));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2453_2454 (.Q(\REG.mem_25_5 ), .C(FIFO_CLK_c), .D(n4548));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2450_2451 (.Q(\REG.mem_25_4 ), .C(FIFO_CLK_c), .D(n4547));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2447_2448 (.Q(\REG.mem_25_3 ), .C(FIFO_CLK_c), .D(n4546));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2444_2445 (.Q(\REG.mem_25_2 ), .C(FIFO_CLK_c), .D(n4545));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2441_2442 (.Q(\REG.mem_25_1 ), .C(FIFO_CLK_c), .D(n4544));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2438_2439 (.Q(\REG.mem_25_0 ), .C(FIFO_CLK_c), .D(n4543));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF wp_sync1_r__i6 (.Q(wp_sync1_r[6]), .C(DEBUG_6_c), .D(n4542));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_DFF wp_sync2_r__i1 (.Q(wp_sync2_r[1]), .C(DEBUG_6_c), .D(n4541));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_DFF wp_sync2_r__i2 (.Q(wp_sync2_r[2]), .C(DEBUG_6_c), .D(n4540));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_DFF wp_sync2_r__i3 (.Q(wp_sync2_r[3]), .C(DEBUG_6_c), .D(n4539));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_DFF wp_sync2_r__i4 (.Q(wp_sync2_r[4]), .C(DEBUG_6_c), .D(n4538));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_DFF wp_sync2_r__i5 (.Q(wp_sync2_r[5]), .C(DEBUG_6_c), .D(n4537));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_DFF wp_sync2_r__i6 (.Q(wp_sync2_r[6]), .C(DEBUG_6_c), .D(n4536));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_DFF i2387_2388 (.Q(\REG.mem_24_15 ), .C(FIFO_CLK_c), .D(n4535));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8139_3_lut (.I0(\REG.mem_16_0 ), .I1(\REG.mem_17_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9681));
    defparam i8139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7842_4_lut (.I0(rd_addr_r[5]), .I1(rd_addr_r[3]), .I2(n3571), 
            .I3(wp_sync_w[3]), .O(n9382));
    defparam i7842_4_lut.LUT_INIT = 16'h7bde;
    SB_DFF i2384_2385 (.Q(\REG.mem_24_14 ), .C(FIFO_CLK_c), .D(n4534));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8140_3_lut (.I0(\REG.mem_18_0 ), .I1(\REG.mem_19_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9682));
    defparam i8140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_28 (.I0(rd_addr_p1_w[4]), .I1(wp_sync_w[4]), .I2(GND_net), 
            .I3(GND_net), .O(n3560));   // src/fifo_dc_32_lut_gen.v(537[38:77])
    defparam i1_2_lut_adj_28.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(rd_addr_p1_w[5]), .I1(rd_addr_p1_w[3]), .I2(n3571), 
            .I3(wp_sync_w[3]), .O(n10_adj_1064));   // src/fifo_dc_32_lut_gen.v(542[28:56])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut (.I0(wp_sync2_r[6]), .I1(rd_addr_p1_w[1]), .I2(rd_addr_p1_w[6]), 
            .I3(wp_sync_w[1]), .O(n8_adj_1065));   // src/fifo_dc_32_lut_gen.v(542[28:56])
    defparam i1_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i8161_3_lut (.I0(\REG.mem_22_0 ), .I1(\REG.mem_23_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9703));
    defparam i8161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut (.I0(rd_addr_p1_w[0]), .I1(n10_adj_1064), .I2(n3560), 
            .I3(wp_sync_w[0]), .O(n12_adj_1066));   // src/fifo_dc_32_lut_gen.v(542[28:56])
    defparam i5_4_lut.LUT_INIT = 16'hfdfe;
    SB_LUT4 i7936_3_lut (.I0(n9378), .I1(n9382), .I2(n9386), .I3(GND_net), 
            .O(n9478));
    defparam i7936_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut (.I0(rd_addr_p1_w[2]), .I1(n12_adj_1066), .I2(n8_adj_1065), 
            .I3(wp_sync_w[2]), .O(n8847));   // src/fifo_dc_32_lut_gen.v(542[28:56])
    defparam i6_4_lut.LUT_INIT = 16'hfdfe;
    SB_LUT4 i8160_3_lut (.I0(\REG.mem_20_0 ), .I1(\REG.mem_21_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9702));
    defparam i8160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 empty_nxt_c_I_10_4_lut (.I0(n8847), .I1(n9478), .I2(DEBUG_1_c), 
            .I3(DEBUG_9_c), .O(empty_nxt_c_N_306));   // src/fifo_dc_32_lut_gen.v(553[46:103])
    defparam empty_nxt_c_I_10_4_lut.LUT_INIT = 16'h3530;
    SB_DFF i2381_2382 (.Q(\REG.mem_24_13 ), .C(FIFO_CLK_c), .D(n4533));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2378_2379 (.Q(\REG.mem_24_12 ), .C(FIFO_CLK_c), .D(n4532));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2375_2376 (.Q(\REG.mem_24_11 ), .C(FIFO_CLK_c), .D(n4531));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2372_2373 (.Q(\REG.mem_24_10 ), .C(FIFO_CLK_c), .D(n4530));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2369_2370 (.Q(\REG.mem_24_9 ), .C(FIFO_CLK_c), .D(n4529));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2366_2367 (.Q(\REG.mem_24_8 ), .C(FIFO_CLK_c), .D(n4528));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2363_2364 (.Q(\REG.mem_24_7 ), .C(FIFO_CLK_c), .D(n4527));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2360_2361 (.Q(\REG.mem_24_6 ), .C(FIFO_CLK_c), .D(n4526));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2357_2358 (.Q(\REG.mem_24_5 ), .C(FIFO_CLK_c), .D(n4525));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2354_2355 (.Q(\REG.mem_24_4 ), .C(FIFO_CLK_c), .D(n4524));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2351_2352 (.Q(\REG.mem_24_3 ), .C(FIFO_CLK_c), .D(n4523));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2348_2349 (.Q(\REG.mem_24_2 ), .C(FIFO_CLK_c), .D(n4522));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2345_2346 (.Q(\REG.mem_24_1 ), .C(FIFO_CLK_c), .D(n4521));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2342_2343 (.Q(\REG.mem_24_0 ), .C(FIFO_CLK_c), .D(n4520));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2291_2292 (.Q(\REG.mem_23_15 ), .C(FIFO_CLK_c), .D(n4519));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2288_2289 (.Q(\REG.mem_23_14 ), .C(FIFO_CLK_c), .D(n4518));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9605 (.I0(rd_addr_r[1]), .I1(n9669), 
            .I2(n9670), .I3(rd_addr_r[2]), .O(n11220));
    defparam rd_addr_r_1__bdd_4_lut_9605.LUT_INIT = 16'he4aa;
    SB_LUT4 n11220_bdd_4_lut (.I0(n11220), .I1(n9667), .I2(n9666), .I3(rd_addr_r[2]), 
            .O(n11223));
    defparam n11220_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2285_2286 (.Q(\REG.mem_23_13 ), .C(FIFO_CLK_c), .D(n4517));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2282_2283 (.Q(\REG.mem_23_12 ), .C(FIFO_CLK_c), .D(n4516));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2279_2280 (.Q(\REG.mem_23_11 ), .C(FIFO_CLK_c), .D(n4515));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2276_2277 (.Q(\REG.mem_23_10 ), .C(FIFO_CLK_c), .D(n4514));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2273_2274 (.Q(\REG.mem_23_9 ), .C(FIFO_CLK_c), .D(n4513));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2270_2271 (.Q(\REG.mem_23_8 ), .C(FIFO_CLK_c), .D(n4512));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2267_2268 (.Q(\REG.mem_23_7 ), .C(FIFO_CLK_c), .D(n4511));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2264_2265 (.Q(\REG.mem_23_6 ), .C(FIFO_CLK_c), .D(n4510));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2261_2262 (.Q(\REG.mem_23_5 ), .C(FIFO_CLK_c), .D(n4509));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2258_2259 (.Q(\REG.mem_23_4 ), .C(FIFO_CLK_c), .D(n4508));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i4064_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_59_8 ), .O(n5153));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4064_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2255_2256 (.Q(\REG.mem_23_3 ), .C(FIFO_CLK_c), .D(n4507));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2252_2253 (.Q(\REG.mem_23_2 ), .C(FIFO_CLK_c), .D(n4506));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2249_2250 (.Q(\REG.mem_23_1 ), .C(FIFO_CLK_c), .D(n4505));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2246_2247 (.Q(\REG.mem_23_0 ), .C(FIFO_CLK_c), .D(n4504));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2195_2196 (.Q(\REG.mem_22_15 ), .C(FIFO_CLK_c), .D(n4503));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2192_2193 (.Q(\REG.mem_22_14 ), .C(FIFO_CLK_c), .D(n4502));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2189_2190 (.Q(\REG.mem_22_13 ), .C(FIFO_CLK_c), .D(n4501));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2186_2187 (.Q(\REG.mem_22_12 ), .C(FIFO_CLK_c), .D(n4500));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2183_2184 (.Q(\REG.mem_22_11 ), .C(FIFO_CLK_c), .D(n4499));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2180_2181 (.Q(\REG.mem_22_10 ), .C(FIFO_CLK_c), .D(n4498));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2177_2178 (.Q(\REG.mem_22_9 ), .C(FIFO_CLK_c), .D(n4497));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2174_2175 (.Q(\REG.mem_22_8 ), .C(FIFO_CLK_c), .D(n4496));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2171_2172 (.Q(\REG.mem_22_7 ), .C(FIFO_CLK_c), .D(n4495));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2168_2169 (.Q(\REG.mem_22_6 ), .C(FIFO_CLK_c), .D(n4494));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2165_2166 (.Q(\REG.mem_22_5 ), .C(FIFO_CLK_c), .D(n4493));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2162_2163 (.Q(\REG.mem_22_4 ), .C(FIFO_CLK_c), .D(n4492));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2159_2160 (.Q(\REG.mem_22_3 ), .C(FIFO_CLK_c), .D(n4491));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2156_2157 (.Q(\REG.mem_22_2 ), .C(FIFO_CLK_c), .D(n4490));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2153_2154 (.Q(\REG.mem_22_1 ), .C(FIFO_CLK_c), .D(n4489));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10104 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_9 ), 
            .I2(\REG.mem_3_9 ), .I3(rd_addr_r[1]), .O(n11826));
    defparam rd_addr_r_0__bdd_4_lut_10104.LUT_INIT = 16'he4aa;
    SB_LUT4 i4063_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_59_7 ), .O(n5152));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4063_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11826_bdd_4_lut (.I0(n11826), .I1(\REG.mem_1_9 ), .I2(\REG.mem_0_9 ), 
            .I3(rd_addr_r[1]), .O(n11829));
    defparam n11826_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4062_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_59_6 ), .O(n5151));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4062_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9590 (.I0(rd_addr_r[1]), .I1(n9648), 
            .I2(n9649), .I3(rd_addr_r[2]), .O(n11214));
    defparam rd_addr_r_1__bdd_4_lut_9590.LUT_INIT = 16'he4aa;
    SB_LUT4 i4061_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_59_5 ), .O(n5150));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4061_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2150_2151 (.Q(\REG.mem_22_0 ), .C(FIFO_CLK_c), .D(n4488));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2099_2100 (.Q(\REG.mem_21_15 ), .C(FIFO_CLK_c), .D(n4487));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2096_2097 (.Q(\REG.mem_21_14 ), .C(FIFO_CLK_c), .D(n4486));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2093_2094 (.Q(\REG.mem_21_13 ), .C(FIFO_CLK_c), .D(n4485));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2090_2091 (.Q(\REG.mem_21_12 ), .C(FIFO_CLK_c), .D(n4484));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2087_2088 (.Q(\REG.mem_21_11 ), .C(FIFO_CLK_c), .D(n4483));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2084_2085 (.Q(\REG.mem_21_10 ), .C(FIFO_CLK_c), .D(n4482));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2081_2082 (.Q(\REG.mem_21_9 ), .C(FIFO_CLK_c), .D(n4481));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2078_2079 (.Q(\REG.mem_21_8 ), .C(FIFO_CLK_c), .D(n4480));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2075_2076 (.Q(\REG.mem_21_7 ), .C(FIFO_CLK_c), .D(n4479));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2072_2073 (.Q(\REG.mem_21_6 ), .C(FIFO_CLK_c), .D(n4478));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2069_2070 (.Q(\REG.mem_21_5 ), .C(FIFO_CLK_c), .D(n4477));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2066_2067 (.Q(\REG.mem_21_4 ), .C(FIFO_CLK_c), .D(n4476));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2063_2064 (.Q(\REG.mem_21_3 ), .C(FIFO_CLK_c), .D(n4475));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2060_2061 (.Q(\REG.mem_21_2 ), .C(FIFO_CLK_c), .D(n4474));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2057_2058 (.Q(\REG.mem_21_1 ), .C(FIFO_CLK_c), .D(n4473));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10095 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_8 ), 
            .I2(\REG.mem_3_8 ), .I3(rd_addr_r[1]), .O(n11820));
    defparam rd_addr_r_0__bdd_4_lut_10095.LUT_INIT = 16'he4aa;
    SB_LUT4 n11214_bdd_4_lut (.I0(n11214), .I1(n9646), .I2(n9645), .I3(rd_addr_r[2]), 
            .O(n11217));
    defparam n11214_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11820_bdd_4_lut (.I0(n11820), .I1(\REG.mem_1_8 ), .I2(\REG.mem_0_8 ), 
            .I3(rd_addr_r[1]), .O(n11823));
    defparam n11820_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8295_3_lut (.I0(\REG.mem_40_7 ), .I1(\REG.mem_41_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9837));
    defparam i8295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8296_3_lut (.I0(\REG.mem_42_7 ), .I1(\REG.mem_43_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9838));
    defparam i8296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10090 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_5 ), 
            .I2(\REG.mem_47_5 ), .I3(rd_addr_r[1]), .O(n11814));
    defparam rd_addr_r_0__bdd_4_lut_10090.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9595 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_12 ), 
            .I2(\REG.mem_7_12 ), .I3(rd_addr_r[1]), .O(n11208));
    defparam rd_addr_r_0__bdd_4_lut_9595.LUT_INIT = 16'he4aa;
    SB_LUT4 i8317_3_lut (.I0(\REG.mem_46_7 ), .I1(\REG.mem_47_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9859));
    defparam i8317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11814_bdd_4_lut (.I0(n11814), .I1(\REG.mem_45_5 ), .I2(\REG.mem_44_5 ), 
            .I3(rd_addr_r[1]), .O(n10454));
    defparam n11814_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8316_3_lut (.I0(\REG.mem_44_7 ), .I1(\REG.mem_45_7 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9858));
    defparam i8316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4060_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_59_4 ), .O(n5149));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4060_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10085 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_12 ), 
            .I2(\REG.mem_63_12 ), .I3(rd_addr_r[1]), .O(n11808));
    defparam rd_addr_r_0__bdd_4_lut_10085.LUT_INIT = 16'he4aa;
    SB_DFF i2054_2055 (.Q(\REG.mem_21_0 ), .C(FIFO_CLK_c), .D(n4472));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2003_2004 (.Q(\REG.mem_20_15 ), .C(FIFO_CLK_c), .D(n4471));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i2000_2001 (.Q(\REG.mem_20_14 ), .C(FIFO_CLK_c), .D(n4470));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1997_1998 (.Q(\REG.mem_20_13 ), .C(FIFO_CLK_c), .D(n4469));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1994_1995 (.Q(\REG.mem_20_12 ), .C(FIFO_CLK_c), .D(n4468));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1991_1992 (.Q(\REG.mem_20_11 ), .C(FIFO_CLK_c), .D(n4467));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1988_1989 (.Q(\REG.mem_20_10 ), .C(FIFO_CLK_c), .D(n4466));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1985_1986 (.Q(\REG.mem_20_9 ), .C(FIFO_CLK_c), .D(n4465));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1982_1983 (.Q(\REG.mem_20_8 ), .C(FIFO_CLK_c), .D(n4464));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1979_1980 (.Q(\REG.mem_20_7 ), .C(FIFO_CLK_c), .D(n4463));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1976_1977 (.Q(\REG.mem_20_6 ), .C(FIFO_CLK_c), .D(n4462));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1973_1974 (.Q(\REG.mem_20_5 ), .C(FIFO_CLK_c), .D(n4461));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1970_1971 (.Q(\REG.mem_20_4 ), .C(FIFO_CLK_c), .D(n4460));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1967_1968 (.Q(\REG.mem_20_3 ), .C(FIFO_CLK_c), .D(n4459));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1964_1965 (.Q(\REG.mem_20_2 ), .C(FIFO_CLK_c), .D(n4458));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1961_1962 (.Q(\REG.mem_20_1 ), .C(FIFO_CLK_c), .D(n4457));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i4059_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_59_3 ), .O(n5148));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4059_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4058_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_59_2 ), .O(n5147));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4058_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i161_162 (.Q(\REG.mem_1_9 ), .C(FIFO_CLK_c), .D(n4147));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFFE \REG.out_raw__i16  (.Q(\REG.out_raw[15] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [15]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFFE \REG.out_raw__i15  (.Q(\REG.out_raw[14] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [14]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_LUT4 i4057_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_59_1 ), .O(n5146));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4057_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE \REG.out_raw__i14  (.Q(\REG.out_raw[13] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [13]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFF i1958_1959 (.Q(\REG.mem_20_0 ), .C(FIFO_CLK_c), .D(n4456));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i4056_3_lut_4_lut (.I0(n59_adj_1060), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_59_0 ), .O(n5145));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4056_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11208_bdd_4_lut (.I0(n11208), .I1(\REG.mem_5_12 ), .I2(\REG.mem_4_12 ), 
            .I3(rd_addr_r[1]), .O(n11211));
    defparam n11208_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i158_159 (.Q(\REG.mem_1_8 ), .C(FIFO_CLK_c), .D(n4146));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_6__I_0_i2_3_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1_w[1]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_176[1] ));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam rd_addr_r_6__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE \REG.out_raw__i13  (.Q(\REG.out_raw[12] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [12]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFFE \REG.out_raw__i12  (.Q(\REG.out_raw[11] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [11]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFFE \REG.out_raw__i11  (.Q(\REG.out_raw[10] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [10]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFF i1907_1908 (.Q(\REG.mem_19_15 ), .C(FIFO_CLK_c), .D(n4455));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1904_1905 (.Q(\REG.mem_19_14 ), .C(FIFO_CLK_c), .D(n4454));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1901_1902 (.Q(\REG.mem_19_13 ), .C(FIFO_CLK_c), .D(n4453));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1898_1899 (.Q(\REG.mem_19_12 ), .C(FIFO_CLK_c), .D(n4452));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1895_1896 (.Q(\REG.mem_19_11 ), .C(FIFO_CLK_c), .D(n4451));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1892_1893 (.Q(\REG.mem_19_10 ), .C(FIFO_CLK_c), .D(n4450));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1889_1890 (.Q(\REG.mem_19_9 ), .C(FIFO_CLK_c), .D(n4449));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1886_1887 (.Q(\REG.mem_19_8 ), .C(FIFO_CLK_c), .D(n4448));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1883_1884 (.Q(\REG.mem_19_7 ), .C(FIFO_CLK_c), .D(n4447));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1880_1881 (.Q(\REG.mem_19_6 ), .C(FIFO_CLK_c), .D(n4446));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1877_1878 (.Q(\REG.mem_19_5 ), .C(FIFO_CLK_c), .D(n4445));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1874_1875 (.Q(\REG.mem_19_4 ), .C(FIFO_CLK_c), .D(n4444));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1871_1872 (.Q(\REG.mem_19_3 ), .C(FIFO_CLK_c), .D(n4443));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1868_1869 (.Q(\REG.mem_19_2 ), .C(FIFO_CLK_c), .D(n4442));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1865_1866 (.Q(\REG.mem_19_1 ), .C(FIFO_CLK_c), .D(n4441));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1862_1863 (.Q(\REG.mem_19_0 ), .C(FIFO_CLK_c), .D(n4440));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFFE \REG.out_raw__i10  (.Q(\REG.out_raw[9] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [9]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFFE \REG.out_raw__i9  (.Q(\REG.out_raw[8] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [8]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFF i1811_1812 (.Q(\REG.mem_18_15 ), .C(FIFO_CLK_c), .D(n4439));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFFE \REG.out_raw__i8  (.Q(\REG.out_raw[7] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [7]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_LUT4 n11808_bdd_4_lut (.I0(n11808), .I1(\REG.mem_61_12 ), .I2(\REG.mem_60_12 ), 
            .I3(rd_addr_r[1]), .O(n10037));
    defparam n11808_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \REG.out_raw__i7  (.Q(\REG.out_raw[6] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [6]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFFE \REG.out_raw__i6  (.Q(\REG.out_raw[5] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [5]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFFE \REG.out_raw__i5  (.Q(\REG.out_raw[4] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [4]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFFE \REG.out_raw__i4  (.Q(\REG.out_raw[3] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [3]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFF i1808_1809 (.Q(\REG.mem_18_14 ), .C(FIFO_CLK_c), .D(n4438));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10080 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_9 ), 
            .I2(\REG.mem_7_9 ), .I3(rd_addr_r[1]), .O(n11802));
    defparam rd_addr_r_0__bdd_4_lut_10080.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i92_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n54));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i92_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 n11802_bdd_4_lut (.I0(n11802), .I1(\REG.mem_5_9 ), .I2(\REG.mem_4_9 ), 
            .I3(rd_addr_r[1]), .O(n11805));
    defparam n11802_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9580 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_2 ), 
            .I2(\REG.mem_39_2 ), .I3(rd_addr_r[1]), .O(n11202));
    defparam rd_addr_r_0__bdd_4_lut_9580.LUT_INIT = 16'he4aa;
    SB_DFF i1805_1806 (.Q(\REG.mem_18_13 ), .C(FIFO_CLK_c), .D(n4437));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1802_1803 (.Q(\REG.mem_18_12 ), .C(FIFO_CLK_c), .D(n4436));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1799_1800 (.Q(\REG.mem_18_11 ), .C(FIFO_CLK_c), .D(n4435));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1796_1797 (.Q(\REG.mem_18_10 ), .C(FIFO_CLK_c), .D(n4434));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1793_1794 (.Q(\REG.mem_18_9 ), .C(FIFO_CLK_c), .D(n4433));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1790_1791 (.Q(\REG.mem_18_8 ), .C(FIFO_CLK_c), .D(n4432));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1787_1788 (.Q(\REG.mem_18_7 ), .C(FIFO_CLK_c), .D(n4431));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1784_1785 (.Q(\REG.mem_18_6 ), .C(FIFO_CLK_c), .D(n4430));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1781_1782 (.Q(\REG.mem_18_5 ), .C(FIFO_CLK_c), .D(n4429));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1778_1779 (.Q(\REG.mem_18_4 ), .C(FIFO_CLK_c), .D(n4428));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1775_1776 (.Q(\REG.mem_18_3 ), .C(FIFO_CLK_c), .D(n4427));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1772_1773 (.Q(\REG.mem_18_2 ), .C(FIFO_CLK_c), .D(n4426));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1769_1770 (.Q(\REG.mem_18_1 ), .C(FIFO_CLK_c), .D(n4425));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1766_1767 (.Q(\REG.mem_18_0 ), .C(FIFO_CLK_c), .D(n4424));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1715_1716 (.Q(\REG.mem_17_15 ), .C(FIFO_CLK_c), .D(n4423));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFFE \REG.out_raw__i3  (.Q(\REG.out_raw[2] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [2]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFF i1712_1713 (.Q(\REG.mem_17_14 ), .C(FIFO_CLK_c), .D(n4422));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11202_bdd_4_lut (.I0(n11202), .I1(\REG.mem_37_2 ), .I2(\REG.mem_36_2 ), 
            .I3(rd_addr_r[1]), .O(n10169));
    defparam n11202_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10139 (.I0(rd_addr_r[1]), .I1(n9927), 
            .I2(n9928), .I3(rd_addr_r[2]), .O(n11796));
    defparam rd_addr_r_1__bdd_4_lut_10139.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i91_2_lut_3_lut_4_lut (.I0(n20_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n22));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i91_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 n11796_bdd_4_lut (.I0(n11796), .I1(n9925), .I2(n9924), .I3(rd_addr_r[2]), 
            .O(n10039));
    defparam n11796_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9575 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_2 ), 
            .I2(\REG.mem_43_2 ), .I3(rd_addr_r[1]), .O(n11196));
    defparam rd_addr_r_0__bdd_4_lut_9575.LUT_INIT = 16'he4aa;
    SB_LUT4 n11196_bdd_4_lut (.I0(n11196), .I1(\REG.mem_41_2 ), .I2(\REG.mem_40_2 ), 
            .I3(rd_addr_r[1]), .O(n10172));
    defparam n11196_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i122_2_lut_3_lut (.I0(n25_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n39));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i122_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10075 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_9 ), 
            .I2(\REG.mem_11_9 ), .I3(rd_addr_r[1]), .O(n11790));
    defparam rd_addr_r_0__bdd_4_lut_10075.LUT_INIT = 16'he4aa;
    SB_DFF i1709_1710 (.Q(\REG.mem_17_13 ), .C(FIFO_CLK_c), .D(n4421));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1706_1707 (.Q(\REG.mem_17_12 ), .C(FIFO_CLK_c), .D(n4420));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1703_1704 (.Q(\REG.mem_17_11 ), .C(FIFO_CLK_c), .D(n4419));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1700_1701 (.Q(\REG.mem_17_10 ), .C(FIFO_CLK_c), .D(n4418));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1697_1698 (.Q(\REG.mem_17_9 ), .C(FIFO_CLK_c), .D(n4417));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1694_1695 (.Q(\REG.mem_17_8 ), .C(FIFO_CLK_c), .D(n4416));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1691_1692 (.Q(\REG.mem_17_7 ), .C(FIFO_CLK_c), .D(n4415));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1688_1689 (.Q(\REG.mem_17_6 ), .C(FIFO_CLK_c), .D(n4414));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1685_1686 (.Q(\REG.mem_17_5 ), .C(FIFO_CLK_c), .D(n4413));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1682_1683 (.Q(\REG.mem_17_4 ), .C(FIFO_CLK_c), .D(n4412));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1679_1680 (.Q(\REG.mem_17_3 ), .C(FIFO_CLK_c), .D(n4411));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1676_1677 (.Q(\REG.mem_17_2 ), .C(FIFO_CLK_c), .D(n4410));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1673_1674 (.Q(\REG.mem_17_1 ), .C(FIFO_CLK_c), .D(n4409));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1670_1671 (.Q(\REG.mem_17_0 ), .C(FIFO_CLK_c), .D(n4408));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1619_1620 (.Q(\REG.mem_16_15 ), .C(FIFO_CLK_c), .D(n4407));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1616_1617 (.Q(\REG.mem_16_14 ), .C(FIFO_CLK_c), .D(n4406));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9189 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_0 ), 
            .I2(\REG.mem_55_0 ), .I3(rd_addr_r[1]), .O(n10722));
    defparam rd_addr_r_0__bdd_4_lut_9189.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9570 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_13 ), 
            .I2(\REG.mem_11_13 ), .I3(rd_addr_r[1]), .O(n11190));
    defparam rd_addr_r_0__bdd_4_lut_9570.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i121_2_lut_3_lut (.I0(n25_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n7));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i121_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i120_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n40));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i120_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 n11790_bdd_4_lut (.I0(n11790), .I1(\REG.mem_9_9 ), .I2(\REG.mem_8_9 ), 
            .I3(rd_addr_r[1]), .O(n11793));
    defparam n11790_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11190_bdd_4_lut (.I0(n11190), .I1(\REG.mem_9_13 ), .I2(\REG.mem_8_13 ), 
            .I3(rd_addr_r[1]), .O(n11193));
    defparam n11190_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i119_2_lut_3_lut (.I0(n23_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n8));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i119_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10065 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_5 ), 
            .I2(\REG.mem_51_5 ), .I3(rd_addr_r[1]), .O(n11784));
    defparam rd_addr_r_0__bdd_4_lut_10065.LUT_INIT = 16'he4aa;
    SB_LUT4 n11784_bdd_4_lut (.I0(n11784), .I1(\REG.mem_49_5 ), .I2(\REG.mem_48_5 ), 
            .I3(rd_addr_r[1]), .O(n10463));
    defparam n11784_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9229 (.I0(rd_addr_r[2]), .I1(n9827), 
            .I2(n10454), .I3(rd_addr_r[3]), .O(n10746));
    defparam rd_addr_r_2__bdd_4_lut_9229.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9204 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_12 ), 
            .I2(\REG.mem_15_12 ), .I3(rd_addr_r[1]), .O(n10740));
    defparam rd_addr_r_0__bdd_4_lut_9204.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i23_2_lut_3_lut (.I0(n12_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n23_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i23_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i1613_1614 (.Q(\REG.mem_16_13 ), .C(FIFO_CLK_c), .D(n4405));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n10722_bdd_4_lut (.I0(n10722), .I1(\REG.mem_53_0 ), .I2(\REG.mem_52_0 ), 
            .I3(rd_addr_r[1]), .O(n10725));
    defparam n10722_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1610_1611 (.Q(\REG.mem_16_12 ), .C(FIFO_CLK_c), .D(n4404));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1607_1608 (.Q(\REG.mem_16_11 ), .C(FIFO_CLK_c), .D(n4403));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1604_1605 (.Q(\REG.mem_16_10 ), .C(FIFO_CLK_c), .D(n4402));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1601_1602 (.Q(\REG.mem_16_9 ), .C(FIFO_CLK_c), .D(n4401));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1598_1599 (.Q(\REG.mem_16_8 ), .C(FIFO_CLK_c), .D(n4400));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1595_1596 (.Q(\REG.mem_16_7 ), .C(FIFO_CLK_c), .D(n4399));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1592_1593 (.Q(\REG.mem_16_6 ), .C(FIFO_CLK_c), .D(n4398));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1589_1590 (.Q(\REG.mem_16_5 ), .C(FIFO_CLK_c), .D(n4397));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1586_1587 (.Q(\REG.mem_16_4 ), .C(FIFO_CLK_c), .D(n4396));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1583_1584 (.Q(\REG.mem_16_3 ), .C(FIFO_CLK_c), .D(n4395));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1580_1581 (.Q(\REG.mem_16_2 ), .C(FIFO_CLK_c), .D(n4394));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1577_1578 (.Q(\REG.mem_16_1 ), .C(FIFO_CLK_c), .D(n4393));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1574_1575 (.Q(\REG.mem_16_0 ), .C(FIFO_CLK_c), .D(n4392));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1523_1524 (.Q(\REG.mem_15_15 ), .C(FIFO_CLK_c), .D(n4391));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFFE \REG.out_raw__i2  (.Q(\REG.out_raw[1] ), .C(DEBUG_6_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_237 [1]));   // src/fifo_dc_32_lut_gen.v(891[25] 897[28])
    SB_DFF i1520_1521 (.Q(\REG.mem_15_14 ), .C(FIFO_CLK_c), .D(n4390));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i40_2_lut_3_lut_4_lut (.I0(n12_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n40_adj_1070));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i40_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9184 (.I0(rd_addr_r[2]), .I1(n10094), 
            .I2(n10118), .I3(rd_addr_r[3]), .O(n10716));
    defparam rd_addr_r_2__bdd_4_lut_9184.LUT_INIT = 16'he4aa;
    SB_LUT4 i3570_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_31_3 ), .O(n4659));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3570_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n10740_bdd_4_lut (.I0(n10740), .I1(\REG.mem_13_12 ), .I2(\REG.mem_12_12 ), 
            .I3(rd_addr_r[1]), .O(n10743));
    defparam n10740_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10734_bdd_4_lut (.I0(n10734), .I1(\REG.mem_25_13 ), .I2(\REG.mem_24_13 ), 
            .I3(rd_addr_r[1]), .O(n10737));
    defparam n10734_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i39_2_lut_3_lut_4_lut (.I0(n12_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n39_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i39_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9194 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_13 ), 
            .I2(\REG.mem_27_13 ), .I3(rd_addr_r[1]), .O(n10734));
    defparam rd_addr_r_0__bdd_4_lut_9194.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_29 (.I0(rp_sync2_r[6]), .I1(rp_sync2_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n3567));   // src/fifo_dc_32_lut_gen.v(286[38:77])
    defparam i1_2_lut_adj_29.LUT_INIT = 16'h6666;
    SB_LUT4 n10716_bdd_4_lut (.I0(n10716), .I1(n10046), .I2(n10025), .I3(rd_addr_r[3]), 
            .O(n10719));
    defparam n10716_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9565 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_0 ), 
            .I2(\REG.mem_39_0 ), .I3(rd_addr_r[1]), .O(n11178));
    defparam rd_addr_r_0__bdd_4_lut_9565.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_30 (.I0(rp_sync2_r[3]), .I1(n3563), .I2(GND_net), 
            .I3(GND_net), .O(n3550));   // src/fifo_dc_32_lut_gen.v(286[38:77])
    defparam i1_2_lut_adj_30.LUT_INIT = 16'h6666;
    SB_LUT4 n11178_bdd_4_lut (.I0(n11178), .I1(\REG.mem_37_0 ), .I2(\REG.mem_36_0 ), 
            .I3(rd_addr_r[1]), .O(n11181));
    defparam n11178_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1517_1518 (.Q(\REG.mem_15_13 ), .C(FIFO_CLK_c), .D(n4389));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1514_1515 (.Q(\REG.mem_15_12 ), .C(FIFO_CLK_c), .D(n4388));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1511_1512 (.Q(\REG.mem_15_11 ), .C(FIFO_CLK_c), .D(n4387));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1508_1509 (.Q(\REG.mem_15_10 ), .C(FIFO_CLK_c), .D(n4386));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1505_1506 (.Q(\REG.mem_15_9 ), .C(FIFO_CLK_c), .D(n4385));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1502_1503 (.Q(\REG.mem_15_8 ), .C(FIFO_CLK_c), .D(n4384));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1499_1500 (.Q(\REG.mem_15_7 ), .C(FIFO_CLK_c), .D(n4383));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1496_1497 (.Q(\REG.mem_15_6 ), .C(FIFO_CLK_c), .D(n4382));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1493_1494 (.Q(\REG.mem_15_5 ), .C(FIFO_CLK_c), .D(n4381));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1490_1491 (.Q(\REG.mem_15_4 ), .C(FIFO_CLK_c), .D(n4380));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1487_1488 (.Q(\REG.mem_15_3 ), .C(FIFO_CLK_c), .D(n4379));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1484_1485 (.Q(\REG.mem_15_2 ), .C(FIFO_CLK_c), .D(n4378));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1481_1482 (.Q(\REG.mem_15_1 ), .C(FIFO_CLK_c), .D(n4377));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1478_1479 (.Q(\REG.mem_15_0 ), .C(FIFO_CLK_c), .D(n4376));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1427_1428 (.Q(\REG.mem_14_15 ), .C(FIFO_CLK_c), .D(n4375));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1424_1425 (.Q(\REG.mem_14_14 ), .C(FIFO_CLK_c), .D(n4374));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9199 (.I0(rd_addr_r[2]), .I1(n9560), 
            .I2(n9569), .I3(rd_addr_r[3]), .O(n10728));
    defparam rd_addr_r_2__bdd_4_lut_9199.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10060 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_8 ), 
            .I2(\REG.mem_7_8 ), .I3(rd_addr_r[1]), .O(n11778));
    defparam rd_addr_r_0__bdd_4_lut_10060.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_31 (.I0(n3597), .I1(rp_sync2_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n9366));   // src/fifo_dc_32_lut_gen.v(286[38:77])
    defparam i1_2_lut_adj_31.LUT_INIT = 16'h6666;
    SB_LUT4 n11778_bdd_4_lut (.I0(n11778), .I1(\REG.mem_5_8 ), .I2(\REG.mem_4_8 ), 
            .I3(rd_addr_r[1]), .O(n11781));
    defparam n11778_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7872_4_lut (.I0(wr_addr_p1_w[4]), .I1(wr_addr_p1_w[1]), .I2(n3563), 
            .I3(n3597), .O(n9412));
    defparam i7872_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i7891_4_lut (.I0(wr_addr_p1_w[5]), .I1(wr_addr_p1_w[3]), .I2(n3567), 
            .I3(n3550), .O(n9432));
    defparam i7891_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut (.I0(wr_addr_p1_w[0]), .I1(wr_addr_p1_w[6]), .I2(n9366), 
            .I3(rp_sync2_r[6]), .O(n9_adj_1071));
    defparam i2_4_lut.LUT_INIT = 16'h2184;
    SB_LUT4 i3569_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_31_2 ), .O(n4658));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3569_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10055 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_10 ), 
            .I2(\REG.mem_55_10 ), .I3(rd_addr_r[1]), .O(n11772));
    defparam rd_addr_r_0__bdd_4_lut_10055.LUT_INIT = 16'he4aa;
    SB_LUT4 n11772_bdd_4_lut (.I0(n11772), .I1(\REG.mem_53_10 ), .I2(\REG.mem_52_10 ), 
            .I3(rd_addr_r[1]), .O(n10046));
    defparam n11772_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_32 (.I0(wr_addr_p1_w[2]), .I1(n3584), .I2(GND_net), 
            .I3(GND_net), .O(n3586));   // src/fifo_dc_32_lut_gen.v(286[38:77])
    defparam i1_2_lut_adj_32.LUT_INIT = 16'h6666;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10050 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_9 ), 
            .I2(\REG.mem_15_9 ), .I3(rd_addr_r[1]), .O(n11766));
    defparam rd_addr_r_0__bdd_4_lut_10050.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9555 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_8 ), 
            .I2(\REG.mem_39_8 ), .I3(rd_addr_r[1]), .O(n11172));
    defparam rd_addr_r_0__bdd_4_lut_9555.LUT_INIT = 16'he4aa;
    SB_LUT4 n11766_bdd_4_lut (.I0(n11766), .I1(\REG.mem_13_9 ), .I2(\REG.mem_12_9 ), 
            .I3(rd_addr_r[1]), .O(n11769));
    defparam n11766_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11172_bdd_4_lut (.I0(n11172), .I1(\REG.mem_37_8 ), .I2(\REG.mem_36_8 ), 
            .I3(rd_addr_r[1]), .O(n11175));
    defparam n11172_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10045 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_15 ), 
            .I2(\REG.mem_39_15 ), .I3(rd_addr_r[1]), .O(n11760));
    defparam rd_addr_r_0__bdd_4_lut_10045.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9550 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_5 ), 
            .I2(\REG.mem_7_5 ), .I3(rd_addr_r[1]), .O(n11166));
    defparam rd_addr_r_0__bdd_4_lut_9550.LUT_INIT = 16'he4aa;
    SB_LUT4 n11760_bdd_4_lut (.I0(n11760), .I1(\REG.mem_37_15 ), .I2(\REG.mem_36_15 ), 
            .I3(rd_addr_r[1]), .O(n11763));
    defparam n11760_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i38_39 (.Q(\REG.mem_0_0 ), .C(FIFO_CLK_c), .D(n4140));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1421_1422 (.Q(\REG.mem_14_13 ), .C(FIFO_CLK_c), .D(n4373));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1418_1419 (.Q(\REG.mem_14_12 ), .C(FIFO_CLK_c), .D(n4372));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1415_1416 (.Q(\REG.mem_14_11 ), .C(FIFO_CLK_c), .D(n4371));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1412_1413 (.Q(\REG.mem_14_10 ), .C(FIFO_CLK_c), .D(n4370));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1409_1410 (.Q(\REG.mem_14_9 ), .C(FIFO_CLK_c), .D(n4369));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1406_1407 (.Q(\REG.mem_14_8 ), .C(FIFO_CLK_c), .D(n4368));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1403_1404 (.Q(\REG.mem_14_7 ), .C(FIFO_CLK_c), .D(n4367));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i7856_4_lut (.I0(wr_addr_r[5]), .I1(wr_addr_r[1]), .I2(n3567), 
            .I3(n3597), .O(n9396));
    defparam i7856_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i7840_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_r[0]), .I2(n3584), 
            .I3(n9366), .O(n9380));
    defparam i7840_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i9046_4_lut (.I0(n3586), .I1(n9_adj_1071), .I2(n9432), .I3(n9412), 
            .O(n10527));   // src/fifo_dc_32_lut_gen.v(298[45:114])
    defparam i9046_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i7938_3_lut (.I0(n9390), .I1(n9380), .I2(n9396), .I3(GND_net), 
            .O(n9480));
    defparam i7938_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 full_nxt_c_I_9_4_lut (.I0(n9480), .I1(n10527), .I2(write_to_dc32_fifo), 
            .I3(dc32_fifo_is_full), .O(full_nxt_c_N_303));   // src/fifo_dc_32_lut_gen.v(298[45:114])
    defparam full_nxt_c_I_9_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 n11166_bdd_4_lut (.I0(n11166), .I1(\REG.mem_5_5 ), .I2(\REG.mem_4_5 ), 
            .I3(rd_addr_r[1]), .O(n11169));
    defparam n11166_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1400_1401 (.Q(\REG.mem_14_6 ), .C(FIFO_CLK_c), .D(n4366));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1397_1398 (.Q(\REG.mem_14_5 ), .C(FIFO_CLK_c), .D(n4365));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1394_1395 (.Q(\REG.mem_14_4 ), .C(FIFO_CLK_c), .D(n4364));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1391_1392 (.Q(\REG.mem_14_3 ), .C(FIFO_CLK_c), .D(n4363));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1388_1389 (.Q(\REG.mem_14_2 ), .C(FIFO_CLK_c), .D(n4362));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1385_1386 (.Q(\REG.mem_14_1 ), .C(FIFO_CLK_c), .D(n4361));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1382_1383 (.Q(\REG.mem_14_0 ), .C(FIFO_CLK_c), .D(n4360));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1331_1332 (.Q(\REG.mem_13_15 ), .C(FIFO_CLK_c), .D(n4359));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8814_3_lut (.I0(\REG.mem_32_14 ), .I1(\REG.mem_33_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10356));
    defparam i8814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8815_3_lut (.I0(\REG.mem_34_14 ), .I1(\REG.mem_35_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10357));
    defparam i8815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7963_3_lut (.I0(n12243), .I1(n12225), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9505));
    defparam i7963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10040 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_9 ), 
            .I2(\REG.mem_19_9 ), .I3(rd_addr_r[1]), .O(n11754));
    defparam rd_addr_r_0__bdd_4_lut_10040.LUT_INIT = 16'he4aa;
    SB_DFF i1328_1329 (.Q(\REG.mem_13_14 ), .C(FIFO_CLK_c), .D(n4358));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i7964_3_lut (.I0(n10965), .I1(n9505), .I2(rd_addr_r[3]), .I3(GND_net), 
            .O(n9506));
    defparam i7964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11754_bdd_4_lut (.I0(n11754), .I1(\REG.mem_17_9 ), .I2(\REG.mem_16_9 ), 
            .I3(rd_addr_r[1]), .O(n11757));
    defparam n11754_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1325_1326 (.Q(\REG.mem_13_13 ), .C(FIFO_CLK_c), .D(n4357));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1322_1323 (.Q(\REG.mem_13_12 ), .C(FIFO_CLK_c), .D(n4356));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1319_1320 (.Q(\REG.mem_13_11 ), .C(FIFO_CLK_c), .D(n4355));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1316_1317 (.Q(\REG.mem_13_10 ), .C(FIFO_CLK_c), .D(n4354));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1313_1314 (.Q(\REG.mem_13_9 ), .C(FIFO_CLK_c), .D(n4353));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1310_1311 (.Q(\REG.mem_13_8 ), .C(FIFO_CLK_c), .D(n4352));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1307_1308 (.Q(\REG.mem_13_7 ), .C(FIFO_CLK_c), .D(n4351));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i41_42 (.Q(\REG.mem_0_1 ), .C(FIFO_CLK_c), .D(n4139));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i44_45 (.Q(\REG.mem_0_2 ), .C(FIFO_CLK_c), .D(n4138));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1304_1305 (.Q(\REG.mem_13_6 ), .C(FIFO_CLK_c), .D(n4350));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i47_48 (.Q(\REG.mem_0_3 ), .C(FIFO_CLK_c), .D(n4136));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8824_3_lut (.I0(\REG.mem_38_14 ), .I1(\REG.mem_39_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10366));
    defparam i8824_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1301_1302 (.Q(\REG.mem_13_5 ), .C(FIFO_CLK_c), .D(n4349));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8823_3_lut (.I0(\REG.mem_36_14 ), .I1(\REG.mem_37_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10365));
    defparam i8823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10159 (.I0(rd_addr_r[4]), .I1(n9632), 
            .I2(n9653), .I3(rd_addr_r[5]), .O(n11748));
    defparam rd_addr_r_4__bdd_4_lut_10159.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9585 (.I0(rd_addr_r[1]), .I1(n10512), 
            .I2(n10513), .I3(rd_addr_r[2]), .O(n11160));
    defparam rd_addr_r_1__bdd_4_lut_9585.LUT_INIT = 16'he4aa;
    SB_DFF i1298_1299 (.Q(\REG.mem_13_4 ), .C(FIFO_CLK_c), .D(n4348));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1295_1296 (.Q(\REG.mem_13_3 ), .C(FIFO_CLK_c), .D(n4347));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1292_1293 (.Q(\REG.mem_13_2 ), .C(FIFO_CLK_c), .D(n4346));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1289_1290 (.Q(\REG.mem_13_1 ), .C(FIFO_CLK_c), .D(n4345));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1286_1287 (.Q(\REG.mem_13_0 ), .C(FIFO_CLK_c), .D(n4344));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1235_1236 (.Q(\REG.mem_12_15 ), .C(FIFO_CLK_c), .D(n4343));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1232_1233 (.Q(\REG.mem_12_14 ), .C(FIFO_CLK_c), .D(n4342));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1229_1230 (.Q(\REG.mem_12_13 ), .C(FIFO_CLK_c), .D(n4341));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11748_bdd_4_lut (.I0(n11748), .I1(n11079), .I2(n9542), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_237 [11]));
    defparam n11748_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7972_3_lut (.I0(n11877), .I1(n11865), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9514));
    defparam i7972_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1226_1227 (.Q(\REG.mem_12_12 ), .C(FIFO_CLK_c), .D(n4340));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1223_1224 (.Q(\REG.mem_12_11 ), .C(FIFO_CLK_c), .D(n4339));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1220_1221 (.Q(\REG.mem_12_10 ), .C(FIFO_CLK_c), .D(n4338));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1217_1218 (.Q(\REG.mem_12_9 ), .C(FIFO_CLK_c), .D(n4337));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1214_1215 (.Q(\REG.mem_12_8 ), .C(FIFO_CLK_c), .D(n4336));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1211_1212 (.Q(\REG.mem_12_7 ), .C(FIFO_CLK_c), .D(n4335));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1208_1209 (.Q(\REG.mem_12_6 ), .C(FIFO_CLK_c), .D(n4334));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1205_1206 (.Q(\REG.mem_12_5 ), .C(FIFO_CLK_c), .D(n4333));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1202_1203 (.Q(\REG.mem_12_4 ), .C(FIFO_CLK_c), .D(n4332));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1199_1200 (.Q(\REG.mem_12_3 ), .C(FIFO_CLK_c), .D(n4331));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1196_1197 (.Q(\REG.mem_12_2 ), .C(FIFO_CLK_c), .D(n4330));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1193_1194 (.Q(\REG.mem_12_1 ), .C(FIFO_CLK_c), .D(n4329));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1190_1191 (.Q(\REG.mem_12_0 ), .C(FIFO_CLK_c), .D(n4328));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1139_1140 (.Q(\REG.mem_11_15 ), .C(FIFO_CLK_c), .D(n4327));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1136_1137 (.Q(\REG.mem_11_14 ), .C(FIFO_CLK_c), .D(n4326));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i7973_3_lut (.I0(n10995), .I1(n9514), .I2(rd_addr_r[3]), .I3(GND_net), 
            .O(n9515));
    defparam i7973_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1133_1134 (.Q(\REG.mem_11_13 ), .C(FIFO_CLK_c), .D(n4325));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1130_1131 (.Q(\REG.mem_11_12 ), .C(FIFO_CLK_c), .D(n4324));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10035 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_5 ), 
            .I2(\REG.mem_55_5 ), .I3(rd_addr_r[1]), .O(n11742));
    defparam rd_addr_r_0__bdd_4_lut_10035.LUT_INIT = 16'he4aa;
    SB_DFF i1127_1128 (.Q(\REG.mem_11_11 ), .C(FIFO_CLK_c), .D(n4323));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i80_2_lut_3_lut (.I0(n32), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n60));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i80_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_DFF i1124_1125 (.Q(\REG.mem_11_10 ), .C(FIFO_CLK_c), .D(n4322));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i79_2_lut_3_lut (.I0(n32), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n28));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i79_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i118_2_lut_3_lut (.I0(n21_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n41));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i118_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i117_2_lut_3_lut (.I0(n21_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n9));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i117_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n11160_bdd_4_lut (.I0(n11160), .I1(n10507), .I2(n10506), .I3(rd_addr_r[2]), 
            .O(n11163));
    defparam n11160_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i21_2_lut_3_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n21_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i21_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i1121_1122 (.Q(\REG.mem_11_9 ), .C(FIFO_CLK_c), .D(n4321));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11742_bdd_4_lut (.I0(n11742), .I1(\REG.mem_53_5 ), .I2(\REG.mem_52_5 ), 
            .I3(rd_addr_r[1]), .O(n10472));
    defparam n11742_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i38_2_lut_3_lut_4_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n38));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i38_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i7969_3_lut (.I0(n12063), .I1(n11919), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9511));
    defparam i7969_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i50_51 (.Q(\REG.mem_0_4 ), .C(FIFO_CLK_c), .D(n4134));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i7970_3_lut (.I0(n10989), .I1(n9511), .I2(rd_addr_r[3]), .I3(GND_net), 
            .O(n9512));
    defparam i7970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i37_2_lut_3_lut_4_lut (.I0(n10_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[4]), .I3(wr_addr_r[3]), .O(n37_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i37_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_DFF i1118_1119 (.Q(\REG.mem_11_8 ), .C(FIFO_CLK_c), .D(n4320));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9224 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_6 ), 
            .I2(\REG.mem_43_6 ), .I3(rd_addr_r[1]), .O(n10770));
    defparam rd_addr_r_0__bdd_4_lut_9224.LUT_INIT = 16'he4aa;
    SB_DFF i1115_1116 (.Q(\REG.mem_11_7 ), .C(FIFO_CLK_c), .D(n4319));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9545 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_2 ), 
            .I2(\REG.mem_47_2 ), .I3(rd_addr_r[1]), .O(n11154));
    defparam rd_addr_r_0__bdd_4_lut_9545.LUT_INIT = 16'he4aa;
    SB_LUT4 n11154_bdd_4_lut (.I0(n11154), .I1(\REG.mem_45_2 ), .I2(\REG.mem_44_2 ), 
            .I3(rd_addr_r[1]), .O(n10181));
    defparam n11154_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i53_54 (.Q(\REG.mem_0_5 ), .C(FIFO_CLK_c), .D(n4133));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1112_1113 (.Q(\REG.mem_11_6 ), .C(FIFO_CLK_c), .D(n4318));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10070 (.I0(rd_addr_r[1]), .I1(n9960), 
            .I2(n9961), .I3(rd_addr_r[2]), .O(n11736));
    defparam rd_addr_r_1__bdd_4_lut_10070.LUT_INIT = 16'he4aa;
    SB_DFF i1109_1110 (.Q(\REG.mem_11_5 ), .C(FIFO_CLK_c), .D(n4317));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9540 (.I0(rd_addr_r[1]), .I1(n10482), 
            .I2(n10483), .I3(rd_addr_r[2]), .O(n11148));
    defparam rd_addr_r_1__bdd_4_lut_9540.LUT_INIT = 16'he4aa;
    SB_DFF i1106_1107 (.Q(\REG.mem_11_4 ), .C(FIFO_CLK_c), .D(n4316));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11736_bdd_4_lut (.I0(n11736), .I1(n9952), .I2(n9951), .I3(rd_addr_r[2]), 
            .O(n10051));
    defparam n11736_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1103_1104 (.Q(\REG.mem_11_3 ), .C(FIFO_CLK_c), .D(n4315));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1100_1101 (.Q(\REG.mem_11_2 ), .C(FIFO_CLK_c), .D(n4314));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1097_1098 (.Q(\REG.mem_11_1 ), .C(FIFO_CLK_c), .D(n4313));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1094_1095 (.Q(\REG.mem_11_0 ), .C(FIFO_CLK_c), .D(n4312));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1043_1044 (.Q(\REG.mem_10_15 ), .C(FIFO_CLK_c), .D(n4311));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i4138_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_63_15 ), .O(n5227));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4138_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i116_2_lut_3_lut (.I0(n36_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n42));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i116_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i1040_1041 (.Q(\REG.mem_10_14 ), .C(FIFO_CLK_c), .D(n4310));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1037_1038 (.Q(\REG.mem_10_13 ), .C(FIFO_CLK_c), .D(n4309));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1034_1035 (.Q(\REG.mem_10_12 ), .C(FIFO_CLK_c), .D(n4308));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3568_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_31_1 ), .O(n4657));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3568_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i115_2_lut_3_lut (.I0(n36_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n10));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i115_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4137_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_63_14 ), .O(n5226));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4137_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1031_1032 (.Q(\REG.mem_10_11 ), .C(FIFO_CLK_c), .D(n4307));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8883_3_lut (.I0(\REG.mem_48_14 ), .I1(\REG.mem_49_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10425));
    defparam i8883_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1028_1029 (.Q(\REG.mem_10_10 ), .C(FIFO_CLK_c), .D(n4306));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i56_57 (.Q(\REG.mem_0_6 ), .C(FIFO_CLK_c), .D(n4132));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3567_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_31_0 ), .O(n4656));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3567_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n10770_bdd_4_lut (.I0(n10770), .I1(\REG.mem_41_6 ), .I2(\REG.mem_40_6 ), 
            .I3(rd_addr_r[1]), .O(n10773));
    defparam n10770_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8884_3_lut (.I0(\REG.mem_50_14 ), .I1(\REG.mem_51_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10426));
    defparam i8884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11148_bdd_4_lut (.I0(n11148), .I1(n10477), .I2(n10476), .I3(rd_addr_r[2]), 
            .O(n11151));
    defparam n11148_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3676_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_36_15 ), .O(n4765));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3676_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1025_1026 (.Q(\REG.mem_10_9 ), .C(FIFO_CLK_c), .D(n4305));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8887_3_lut (.I0(\REG.mem_54_14 ), .I1(\REG.mem_55_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10429));
    defparam i8887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10025 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_9 ), 
            .I2(\REG.mem_23_9 ), .I3(rd_addr_r[1]), .O(n11730));
    defparam rd_addr_r_0__bdd_4_lut_10025.LUT_INIT = 16'he4aa;
    SB_DFF i1022_1023 (.Q(\REG.mem_10_8 ), .C(FIFO_CLK_c), .D(n4304));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i4136_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_63_13 ), .O(n5225));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4136_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8886_3_lut (.I0(\REG.mem_52_14 ), .I1(\REG.mem_53_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10428));
    defparam i8886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11730_bdd_4_lut (.I0(n11730), .I1(\REG.mem_21_9 ), .I2(\REG.mem_20_9 ), 
            .I3(rd_addr_r[1]), .O(n11733));
    defparam n11730_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1019_1020 (.Q(\REG.mem_10_7 ), .C(FIFO_CLK_c), .D(n4303));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3675_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_36_14 ), .O(n4764));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3675_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1016_1017 (.Q(\REG.mem_10_6 ), .C(FIFO_CLK_c), .D(n4302));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1013_1014 (.Q(\REG.mem_10_5 ), .C(FIFO_CLK_c), .D(n4301));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9535 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_5 ), 
            .I2(\REG.mem_11_5 ), .I3(rd_addr_r[1]), .O(n11142));
    defparam rd_addr_r_0__bdd_4_lut_9535.LUT_INIT = 16'he4aa;
    SB_LUT4 i3674_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_36_13 ), .O(n4763));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3674_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1010_1011 (.Q(\REG.mem_10_4 ), .C(FIFO_CLK_c), .D(n4300));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3673_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_36_12 ), .O(n4762));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3673_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1007_1008 (.Q(\REG.mem_10_3 ), .C(FIFO_CLK_c), .D(n4299));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i1004_1005 (.Q(\REG.mem_10_2 ), .C(FIFO_CLK_c), .D(n4298));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i4135_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_63_12 ), .O(n5224));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4135_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3672_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_36_11 ), .O(n4761));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3672_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1001_1002 (.Q(\REG.mem_10_1 ), .C(FIFO_CLK_c), .D(n4297));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3671_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_36_10 ), .O(n4760));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3671_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i998_999 (.Q(\REG.mem_10_0 ), .C(FIFO_CLK_c), .D(n4296));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i59_60 (.Q(\REG.mem_0_7 ), .C(FIFO_CLK_c), .D(n4131));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF \genblk16.rd_prev_r_111  (.Q(\genblk16.rd_prev_r ), .C(DEBUG_6_c), 
           .D(n4130));   // src/fifo_dc_32_lut_gen.v(749[29] 759[32])
    SB_LUT4 i3670_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_36_9 ), .O(n4759));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3670_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i86_2_lut_3_lut (.I0(n21_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n57));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i86_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i4134_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_63_11 ), .O(n5223));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4134_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3669_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_36_8 ), .O(n4758));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3669_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3668_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_36_7 ), .O(n4757));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3668_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11142_bdd_4_lut (.I0(n11142), .I1(\REG.mem_9_5 ), .I2(\REG.mem_8_5 ), 
            .I3(rd_addr_r[1]), .O(n11145));
    defparam n11142_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3667_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_36_6 ), .O(n4756));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3667_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3666_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_36_5 ), .O(n4755));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3666_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i62_63 (.Q(\REG.mem_0_8 ), .C(FIFO_CLK_c), .D(n4126));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10299 (.I0(rd_addr_r[2]), .I1(n11115), 
            .I2(n9842), .I3(rd_addr_r[3]), .O(n11724));
    defparam rd_addr_r_2__bdd_4_lut_10299.LUT_INIT = 16'he4aa;
    SB_DFF i65_66 (.Q(\REG.mem_0_9 ), .C(FIFO_CLK_c), .D(n4125));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i68_69 (.Q(\REG.mem_0_10 ), .C(FIFO_CLK_c), .D(n4124));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3665_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_36_4 ), .O(n4754));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3665_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9525 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_3 ), 
            .I2(\REG.mem_39_3 ), .I3(rd_addr_r[1]), .O(n11136));
    defparam rd_addr_r_0__bdd_4_lut_9525.LUT_INIT = 16'he4aa;
    SB_LUT4 n11724_bdd_4_lut (.I0(n11724), .I1(n10472), .I2(n10463), .I3(rd_addr_r[3]), 
            .O(n10481));
    defparam n11724_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i947_948 (.Q(\REG.mem_9_15 ), .C(FIFO_CLK_c), .D(n4288));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(FIFO_CLK_c), .D(n4287));   // src/fifo_dc_32_lut_gen.v(308[21] 324[24])
    SB_DFF i944_945 (.Q(\REG.mem_9_14 ), .C(FIFO_CLK_c), .D(n4286));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i941_942 (.Q(\REG.mem_9_13 ), .C(FIFO_CLK_c), .D(n4285));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i938_939 (.Q(\REG.mem_9_12 ), .C(FIFO_CLK_c), .D(n4284));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i935_936 (.Q(\REG.mem_9_11 ), .C(FIFO_CLK_c), .D(n4283));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i932_933 (.Q(\REG.mem_9_10 ), .C(FIFO_CLK_c), .D(n4282));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i929_930 (.Q(\REG.mem_9_9 ), .C(FIFO_CLK_c), .D(n4281));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i71_72 (.Q(\REG.mem_0_11 ), .C(FIFO_CLK_c), .D(n4120));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i74_75 (.Q(\REG.mem_0_12 ), .C(FIFO_CLK_c), .D(n4119));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i143_144 (.Q(\REG.mem_1_3 ), .C(FIFO_CLK_c), .D(n4118));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(FIFO_CLK_c), .D(n4117));   // src/fifo_dc_32_lut_gen.v(308[21] 324[24])
    SB_DFF i77_78 (.Q(\REG.mem_0_13 ), .C(FIFO_CLK_c), .D(n4114));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i80_81 (.Q(\REG.mem_0_14 ), .C(FIFO_CLK_c), .D(n4113));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i83_84 (.Q(\REG.mem_0_15 ), .C(FIFO_CLK_c), .D(n4112));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i926_927 (.Q(\REG.mem_9_8 ), .C(FIFO_CLK_c), .D(n4280));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9179 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_13 ), 
            .I2(\REG.mem_31_13 ), .I3(rd_addr_r[1]), .O(n10710));
    defparam rd_addr_r_0__bdd_4_lut_9179.LUT_INIT = 16'he4aa;
    SB_LUT4 i3664_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_36_3 ), .O(n4753));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3664_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3663_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_36_2 ), .O(n4752));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3663_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i923_924 (.Q(\REG.mem_9_7 ), .C(FIFO_CLK_c), .D(n4279));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11136_bdd_4_lut (.I0(n11136), .I1(\REG.mem_37_3 ), .I2(\REG.mem_36_3 ), 
            .I3(rd_addr_r[1]), .O(n11139));
    defparam n11136_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3662_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_36_1 ), .O(n4751));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3662_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3661_3_lut_4_lut (.I0(n46_c), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_36_0 ), .O(n4750));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3661_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3660_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_35_15 ), .O(n4749));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3660_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i920_921 (.Q(\REG.mem_9_6 ), .C(FIFO_CLK_c), .D(n4278));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8319_3_lut (.I0(n10821), .I1(n12201), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9861));
    defparam i8319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10020 (.I0(rd_addr_r[1]), .I1(n9993), 
            .I2(n9994), .I3(rd_addr_r[2]), .O(n11718));
    defparam rd_addr_r_1__bdd_4_lut_10020.LUT_INIT = 16'he4aa;
    SB_LUT4 i3659_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_35_14 ), .O(n4748));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3659_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8320_3_lut (.I0(n12159), .I1(n12069), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9862));
    defparam i8320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11718_bdd_4_lut (.I0(n11718), .I1(n9988), .I2(n9987), .I3(rd_addr_r[2]), 
            .O(n10054));
    defparam n11718_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3658_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_35_13 ), .O(n4747));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3658_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4133_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_63_10 ), .O(n5222));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4133_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4132_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_63_9 ), .O(n5221));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4132_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i917_918 (.Q(\REG.mem_9_5 ), .C(FIFO_CLK_c), .D(n4277));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3657_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_35_12 ), .O(n4746));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3657_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3656_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_35_11 ), .O(n4745));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3656_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4131_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_63_8 ), .O(n5220));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4131_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9520 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_0 ), 
            .I2(\REG.mem_43_0 ), .I3(rd_addr_r[1]), .O(n11130));
    defparam rd_addr_r_0__bdd_4_lut_9520.LUT_INIT = 16'he4aa;
    SB_LUT4 n11130_bdd_4_lut (.I0(n11130), .I1(\REG.mem_41_0 ), .I2(\REG.mem_40_0 ), 
            .I3(rd_addr_r[1]), .O(n11133));
    defparam n11130_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3655_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_35_10 ), .O(n4744));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3655_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF wp_sync2_r__i0 (.Q(wp_sync2_r[0]), .C(DEBUG_6_c), .D(n4108));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10010 (.I0(rd_addr_r[2]), .I1(n9932), 
            .I2(n9977), .I3(rd_addr_r[3]), .O(n11712));
    defparam rd_addr_r_2__bdd_4_lut_10010.LUT_INIT = 16'he4aa;
    SB_LUT4 i3654_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_35_9 ), .O(n4743));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3654_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3653_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_35_8 ), .O(n4742));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3653_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11712_bdd_4_lut (.I0(n11712), .I1(n9887), .I2(n11283), .I3(rd_addr_r[3]), 
            .O(n10487));
    defparam n11712_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3652_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_35_7 ), .O(n4741));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3652_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3651_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_35_6 ), .O(n4740));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3651_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3650_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_35_5 ), .O(n4739));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3650_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3649_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_35_4 ), .O(n4738));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3649_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i85_2_lut_3_lut (.I0(n21_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n25));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i85_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_10015 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_11 ), 
            .I2(\REG.mem_63_11 ), .I3(rd_addr_r[1]), .O(n11706));
    defparam rd_addr_r_0__bdd_4_lut_10015.LUT_INIT = 16'he4aa;
    SB_LUT4 n11706_bdd_4_lut (.I0(n11706), .I1(\REG.mem_61_11 ), .I2(\REG.mem_60_11 ), 
            .I3(rd_addr_r[1]), .O(n11709));
    defparam n11706_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3648_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_35_3 ), .O(n4737));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3648_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3647_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_35_2 ), .O(n4736));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3647_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i914_915 (.Q(\REG.mem_9_4 ), .C(FIFO_CLK_c), .D(n4276));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i4130_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_63_7 ), .O(n5219));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4130_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3646_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_35_1 ), .O(n4735));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3646_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3645_3_lut_4_lut (.I0(n44_c), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_35_0 ), .O(n4734));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3645_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9995 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_11 ), 
            .I2(\REG.mem_43_11 ), .I3(rd_addr_r[1]), .O(n11700));
    defparam rd_addr_r_0__bdd_4_lut_9995.LUT_INIT = 16'he4aa;
    SB_LUT4 n11700_bdd_4_lut (.I0(n11700), .I1(\REG.mem_41_11 ), .I2(\REG.mem_40_11 ), 
            .I3(rd_addr_r[1]), .O(n11703));
    defparam n11700_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i114_2_lut_3_lut (.I0(n34), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n43));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i114_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i4129_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_63_6 ), .O(n5218));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4129_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i113_2_lut_3_lut (.I0(n34), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n11));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i113_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i112_2_lut_3_lut (.I0(n32), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n44));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i112_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i111_2_lut_3_lut (.I0(n32), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n12));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i111_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9515 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_3 ), 
            .I2(\REG.mem_43_3 ), .I3(rd_addr_r[1]), .O(n11124));
    defparam rd_addr_r_0__bdd_4_lut_9515.LUT_INIT = 16'he4aa;
    SB_DFF i911_912 (.Q(\REG.mem_9_3 ), .C(FIFO_CLK_c), .D(n4275));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11124_bdd_4_lut (.I0(n11124), .I1(\REG.mem_41_3 ), .I2(\REG.mem_40_3 ), 
            .I3(rd_addr_r[1]), .O(n11127));
    defparam n11124_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i908_909 (.Q(\REG.mem_9_2 ), .C(FIFO_CLK_c), .D(n4274));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3951_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_52_15 ), .O(n5040));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3951_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4128_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_63_5 ), .O(n5217));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4128_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i905_906 (.Q(\REG.mem_9_1 ), .C(FIFO_CLK_c), .D(n4273));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3950_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_52_14 ), .O(n5039));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3950_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_10000 (.I0(rd_addr_r[2]), .I1(n11271), 
            .I2(n10779), .I3(rd_addr_r[3]), .O(n11694));
    defparam rd_addr_r_2__bdd_4_lut_10000.LUT_INIT = 16'he4aa;
    SB_LUT4 n11694_bdd_4_lut (.I0(n11694), .I1(n11409), .I2(n10022), .I3(rd_addr_r[3]), 
            .O(n10493));
    defparam n11694_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3949_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_52_13 ), .O(n5038));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3949_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i902_903 (.Q(\REG.mem_9_0 ), .C(FIFO_CLK_c), .D(n4272));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i8332_3_lut (.I0(n11679), .I1(n11505), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9874));
    defparam i8332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3948_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_52_12 ), .O(n5037));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3948_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4127_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_63_4 ), .O(n5216));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4127_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4126_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_63_3 ), .O(n5215));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4126_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3947_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_52_11 ), .O(n5036));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3947_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(FIFO_CLK_c), .D(n4271));   // src/fifo_dc_32_lut_gen.v(308[21] 324[24])
    SB_LUT4 i3946_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_52_10 ), .O(n5035));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3946_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9510 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_15 ), 
            .I2(\REG.mem_55_15 ), .I3(rd_addr_r[1]), .O(n11118));
    defparam rd_addr_r_0__bdd_4_lut_9510.LUT_INIT = 16'he4aa;
    SB_LUT4 i4125_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_63_2 ), .O(n5214));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4125_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8595_3_lut (.I0(\REG.mem_32_6 ), .I1(\REG.mem_33_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10137));
    defparam i8595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4124_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_63_1 ), .O(n5213));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4124_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8596_3_lut (.I0(\REG.mem_34_6 ), .I1(\REG.mem_35_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10138));
    defparam i8596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_10144 (.I0(rd_addr_r[3]), .I1(n10422), 
            .I2(n10423), .I3(rd_addr_r[4]), .O(n11688));
    defparam rd_addr_r_3__bdd_4_lut_10144.LUT_INIT = 16'he4aa;
    SB_DFF wr_addr_r__i3 (.Q(wr_addr_r[3]), .C(FIFO_CLK_c), .D(n4270));   // src/fifo_dc_32_lut_gen.v(308[21] 324[24])
    SB_LUT4 n11118_bdd_4_lut (.I0(n11118), .I1(\REG.mem_53_15 ), .I2(\REG.mem_52_15 ), 
            .I3(rd_addr_r[1]), .O(n11121));
    defparam n11118_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3945_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_52_9 ), .O(n5034));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3945_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9505 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_5 ), 
            .I2(\REG.mem_59_5 ), .I3(rd_addr_r[1]), .O(n11112));
    defparam rd_addr_r_0__bdd_4_lut_9505.LUT_INIT = 16'he4aa;
    SB_LUT4 i3944_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_52_8 ), .O(n5033));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3944_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11112_bdd_4_lut (.I0(n11112), .I1(\REG.mem_57_5 ), .I2(\REG.mem_56_5 ), 
            .I3(rd_addr_r[1]), .O(n11115));
    defparam n11112_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF wr_addr_r__i4 (.Q(wr_addr_r[4]), .C(FIFO_CLK_c), .D(n4269));   // src/fifo_dc_32_lut_gen.v(308[21] 324[24])
    SB_LUT4 i3943_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_52_7 ), .O(n5032));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3943_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3942_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_52_6 ), .O(n5031));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3942_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11688_bdd_4_lut (.I0(n11688), .I1(n10351), .I2(n10350), .I3(rd_addr_r[4]), 
            .O(n11691));
    defparam n11688_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3941_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_52_5 ), .O(n5030));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3941_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8641_3_lut (.I0(\REG.mem_38_6 ), .I1(\REG.mem_39_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10183));
    defparam i8641_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF wr_addr_r__i5 (.Q(wr_addr_r[5]), .C(FIFO_CLK_c), .D(n4268));   // src/fifo_dc_32_lut_gen.v(308[21] 324[24])
    SB_DFF wp_sync1_r__i0 (.Q(wp_sync1_r[0]), .C(DEBUG_6_c), .D(n4107));   // src/fifo_dc_32_lut_gen.v(602[21] 614[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9990 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_7 ), 
            .I2(\REG.mem_11_7 ), .I3(rd_addr_r[1]), .O(n11682));
    defparam rd_addr_r_0__bdd_4_lut_9990.LUT_INIT = 16'he4aa;
    SB_LUT4 n11682_bdd_4_lut (.I0(n11682), .I1(\REG.mem_9_7 ), .I2(\REG.mem_8_7 ), 
            .I3(rd_addr_r[1]), .O(n11685));
    defparam n11682_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8640_3_lut (.I0(\REG.mem_36_6 ), .I1(\REG.mem_37_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10182));
    defparam i8640_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF wr_addr_r__i6 (.Q(\wr_addr_r[6] ), .C(FIFO_CLK_c), .D(n4266));   // src/fifo_dc_32_lut_gen.v(308[21] 324[24])
    SB_LUT4 i8724_3_lut (.I0(\REG.mem_32_13 ), .I1(\REG.mem_33_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10266));
    defparam i8724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9975 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_0 ), 
            .I2(\REG.mem_27_0 ), .I3(rd_addr_r[1]), .O(n11676));
    defparam rd_addr_r_0__bdd_4_lut_9975.LUT_INIT = 16'he4aa;
    SB_LUT4 i3940_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_52_4 ), .O(n5029));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3940_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8725_3_lut (.I0(\REG.mem_34_13 ), .I1(\REG.mem_35_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10267));
    defparam i8725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_en_i_I_0_2_lut (.I0(DEBUG_9_c), .I1(DEBUG_1_c), .I2(GND_net), 
            .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(239[29:51])
    defparam rd_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9500 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_10 ), 
            .I2(\REG.mem_15_10 ), .I3(rd_addr_r[1]), .O(n11106));
    defparam rd_addr_r_0__bdd_4_lut_9500.LUT_INIT = 16'he4aa;
    SB_LUT4 i3939_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_52_3 ), .O(n5028));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3939_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11106_bdd_4_lut (.I0(n11106), .I1(\REG.mem_13_10 ), .I2(\REG.mem_12_10 ), 
            .I3(rd_addr_r[1]), .O(n11109));
    defparam n11106_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4120_3_lut_4_lut (.I0(n67), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_63_0 ), .O(n5209));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i4120_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i851_852 (.Q(\REG.mem_8_15 ), .C(FIFO_CLK_c), .D(n4265));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11676_bdd_4_lut (.I0(n11676), .I1(\REG.mem_25_0 ), .I2(\REG.mem_24_0 ), 
            .I3(rd_addr_r[1]), .O(n11679));
    defparam n11676_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8534_3_lut (.I0(n11535), .I1(n11607), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n10076));
    defparam i8534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9970 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_11 ), 
            .I2(\REG.mem_47_11 ), .I3(rd_addr_r[1]), .O(n11670));
    defparam rd_addr_r_0__bdd_4_lut_9970.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9495 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_2 ), 
            .I2(\REG.mem_51_2 ), .I3(rd_addr_r[1]), .O(n11100));
    defparam rd_addr_r_0__bdd_4_lut_9495.LUT_INIT = 16'he4aa;
    SB_LUT4 i3938_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_52_2 ), .O(n5027));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3938_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11100_bdd_4_lut (.I0(n11100), .I1(\REG.mem_49_2 ), .I2(\REG.mem_48_2 ), 
            .I3(rd_addr_r[1]), .O(n10190));
    defparam n11100_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11670_bdd_4_lut (.I0(n11670), .I1(\REG.mem_45_11 ), .I2(\REG.mem_44_11 ), 
            .I3(rd_addr_r[1]), .O(n11673));
    defparam n11670_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i848_849 (.Q(\REG.mem_8_14 ), .C(FIFO_CLK_c), .D(n4264));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3937_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_52_1 ), .O(n5026));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3937_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3936_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_52_0 ), .O(n5025));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3936_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9490 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_5 ), 
            .I2(\REG.mem_15_5 ), .I3(rd_addr_r[1]), .O(n11094));
    defparam rd_addr_r_0__bdd_4_lut_9490.LUT_INIT = 16'he4aa;
    SB_LUT4 i8357_3_lut (.I0(n11349), .I1(n12279), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_237 [0]));
    defparam i8357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n11094_bdd_4_lut (.I0(n11094), .I1(\REG.mem_13_5 ), .I2(\REG.mem_12_5 ), 
            .I3(rd_addr_r[1]), .O(n11097));
    defparam n11094_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8734_3_lut (.I0(\REG.mem_38_13 ), .I1(\REG.mem_39_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10276));
    defparam i8734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8733_3_lut (.I0(\REG.mem_36_13 ), .I1(\REG.mem_37_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10275));
    defparam i8733_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i845_846 (.Q(\REG.mem_8_13 ), .C(FIFO_CLK_c), .D(n4263));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_4__bdd_4_lut_10030 (.I0(rd_addr_r[4]), .I1(n10749), 
            .I2(n10481), .I3(rd_addr_r[5]), .O(n11664));
    defparam rd_addr_r_4__bdd_4_lut_10030.LUT_INIT = 16'he4aa;
    SB_LUT4 n11664_bdd_4_lut (.I0(n11664), .I1(n11025), .I2(n11625), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_237 [5]));
    defparam n11664_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9530 (.I0(rd_addr_r[1]), .I1(n10392), 
            .I2(n10393), .I3(rd_addr_r[2]), .O(n11088));
    defparam rd_addr_r_1__bdd_4_lut_9530.LUT_INIT = 16'he4aa;
    SB_LUT4 n11088_bdd_4_lut (.I0(n11088), .I1(n10375), .I2(n10374), .I3(rd_addr_r[2]), 
            .O(n11091));
    defparam n11088_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i842_843 (.Q(\REG.mem_8_12 ), .C(FIFO_CLK_c), .D(n4262));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i36_2_lut_3_lut (.I0(n11_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n36_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i36_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_9620 (.I0(rd_addr_r[3]), .I1(n9507), 
            .I2(n9508), .I3(rd_addr_r[4]), .O(n11082));
    defparam rd_addr_r_3__bdd_4_lut_9620.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9985 (.I0(rd_addr_r[2]), .I1(n10983), 
            .I2(n10743), .I3(rd_addr_r[3]), .O(n11658));
    defparam rd_addr_r_2__bdd_4_lut_9985.LUT_INIT = 16'he4aa;
    SB_DFF i146_147 (.Q(\REG.mem_1_4 ), .C(FIFO_CLK_c), .D(n4106));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3015_2_lut_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_p1_w[0]), 
            .I2(rd_fifo_en_w), .I3(reset_all), .O(n4104));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam i3015_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 EnabledDecoder_2_i35_2_lut_3_lut (.I0(n11_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n35_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i35_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_nxt_c_6__I_0_130_i1_2_lut_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_p1_w[0]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_176[1] ), .O(rd_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(548[59:99])
    defparam rd_addr_nxt_c_6__I_0_130_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_DFF i839_840 (.Q(\REG.mem_8_11 ), .C(FIFO_CLK_c), .D(n4261));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9219 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_5 ), 
            .I2(\REG.mem_43_5 ), .I3(rd_addr_r[1]), .O(n10764));
    defparam rd_addr_r_0__bdd_4_lut_9219.LUT_INIT = 16'he4aa;
    SB_LUT4 n10746_bdd_4_lut (.I0(n10746), .I1(n9824), .I2(n9812), .I3(rd_addr_r[3]), 
            .O(n10749));
    defparam n10746_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n10764_bdd_4_lut (.I0(n10764), .I1(\REG.mem_41_5 ), .I2(\REG.mem_40_5 ), 
            .I3(rd_addr_r[1]), .O(n9827));
    defparam n10764_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i96_2_lut_3_lut (.I0(n31_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n52));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i96_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_DFF i149_150 (.Q(\REG.mem_1_5 ), .C(FIFO_CLK_c), .D(n4105));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11658_bdd_4_lut (.I0(n11658), .I1(n11211), .I2(n11619), .I3(rd_addr_r[3]), 
            .O(n10061));
    defparam n11658_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3064_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_1_15 ), .O(n4153));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3064_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(DEBUG_6_c), .D(n4104));   // src/fifo_dc_32_lut_gen.v(558[21] 574[24])
    SB_LUT4 i3063_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_1_14 ), .O(n4152));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3063_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3062_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_1_13 ), .O(n4151));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3062_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3061_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_1_12 ), .O(n4150));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3061_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3060_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_1_11 ), .O(n4149));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3060_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3059_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_1_10 ), .O(n4148));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3059_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3058_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_1_9 ), .O(n4147));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3058_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2986_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_1_0 ), .O(n4075));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i2986_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3013_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_1_6 ), .O(n4102));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3013_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n10710_bdd_4_lut (.I0(n10710), .I1(\REG.mem_29_13 ), .I2(\REG.mem_28_13 ), 
            .I3(rd_addr_r[1]), .O(n10713));
    defparam n10710_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i836_837 (.Q(\REG.mem_8_10 ), .C(FIFO_CLK_c), .D(n4260));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3017_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_1_4 ), .O(n4106));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3017_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3057_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_1_8 ), .O(n4146));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3057_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9965 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_8 ), 
            .I2(\REG.mem_11_8 ), .I3(rd_addr_r[1]), .O(n11652));
    defparam rd_addr_r_0__bdd_4_lut_9965.LUT_INIT = 16'he4aa;
    SB_LUT4 i2981_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_1_2 ), .O(n4070));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i2981_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n11652_bdd_4_lut (.I0(n11652), .I1(\REG.mem_9_8 ), .I2(\REG.mem_8_8 ), 
            .I3(rd_addr_r[1]), .O(n11655));
    defparam n11652_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11082_bdd_4_lut (.I0(n11082), .I1(n10432), .I2(n10431), .I3(rd_addr_r[4]), 
            .O(n11085));
    defparam n11082_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i833_834 (.Q(\REG.mem_8_9 ), .C(FIFO_CLK_c), .D(n4259));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i2985_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_1_1 ), .O(n4074));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i2985_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i830_831 (.Q(\REG.mem_8_8 ), .C(FIFO_CLK_c), .D(n4258));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i827_828 (.Q(\REG.mem_8_7 ), .C(FIFO_CLK_c), .D(n4257));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i824_825 (.Q(\REG.mem_8_6 ), .C(FIFO_CLK_c), .D(n4256));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i821_822 (.Q(\REG.mem_8_5 ), .C(FIFO_CLK_c), .D(n4255));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i818_819 (.Q(\REG.mem_8_4 ), .C(FIFO_CLK_c), .D(n4254));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i815_816 (.Q(\REG.mem_8_3 ), .C(FIFO_CLK_c), .D(n4253));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i812_813 (.Q(\REG.mem_8_2 ), .C(FIFO_CLK_c), .D(n4252));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i809_810 (.Q(\REG.mem_8_1 ), .C(FIFO_CLK_c), .D(n4251));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i806_807 (.Q(\REG.mem_8_0 ), .C(FIFO_CLK_c), .D(n4250));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i755_756 (.Q(\REG.mem_7_15 ), .C(FIFO_CLK_c), .D(n4249));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i752_753 (.Q(\REG.mem_7_14 ), .C(FIFO_CLK_c), .D(n4248));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i749_750 (.Q(\REG.mem_7_13 ), .C(FIFO_CLK_c), .D(n4247));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i746_747 (.Q(\REG.mem_7_12 ), .C(FIFO_CLK_c), .D(n4246));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i743_744 (.Q(\REG.mem_7_11 ), .C(FIFO_CLK_c), .D(n4245));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i740_741 (.Q(\REG.mem_7_10 ), .C(FIFO_CLK_c), .D(n4244));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i737_738 (.Q(\REG.mem_7_9 ), .C(FIFO_CLK_c), .D(n4243));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i734_735 (.Q(\REG.mem_7_8 ), .C(FIFO_CLK_c), .D(n4242));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i731_732 (.Q(\REG.mem_7_7 ), .C(FIFO_CLK_c), .D(n4241));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i728_729 (.Q(\REG.mem_7_6 ), .C(FIFO_CLK_c), .D(n4240));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i725_726 (.Q(\REG.mem_7_5 ), .C(FIFO_CLK_c), .D(n4239));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i722_723 (.Q(\REG.mem_7_4 ), .C(FIFO_CLK_c), .D(n4238));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i719_720 (.Q(\REG.mem_7_3 ), .C(FIFO_CLK_c), .D(n4237));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i716_717 (.Q(\REG.mem_7_2 ), .C(FIFO_CLK_c), .D(n4236));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i713_714 (.Q(\REG.mem_7_1 ), .C(FIFO_CLK_c), .D(n4235));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i710_711 (.Q(\REG.mem_7_0 ), .C(FIFO_CLK_c), .D(n4234));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i659_660 (.Q(\REG.mem_6_15 ), .C(FIFO_CLK_c), .D(n4233));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i656_657 (.Q(\REG.mem_6_14 ), .C(FIFO_CLK_c), .D(n4232));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i653_654 (.Q(\REG.mem_6_13 ), .C(FIFO_CLK_c), .D(n4231));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i650_651 (.Q(\REG.mem_6_12 ), .C(FIFO_CLK_c), .D(n4230));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i647_648 (.Q(\REG.mem_6_11 ), .C(FIFO_CLK_c), .D(n4229));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i644_645 (.Q(\REG.mem_6_10 ), .C(FIFO_CLK_c), .D(n4228));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i641_642 (.Q(\REG.mem_6_9 ), .C(FIFO_CLK_c), .D(n4227));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i638_639 (.Q(\REG.mem_6_8 ), .C(FIFO_CLK_c), .D(n4226));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i635_636 (.Q(\REG.mem_6_7 ), .C(FIFO_CLK_c), .D(n4225));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i632_633 (.Q(\REG.mem_6_6 ), .C(FIFO_CLK_c), .D(n4224));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i629_630 (.Q(\REG.mem_6_5 ), .C(FIFO_CLK_c), .D(n4223));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i626_627 (.Q(\REG.mem_6_4 ), .C(FIFO_CLK_c), .D(n4222));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i623_624 (.Q(\REG.mem_6_3 ), .C(FIFO_CLK_c), .D(n4221));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i620_621 (.Q(\REG.mem_6_2 ), .C(FIFO_CLK_c), .D(n4220));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i617_618 (.Q(\REG.mem_6_1 ), .C(FIFO_CLK_c), .D(n4219));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i614_615 (.Q(\REG.mem_6_0 ), .C(FIFO_CLK_c), .D(n4218));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i563_564 (.Q(\REG.mem_5_15 ), .C(FIFO_CLK_c), .D(n4217));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i560_561 (.Q(\REG.mem_5_14 ), .C(FIFO_CLK_c), .D(n4216));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i557_558 (.Q(\REG.mem_5_13 ), .C(FIFO_CLK_c), .D(n4215));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i554_555 (.Q(\REG.mem_5_12 ), .C(FIFO_CLK_c), .D(n4214));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i551_552 (.Q(\REG.mem_5_11 ), .C(FIFO_CLK_c), .D(n4213));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i548_549 (.Q(\REG.mem_5_10 ), .C(FIFO_CLK_c), .D(n4212));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i545_546 (.Q(\REG.mem_5_9 ), .C(FIFO_CLK_c), .D(n4211));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i542_543 (.Q(\REG.mem_5_8 ), .C(FIFO_CLK_c), .D(n4210));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i539_540 (.Q(\REG.mem_5_7 ), .C(FIFO_CLK_c), .D(n4209));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i536_537 (.Q(\REG.mem_5_6 ), .C(FIFO_CLK_c), .D(n4208));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i533_534 (.Q(\REG.mem_5_5 ), .C(FIFO_CLK_c), .D(n4207));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i530_531 (.Q(\REG.mem_5_4 ), .C(FIFO_CLK_c), .D(n4206));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i527_528 (.Q(\REG.mem_5_3 ), .C(FIFO_CLK_c), .D(n4205));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i524_525 (.Q(\REG.mem_5_2 ), .C(FIFO_CLK_c), .D(n4204));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i521_522 (.Q(\REG.mem_5_1 ), .C(FIFO_CLK_c), .D(n4203));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i518_519 (.Q(\REG.mem_5_0 ), .C(FIFO_CLK_c), .D(n4202));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF rp_sync2_r__i0 (.Q(rp_sync2_r[0]), .C(FIFO_CLK_c), .D(n4103));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_LUT4 EnabledDecoder_2_i95_2_lut_3_lut (.I0(n31_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n20));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i95_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i3003_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_1_7 ), .O(n4092));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3003_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3177_2_lut_4_lut (.I0(\wr_addr_r[6] ), .I1(wr_addr_p1_w[6]), 
            .I2(write_to_dc32_fifo), .I3(reset_all), .O(n4266));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam i3177_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i3016_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_1_5 ), .O(n4105));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3016_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3029_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_1_3 ), .O(n4118));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3029_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n10728_bdd_4_lut (.I0(n10728), .I1(n9557), .I2(n9551), .I3(rd_addr_r[3]), 
            .O(n10731));
    defparam n10728_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_10005 (.I0(rd_addr_r[1]), .I1(n10029), 
            .I2(n10030), .I3(rd_addr_r[2]), .O(n11646));
    defparam rd_addr_r_1__bdd_4_lut_10005.LUT_INIT = 16'he4aa;
    SB_DFF i467_468 (.Q(\REG.mem_4_15 ), .C(FIFO_CLK_c), .D(n4201));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 wr_addr_nxt_c_6__I_0_128_i6_2_lut_4_lut (.I0(\wr_addr_r[6] ), 
            .I1(wr_addr_p1_w[6]), .I2(write_to_dc32_fifo), .I3(\wr_addr_nxt_c[5] ), 
            .O(wr_grey_w[5]));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam wr_addr_nxt_c_6__I_0_128_i6_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 EnabledDecoder_2_i94_2_lut_3_lut (.I0(n29), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n53));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i94_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_DFF i152_153 (.Q(\REG.mem_1_6 ), .C(FIFO_CLK_c), .D(n4102));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF rp_sync1_r__i0 (.Q(rp_sync1_r[0]), .C(FIFO_CLK_c), .D(n4101));   // src/fifo_dc_32_lut_gen.v(352[21] 364[24])
    SB_LUT4 n11646_bdd_4_lut (.I0(n11646), .I1(n10018), .I2(n10017), .I3(rd_addr_r[2]), 
            .O(n10066));
    defparam n11646_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9615 (.I0(rd_addr_r[2]), .I1(n10406), 
            .I2(n10409), .I3(rd_addr_r[3]), .O(n11076));
    defparam rd_addr_r_2__bdd_4_lut_9615.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9955 (.I0(rd_addr_r[2]), .I1(n9677), 
            .I2(n10851), .I3(rd_addr_r[3]), .O(n11640));
    defparam rd_addr_r_2__bdd_4_lut_9955.LUT_INIT = 16'he4aa;
    SB_LUT4 n11076_bdd_4_lut (.I0(n11076), .I1(n10400), .I2(n10397), .I3(rd_addr_r[3]), 
            .O(n11079));
    defparam n11076_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11640_bdd_4_lut (.I0(n11640), .I1(n9539), .I2(n11583), .I3(rd_addr_r[3]), 
            .O(n10502));
    defparam n11640_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3628_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_33_15 ), .O(n4717));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3628_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_9960 (.I0(rd_addr_r[4]), .I1(n10487), 
            .I2(n10493), .I3(rd_addr_r[5]), .O(n11634));
    defparam rd_addr_r_4__bdd_4_lut_9960.LUT_INIT = 16'he4aa;
    SB_LUT4 n11634_bdd_4_lut (.I0(n11634), .I1(n10373), .I2(n10313), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_237 [9]));
    defparam n11634_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9485 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_8 ), 
            .I2(\REG.mem_43_8 ), .I3(rd_addr_r[1]), .O(n11070));
    defparam rd_addr_r_0__bdd_4_lut_9485.LUT_INIT = 16'he4aa;
    SB_LUT4 i3627_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_33_14 ), .O(n4716));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3627_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3626_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_33_13 ), .O(n4715));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3626_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3625_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_33_12 ), .O(n4714));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3625_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i464_465 (.Q(\REG.mem_4_14 ), .C(FIFO_CLK_c), .D(n4200));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3624_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_33_11 ), .O(n4713));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3624_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9950 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_10 ), 
            .I2(\REG.mem_23_10 ), .I3(rd_addr_r[1]), .O(n11628));
    defparam rd_addr_r_0__bdd_4_lut_9950.LUT_INIT = 16'he4aa;
    SB_LUT4 n11628_bdd_4_lut (.I0(n11628), .I1(\REG.mem_21_10 ), .I2(\REG.mem_20_10 ), 
            .I3(rd_addr_r[1]), .O(n9722));
    defparam n11628_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i93_2_lut_3_lut (.I0(n29), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n21));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i93_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i3623_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_33_10 ), .O(n4712));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3623_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3622_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_33_9 ), .O(n4711));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3622_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11070_bdd_4_lut (.I0(n11070), .I1(\REG.mem_41_8 ), .I2(\REG.mem_40_8 ), 
            .I3(rd_addr_r[1]), .O(n11073));
    defparam n11070_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3621_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_33_8 ), .O(n4710));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3621_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3180_2_lut_4_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(write_to_dc32_fifo), .I3(reset_all), .O(n4269));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam i3180_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_DFF i461_462 (.Q(\REG.mem_4_13 ), .C(FIFO_CLK_c), .D(n4199));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3620_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_33_7 ), .O(n4709));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3620_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_9940 (.I0(rd_addr_r[2]), .I1(n11145), 
            .I2(n11097), .I3(rd_addr_r[3]), .O(n11622));
    defparam rd_addr_r_2__bdd_4_lut_9940.LUT_INIT = 16'he4aa;
    SB_LUT4 n11622_bdd_4_lut (.I0(n11622), .I1(n11169), .I2(n11319), .I3(rd_addr_r[3]), 
            .O(n11625));
    defparam n11622_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_nxt_c_6__I_0_128_i4_2_lut_4_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(write_to_dc32_fifo), .I3(\wr_addr_nxt_c[3] ), .O(wr_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam wr_addr_nxt_c_6__I_0_128_i4_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i3619_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_33_6 ), .O(n4708));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3619_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9214 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_7 ), 
            .I2(\REG.mem_15_7 ), .I3(rd_addr_r[1]), .O(n10758));
    defparam rd_addr_r_0__bdd_4_lut_9214.LUT_INIT = 16'he4aa;
    SB_LUT4 i3618_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_33_5 ), .O(n4707));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3618_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9930 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_12 ), 
            .I2(\REG.mem_3_12 ), .I3(rd_addr_r[1]), .O(n11616));
    defparam rd_addr_r_0__bdd_4_lut_9930.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_nxt_c_6__I_0_128_i5_2_lut_4_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(write_to_dc32_fifo), .I3(\wr_addr_nxt_c[5] ), .O(wr_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam wr_addr_nxt_c_6__I_0_128_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i3617_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_33_4 ), .O(n4706));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3617_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n10758_bdd_4_lut (.I0(n10758), .I1(\REG.mem_13_7 ), .I2(\REG.mem_12_7 ), 
            .I3(rd_addr_r[1]), .O(n10761));
    defparam n10758_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i458_459 (.Q(\REG.mem_4_12 ), .C(FIFO_CLK_c), .D(n4198));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i455_456 (.Q(\REG.mem_4_11 ), .C(FIFO_CLK_c), .D(n4197));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i452_453 (.Q(\REG.mem_4_10 ), .C(FIFO_CLK_c), .D(n4196));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i449_450 (.Q(\REG.mem_4_9 ), .C(FIFO_CLK_c), .D(n4195));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3616_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_33_3 ), .O(n4705));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3616_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11616_bdd_4_lut (.I0(n11616), .I1(\REG.mem_1_12 ), .I2(\REG.mem_0_12 ), 
            .I3(rd_addr_r[1]), .O(n11619));
    defparam n11616_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i130_2_lut_3_lut (.I0(n33), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n35));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i130_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i446_447 (.Q(\REG.mem_4_8 ), .C(FIFO_CLK_c), .D(n4194));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i443_444 (.Q(\REG.mem_4_7 ), .C(FIFO_CLK_c), .D(n4193));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9920 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_6 ), 
            .I2(\REG.mem_31_6 ), .I3(rd_addr_r[1]), .O(n11610));
    defparam rd_addr_r_0__bdd_4_lut_9920.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9465 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_3 ), 
            .I2(\REG.mem_47_3 ), .I3(rd_addr_r[1]), .O(n11058));
    defparam rd_addr_r_0__bdd_4_lut_9465.LUT_INIT = 16'he4aa;
    SB_LUT4 n11058_bdd_4_lut (.I0(n11058), .I1(\REG.mem_45_3 ), .I2(\REG.mem_44_3 ), 
            .I3(rd_addr_r[1]), .O(n11061));
    defparam n11058_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i440_441 (.Q(\REG.mem_4_6 ), .C(FIFO_CLK_c), .D(n4192));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i155_156 (.Q(\REG.mem_1_7 ), .C(FIFO_CLK_c), .D(n4092));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 i3615_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_33_2 ), .O(n4704));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3615_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n11610_bdd_4_lut (.I0(n11610), .I1(\REG.mem_29_6 ), .I2(\REG.mem_28_6 ), 
            .I3(rd_addr_r[1]), .O(n10073));
    defparam n11610_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3614_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_33_1 ), .O(n4703));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3614_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3613_3_lut_4_lut (.I0(n40_adj_1070), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_33_0 ), .O(n4702));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3613_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9480 (.I0(rd_addr_r[1]), .I1(n10338), 
            .I2(n10339), .I3(rd_addr_r[2]), .O(n11052));
    defparam rd_addr_r_1__bdd_4_lut_9480.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9945 (.I0(rd_addr_r[1]), .I1(n9900), 
            .I2(n9901), .I3(rd_addr_r[2]), .O(n11604));
    defparam rd_addr_r_1__bdd_4_lut_9945.LUT_INIT = 16'he4aa;
    SB_DFF i134_135 (.Q(\REG.mem_1_0 ), .C(FIFO_CLK_c), .D(n4075));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11604_bdd_4_lut (.I0(n11604), .I1(n9877), .I2(n9876), .I3(rd_addr_r[2]), 
            .O(n11607));
    defparam n11604_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9915 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_10 ), 
            .I2(\REG.mem_3_10 ), .I3(rd_addr_r[1]), .O(n11598));
    defparam rd_addr_r_0__bdd_4_lut_9915.LUT_INIT = 16'he4aa;
    SB_LUT4 n11052_bdd_4_lut (.I0(n11052), .I1(n10327), .I2(n10326), .I3(rd_addr_r[2]), 
            .O(n11055));
    defparam n11052_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11598_bdd_4_lut (.I0(n11598), .I1(\REG.mem_1_10 ), .I2(\REG.mem_0_10 ), 
            .I3(rd_addr_r[1]), .O(n10511));
    defparam n11598_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i137_138 (.Q(\REG.mem_1_1 ), .C(FIFO_CLK_c), .D(n4074));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i20_2_lut (.I0(n11_c), .I1(wr_addr_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n20_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i20_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_9451 (.I0(rd_addr_r[1]), .I1(n10335), 
            .I2(n10336), .I3(rd_addr_r[2]), .O(n11046));
    defparam rd_addr_r_1__bdd_4_lut_9451.LUT_INIT = 16'he4aa;
    SB_DFF i437_438 (.Q(\REG.mem_4_5 ), .C(FIFO_CLK_c), .D(n4191));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i129_2_lut_3_lut (.I0(n33), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n3));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i129_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3028_2_lut_4_lut (.I0(wr_addr_r[0]), .I1(wr_addr_p1_w[0]), 
            .I2(write_to_dc32_fifo), .I3(reset_all), .O(n4117));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam i3028_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 wr_addr_nxt_c_6__I_0_128_i1_2_lut_4_lut (.I0(wr_addr_r[0]), .I1(wr_addr_p1_w[0]), 
            .I2(write_to_dc32_fifo), .I3(\wr_addr_nxt_c[1] ), .O(wr_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(303[33:89])
    defparam wr_addr_nxt_c_6__I_0_128_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 n11046_bdd_4_lut (.I0(n11046), .I1(n10315), .I2(n10314), .I3(rd_addr_r[2]), 
            .O(n11049));
    defparam n11046_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9456 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_13 ), 
            .I2(\REG.mem_15_13 ), .I3(rd_addr_r[1]), .O(n11040));
    defparam rd_addr_r_0__bdd_4_lut_9456.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i128_2_lut_3_lut (.I0(n31_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n36));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i128_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i90_2_lut_3_lut (.I0(n25_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n55));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i90_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9905 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_7 ), 
            .I2(\REG.mem_27_7 ), .I3(rd_addr_r[1]), .O(n11592));
    defparam rd_addr_r_0__bdd_4_lut_9905.LUT_INIT = 16'he4aa;
    SB_LUT4 n11592_bdd_4_lut (.I0(n11592), .I1(\REG.mem_25_7 ), .I2(\REG.mem_24_7 ), 
            .I3(rd_addr_r[1]), .O(n11595));
    defparam n11592_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i434_435 (.Q(\REG.mem_4_4 ), .C(FIFO_CLK_c), .D(n4190));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i431_432 (.Q(\REG.mem_4_3 ), .C(FIFO_CLK_c), .D(n4189));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i428_429 (.Q(\REG.mem_4_2 ), .C(FIFO_CLK_c), .D(n4188));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11040_bdd_4_lut (.I0(n11040), .I1(\REG.mem_13_13 ), .I2(\REG.mem_12_13 ), 
            .I3(rd_addr_r[1]), .O(n11043));
    defparam n11040_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i425_426 (.Q(\REG.mem_4_1 ), .C(FIFO_CLK_c), .D(n4187));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i422_423 (.Q(\REG.mem_4_0 ), .C(FIFO_CLK_c), .D(n4186));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9209 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_0 ), 
            .I2(\REG.mem_51_0 ), .I3(rd_addr_r[1]), .O(n10752));
    defparam rd_addr_r_0__bdd_4_lut_9209.LUT_INIT = 16'he4aa;
    SB_DFF i371_372 (.Q(\REG.mem_3_15 ), .C(FIFO_CLK_c), .D(n4185));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9900 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_8 ), 
            .I2(\REG.mem_15_8 ), .I3(rd_addr_r[1]), .O(n11586));
    defparam rd_addr_r_0__bdd_4_lut_9900.LUT_INIT = 16'he4aa;
    SB_DFF i368_369 (.Q(\REG.mem_3_14 ), .C(FIFO_CLK_c), .D(n4184));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i365_366 (.Q(\REG.mem_3_13 ), .C(FIFO_CLK_c), .D(n4183));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 n11586_bdd_4_lut (.I0(n11586), .I1(\REG.mem_13_8 ), .I2(\REG.mem_12_8 ), 
            .I3(rd_addr_r[1]), .O(n11589));
    defparam n11586_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9441 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_2 ), 
            .I2(\REG.mem_55_2 ), .I3(rd_addr_r[1]), .O(n11034));
    defparam rd_addr_r_0__bdd_4_lut_9441.LUT_INIT = 16'he4aa;
    SB_LUT4 n11034_bdd_4_lut (.I0(n11034), .I1(\REG.mem_53_2 ), .I2(\REG.mem_52_2 ), 
            .I3(rd_addr_r[1]), .O(n10199));
    defparam n11034_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9895 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_6 ), 
            .I2(\REG.mem_3_6 ), .I3(rd_addr_r[1]), .O(n11580));
    defparam rd_addr_r_0__bdd_4_lut_9895.LUT_INIT = 16'he4aa;
    SB_LUT4 n11580_bdd_4_lut (.I0(n11580), .I1(\REG.mem_1_6 ), .I2(\REG.mem_0_6 ), 
            .I3(rd_addr_r[1]), .O(n11583));
    defparam n11580_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_9980 (.I0(rd_addr_r[3]), .I1(n11529), 
            .I2(n10066), .I3(rd_addr_r[4]), .O(n11574));
    defparam rd_addr_r_3__bdd_4_lut_9980.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i89_2_lut_3_lut (.I0(n25_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n23));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i89_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF i140_141 (.Q(\REG.mem_1_2 ), .C(FIFO_CLK_c), .D(n4070));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i127_2_lut_3_lut (.I0(n31_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n4));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i127_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n11574_bdd_4_lut (.I0(n11574), .I1(n10054), .I2(n11523), .I3(rd_addr_r[4]), 
            .O(n11577));
    defparam n11574_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i362_363 (.Q(\REG.mem_3_12 ), .C(FIFO_CLK_c), .D(n4182));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i359_360 (.Q(\REG.mem_3_11 ), .C(FIFO_CLK_c), .D(n4181));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_DFF i356_357 (.Q(\REG.mem_3_10 ), .C(FIFO_CLK_c), .D(n4180));   // src/fifo_dc_32_lut_gen.v(876[78:81])
    SB_LUT4 EnabledDecoder_2_i34_2_lut_3_lut (.I0(n9_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n34));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i34_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i32_2_lut_3_lut (.I0(n12_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n32));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i32_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_9436 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_2 ), 
            .I2(\REG.mem_59_2 ), .I3(rd_addr_r[1]), .O(n11028));
    defparam rd_addr_r_0__bdd_4_lut_9436.LUT_INIT = 16'he4aa;
    SB_LUT4 n11028_bdd_4_lut (.I0(n11028), .I1(\REG.mem_57_2 ), .I2(\REG.mem_56_2 ), 
            .I3(rd_addr_r[1]), .O(n10202));
    defparam n11028_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3611_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_32_15 ), .O(n4700));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3611_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3609_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_32_14 ), .O(n4698));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3609_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3608_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_32_13 ), .O(n4697));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3608_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3607_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_32_12 ), .O(n4696));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3607_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3606_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_32_11 ), .O(n4695));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3606_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3605_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_32_10 ), .O(n4694));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3605_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3604_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_32_9 ), .O(n4693));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3604_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3603_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_32_8 ), .O(n4692));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3603_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8442_3_lut (.I0(n10977), .I1(n10809), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9984));
    defparam i8442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8379_3_lut (.I0(\REG.mem_20_15 ), .I1(\REG.mem_21_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9921));
    defparam i8379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8380_3_lut (.I0(\REG.mem_22_15 ), .I1(\REG.mem_23_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9922));
    defparam i8380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3602_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_32_7 ), .O(n4691));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3602_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8350_3_lut (.I0(\REG.mem_18_15 ), .I1(\REG.mem_19_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9892));
    defparam i8350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8349_3_lut (.I0(\REG.mem_16_15 ), .I1(\REG.mem_17_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9891));
    defparam i8349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8175_3_lut (.I0(\REG.mem_52_4 ), .I1(\REG.mem_53_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9717));
    defparam i8175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8176_3_lut (.I0(\REG.mem_54_4 ), .I1(\REG.mem_55_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9718));
    defparam i8176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8173_3_lut (.I0(\REG.mem_50_4 ), .I1(\REG.mem_51_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9715));
    defparam i8173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8172_3_lut (.I0(\REG.mem_48_4 ), .I1(\REG.mem_49_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9714));
    defparam i8172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3601_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_32_6 ), .O(n4690));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3601_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8154_3_lut (.I0(\REG.mem_36_4 ), .I1(\REG.mem_37_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9696));
    defparam i8154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8155_3_lut (.I0(\REG.mem_38_4 ), .I1(\REG.mem_39_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9697));
    defparam i8155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8152_3_lut (.I0(\REG.mem_34_4 ), .I1(\REG.mem_35_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9694));
    defparam i8152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8151_3_lut (.I0(\REG.mem_32_4 ), .I1(\REG.mem_33_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9693));
    defparam i8151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3600_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_32_5 ), .O(n4689));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3600_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3599_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_32_4 ), .O(n4688));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3599_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3598_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_32_3 ), .O(n4687));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3598_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3597_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_32_2 ), .O(n4686));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3597_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3596_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_32_1 ), .O(n4685));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3596_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3595_3_lut_4_lut (.I0(n38), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_32_0 ), .O(n4684));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3595_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i106_2_lut_3_lut (.I0(n26_adj_1085), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n47));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i106_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i105_2_lut_3_lut (.I0(n26_adj_1085), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n15));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i105_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 EnabledDecoder_2_i73_2_lut_3_lut (.I0(n26_adj_1085), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n31));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i73_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i74_2_lut_3_lut (.I0(n26_adj_1085), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n63));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i74_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i25_2_lut_3_lut (.I0(n9_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n25_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i25_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i26_2_lut_3_lut (.I0(n9_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n26_adj_1085));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i26_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i10_2_lut_3_lut (.I0(write_to_dc32_fifo), .I1(wr_addr_r[0]), 
            .I2(wr_addr_r[1]), .I3(GND_net), .O(n10_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i10_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 EnabledDecoder_2_i9_2_lut_3_lut (.I0(write_to_dc32_fifo), .I1(wr_addr_r[0]), 
            .I2(wr_addr_r[1]), .I3(GND_net), .O(n9_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i9_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i8127_3_lut (.I0(\REG.mem_20_4 ), .I1(\REG.mem_21_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9669));
    defparam i8127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8128_3_lut (.I0(\REG.mem_22_4 ), .I1(\REG.mem_23_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9670));
    defparam i8128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8125_3_lut (.I0(\REG.mem_18_4 ), .I1(\REG.mem_19_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9667));
    defparam i8125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8124_3_lut (.I0(\REG.mem_16_4 ), .I1(\REG.mem_17_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9666));
    defparam i8124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8106_3_lut (.I0(\REG.mem_4_4 ), .I1(\REG.mem_5_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9648));
    defparam i8106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8107_3_lut (.I0(\REG.mem_6_4 ), .I1(\REG.mem_7_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9649));
    defparam i8107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8104_3_lut (.I0(\REG.mem_2_4 ), .I1(\REG.mem_3_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9646));
    defparam i8104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8103_3_lut (.I0(\REG.mem_0_4 ), .I1(\REG.mem_1_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9645));
    defparam i8103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7958_3_lut (.I0(n10875), .I1(n11691), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_237 [15]));
    defparam i7958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8012_3_lut (.I0(n11085), .I1(n12033), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_237 [13]));
    defparam i8012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8474_3_lut (.I0(n11481), .I1(n11889), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_237 [7]));
    defparam i8474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8219_3_lut (.I0(n11259), .I1(n11337), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_237 [4]));
    defparam i8219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3901_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_49_15 ), .O(n4990));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3901_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8385_3_lut (.I0(\REG.mem_12_1 ), .I1(\REG.mem_13_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9927));
    defparam i8385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8386_3_lut (.I0(\REG.mem_14_1 ), .I1(\REG.mem_15_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9928));
    defparam i8386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8383_3_lut (.I0(\REG.mem_10_1 ), .I1(\REG.mem_11_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9925));
    defparam i8383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8382_3_lut (.I0(\REG.mem_8_1 ), .I1(\REG.mem_9_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9924));
    defparam i8382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3900_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_49_14 ), .O(n4989));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3900_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3899_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_49_13 ), .O(n4988));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3899_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8540_3_lut (.I0(n11541), .I1(n11577), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_237 [1]));
    defparam i8540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3898_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_49_12 ), .O(n4987));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3898_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3897_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_49_11 ), .O(n4986));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3897_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3896_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_49_10 ), .O(n4985));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3896_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8090_3_lut (.I0(n11151), .I1(n9631), .I2(rd_addr_r[3]), .I3(GND_net), 
            .O(n9632));
    defparam i8090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8089_3_lut (.I0(n11703), .I1(n11673), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9631));
    defparam i8089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8111_3_lut (.I0(n11163), .I1(n9652), .I2(rd_addr_r[3]), .I3(GND_net), 
            .O(n9653));
    defparam i8111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8110_3_lut (.I0(n12339), .I1(n11709), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9652));
    defparam i8110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8970_3_lut (.I0(\REG.mem_52_11 ), .I1(\REG.mem_53_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10512));
    defparam i8970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8971_3_lut (.I0(\REG.mem_54_11 ), .I1(\REG.mem_55_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10513));
    defparam i8971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3895_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_49_9 ), .O(n4984));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3895_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8000_3_lut (.I0(n11049), .I1(n9541), .I2(rd_addr_r[3]), .I3(GND_net), 
            .O(n9542));
    defparam i8000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7999_3_lut (.I0(n12057), .I1(n12039), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9541));
    defparam i7999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3894_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_49_8 ), .O(n4983));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3894_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3893_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_49_7 ), .O(n4982));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3893_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8965_3_lut (.I0(\REG.mem_50_11 ), .I1(\REG.mem_51_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10507));
    defparam i8965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8964_3_lut (.I0(\REG.mem_48_11 ), .I1(\REG.mem_49_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10506));
    defparam i8964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8418_3_lut (.I0(\REG.mem_28_1 ), .I1(\REG.mem_29_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9960));
    defparam i8418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8419_3_lut (.I0(\REG.mem_30_1 ), .I1(\REG.mem_31_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9961));
    defparam i8419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8940_3_lut (.I0(\REG.mem_36_11 ), .I1(\REG.mem_37_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10482));
    defparam i8940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8941_3_lut (.I0(\REG.mem_38_11 ), .I1(\REG.mem_39_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10483));
    defparam i8941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8410_3_lut (.I0(\REG.mem_26_1 ), .I1(\REG.mem_27_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9952));
    defparam i8410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8409_3_lut (.I0(\REG.mem_24_1 ), .I1(\REG.mem_25_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9951));
    defparam i8409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3892_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D6_c_6), 
            .I3(\REG.mem_49_6 ), .O(n4981));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3892_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(wp_sync2_r[3]), .I1(wp_sync2_r[4]), 
            .I2(wp_sync2_r[6]), .I3(wp_sync2_r[5]), .O(wp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(537[38:77])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8935_3_lut (.I0(\REG.mem_34_11 ), .I1(\REG.mem_35_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10477));
    defparam i8935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8934_3_lut (.I0(\REG.mem_32_11 ), .I1(\REG.mem_33_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10476));
    defparam i8934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_33 (.I0(rp_sync2_r[1]), .I1(rp_sync2_r[2]), 
            .I2(rp_sync2_r[3]), .I3(n3563), .O(n3597));   // src/fifo_dc_32_lut_gen.v(286[38:77])
    defparam i1_2_lut_3_lut_4_lut_adj_33.LUT_INIT = 16'h6996;
    SB_LUT4 i3891_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D5_c_5), 
            .I3(\REG.mem_49_5 ), .O(n4980));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3891_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3890_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D4_c_4), 
            .I3(\REG.mem_49_4 ), .O(n4979));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3890_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3889_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D3_c_3), 
            .I3(\REG.mem_49_3 ), .O(n4978));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3889_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3888_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D2_c_2), 
            .I3(\REG.mem_49_2 ), .O(n4977));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3888_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8451_3_lut (.I0(\REG.mem_44_1 ), .I1(\REG.mem_45_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9993));
    defparam i8451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8452_3_lut (.I0(\REG.mem_46_1 ), .I1(\REG.mem_47_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9994));
    defparam i8452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8446_3_lut (.I0(\REG.mem_42_1 ), .I1(\REG.mem_43_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9988));
    defparam i8446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8445_3_lut (.I0(\REG.mem_40_1 ), .I1(\REG.mem_41_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9987));
    defparam i8445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3887_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D1_c_1), 
            .I3(\REG.mem_49_1 ), .O(n4976));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3887_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3886_3_lut_4_lut (.I0(n39_c), .I1(wr_addr_r[5]), .I2(FIFO_D0_c_0), 
            .I3(\REG.mem_49_0 ), .O(n4975));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3886_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8880_3_lut (.I0(n11295), .I1(n11121), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10422));
    defparam i8880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8881_3_lut (.I0(n10935), .I1(n10845), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10423));
    defparam i8881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_fifo_en_w_I_0_133_2_lut_3_lut (.I0(DEBUG_9_c), .I1(DEBUG_1_c), 
            .I2(\genblk16.rd_prev_r ), .I3(GND_net), .O(t_rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(745[41:67])
    defparam rd_fifo_en_w_I_0_133_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i8809_3_lut (.I0(n11571), .I1(n11385), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10351));
    defparam i8809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8808_3_lut (.I0(n11841), .I1(n11763), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10350));
    defparam i8808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3879_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D15_c_15), 
            .I3(\REG.mem_48_15 ), .O(n4968));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3879_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3877_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D14_c_14), 
            .I3(\REG.mem_48_14 ), .O(n4966));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3877_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3876_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D13_c_13), 
            .I3(\REG.mem_48_13 ), .O(n4965));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3876_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3875_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D12_c_12), 
            .I3(\REG.mem_48_12 ), .O(n4964));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3875_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8850_3_lut (.I0(\REG.mem_52_6 ), .I1(\REG.mem_53_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10392));
    defparam i8850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8851_3_lut (.I0(\REG.mem_54_6 ), .I1(\REG.mem_55_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10393));
    defparam i8851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8833_3_lut (.I0(\REG.mem_50_6 ), .I1(\REG.mem_51_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10375));
    defparam i8833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8832_3_lut (.I0(\REG.mem_48_6 ), .I1(\REG.mem_49_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10374));
    defparam i8832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7965_3_lut (.I0(n10959), .I1(n10899), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9507));
    defparam i7965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7966_3_lut (.I0(n10737), .I1(n10713), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n9508));
    defparam i7966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7850_4_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_r[4]), .I2(rp_sync2_r[3]), 
            .I3(n3563), .O(n9390));
    defparam i7850_4_lut_4_lut.LUT_INIT = 16'hb7de;
    SB_LUT4 i3874_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D11_c_11), 
            .I3(\REG.mem_48_11 ), .O(n4963));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3874_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut (.I0(rp_sync2_r[2]), .I1(rp_sync2_r[3]), .I2(n3563), 
            .I3(GND_net), .O(n3584));   // src/fifo_dc_32_lut_gen.v(286[38:77])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i8890_3_lut (.I0(n11193), .I1(n11043), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10432));
    defparam i8890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8889_3_lut (.I0(n11313), .I1(n11235), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n10431));
    defparam i8889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3873_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D10_c_10), 
            .I3(\REG.mem_48_10 ), .O(n4962));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3873_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_34 (.I0(rp_sync2_r[4]), .I1(rp_sync2_r[6]), 
            .I2(rp_sync2_r[5]), .I3(GND_net), .O(n3563));   // src/fifo_dc_32_lut_gen.v(286[38:77])
    defparam i1_2_lut_3_lut_adj_34.LUT_INIT = 16'h9696;
    SB_LUT4 i3872_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D9_c_9), 
            .I3(\REG.mem_48_9 ), .O(n4961));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3872_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3871_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D8_c_8), 
            .I3(\REG.mem_48_8 ), .O(n4960));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3871_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3870_3_lut_4_lut (.I0(n37_c), .I1(wr_addr_r[5]), .I2(FIFO_D7_c_7), 
            .I3(\REG.mem_48_7 ), .O(n4959));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam i3870_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i8487_3_lut (.I0(\REG.mem_60_1 ), .I1(\REG.mem_61_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10029));
    defparam i8487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8488_3_lut (.I0(\REG.mem_62_1 ), .I1(\REG.mem_63_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10030));
    defparam i8488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i59_2_lut_3_lut_4_lut (.I0(n11_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n59_adj_1060));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i59_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i8476_3_lut (.I0(\REG.mem_58_1 ), .I1(\REG.mem_59_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10018));
    defparam i8476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8475_3_lut (.I0(\REG.mem_56_1 ), .I1(\REG.mem_57_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10017));
    defparam i8475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7838_4_lut_4_lut (.I0(rd_addr_r[1]), .I1(rd_addr_r[2]), .I2(wp_sync2_r[1]), 
            .I3(wp_sync_w[2]), .O(n9378));
    defparam i7838_4_lut_4_lut.LUT_INIT = 16'hb7de;
    SB_LUT4 i1_2_lut_3_lut_adj_35 (.I0(wp_sync2_r[0]), .I1(wp_sync2_r[1]), 
            .I2(wp_sync_w[2]), .I3(GND_net), .O(wp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(537[38:77])
    defparam i1_2_lut_3_lut_adj_35.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_36 (.I0(wp_sync2_r[4]), .I1(wp_sync2_r[6]), 
            .I2(wp_sync2_r[5]), .I3(GND_net), .O(wp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(537[38:77])
    defparam i1_2_lut_3_lut_adj_36.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_37 (.I0(wp_sync2_r[2]), .I1(wp_sync2_r[3]), 
            .I2(wp_sync_w[4]), .I3(GND_net), .O(wp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(537[38:77])
    defparam i1_2_lut_3_lut_adj_37.LUT_INIT = 16'h9696;
    SB_LUT4 EnabledDecoder_2_i44_2_lut_3_lut_4_lut (.I0(n11_c), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n44_c));   // src/fifo_dc_32_lut_gen.v(887[37:55])
    defparam EnabledDecoder_2_i44_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i8796_3_lut (.I0(\REG.mem_52_13 ), .I1(\REG.mem_53_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10338));
    defparam i8796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8797_3_lut (.I0(\REG.mem_54_13 ), .I1(\REG.mem_55_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10339));
    defparam i8797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8358_3_lut (.I0(\REG.mem_28_12 ), .I1(\REG.mem_29_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9900));
    defparam i8358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8359_3_lut (.I0(\REG.mem_30_12 ), .I1(\REG.mem_31_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9901));
    defparam i8359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8335_3_lut (.I0(\REG.mem_26_12 ), .I1(\REG.mem_27_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9877));
    defparam i8335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8334_3_lut (.I0(\REG.mem_24_12 ), .I1(\REG.mem_25_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n9876));
    defparam i8334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8785_3_lut (.I0(\REG.mem_50_13 ), .I1(\REG.mem_51_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10327));
    defparam i8785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8784_3_lut (.I0(\REG.mem_48_13 ), .I1(\REG.mem_49_13 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10326));
    defparam i8784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8793_3_lut (.I0(\REG.mem_4_11 ), .I1(\REG.mem_5_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10335));
    defparam i8793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8794_3_lut (.I0(\REG.mem_6_11 ), .I1(\REG.mem_7_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10336));
    defparam i8794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8773_3_lut (.I0(\REG.mem_2_11 ), .I1(\REG.mem_3_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10315));
    defparam i8773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8772_3_lut (.I0(\REG.mem_0_11 ), .I1(\REG.mem_1_11 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n10314));
    defparam i8772_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module spi
//

module spi (SEN_c_1, DEBUG_6_c, SOUT_c, n3629, \rx_shift_reg[0] , 
            GND_net, multi_byte_spi_trans_flag_r, n9073, VCC_net, \tx_shift_reg[0] , 
            spi_start_transfer_r, n1638, spi_rx_byte_ready, n4701, \rx_shift_reg[1] , 
            n4699, rx_buf_byte, n4683, n4682, n4681, n4680, n4679, 
            n4678, n4145, \rx_shift_reg[2] , n4144, \rx_shift_reg[3] , 
            n4137, \rx_shift_reg[4] , n3626, SCK_c_0, SDAT_c_15, n4099, 
            n4081, \rx_shift_reg[5] , n4080, \rx_shift_reg[6] , n4079, 
            \rx_shift_reg[7] , tx_addr_byte, \tx_data_byte[7] , \tx_data_byte[6] , 
            \tx_data_byte[5] , \tx_data_byte[4] , \tx_data_byte[3] , \tx_data_byte[2] , 
            \tx_data_byte[1] , n2851) /* synthesis syn_module_defined=1 */ ;
    output SEN_c_1;
    input DEBUG_6_c;
    input SOUT_c;
    output n3629;
    output \rx_shift_reg[0] ;
    input GND_net;
    input multi_byte_spi_trans_flag_r;
    input n9073;
    input VCC_net;
    output \tx_shift_reg[0] ;
    input spi_start_transfer_r;
    output n1638;
    output spi_rx_byte_ready;
    input n4701;
    output \rx_shift_reg[1] ;
    input n4699;
    output [7:0]rx_buf_byte;
    input n4683;
    input n4682;
    input n4681;
    input n4680;
    input n4679;
    input n4678;
    input n4145;
    output \rx_shift_reg[2] ;
    input n4144;
    output \rx_shift_reg[3] ;
    input n4137;
    output \rx_shift_reg[4] ;
    output n3626;
    output SCK_c_0;
    output SDAT_c_15;
    input n4099;
    input n4081;
    output \rx_shift_reg[5] ;
    input n4080;
    output \rx_shift_reg[6] ;
    input n4079;
    output \rx_shift_reg[7] ;
    input [7:0]tx_addr_byte;
    input \tx_data_byte[7] ;
    input \tx_data_byte[6] ;
    input \tx_data_byte[5] ;
    input \tx_data_byte[4] ;
    input \tx_data_byte[3] ;
    input \tx_data_byte[2] ;
    input \tx_data_byte[1] ;
    output n2851;
    
    wire DEBUG_6_c /* synthesis SET_AS_NETWORK=DEBUG_6_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [2:0]n598;
    wire [3:0]state_3__N_822;
    
    wire n9321;
    wire [3:0]state;   // src/spi.v(71[11:16])
    
    wire n9331, n9476, n9332, n19, n10584, n3, n7, n3747, n9285, 
        n3_adj_1054, n21, n22, n9472, n19_adj_1055, n6394, n10579;
    wire [7:0]n1688;
    
    wire n10537, n10532, n34, n37, n9434, n3955, n12, n3683, 
        n9333, n9294;
    wire [9:0]counter;   // src/spi.v(69[11:18])
    
    wire n16, n24, n4;
    wire [7:0]n315;
    wire [7:0]multi_byte_counter;   // src/spi.v(68[11:29])
    
    wire n8736, n8735, n8734, n8733, n8732, n8731, n8730;
    wire [9:0]n45;
    
    wire n3766, n3926, n2505, n3745, n9416, n3340, n8785, n8784;
    wire [15:0]n1639;
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    
    wire n3471, n10, n14, n10_adj_1056, n14_adj_1057, n10577, n7_adj_1058, 
        n8783, n3_adj_1059, n8782, n8781, n8780, n8779, n8778, 
        n8777, n10538, n10539, n10540, n8;
    
    SB_DFF byte_recv_92_i2 (.Q(SEN_c_1), .C(DEBUG_6_c), .D(n598[1]));   // src/spi.v(88[9] 219[16])
    SB_DFFE rx_shift_reg_i0 (.Q(\rx_shift_reg[0] ), .C(DEBUG_6_c), .E(n3629), 
            .D(SOUT_c));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i0 (.Q(state[0]), .C(DEBUG_6_c), .E(n9321), .D(state_3__N_822[0]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_3_lut (.I0(state[3]), .I1(n9331), .I2(n9476), .I3(GND_net), 
            .O(n9332));
    defparam i1_3_lut.LUT_INIT = 16'h4c4c;
    SB_LUT4 i9099_2_lut (.I0(n19), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n10584));   // src/spi.v(88[9] 219[16])
    defparam i9099_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 mux_56_Mux_1_i7_4_lut (.I0(n3), .I1(n10584), .I2(state[2]), 
            .I3(state[1]), .O(n7));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i7_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_3_lut_adj_16 (.I0(n3747), .I1(state[2]), .I2(n9285), .I3(GND_net), 
            .O(n9331));
    defparam i1_3_lut_adj_16.LUT_INIT = 16'ha8a8;
    SB_LUT4 mux_56_Mux_2_i3_3_lut (.I0(multi_byte_spi_trans_flag_r), .I1(state[0]), 
            .I2(state[1]), .I3(GND_net), .O(n3_adj_1054));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i3_3_lut.LUT_INIT = 16'hc2c2;
    SB_LUT4 mux_56_Mux_2_i15_4_lut (.I0(n3_adj_1054), .I1(state[2]), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_822[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 i1_2_lut (.I0(n19), .I1(n21), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9133_4_lut (.I0(n22), .I1(n9472), .I2(n9476), .I3(state[3]), 
            .O(n19_adj_1055));
    defparam i9133_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i5312_2_lut (.I0(state[3]), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n6394));
    defparam i5312_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mux_56_Mux_3_i15_4_lut (.I0(n10579), .I1(state[1]), .I2(state[3]), 
            .I3(n1688[5]), .O(state_3__N_822[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_3_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i9062_3_lut (.I0(state[0]), .I1(state[2]), .I2(n19), .I3(GND_net), 
            .O(n10537));
    defparam i9062_3_lut.LUT_INIT = 16'h4d4d;
    SB_DFFE tx_shift_reg_i0_i0 (.Q(\tx_shift_reg[0] ), .C(DEBUG_6_c), .E(VCC_net), 
            .D(n9073));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i9049_3_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), 
            .I3(GND_net), .O(n10532));
    defparam i9049_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i65_4_lut (.I0(n6394), .I1(n10537), .I2(state[1]), .I3(state[2]), 
            .O(n34));
    defparam i65_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i66_4_lut (.I0(n10532), .I1(n1688[5]), .I2(state[1]), .I3(state[3]), 
            .O(n37));
    defparam i66_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut (.I0(state[3]), .I1(n37), .I2(n34), .I3(n9434), 
            .O(n3955));
    defparam i1_4_lut.LUT_INIT = 16'h50dc;
    SB_LUT4 i1_4_lut_adj_17 (.I0(state[3]), .I1(n1688[5]), .I2(n9434), 
            .I3(state[1]), .O(n12));   // src/spi.v(88[9] 219[16])
    defparam i1_4_lut_adj_17.LUT_INIT = 16'ha2a0;
    SB_LUT4 i9156_4_lut (.I0(n12), .I1(state[1]), .I2(n6394), .I3(state[2]), 
            .O(n3683));   // src/spi.v(88[9] 219[16])
    defparam i9156_4_lut.LUT_INIT = 16'h4454;
    SB_DFFE state_i3 (.Q(state[3]), .C(DEBUG_6_c), .E(n19_adj_1055), .D(state_3__N_822[3]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i2 (.Q(state[2]), .C(DEBUG_6_c), .E(n9333), .D(state_3__N_822[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(DEBUG_6_c), .E(n9332), .D(state_3__N_822[1]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_4_lut_adj_18 (.I0(n9294), .I1(state[3]), .I2(counter[4]), 
            .I3(state[1]), .O(n16));   // src/spi.v(88[9] 219[16])
    defparam i1_4_lut_adj_18.LUT_INIT = 16'hf5c4;
    SB_LUT4 i30_4_lut (.I0(spi_start_transfer_r), .I1(state[3]), .I2(state[1]), 
            .I3(state[0]), .O(n24));   // src/spi.v(88[9] 219[16])
    defparam i30_4_lut.LUT_INIT = 16'hcfc1;
    SB_LUT4 i1_4_lut_adj_19 (.I0(state[0]), .I1(state[3]), .I2(state[1]), 
            .I3(state[2]), .O(n4));
    defparam i1_4_lut_adj_19.LUT_INIT = 16'h2034;
    SB_LUT4 i1_3_lut_adj_20 (.I0(counter[4]), .I1(n4), .I2(n9294), .I3(GND_net), 
            .O(n1638));
    defparam i1_3_lut_adj_20.LUT_INIT = 16'h4040;
    SB_LUT4 add_794_9_lut (.I0(GND_net), .I1(multi_byte_counter[7]), .I2(n1688[5]), 
            .I3(n8736), .O(n315[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_794_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_794_8_lut (.I0(GND_net), .I1(multi_byte_counter[6]), .I2(n1688[5]), 
            .I3(n8735), .O(n315[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_794_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_794_8 (.CI(n8735), .I0(multi_byte_counter[6]), .I1(n1688[5]), 
            .CO(n8736));
    SB_LUT4 add_794_7_lut (.I0(GND_net), .I1(multi_byte_counter[5]), .I2(n1688[5]), 
            .I3(n8734), .O(n315[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_794_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_794_7 (.CI(n8734), .I0(multi_byte_counter[5]), .I1(n1688[5]), 
            .CO(n8735));
    SB_LUT4 add_794_6_lut (.I0(GND_net), .I1(multi_byte_counter[4]), .I2(n1688[5]), 
            .I3(n8733), .O(n315[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_794_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_794_6 (.CI(n8733), .I0(multi_byte_counter[4]), .I1(n1688[5]), 
            .CO(n8734));
    SB_DFF byte_recv_92_i3 (.Q(spi_rx_byte_ready), .C(DEBUG_6_c), .D(n598[2]));   // src/spi.v(88[9] 219[16])
    SB_LUT4 add_794_5_lut (.I0(GND_net), .I1(multi_byte_counter[3]), .I2(n1688[5]), 
            .I3(n8732), .O(n315[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_794_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_794_5 (.CI(n8732), .I0(multi_byte_counter[3]), .I1(n1688[5]), 
            .CO(n8733));
    SB_LUT4 add_794_4_lut (.I0(GND_net), .I1(multi_byte_counter[2]), .I2(n1688[5]), 
            .I3(n8731), .O(n315[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_794_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_794_4 (.CI(n8731), .I0(multi_byte_counter[2]), .I1(n1688[5]), 
            .CO(n8732));
    SB_LUT4 add_794_3_lut (.I0(GND_net), .I1(multi_byte_counter[1]), .I2(n1688[5]), 
            .I3(n8730), .O(n315[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_794_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_794_3 (.CI(n8730), .I0(multi_byte_counter[1]), .I1(n1688[5]), 
            .CO(n8731));
    SB_LUT4 add_794_2_lut (.I0(GND_net), .I1(multi_byte_counter[0]), .I2(n1688[5]), 
            .I3(GND_net), .O(n315[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_794_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF rx_shift_reg_i1 (.Q(\rx_shift_reg[1] ), .C(DEBUG_6_c), .D(n4701));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i1 (.Q(rx_buf_byte[1]), .C(DEBUG_6_c), .D(n4699));   // src/spi.v(76[8] 221[4])
    SB_CARRY add_794_2 (.CI(GND_net), .I0(multi_byte_counter[0]), .I1(n1688[5]), 
            .CO(n8730));
    SB_DFF Rx_Recv_Byte_i2 (.Q(rx_buf_byte[2]), .C(DEBUG_6_c), .D(n4683));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i3 (.Q(rx_buf_byte[3]), .C(DEBUG_6_c), .D(n4682));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i4 (.Q(rx_buf_byte[4]), .C(DEBUG_6_c), .D(n4681));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i5 (.Q(rx_buf_byte[5]), .C(DEBUG_6_c), .D(n4680));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i6 (.Q(rx_buf_byte[6]), .C(DEBUG_6_c), .D(n4679));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i7 (.Q(rx_buf_byte[7]), .C(DEBUG_6_c), .D(n4678));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_939__i0 (.Q(counter[0]), .C(DEBUG_6_c), .E(n3683), 
            .D(n45[0]), .R(n3955));   // src/spi.v(183[28:41])
    SB_DFFESR multi_byte_counter_i4 (.Q(multi_byte_counter[4]), .C(DEBUG_6_c), 
            .E(n3766), .D(n315[4]), .R(n3926));   // src/spi.v(76[8] 221[4])
    SB_DFFESS multi_byte_counter_i5 (.Q(multi_byte_counter[5]), .C(DEBUG_6_c), 
            .E(n3766), .D(n315[5]), .S(n3926));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i2 (.Q(\rx_shift_reg[2] ), .C(DEBUG_6_c), .D(n4145));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i2_3_lut (.I0(state[3]), .I1(n19), .I2(state[1]), .I3(GND_net), 
            .O(n9285));
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i4_4_lut (.I0(n2505), .I1(state[3]), .I2(spi_start_transfer_r), 
            .I3(state[0]), .O(n3747));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1430_2_lut (.I0(state[1]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n2505));   // src/spi.v(88[9] 219[16])
    defparam i1430_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(state[3]), .I1(n3745), .I2(n9416), .I3(n3747), 
            .O(n9321));
    defparam i2_4_lut.LUT_INIT = 16'hc400;
    SB_LUT4 i7893_2_lut (.I0(state[0]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n9434));
    defparam i7893_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mux_56_Mux_1_i15_3_lut_4_lut (.I0(state[1]), .I1(state[0]), 
            .I2(state[3]), .I3(n7), .O(state_3__N_822[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_1_i15_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i3_4_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[3]), 
            .I3(counter[1]), .O(n9294));
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i9159_3_lut (.I0(counter[4]), .I1(n9294), .I2(n3340), .I3(GND_net), 
            .O(n3629));   // src/spi.v(88[9] 219[16])
    defparam i9159_3_lut.LUT_INIT = 16'h0808;
    SB_DFF rx_shift_reg_i3 (.Q(\rx_shift_reg[3] ), .C(DEBUG_6_c), .D(n4144));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i4 (.Q(\rx_shift_reg[4] ), .C(DEBUG_6_c), .D(n4137));   // src/spi.v(76[8] 221[4])
    SB_LUT4 counter_939_add_4_11_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[9]), 
            .I3(n8785), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_939_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_939_add_4_10_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[8]), 
            .I3(n8784), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_939_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_939_add_4_10 (.CI(n8784), .I0(VCC_net), .I1(counter[8]), 
            .CO(n8785));
    SB_DFFE tx_shift_reg_i0_i14 (.Q(tx_shift_reg[14]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[14]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i13 (.Q(tx_shift_reg[13]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[13]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i12 (.Q(tx_shift_reg[12]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[12]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i11 (.Q(tx_shift_reg[11]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[11]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i10 (.Q(tx_shift_reg[10]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[10]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i9 (.Q(tx_shift_reg[9]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[9]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i8 (.Q(tx_shift_reg[8]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[8]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i7 (.Q(tx_shift_reg[7]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[7]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i6 (.Q(tx_shift_reg[6]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[6]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i5 (.Q(tx_shift_reg[5]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[5]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i4 (.Q(tx_shift_reg[4]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[4]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i3 (.Q(tx_shift_reg[3]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[3]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i2 (.Q(tx_shift_reg[2]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i1 (.Q(tx_shift_reg[1]), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[1]));   // src/spi.v(76[8] 221[4])
    SB_DFF byte_recv_92_i1 (.Q(SCK_c_0), .C(DEBUG_6_c), .D(n598[0]));   // src/spi.v(88[9] 219[16])
    SB_LUT4 i2_3_lut_adj_21 (.I0(counter[1]), .I1(counter[3]), .I2(counter[2]), 
            .I3(GND_net), .O(n3471));
    defparam i2_3_lut_adj_21.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut (.I0(counter[7]), .I1(counter[5]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // src/spi.v(141[21:41])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(counter[4]), .I1(counter[6]), .I2(counter[8]), 
            .I3(counter[9]), .O(n14));   // src/spi.v(141[21:41])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(counter[0]), .I1(n14), .I2(n10), .I3(n3471), 
            .O(n19));   // src/spi.v(141[21:41])
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_2_lut_adj_22 (.I0(multi_byte_counter[2]), .I1(multi_byte_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_1056));   // src/spi.v(208[21:52])
    defparam i2_2_lut_adj_22.LUT_INIT = 16'heeee;
    SB_LUT4 i7913_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n9476));
    defparam i7913_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i6_4_lut_adj_23 (.I0(multi_byte_counter[3]), .I1(multi_byte_counter[1]), 
            .I2(multi_byte_counter[5]), .I3(multi_byte_counter[7]), .O(n14_adj_1057));   // src/spi.v(208[21:52])
    defparam i6_4_lut_adj_23.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_24 (.I0(multi_byte_counter[0]), .I1(n14_adj_1057), 
            .I2(n10_adj_1056), .I3(multi_byte_counter[6]), .O(n1688[5]));   // src/spi.v(208[21:52])
    defparam i7_4_lut_adj_24.LUT_INIT = 16'hfffd;
    SB_LUT4 i9092_3_lut (.I0(n1688[5]), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n10577));   // src/spi.v(88[9] 219[16])
    defparam i9092_3_lut.LUT_INIT = 16'hc4c4;
    SB_DFFESR counter_939__i1 (.Q(counter[1]), .C(DEBUG_6_c), .E(n3683), 
            .D(n45[1]), .R(n3955));   // src/spi.v(183[28:41])
    SB_LUT4 mux_188_Mux_1_i7_4_lut (.I0(state[0]), .I1(state[2]), .I2(n19), 
            .I3(state[1]), .O(n7_adj_1058));   // src/spi.v(88[9] 219[16])
    defparam mux_188_Mux_1_i7_4_lut.LUT_INIT = 16'h02dd;
    SB_DFFESR counter_939__i2 (.Q(counter[2]), .C(DEBUG_6_c), .E(n3683), 
            .D(n45[2]), .R(n3955));   // src/spi.v(183[28:41])
    SB_LUT4 mux_188_Mux_1_i15_4_lut (.I0(n7_adj_1058), .I1(n10577), .I2(state[3]), 
            .I3(state[2]), .O(n598[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_188_Mux_1_i15_4_lut.LUT_INIT = 16'hfaca;
    SB_DFFESR counter_939__i3 (.Q(counter[3]), .C(DEBUG_6_c), .E(n3683), 
            .D(n45[3]), .R(n3955));   // src/spi.v(183[28:41])
    SB_LUT4 i9090_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n10579));
    defparam i9090_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFFESR counter_939__i4 (.Q(counter[4]), .C(DEBUG_6_c), .E(n3683), 
            .D(n45[4]), .R(n3955));   // src/spi.v(183[28:41])
    SB_DFFESR counter_939__i5 (.Q(counter[5]), .C(DEBUG_6_c), .E(n3683), 
            .D(n45[5]), .R(n3955));   // src/spi.v(183[28:41])
    SB_DFFESR counter_939__i6 (.Q(counter[6]), .C(DEBUG_6_c), .E(n3683), 
            .D(n45[6]), .R(n3955));   // src/spi.v(183[28:41])
    SB_DFFESR counter_939__i7 (.Q(counter[7]), .C(DEBUG_6_c), .E(n3683), 
            .D(n45[7]), .R(n3955));   // src/spi.v(183[28:41])
    SB_DFFESS counter_939__i8 (.Q(counter[8]), .C(DEBUG_6_c), .E(n3683), 
            .D(n45[8]), .S(n3955));   // src/spi.v(183[28:41])
    SB_DFFE tx_shift_reg_i0_i15 (.Q(SDAT_c_15), .C(DEBUG_6_c), .E(n3626), 
            .D(n1639[15]));   // src/spi.v(76[8] 221[4])
    SB_DFFESR counter_939__i9 (.Q(counter[9]), .C(DEBUG_6_c), .E(n3683), 
            .D(n45[9]), .R(n3955));   // src/spi.v(183[28:41])
    SB_DFFESR multi_byte_counter_i0 (.Q(multi_byte_counter[0]), .C(DEBUG_6_c), 
            .E(n3766), .D(n315[0]), .R(n3926));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_56_Mux_1_i3_3_lut_3_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(GND_net), .O(n3));
    defparam mux_56_Mux_1_i3_3_lut_3_lut.LUT_INIT = 16'h3e3e;
    SB_LUT4 counter_939_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[7]), 
            .I3(n8783), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_939_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_56_Mux_0_i3_4_lut_4_lut (.I0(multi_byte_spi_trans_flag_r), 
            .I1(state[0]), .I2(state[1]), .I3(n19), .O(n3_adj_1059));
    defparam mux_56_Mux_0_i3_4_lut_4_lut.LUT_INIT = 16'hc131;
    SB_LUT4 i43_4_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(state[1]), 
            .I3(state[0]), .O(n21));
    defparam i43_4_lut_4_lut.LUT_INIT = 16'hf01a;
    SB_LUT4 i2833_3_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(state[0]), 
            .I3(n3_adj_1059), .O(state_3__N_822[0]));
    defparam i2833_3_lut_4_lut.LUT_INIT = 16'h1f0e;
    SB_CARRY counter_939_add_4_9 (.CI(n8783), .I0(VCC_net), .I1(counter[7]), 
            .CO(n8784));
    SB_LUT4 counter_939_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[6]), 
            .I3(n8782), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_939_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_939_add_4_8 (.CI(n8782), .I0(VCC_net), .I1(counter[6]), 
            .CO(n8783));
    SB_LUT4 counter_939_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[5]), 
            .I3(n8781), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_939_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_939_add_4_7 (.CI(n8781), .I0(VCC_net), .I1(counter[5]), 
            .CO(n8782));
    SB_LUT4 counter_939_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[4]), 
            .I3(n8780), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_939_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_939_add_4_6 (.CI(n8780), .I0(VCC_net), .I1(counter[4]), 
            .CO(n8781));
    SB_LUT4 counter_939_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[3]), 
            .I3(n8779), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_939_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF Rx_Recv_Byte_i0 (.Q(rx_buf_byte[0]), .C(DEBUG_6_c), .D(n4099));   // src/spi.v(76[8] 221[4])
    SB_CARRY counter_939_add_4_5 (.CI(n8779), .I0(VCC_net), .I1(counter[3]), 
            .CO(n8780));
    SB_LUT4 counter_939_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[2]), 
            .I3(n8778), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_939_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_939_add_4_4 (.CI(n8778), .I0(VCC_net), .I1(counter[2]), 
            .CO(n8779));
    SB_LUT4 counter_939_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[1]), 
            .I3(n8777), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_939_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_939_add_4_3 (.CI(n8777), .I0(VCC_net), .I1(counter[1]), 
            .CO(n8778));
    SB_LUT4 counter_939_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_939_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF rx_shift_reg_i5 (.Q(\rx_shift_reg[5] ), .C(DEBUG_6_c), .D(n4081));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i6 (.Q(\rx_shift_reg[6] ), .C(DEBUG_6_c), .D(n4080));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i7 (.Q(\rx_shift_reg[7] ), .C(DEBUG_6_c), .D(n4079));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i6 (.Q(multi_byte_counter[6]), .C(DEBUG_6_c), 
            .E(n3766), .D(n315[6]), .R(n3926));   // src/spi.v(76[8] 221[4])
    SB_DFFESS multi_byte_counter_i7 (.Q(multi_byte_counter[7]), .C(DEBUG_6_c), 
            .E(n3766), .D(n315[7]), .S(n3926));   // src/spi.v(76[8] 221[4])
    SB_CARRY counter_939_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n8777));
    SB_DFFESR multi_byte_counter_i1 (.Q(multi_byte_counter[1]), .C(DEBUG_6_c), 
            .E(n3766), .D(n315[1]), .R(n3926));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i2 (.Q(multi_byte_counter[2]), .C(DEBUG_6_c), 
            .E(n3766), .D(n315[2]), .R(n3926));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i3 (.Q(multi_byte_counter[3]), .C(DEBUG_6_c), 
            .E(n3766), .D(n315[3]), .R(n3926));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_4_lut_adj_25 (.I0(state[1]), .I1(n10538), .I2(n9434), .I3(state[3]), 
            .O(n3766));
    defparam i1_4_lut_adj_25.LUT_INIT = 16'h0a88;
    SB_LUT4 i2921_2_lut (.I0(n3766), .I1(state[3]), .I2(GND_net), .I3(GND_net), 
            .O(n3926));   // src/spi.v(76[8] 221[4])
    defparam i2921_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_784_i15_3_lut (.I0(tx_addr_byte[6]), .I1(tx_shift_reg[13]), 
            .I2(n1638), .I3(GND_net), .O(n1639[14]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i14_3_lut (.I0(tx_addr_byte[5]), .I1(tx_shift_reg[12]), 
            .I2(n1638), .I3(GND_net), .O(n1639[13]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i13_3_lut (.I0(tx_addr_byte[4]), .I1(tx_shift_reg[11]), 
            .I2(n1638), .I3(GND_net), .O(n1639[12]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i12_3_lut (.I0(tx_addr_byte[3]), .I1(tx_shift_reg[10]), 
            .I2(n1638), .I3(GND_net), .O(n1639[11]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i11_3_lut (.I0(tx_addr_byte[2]), .I1(tx_shift_reg[9]), 
            .I2(n1638), .I3(GND_net), .O(n1639[10]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i10_3_lut (.I0(tx_addr_byte[1]), .I1(tx_shift_reg[8]), 
            .I2(n1638), .I3(GND_net), .O(n1639[9]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i9_3_lut (.I0(tx_addr_byte[0]), .I1(tx_shift_reg[7]), 
            .I2(n1638), .I3(GND_net), .O(n1639[8]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i8_3_lut (.I0(\tx_data_byte[7] ), .I1(tx_shift_reg[6]), 
            .I2(n1638), .I3(GND_net), .O(n1639[7]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i7_3_lut (.I0(\tx_data_byte[6] ), .I1(tx_shift_reg[5]), 
            .I2(n1638), .I3(GND_net), .O(n1639[6]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i6_3_lut (.I0(\tx_data_byte[5] ), .I1(tx_shift_reg[4]), 
            .I2(n1638), .I3(GND_net), .O(n1639[5]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i5_3_lut (.I0(\tx_data_byte[4] ), .I1(tx_shift_reg[3]), 
            .I2(n1638), .I3(GND_net), .O(n1639[4]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i4_3_lut (.I0(\tx_data_byte[3] ), .I1(tx_shift_reg[2]), 
            .I2(n1638), .I3(GND_net), .O(n1639[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i3_3_lut (.I0(\tx_data_byte[2] ), .I1(tx_shift_reg[1]), 
            .I2(n1638), .I3(GND_net), .O(n1639[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_784_i2_3_lut (.I0(\tx_data_byte[1] ), .I1(\tx_shift_reg[0] ), 
            .I2(n1638), .I3(GND_net), .O(n1639[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(n9285), .I1(state[0]), .I2(state[2]), 
            .I3(n3747), .O(n9333));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'hba00;
    SB_LUT4 i1_4_lut_adj_26 (.I0(counter[4]), .I1(n10539), .I2(n10540), 
            .I3(state[3]), .O(n598[0]));   // src/spi.v(88[9] 219[16])
    defparam i1_4_lut_adj_26.LUT_INIT = 16'ha088;
    SB_LUT4 i9088_4_lut (.I0(n8), .I1(state[1]), .I2(state[0]), .I3(state[2]), 
            .O(n10539));   // src/spi.v(88[9] 219[16])
    defparam i9088_4_lut.LUT_INIT = 16'hc08c;
    SB_LUT4 mux_784_i16_3_lut (.I0(tx_addr_byte[7]), .I1(tx_shift_reg[14]), 
            .I2(n1638), .I3(GND_net), .O(n1639[15]));   // src/spi.v(88[9] 219[16])
    defparam mux_784_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(counter[0]), .I1(counter[1]), .I2(counter[3]), 
            .I3(counter[2]), .O(n8));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9061_2_lut_3_lut (.I0(n19), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n10538));
    defparam i9061_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 mux_188_Mux_2_i15_4_lut_4_lut (.I0(state[0]), .I1(state[2]), 
            .I2(state[3]), .I3(state[1]), .O(n598[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_188_Mux_2_i15_4_lut_4_lut.LUT_INIT = 16'h1008;
    SB_LUT4 i2253_4_lut_4_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(state[3]), .O(n3340));   // src/spi.v(88[9] 219[16])
    defparam i2253_4_lut_4_lut_4_lut.LUT_INIT = 16'hfe75;
    SB_LUT4 i9101_2_lut_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(n8), .O(n10540));   // src/spi.v(88[9] 219[16])
    defparam i9101_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_3_lut_4_lut (.I0(state[1]), .I1(state[2]), .I2(n19), .I3(state[0]), 
            .O(n9416));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i2_2_lut_3_lut (.I0(n9285), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n3745));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i1752_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(state[3]), .O(n2851));   // src/spi.v(88[9] 219[16])
    defparam i1752_4_lut_4_lut.LUT_INIT = 16'hfdef;
    SB_LUT4 i9162_3_lut_4_lut (.I0(state[2]), .I1(state[0]), .I2(n24), 
            .I3(n16), .O(n3626));   // src/spi.v(88[9] 219[16])
    defparam i9162_3_lut_4_lut.LUT_INIT = 16'h000d;
    SB_LUT4 i7931_3_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(spi_start_transfer_r), 
            .I3(state[1]), .O(n9472));
    defparam i7931_3_lut_4_lut.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module clock
//

module clock (GND_net, VCC_net, ICE_SYSCLK_c, pll_clk_unbuf) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    input ICE_SYSCLK_c;
    output pll_clk_unbuf;
    
    
    SB_PLL40_CORE pll_config (.REFERENCECLK(ICE_SYSCLK_c), .PLLOUTGLOBAL(pll_clk_unbuf), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=14, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/top.v(222[7] 228[3])
    defparam pll_config.FEEDBACK_PATH = "SIMPLE";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll_config.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll_config.FDA_FEEDBACK = 0;
    defparam pll_config.FDA_RELATIVE = 0;
    defparam pll_config.PLLOUT_SELECT = "GENCLK";
    defparam pll_config.DIVR = 4'b0001;
    defparam pll_config.DIVF = 7'b1010010;
    defparam pll_config.DIVQ = 3'b100;
    defparam pll_config.FILTER_RANGE = 3'b001;
    defparam pll_config.ENABLE_ICEGATE = 1'b0;
    defparam pll_config.TEST_MODE = 1'b0;
    defparam pll_config.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \uart_tx(CLKS_PER_BIT=20) 
//

module \uart_tx(CLKS_PER_BIT=20)  (DEBUG_6_c, UART_TX_c, r_SM_Main, VCC_net, 
            n4974, r_Tx_Data, n4973, n4972, n4971, n4970, n4969, 
            n4967, GND_net, \r_SM_Main_2__N_728[0] , \r_SM_Main_2__N_725[1] , 
            n3151, n4091, n4090, tx_uart_active_flag, n12410, n4) /* synthesis syn_module_defined=1 */ ;
    input DEBUG_6_c;
    output UART_TX_c;
    output [2:0]r_SM_Main;
    input VCC_net;
    input n4974;
    output [7:0]r_Tx_Data;
    input n4973;
    input n4972;
    input n4971;
    input n4970;
    input n4969;
    input n4967;
    input GND_net;
    input \r_SM_Main_2__N_728[0] ;
    output \r_SM_Main_2__N_725[1] ;
    output n3151;
    input n4091;
    input n4090;
    output tx_uart_active_flag;
    input n12410;
    output n4;
    
    wire DEBUG_6_c /* synthesis SET_AS_NETWORK=DEBUG_6_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [9:0]n45;
    
    wire n1;
    wire [9:0]r_Clock_Count;   // src/uart_tx.v(32[16:29])
    
    wire n4044;
    wire [2:0]n312;
    
    wire n9466;
    wire [2:0]r_Bit_Index;   // src/uart_tx.v(33[16:27])
    
    wire n9468, n3, n2521, n5333, n3_adj_1052, n11184, n11187, 
        n8803, n8802, n8801, n8800, n8799, n8798, n8797, n8796, 
        n8795, n6582, n2520, n11067, o_Tx_Serial_N_757, n4_c, n8, 
        n7, n11064;
    
    SB_DFFESR r_Clock_Count_943__i8 (.Q(r_Clock_Count[8]), .C(DEBUG_6_c), 
            .E(n1), .D(n45[8]), .R(n4044));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_943__i7 (.Q(r_Clock_Count[7]), .C(DEBUG_6_c), 
            .E(n1), .D(n45[7]), .R(n4044));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_943__i6 (.Q(r_Clock_Count[6]), .C(DEBUG_6_c), 
            .E(n1), .D(n45[6]), .R(n4044));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_943__i5 (.Q(r_Clock_Count[5]), .C(DEBUG_6_c), 
            .E(n1), .D(n45[5]), .R(n4044));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_943__i4 (.Q(r_Clock_Count[4]), .C(DEBUG_6_c), 
            .E(n1), .D(n45[4]), .R(n4044));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_943__i3 (.Q(r_Clock_Count[3]), .C(DEBUG_6_c), 
            .E(n1), .D(n45[3]), .R(n4044));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_943__i2 (.Q(r_Clock_Count[2]), .C(DEBUG_6_c), 
            .E(n1), .D(n45[2]), .R(n4044));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_943__i1 (.Q(r_Clock_Count[1]), .C(DEBUG_6_c), 
            .E(n1), .D(n45[1]), .R(n4044));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(DEBUG_6_c), .E(n9466), 
            .D(n312[2]), .R(n9468));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFE o_Tx_Serial_44 (.Q(UART_TX_c), .C(DEBUG_6_c), .E(n1), .D(n3));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(DEBUG_6_c), .D(n2521), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Clock_Count_943__i0 (.Q(r_Clock_Count[0]), .C(DEBUG_6_c), 
            .E(n1), .D(n45[0]), .R(n4044));   // src/uart_tx.v(116[34:51])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(DEBUG_6_c), .E(VCC_net), 
            .D(n5333));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(DEBUG_6_c), .D(n4974));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(DEBUG_6_c), .D(n4973));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(DEBUG_6_c), .D(n4972));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(DEBUG_6_c), .D(n4971));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(DEBUG_6_c), .D(n4970));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(DEBUG_6_c), .D(n4969));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(DEBUG_6_c), .D(n4967));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(DEBUG_6_c), .D(n3_adj_1052), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n11184));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n11184_bdd_4_lut (.I0(n11184), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n11187));
    defparam n11184_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 r_Clock_Count_943_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n8803), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_943_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_943_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n8802), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_943_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_943_add_4_10 (.CI(n8802), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n8803));
    SB_LUT4 r_Clock_Count_943_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[7]), 
            .I3(n8801), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_943_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_943_add_4_9 (.CI(n8801), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n8802));
    SB_LUT4 r_Clock_Count_943_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[6]), 
            .I3(n8800), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_943_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_943_add_4_8 (.CI(n8800), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n8801));
    SB_LUT4 r_Clock_Count_943_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[5]), 
            .I3(n8799), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_943_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_943_add_4_7 (.CI(n8799), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n8800));
    SB_LUT4 r_Clock_Count_943_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[4]), 
            .I3(n8798), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_943_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_943_add_4_6 (.CI(n8798), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n8799));
    SB_LUT4 r_Clock_Count_943_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[3]), 
            .I3(n8797), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_943_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_943_add_4_5 (.CI(n8797), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n8798));
    SB_LUT4 r_Clock_Count_943_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[2]), 
            .I3(n8796), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_943_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_943_add_4_4 (.CI(n8796), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n8797));
    SB_LUT4 r_Clock_Count_943_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[1]), 
            .I3(n8795), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_943_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_943_add_4_3 (.CI(n8795), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n8796));
    SB_LUT4 r_Clock_Count_943_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(r_Clock_Count[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_943_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_943_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n8795));
    SB_LUT4 i1445_4_lut (.I0(\r_SM_Main_2__N_728[0] ), .I1(n6582), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_725[1] ), .O(n2520));   // src/uart_tx.v(41[7] 140[14])
    defparam i1445_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1446_3_lut (.I0(n2520), .I1(\r_SM_Main_2__N_725[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n2521));   // src/uart_tx.v(41[7] 140[14])
    defparam i1446_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i9146_2_lut_3_lut (.I0(n6582), .I1(r_SM_Main[1]), .I2(n9466), 
            .I3(GND_net), .O(n9468));   // src/uart_tx.v(41[7] 140[14])
    defparam i9146_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i4244_3_lut_4_lut (.I0(n6582), .I1(r_SM_Main[1]), .I2(r_Bit_Index[0]), 
            .I3(n9466), .O(n5333));   // src/uart_tx.v(41[7] 140[14])
    defparam i4244_3_lut_4_lut.LUT_INIT = 16'h04f0;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n6582));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1090_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n312[2]));
    defparam i1090_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_728[0] ), .O(n3151));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_725[1] ), .O(n9466));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i5796138_i1_3_lut (.I0(n11187), .I1(n11067), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_757));
    defparam i5796138_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_55_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_757), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // src/uart_tx.v(41[7] 140[14])
    defparam r_SM_Main_2__I_0_55_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n4_c));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[9]), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(GND_net), .O(n8));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[8]), .I2(r_Clock_Count[4]), 
            .I3(n4_c), .O(n7));
    defparam i1_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i5_4_lut (.I0(r_Clock_Count[5]), .I1(n7), .I2(r_Clock_Count[6]), 
            .I3(n8), .O(\r_SM_Main_2__N_725[1] ));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_9560 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n11064));
    defparam r_Bit_Index_0__bdd_4_lut_9560.LUT_INIT = 16'he4aa;
    SB_LUT4 n11064_bdd_4_lut (.I0(n11064), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n11067));
    defparam n11064_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(DEBUG_6_c), .D(n4091));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Active_46 (.Q(tx_uart_active_flag), .C(DEBUG_6_c), .D(n4090));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(DEBUG_6_c), .D(n12410));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i9107_4_lut_4_lut (.I0(\r_SM_Main_2__N_725[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_728[0] ), .O(n4));   // src/uart_tx.v(41[7] 140[14])
    defparam i9107_4_lut_4_lut.LUT_INIT = 16'h8380;
    SB_LUT4 i2032_2_lut_3_lut (.I0(\r_SM_Main_2__N_725[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_1052));   // src/uart_tx.v(41[7] 140[14])
    defparam i2032_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(DEBUG_6_c), .E(n9466), 
            .D(n312[1]), .R(n9468));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Clock_Count_943__i9 (.Q(r_Clock_Count[9]), .C(DEBUG_6_c), 
            .E(n1), .D(n45[9]), .R(n4044));   // src/uart_tx.v(116[34:51])
    SB_LUT4 i9136_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_725[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n4044));
    defparam i9136_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1083_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n312[1]));   // src/uart_tx.v(96[36:51])
    defparam i1083_2_lut.LUT_INIT = 16'h6666;
    
endmodule

// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Jun 15 2020 23:04:52

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    SOUT,
    SCK,
    FIFO_D31,
    FIFO_D20,
    FIFO_D13,
    FIFO_D1,
    FIFO_CLK,
    FIFO_BE2,
    DATA15,
    DATA4,
    DATA23,
    RST,
    FIFO_D4,
    FIFO_D14,
    UART_TX,
    DATA10,
    DATA28,
    DATA19,
    SDAT,
    FT_SIWU,
    DATA0,
    FT_WR,
    FIFO_D27,
    FIFO_D10,
    FIFO_D0,
    FIFO_BE3,
    DEBUG_0,
    FIFO_D9,
    DATA14,
    UPDATE,
    RESET,
    FIFO_D21,
    FIFO_D12,
    FIFO_BE1,
    DEBUG_6,
    DATA5,
    DATA24,
    SEN,
    FIFO_D7,
    FIFO_D15,
    ICE_CREST,
    FIFO_D23,
    DATA3,
    DATA22,
    DATA13,
    INVERT,
    FT_RD,
    FIFO_D5,
    FIFO_D24,
    FIFO_D17,
    DSR,
    DEBUG_3,
    DATA29,
    DATA18,
    ICE_SYSCLK,
    ICE_CLK,
    DATA20,
    DATA11,
    DATA1,
    VALID,
    SYNC,
    FIFO_D3,
    FIFO_D26,
    FIFO_D11,
    DEBUG_1,
    DATA8,
    DATA31,
    DATA27,
    CTS,
    FIFO_D8,
    FIFO_D18,
    DEBUG_8,
    DCD,
    DATA17,
    SLM_CLK,
    DATA6,
    DATA25,
    ICE_CDONE,
    FIFO_D6,
    FIFO_D29,
    UART_RX,
    FIFO_D22,
    FIFO_BE0,
    DEBUG_5,
    DATA12,
    DTR,
    DATA21,
    DATA2,
    FIFO_D25,
    FIFO_D2,
    FIFO_D16,
    DEBUG_2,
    DATA9,
    DATA30,
    FT_TXE,
    FR_RXF,
    FIFO_D19,
    DEBUG_9,
    DATA16,
    FT_OE,
    DATA7,
    DATA26,
    FIFO_D30,
    FIFO_D28);

    input SOUT;
    output SCK;
    input FIFO_D31;
    input FIFO_D20;
    input FIFO_D13;
    input FIFO_D1;
    input FIFO_CLK;
    input FIFO_BE2;
    output DATA15;
    output DATA4;
    output DATA23;
    output RST;
    input FIFO_D4;
    input FIFO_D14;
    output UART_TX;
    output DATA10;
    output DATA28;
    output DATA19;
    output SDAT;
    output FT_SIWU;
    output DATA0;
    output FT_WR;
    input FIFO_D27;
    input FIFO_D10;
    input FIFO_D0;
    input FIFO_BE3;
    output DEBUG_0;
    input FIFO_D9;
    output DATA14;
    output UPDATE;
    output RESET;
    input FIFO_D21;
    input FIFO_D12;
    input FIFO_BE1;
    output DEBUG_6;
    output DATA5;
    output DATA24;
    output SEN;
    input FIFO_D7;
    input FIFO_D15;
    output ICE_CREST;
    input FIFO_D23;
    output DATA3;
    output DATA22;
    output DATA13;
    output INVERT;
    output FT_RD;
    input FIFO_D5;
    input FIFO_D24;
    input FIFO_D17;
    output DSR;
    output DEBUG_3;
    output DATA29;
    output DATA18;
    input ICE_SYSCLK;
    output ICE_CLK;
    output DATA20;
    output DATA11;
    output DATA1;
    output VALID;
    output SYNC;
    input FIFO_D3;
    input FIFO_D26;
    input FIFO_D11;
    output DEBUG_1;
    output DATA8;
    output DATA31;
    output DATA27;
    output CTS;
    input FIFO_D8;
    input FIFO_D18;
    output DEBUG_8;
    output DCD;
    output DATA17;
    output SLM_CLK;
    output DATA6;
    output DATA25;
    output ICE_CDONE;
    input FIFO_D6;
    input FIFO_D29;
    input UART_RX;
    input FIFO_D22;
    input FIFO_BE0;
    output DEBUG_5;
    output DATA12;
    output DTR;
    output DATA21;
    output DATA2;
    input FIFO_D25;
    input FIFO_D2;
    input FIFO_D16;
    output DEBUG_2;
    output DATA9;
    output DATA30;
    input FT_TXE;
    input FR_RXF;
    input FIFO_D19;
    output DEBUG_9;
    output DATA16;
    output FT_OE;
    output DATA7;
    output DATA26;
    input FIFO_D30;
    input FIFO_D28;

    wire N__98338;
    wire N__98337;
    wire N__98336;
    wire N__98327;
    wire N__98326;
    wire N__98325;
    wire N__98318;
    wire N__98317;
    wire N__98316;
    wire N__98309;
    wire N__98308;
    wire N__98307;
    wire N__98300;
    wire N__98299;
    wire N__98298;
    wire N__98291;
    wire N__98290;
    wire N__98289;
    wire N__98282;
    wire N__98281;
    wire N__98280;
    wire N__98273;
    wire N__98272;
    wire N__98271;
    wire N__98264;
    wire N__98263;
    wire N__98262;
    wire N__98255;
    wire N__98254;
    wire N__98253;
    wire N__98246;
    wire N__98245;
    wire N__98244;
    wire N__98237;
    wire N__98236;
    wire N__98235;
    wire N__98228;
    wire N__98227;
    wire N__98226;
    wire N__98219;
    wire N__98218;
    wire N__98217;
    wire N__98210;
    wire N__98209;
    wire N__98208;
    wire N__98201;
    wire N__98200;
    wire N__98199;
    wire N__98192;
    wire N__98191;
    wire N__98190;
    wire N__98183;
    wire N__98182;
    wire N__98181;
    wire N__98174;
    wire N__98173;
    wire N__98172;
    wire N__98165;
    wire N__98164;
    wire N__98163;
    wire N__98156;
    wire N__98155;
    wire N__98154;
    wire N__98147;
    wire N__98146;
    wire N__98145;
    wire N__98138;
    wire N__98137;
    wire N__98136;
    wire N__98129;
    wire N__98128;
    wire N__98127;
    wire N__98120;
    wire N__98119;
    wire N__98118;
    wire N__98111;
    wire N__98110;
    wire N__98109;
    wire N__98102;
    wire N__98101;
    wire N__98100;
    wire N__98093;
    wire N__98092;
    wire N__98091;
    wire N__98084;
    wire N__98083;
    wire N__98082;
    wire N__98075;
    wire N__98074;
    wire N__98073;
    wire N__98066;
    wire N__98065;
    wire N__98064;
    wire N__98057;
    wire N__98056;
    wire N__98055;
    wire N__98048;
    wire N__98047;
    wire N__98046;
    wire N__98039;
    wire N__98038;
    wire N__98037;
    wire N__98030;
    wire N__98029;
    wire N__98028;
    wire N__98021;
    wire N__98020;
    wire N__98019;
    wire N__98012;
    wire N__98011;
    wire N__98010;
    wire N__98003;
    wire N__98002;
    wire N__98001;
    wire N__97994;
    wire N__97993;
    wire N__97992;
    wire N__97985;
    wire N__97984;
    wire N__97983;
    wire N__97976;
    wire N__97975;
    wire N__97974;
    wire N__97967;
    wire N__97966;
    wire N__97965;
    wire N__97958;
    wire N__97957;
    wire N__97956;
    wire N__97949;
    wire N__97948;
    wire N__97947;
    wire N__97940;
    wire N__97939;
    wire N__97938;
    wire N__97931;
    wire N__97930;
    wire N__97929;
    wire N__97922;
    wire N__97921;
    wire N__97920;
    wire N__97913;
    wire N__97912;
    wire N__97911;
    wire N__97904;
    wire N__97903;
    wire N__97902;
    wire N__97895;
    wire N__97894;
    wire N__97893;
    wire N__97886;
    wire N__97885;
    wire N__97884;
    wire N__97877;
    wire N__97876;
    wire N__97875;
    wire N__97868;
    wire N__97867;
    wire N__97866;
    wire N__97859;
    wire N__97858;
    wire N__97857;
    wire N__97850;
    wire N__97849;
    wire N__97848;
    wire N__97841;
    wire N__97840;
    wire N__97839;
    wire N__97832;
    wire N__97831;
    wire N__97830;
    wire N__97823;
    wire N__97822;
    wire N__97821;
    wire N__97814;
    wire N__97813;
    wire N__97812;
    wire N__97805;
    wire N__97804;
    wire N__97803;
    wire N__97796;
    wire N__97795;
    wire N__97794;
    wire N__97787;
    wire N__97786;
    wire N__97785;
    wire N__97778;
    wire N__97777;
    wire N__97776;
    wire N__97769;
    wire N__97768;
    wire N__97767;
    wire N__97760;
    wire N__97759;
    wire N__97758;
    wire N__97751;
    wire N__97750;
    wire N__97749;
    wire N__97742;
    wire N__97741;
    wire N__97740;
    wire N__97733;
    wire N__97732;
    wire N__97731;
    wire N__97724;
    wire N__97723;
    wire N__97722;
    wire N__97715;
    wire N__97714;
    wire N__97713;
    wire N__97706;
    wire N__97705;
    wire N__97704;
    wire N__97697;
    wire N__97696;
    wire N__97695;
    wire N__97688;
    wire N__97687;
    wire N__97686;
    wire N__97679;
    wire N__97678;
    wire N__97677;
    wire N__97670;
    wire N__97669;
    wire N__97668;
    wire N__97661;
    wire N__97660;
    wire N__97659;
    wire N__97652;
    wire N__97651;
    wire N__97650;
    wire N__97643;
    wire N__97642;
    wire N__97641;
    wire N__97634;
    wire N__97633;
    wire N__97632;
    wire N__97625;
    wire N__97624;
    wire N__97623;
    wire N__97616;
    wire N__97615;
    wire N__97614;
    wire N__97607;
    wire N__97606;
    wire N__97605;
    wire N__97598;
    wire N__97597;
    wire N__97596;
    wire N__97579;
    wire N__97578;
    wire N__97575;
    wire N__97572;
    wire N__97567;
    wire N__97564;
    wire N__97563;
    wire N__97560;
    wire N__97557;
    wire N__97552;
    wire N__97549;
    wire N__97548;
    wire N__97545;
    wire N__97542;
    wire N__97537;
    wire N__97534;
    wire N__97531;
    wire N__97530;
    wire N__97527;
    wire N__97524;
    wire N__97519;
    wire N__97516;
    wire N__97515;
    wire N__97512;
    wire N__97509;
    wire N__97504;
    wire N__97501;
    wire N__97500;
    wire N__97497;
    wire N__97494;
    wire N__97489;
    wire N__97486;
    wire N__97485;
    wire N__97482;
    wire N__97479;
    wire N__97474;
    wire N__97471;
    wire N__97468;
    wire N__97467;
    wire N__97464;
    wire N__97461;
    wire N__97456;
    wire N__97453;
    wire N__97452;
    wire N__97451;
    wire N__97450;
    wire N__97449;
    wire N__97448;
    wire N__97447;
    wire N__97446;
    wire N__97445;
    wire N__97444;
    wire N__97443;
    wire N__97442;
    wire N__97441;
    wire N__97440;
    wire N__97439;
    wire N__97438;
    wire N__97437;
    wire N__97436;
    wire N__97435;
    wire N__97434;
    wire N__97433;
    wire N__97432;
    wire N__97431;
    wire N__97430;
    wire N__97429;
    wire N__97428;
    wire N__97427;
    wire N__97426;
    wire N__97425;
    wire N__97424;
    wire N__97423;
    wire N__97422;
    wire N__97421;
    wire N__97420;
    wire N__97419;
    wire N__97418;
    wire N__97417;
    wire N__97414;
    wire N__97413;
    wire N__97412;
    wire N__97411;
    wire N__97410;
    wire N__97409;
    wire N__97408;
    wire N__97407;
    wire N__97406;
    wire N__97405;
    wire N__97404;
    wire N__97403;
    wire N__97402;
    wire N__97401;
    wire N__97400;
    wire N__97399;
    wire N__97398;
    wire N__97397;
    wire N__97396;
    wire N__97395;
    wire N__97394;
    wire N__97393;
    wire N__97392;
    wire N__97391;
    wire N__97390;
    wire N__97389;
    wire N__97388;
    wire N__97387;
    wire N__97386;
    wire N__97385;
    wire N__97384;
    wire N__97383;
    wire N__97382;
    wire N__97381;
    wire N__97380;
    wire N__97379;
    wire N__97378;
    wire N__97377;
    wire N__97376;
    wire N__97375;
    wire N__97374;
    wire N__97373;
    wire N__97372;
    wire N__97371;
    wire N__97370;
    wire N__97369;
    wire N__97368;
    wire N__97367;
    wire N__97366;
    wire N__97365;
    wire N__97364;
    wire N__97363;
    wire N__97362;
    wire N__97361;
    wire N__97360;
    wire N__97359;
    wire N__97358;
    wire N__97357;
    wire N__97356;
    wire N__97355;
    wire N__97354;
    wire N__97353;
    wire N__97352;
    wire N__97351;
    wire N__97350;
    wire N__97349;
    wire N__97348;
    wire N__97347;
    wire N__97346;
    wire N__97345;
    wire N__97344;
    wire N__97343;
    wire N__97342;
    wire N__97123;
    wire N__97120;
    wire N__97117;
    wire N__97114;
    wire N__97111;
    wire N__97110;
    wire N__97107;
    wire N__97104;
    wire N__97099;
    wire N__97098;
    wire N__97095;
    wire N__97092;
    wire N__97087;
    wire N__97084;
    wire N__97081;
    wire N__97078;
    wire N__97077;
    wire N__97074;
    wire N__97071;
    wire N__97066;
    wire N__97063;
    wire N__97060;
    wire N__97059;
    wire N__97056;
    wire N__97055;
    wire N__97054;
    wire N__97053;
    wire N__97050;
    wire N__97049;
    wire N__97048;
    wire N__97047;
    wire N__97046;
    wire N__97045;
    wire N__97042;
    wire N__97041;
    wire N__97040;
    wire N__97039;
    wire N__97038;
    wire N__97037;
    wire N__97036;
    wire N__97035;
    wire N__97034;
    wire N__97031;
    wire N__97026;
    wire N__97025;
    wire N__97024;
    wire N__97023;
    wire N__97022;
    wire N__97021;
    wire N__97018;
    wire N__97013;
    wire N__97010;
    wire N__97005;
    wire N__97002;
    wire N__96991;
    wire N__96990;
    wire N__96989;
    wire N__96988;
    wire N__96985;
    wire N__96982;
    wire N__96981;
    wire N__96980;
    wire N__96977;
    wire N__96974;
    wire N__96971;
    wire N__96964;
    wire N__96959;
    wire N__96954;
    wire N__96949;
    wire N__96944;
    wire N__96943;
    wire N__96942;
    wire N__96941;
    wire N__96938;
    wire N__96935;
    wire N__96934;
    wire N__96931;
    wire N__96928;
    wire N__96925;
    wire N__96920;
    wire N__96917;
    wire N__96910;
    wire N__96905;
    wire N__96900;
    wire N__96895;
    wire N__96892;
    wire N__96889;
    wire N__96886;
    wire N__96883;
    wire N__96880;
    wire N__96877;
    wire N__96874;
    wire N__96871;
    wire N__96868;
    wire N__96863;
    wire N__96860;
    wire N__96857;
    wire N__96852;
    wire N__96849;
    wire N__96842;
    wire N__96837;
    wire N__96830;
    wire N__96817;
    wire N__96816;
    wire N__96815;
    wire N__96814;
    wire N__96813;
    wire N__96812;
    wire N__96811;
    wire N__96808;
    wire N__96807;
    wire N__96806;
    wire N__96801;
    wire N__96794;
    wire N__96791;
    wire N__96788;
    wire N__96785;
    wire N__96784;
    wire N__96783;
    wire N__96782;
    wire N__96779;
    wire N__96778;
    wire N__96777;
    wire N__96776;
    wire N__96775;
    wire N__96774;
    wire N__96773;
    wire N__96772;
    wire N__96771;
    wire N__96770;
    wire N__96769;
    wire N__96764;
    wire N__96757;
    wire N__96754;
    wire N__96751;
    wire N__96750;
    wire N__96747;
    wire N__96744;
    wire N__96741;
    wire N__96740;
    wire N__96739;
    wire N__96738;
    wire N__96737;
    wire N__96736;
    wire N__96735;
    wire N__96734;
    wire N__96733;
    wire N__96732;
    wire N__96731;
    wire N__96730;
    wire N__96729;
    wire N__96728;
    wire N__96727;
    wire N__96724;
    wire N__96721;
    wire N__96718;
    wire N__96713;
    wire N__96712;
    wire N__96711;
    wire N__96710;
    wire N__96709;
    wire N__96706;
    wire N__96703;
    wire N__96700;
    wire N__96699;
    wire N__96698;
    wire N__96697;
    wire N__96696;
    wire N__96695;
    wire N__96694;
    wire N__96691;
    wire N__96682;
    wire N__96679;
    wire N__96676;
    wire N__96671;
    wire N__96666;
    wire N__96665;
    wire N__96664;
    wire N__96661;
    wire N__96654;
    wire N__96651;
    wire N__96646;
    wire N__96643;
    wire N__96640;
    wire N__96639;
    wire N__96638;
    wire N__96637;
    wire N__96636;
    wire N__96635;
    wire N__96632;
    wire N__96629;
    wire N__96626;
    wire N__96623;
    wire N__96616;
    wire N__96607;
    wire N__96604;
    wire N__96599;
    wire N__96588;
    wire N__96585;
    wire N__96584;
    wire N__96583;
    wire N__96582;
    wire N__96581;
    wire N__96580;
    wire N__96577;
    wire N__96576;
    wire N__96575;
    wire N__96574;
    wire N__96573;
    wire N__96568;
    wire N__96561;
    wire N__96558;
    wire N__96555;
    wire N__96548;
    wire N__96541;
    wire N__96538;
    wire N__96529;
    wire N__96528;
    wire N__96525;
    wire N__96520;
    wire N__96513;
    wire N__96504;
    wire N__96493;
    wire N__96490;
    wire N__96485;
    wire N__96480;
    wire N__96477;
    wire N__96472;
    wire N__96461;
    wire N__96458;
    wire N__96447;
    wire N__96430;
    wire N__96429;
    wire N__96426;
    wire N__96423;
    wire N__96420;
    wire N__96415;
    wire N__96412;
    wire N__96409;
    wire N__96408;
    wire N__96405;
    wire N__96402;
    wire N__96399;
    wire N__96396;
    wire N__96391;
    wire N__96390;
    wire N__96389;
    wire N__96388;
    wire N__96387;
    wire N__96386;
    wire N__96383;
    wire N__96382;
    wire N__96371;
    wire N__96370;
    wire N__96369;
    wire N__96368;
    wire N__96367;
    wire N__96366;
    wire N__96365;
    wire N__96362;
    wire N__96359;
    wire N__96358;
    wire N__96357;
    wire N__96356;
    wire N__96355;
    wire N__96354;
    wire N__96353;
    wire N__96352;
    wire N__96351;
    wire N__96350;
    wire N__96349;
    wire N__96346;
    wire N__96345;
    wire N__96344;
    wire N__96343;
    wire N__96342;
    wire N__96341;
    wire N__96340;
    wire N__96337;
    wire N__96328;
    wire N__96325;
    wire N__96324;
    wire N__96323;
    wire N__96322;
    wire N__96321;
    wire N__96316;
    wire N__96315;
    wire N__96314;
    wire N__96313;
    wire N__96312;
    wire N__96299;
    wire N__96296;
    wire N__96289;
    wire N__96286;
    wire N__96281;
    wire N__96276;
    wire N__96273;
    wire N__96270;
    wire N__96269;
    wire N__96264;
    wire N__96261;
    wire N__96260;
    wire N__96257;
    wire N__96252;
    wire N__96251;
    wire N__96248;
    wire N__96247;
    wire N__96246;
    wire N__96245;
    wire N__96244;
    wire N__96243;
    wire N__96240;
    wire N__96237;
    wire N__96232;
    wire N__96231;
    wire N__96230;
    wire N__96229;
    wire N__96228;
    wire N__96227;
    wire N__96226;
    wire N__96225;
    wire N__96222;
    wire N__96215;
    wire N__96210;
    wire N__96209;
    wire N__96206;
    wire N__96199;
    wire N__96194;
    wire N__96193;
    wire N__96192;
    wire N__96191;
    wire N__96190;
    wire N__96189;
    wire N__96186;
    wire N__96183;
    wire N__96180;
    wire N__96177;
    wire N__96174;
    wire N__96163;
    wire N__96158;
    wire N__96157;
    wire N__96156;
    wire N__96155;
    wire N__96154;
    wire N__96153;
    wire N__96152;
    wire N__96149;
    wire N__96144;
    wire N__96141;
    wire N__96132;
    wire N__96125;
    wire N__96122;
    wire N__96115;
    wire N__96106;
    wire N__96103;
    wire N__96100;
    wire N__96089;
    wire N__96086;
    wire N__96083;
    wire N__96072;
    wire N__96067;
    wire N__96064;
    wire N__96053;
    wire N__96048;
    wire N__96045;
    wire N__96040;
    wire N__96037;
    wire N__96032;
    wire N__96029;
    wire N__96022;
    wire N__96013;
    wire N__96012;
    wire N__96011;
    wire N__96010;
    wire N__96009;
    wire N__96008;
    wire N__96007;
    wire N__96006;
    wire N__96005;
    wire N__96004;
    wire N__96003;
    wire N__96000;
    wire N__95999;
    wire N__95998;
    wire N__95997;
    wire N__95994;
    wire N__95991;
    wire N__95990;
    wire N__95989;
    wire N__95986;
    wire N__95985;
    wire N__95984;
    wire N__95983;
    wire N__95982;
    wire N__95981;
    wire N__95980;
    wire N__95979;
    wire N__95978;
    wire N__95973;
    wire N__95970;
    wire N__95967;
    wire N__95962;
    wire N__95959;
    wire N__95956;
    wire N__95955;
    wire N__95950;
    wire N__95947;
    wire N__95944;
    wire N__95941;
    wire N__95938;
    wire N__95937;
    wire N__95934;
    wire N__95931;
    wire N__95930;
    wire N__95925;
    wire N__95922;
    wire N__95915;
    wire N__95910;
    wire N__95907;
    wire N__95902;
    wire N__95899;
    wire N__95894;
    wire N__95893;
    wire N__95892;
    wire N__95891;
    wire N__95890;
    wire N__95887;
    wire N__95884;
    wire N__95881;
    wire N__95876;
    wire N__95873;
    wire N__95870;
    wire N__95867;
    wire N__95864;
    wire N__95861;
    wire N__95858;
    wire N__95851;
    wire N__95844;
    wire N__95841;
    wire N__95836;
    wire N__95833;
    wire N__95830;
    wire N__95827;
    wire N__95824;
    wire N__95819;
    wire N__95810;
    wire N__95803;
    wire N__95798;
    wire N__95779;
    wire N__95776;
    wire N__95775;
    wire N__95774;
    wire N__95773;
    wire N__95772;
    wire N__95771;
    wire N__95770;
    wire N__95763;
    wire N__95762;
    wire N__95761;
    wire N__95760;
    wire N__95759;
    wire N__95756;
    wire N__95753;
    wire N__95752;
    wire N__95751;
    wire N__95750;
    wire N__95749;
    wire N__95748;
    wire N__95747;
    wire N__95746;
    wire N__95745;
    wire N__95744;
    wire N__95743;
    wire N__95742;
    wire N__95741;
    wire N__95740;
    wire N__95737;
    wire N__95736;
    wire N__95735;
    wire N__95732;
    wire N__95731;
    wire N__95730;
    wire N__95729;
    wire N__95728;
    wire N__95727;
    wire N__95726;
    wire N__95725;
    wire N__95724;
    wire N__95723;
    wire N__95722;
    wire N__95721;
    wire N__95720;
    wire N__95719;
    wire N__95718;
    wire N__95717;
    wire N__95714;
    wire N__95709;
    wire N__95708;
    wire N__95707;
    wire N__95706;
    wire N__95705;
    wire N__95704;
    wire N__95703;
    wire N__95702;
    wire N__95701;
    wire N__95700;
    wire N__95699;
    wire N__95698;
    wire N__95695;
    wire N__95692;
    wire N__95691;
    wire N__95690;
    wire N__95689;
    wire N__95688;
    wire N__95687;
    wire N__95686;
    wire N__95685;
    wire N__95684;
    wire N__95683;
    wire N__95682;
    wire N__95677;
    wire N__95672;
    wire N__95669;
    wire N__95658;
    wire N__95651;
    wire N__95650;
    wire N__95645;
    wire N__95644;
    wire N__95643;
    wire N__95642;
    wire N__95635;
    wire N__95634;
    wire N__95633;
    wire N__95632;
    wire N__95631;
    wire N__95630;
    wire N__95629;
    wire N__95628;
    wire N__95627;
    wire N__95626;
    wire N__95625;
    wire N__95624;
    wire N__95623;
    wire N__95622;
    wire N__95621;
    wire N__95620;
    wire N__95619;
    wire N__95618;
    wire N__95617;
    wire N__95616;
    wire N__95613;
    wire N__95608;
    wire N__95595;
    wire N__95594;
    wire N__95591;
    wire N__95588;
    wire N__95585;
    wire N__95584;
    wire N__95583;
    wire N__95582;
    wire N__95579;
    wire N__95572;
    wire N__95567;
    wire N__95562;
    wire N__95559;
    wire N__95556;
    wire N__95555;
    wire N__95554;
    wire N__95553;
    wire N__95550;
    wire N__95549;
    wire N__95548;
    wire N__95547;
    wire N__95546;
    wire N__95545;
    wire N__95542;
    wire N__95541;
    wire N__95540;
    wire N__95539;
    wire N__95538;
    wire N__95537;
    wire N__95536;
    wire N__95535;
    wire N__95534;
    wire N__95533;
    wire N__95532;
    wire N__95531;
    wire N__95530;
    wire N__95529;
    wire N__95528;
    wire N__95517;
    wire N__95504;
    wire N__95503;
    wire N__95502;
    wire N__95501;
    wire N__95498;
    wire N__95497;
    wire N__95496;
    wire N__95495;
    wire N__95494;
    wire N__95493;
    wire N__95492;
    wire N__95481;
    wire N__95478;
    wire N__95475;
    wire N__95470;
    wire N__95467;
    wire N__95466;
    wire N__95465;
    wire N__95464;
    wire N__95463;
    wire N__95462;
    wire N__95461;
    wire N__95460;
    wire N__95459;
    wire N__95458;
    wire N__95457;
    wire N__95456;
    wire N__95453;
    wire N__95452;
    wire N__95451;
    wire N__95450;
    wire N__95449;
    wire N__95448;
    wire N__95447;
    wire N__95446;
    wire N__95445;
    wire N__95444;
    wire N__95443;
    wire N__95442;
    wire N__95439;
    wire N__95436;
    wire N__95431;
    wire N__95428;
    wire N__95427;
    wire N__95426;
    wire N__95425;
    wire N__95424;
    wire N__95423;
    wire N__95422;
    wire N__95421;
    wire N__95420;
    wire N__95419;
    wire N__95418;
    wire N__95417;
    wire N__95416;
    wire N__95415;
    wire N__95414;
    wire N__95413;
    wire N__95412;
    wire N__95411;
    wire N__95410;
    wire N__95409;
    wire N__95408;
    wire N__95407;
    wire N__95404;
    wire N__95403;
    wire N__95402;
    wire N__95401;
    wire N__95400;
    wire N__95399;
    wire N__95398;
    wire N__95397;
    wire N__95396;
    wire N__95395;
    wire N__95394;
    wire N__95393;
    wire N__95392;
    wire N__95391;
    wire N__95390;
    wire N__95389;
    wire N__95388;
    wire N__95387;
    wire N__95386;
    wire N__95385;
    wire N__95384;
    wire N__95383;
    wire N__95382;
    wire N__95381;
    wire N__95380;
    wire N__95379;
    wire N__95378;
    wire N__95377;
    wire N__95376;
    wire N__95375;
    wire N__95374;
    wire N__95373;
    wire N__95372;
    wire N__95371;
    wire N__95370;
    wire N__95369;
    wire N__95368;
    wire N__95367;
    wire N__95364;
    wire N__95359;
    wire N__95356;
    wire N__95349;
    wire N__95348;
    wire N__95347;
    wire N__95346;
    wire N__95345;
    wire N__95344;
    wire N__95343;
    wire N__95342;
    wire N__95339;
    wire N__95338;
    wire N__95337;
    wire N__95336;
    wire N__95335;
    wire N__95334;
    wire N__95333;
    wire N__95330;
    wire N__95327;
    wire N__95326;
    wire N__95325;
    wire N__95324;
    wire N__95323;
    wire N__95322;
    wire N__95321;
    wire N__95320;
    wire N__95319;
    wire N__95318;
    wire N__95317;
    wire N__95316;
    wire N__95315;
    wire N__95314;
    wire N__95305;
    wire N__95300;
    wire N__95299;
    wire N__95298;
    wire N__95295;
    wire N__95294;
    wire N__95291;
    wire N__95290;
    wire N__95289;
    wire N__95288;
    wire N__95287;
    wire N__95286;
    wire N__95285;
    wire N__95284;
    wire N__95283;
    wire N__95276;
    wire N__95273;
    wire N__95262;
    wire N__95259;
    wire N__95254;
    wire N__95249;
    wire N__95238;
    wire N__95225;
    wire N__95224;
    wire N__95223;
    wire N__95222;
    wire N__95221;
    wire N__95220;
    wire N__95219;
    wire N__95218;
    wire N__95211;
    wire N__95206;
    wire N__95197;
    wire N__95186;
    wire N__95183;
    wire N__95178;
    wire N__95177;
    wire N__95176;
    wire N__95175;
    wire N__95174;
    wire N__95173;
    wire N__95166;
    wire N__95157;
    wire N__95156;
    wire N__95155;
    wire N__95154;
    wire N__95153;
    wire N__95152;
    wire N__95151;
    wire N__95150;
    wire N__95149;
    wire N__95148;
    wire N__95147;
    wire N__95146;
    wire N__95139;
    wire N__95132;
    wire N__95127;
    wire N__95122;
    wire N__95119;
    wire N__95106;
    wire N__95105;
    wire N__95104;
    wire N__95103;
    wire N__95102;
    wire N__95101;
    wire N__95100;
    wire N__95099;
    wire N__95098;
    wire N__95097;
    wire N__95096;
    wire N__95095;
    wire N__95094;
    wire N__95093;
    wire N__95092;
    wire N__95091;
    wire N__95090;
    wire N__95089;
    wire N__95088;
    wire N__95087;
    wire N__95084;
    wire N__95081;
    wire N__95080;
    wire N__95079;
    wire N__95078;
    wire N__95077;
    wire N__95076;
    wire N__95075;
    wire N__95070;
    wire N__95067;
    wire N__95058;
    wire N__95055;
    wire N__95054;
    wire N__95053;
    wire N__95052;
    wire N__95051;
    wire N__95050;
    wire N__95049;
    wire N__95048;
    wire N__95039;
    wire N__95030;
    wire N__95019;
    wire N__95010;
    wire N__95009;
    wire N__95008;
    wire N__95007;
    wire N__95006;
    wire N__95005;
    wire N__95002;
    wire N__94993;
    wire N__94990;
    wire N__94987;
    wire N__94984;
    wire N__94981;
    wire N__94980;
    wire N__94979;
    wire N__94978;
    wire N__94975;
    wire N__94974;
    wire N__94973;
    wire N__94972;
    wire N__94971;
    wire N__94970;
    wire N__94967;
    wire N__94964;
    wire N__94957;
    wire N__94944;
    wire N__94931;
    wire N__94920;
    wire N__94915;
    wire N__94904;
    wire N__94899;
    wire N__94894;
    wire N__94889;
    wire N__94878;
    wire N__94877;
    wire N__94876;
    wire N__94875;
    wire N__94874;
    wire N__94871;
    wire N__94868;
    wire N__94863;
    wire N__94858;
    wire N__94849;
    wire N__94846;
    wire N__94835;
    wire N__94832;
    wire N__94831;
    wire N__94830;
    wire N__94829;
    wire N__94828;
    wire N__94827;
    wire N__94826;
    wire N__94825;
    wire N__94824;
    wire N__94823;
    wire N__94822;
    wire N__94819;
    wire N__94810;
    wire N__94805;
    wire N__94794;
    wire N__94785;
    wire N__94780;
    wire N__94777;
    wire N__94776;
    wire N__94773;
    wire N__94772;
    wire N__94771;
    wire N__94770;
    wire N__94769;
    wire N__94768;
    wire N__94767;
    wire N__94766;
    wire N__94765;
    wire N__94764;
    wire N__94763;
    wire N__94760;
    wire N__94757;
    wire N__94752;
    wire N__94743;
    wire N__94736;
    wire N__94723;
    wire N__94720;
    wire N__94717;
    wire N__94712;
    wire N__94701;
    wire N__94692;
    wire N__94687;
    wire N__94686;
    wire N__94685;
    wire N__94682;
    wire N__94681;
    wire N__94678;
    wire N__94675;
    wire N__94672;
    wire N__94671;
    wire N__94670;
    wire N__94669;
    wire N__94668;
    wire N__94667;
    wire N__94666;
    wire N__94665;
    wire N__94664;
    wire N__94663;
    wire N__94662;
    wire N__94661;
    wire N__94660;
    wire N__94657;
    wire N__94654;
    wire N__94651;
    wire N__94648;
    wire N__94645;
    wire N__94636;
    wire N__94633;
    wire N__94624;
    wire N__94613;
    wire N__94610;
    wire N__94605;
    wire N__94604;
    wire N__94603;
    wire N__94602;
    wire N__94601;
    wire N__94600;
    wire N__94599;
    wire N__94598;
    wire N__94597;
    wire N__94596;
    wire N__94595;
    wire N__94594;
    wire N__94593;
    wire N__94592;
    wire N__94591;
    wire N__94590;
    wire N__94585;
    wire N__94584;
    wire N__94583;
    wire N__94582;
    wire N__94581;
    wire N__94580;
    wire N__94579;
    wire N__94578;
    wire N__94577;
    wire N__94574;
    wire N__94565;
    wire N__94556;
    wire N__94553;
    wire N__94542;
    wire N__94531;
    wire N__94524;
    wire N__94521;
    wire N__94516;
    wire N__94513;
    wire N__94510;
    wire N__94505;
    wire N__94496;
    wire N__94493;
    wire N__94486;
    wire N__94485;
    wire N__94484;
    wire N__94483;
    wire N__94482;
    wire N__94481;
    wire N__94480;
    wire N__94477;
    wire N__94474;
    wire N__94473;
    wire N__94472;
    wire N__94471;
    wire N__94464;
    wire N__94459;
    wire N__94458;
    wire N__94457;
    wire N__94456;
    wire N__94441;
    wire N__94438;
    wire N__94433;
    wire N__94426;
    wire N__94411;
    wire N__94406;
    wire N__94399;
    wire N__94396;
    wire N__94393;
    wire N__94390;
    wire N__94387;
    wire N__94376;
    wire N__94369;
    wire N__94364;
    wire N__94359;
    wire N__94354;
    wire N__94351;
    wire N__94344;
    wire N__94337;
    wire N__94330;
    wire N__94329;
    wire N__94328;
    wire N__94325;
    wire N__94318;
    wire N__94315;
    wire N__94308;
    wire N__94297;
    wire N__94296;
    wire N__94279;
    wire N__94270;
    wire N__94259;
    wire N__94252;
    wire N__94245;
    wire N__94244;
    wire N__94243;
    wire N__94242;
    wire N__94241;
    wire N__94240;
    wire N__94239;
    wire N__94238;
    wire N__94237;
    wire N__94236;
    wire N__94235;
    wire N__94234;
    wire N__94233;
    wire N__94224;
    wire N__94223;
    wire N__94222;
    wire N__94221;
    wire N__94212;
    wire N__94203;
    wire N__94192;
    wire N__94187;
    wire N__94182;
    wire N__94181;
    wire N__94180;
    wire N__94179;
    wire N__94178;
    wire N__94177;
    wire N__94176;
    wire N__94173;
    wire N__94172;
    wire N__94171;
    wire N__94170;
    wire N__94169;
    wire N__94168;
    wire N__94163;
    wire N__94162;
    wire N__94161;
    wire N__94160;
    wire N__94157;
    wire N__94154;
    wire N__94151;
    wire N__94150;
    wire N__94149;
    wire N__94146;
    wire N__94143;
    wire N__94142;
    wire N__94141;
    wire N__94140;
    wire N__94139;
    wire N__94132;
    wire N__94129;
    wire N__94126;
    wire N__94123;
    wire N__94122;
    wire N__94121;
    wire N__94120;
    wire N__94109;
    wire N__94104;
    wire N__94103;
    wire N__94102;
    wire N__94101;
    wire N__94100;
    wire N__94097;
    wire N__94090;
    wire N__94085;
    wire N__94074;
    wire N__94069;
    wire N__94062;
    wire N__94055;
    wire N__94052;
    wire N__94051;
    wire N__94050;
    wire N__94049;
    wire N__94048;
    wire N__94045;
    wire N__94042;
    wire N__94037;
    wire N__94034;
    wire N__94029;
    wire N__94024;
    wire N__94021;
    wire N__94016;
    wire N__94013;
    wire N__94010;
    wire N__93999;
    wire N__93990;
    wire N__93983;
    wire N__93972;
    wire N__93969;
    wire N__93968;
    wire N__93967;
    wire N__93966;
    wire N__93965;
    wire N__93964;
    wire N__93961;
    wire N__93958;
    wire N__93947;
    wire N__93944;
    wire N__93933;
    wire N__93932;
    wire N__93931;
    wire N__93930;
    wire N__93929;
    wire N__93928;
    wire N__93927;
    wire N__93926;
    wire N__93925;
    wire N__93924;
    wire N__93923;
    wire N__93920;
    wire N__93909;
    wire N__93906;
    wire N__93899;
    wire N__93894;
    wire N__93891;
    wire N__93886;
    wire N__93883;
    wire N__93872;
    wire N__93865;
    wire N__93858;
    wire N__93845;
    wire N__93842;
    wire N__93829;
    wire N__93816;
    wire N__93815;
    wire N__93812;
    wire N__93811;
    wire N__93810;
    wire N__93809;
    wire N__93808;
    wire N__93807;
    wire N__93806;
    wire N__93805;
    wire N__93804;
    wire N__93801;
    wire N__93798;
    wire N__93795;
    wire N__93792;
    wire N__93789;
    wire N__93782;
    wire N__93777;
    wire N__93774;
    wire N__93773;
    wire N__93772;
    wire N__93771;
    wire N__93770;
    wire N__93769;
    wire N__93768;
    wire N__93765;
    wire N__93760;
    wire N__93753;
    wire N__93744;
    wire N__93729;
    wire N__93722;
    wire N__93717;
    wire N__93704;
    wire N__93699;
    wire N__93696;
    wire N__93687;
    wire N__93676;
    wire N__93665;
    wire N__93654;
    wire N__93643;
    wire N__93638;
    wire N__93635;
    wire N__93632;
    wire N__93619;
    wire N__93618;
    wire N__93615;
    wire N__93608;
    wire N__93599;
    wire N__93594;
    wire N__93591;
    wire N__93588;
    wire N__93585;
    wire N__93580;
    wire N__93575;
    wire N__93564;
    wire N__93559;
    wire N__93556;
    wire N__93547;
    wire N__93532;
    wire N__93517;
    wire N__93514;
    wire N__93481;
    wire N__93478;
    wire N__93477;
    wire N__93474;
    wire N__93471;
    wire N__93468;
    wire N__93465;
    wire N__93460;
    wire N__93457;
    wire N__93456;
    wire N__93455;
    wire N__93454;
    wire N__93453;
    wire N__93452;
    wire N__93451;
    wire N__93450;
    wire N__93449;
    wire N__93448;
    wire N__93447;
    wire N__93446;
    wire N__93443;
    wire N__93442;
    wire N__93441;
    wire N__93440;
    wire N__93439;
    wire N__93438;
    wire N__93437;
    wire N__93436;
    wire N__93435;
    wire N__93434;
    wire N__93433;
    wire N__93432;
    wire N__93431;
    wire N__93430;
    wire N__93429;
    wire N__93428;
    wire N__93427;
    wire N__93426;
    wire N__93425;
    wire N__93424;
    wire N__93423;
    wire N__93422;
    wire N__93421;
    wire N__93420;
    wire N__93419;
    wire N__93418;
    wire N__93417;
    wire N__93416;
    wire N__93415;
    wire N__93414;
    wire N__93413;
    wire N__93412;
    wire N__93411;
    wire N__93410;
    wire N__93409;
    wire N__93408;
    wire N__93407;
    wire N__93406;
    wire N__93405;
    wire N__93404;
    wire N__93403;
    wire N__93402;
    wire N__93401;
    wire N__93400;
    wire N__93399;
    wire N__93398;
    wire N__93397;
    wire N__93396;
    wire N__93395;
    wire N__93394;
    wire N__93393;
    wire N__93392;
    wire N__93391;
    wire N__93390;
    wire N__93389;
    wire N__93388;
    wire N__93387;
    wire N__93386;
    wire N__93385;
    wire N__93384;
    wire N__93383;
    wire N__93382;
    wire N__93381;
    wire N__93380;
    wire N__93379;
    wire N__93378;
    wire N__93377;
    wire N__93376;
    wire N__93375;
    wire N__93374;
    wire N__93373;
    wire N__93372;
    wire N__93371;
    wire N__93370;
    wire N__93369;
    wire N__93368;
    wire N__93367;
    wire N__93366;
    wire N__93365;
    wire N__93364;
    wire N__93363;
    wire N__93362;
    wire N__93361;
    wire N__93360;
    wire N__93359;
    wire N__93358;
    wire N__93357;
    wire N__93356;
    wire N__93355;
    wire N__93354;
    wire N__93353;
    wire N__93352;
    wire N__93351;
    wire N__93350;
    wire N__93349;
    wire N__93348;
    wire N__93347;
    wire N__93346;
    wire N__93345;
    wire N__93344;
    wire N__93343;
    wire N__93342;
    wire N__93341;
    wire N__93340;
    wire N__93339;
    wire N__93338;
    wire N__93337;
    wire N__93336;
    wire N__93335;
    wire N__93334;
    wire N__93333;
    wire N__93332;
    wire N__93331;
    wire N__93330;
    wire N__93329;
    wire N__93328;
    wire N__93327;
    wire N__93326;
    wire N__93325;
    wire N__93324;
    wire N__93323;
    wire N__93322;
    wire N__93321;
    wire N__93320;
    wire N__93319;
    wire N__93318;
    wire N__93317;
    wire N__93316;
    wire N__93315;
    wire N__93314;
    wire N__93313;
    wire N__93312;
    wire N__93311;
    wire N__93310;
    wire N__93309;
    wire N__93308;
    wire N__93307;
    wire N__93306;
    wire N__93305;
    wire N__93304;
    wire N__93303;
    wire N__93302;
    wire N__93301;
    wire N__93300;
    wire N__93299;
    wire N__93298;
    wire N__93297;
    wire N__93296;
    wire N__93295;
    wire N__93294;
    wire N__93293;
    wire N__93292;
    wire N__93291;
    wire N__93290;
    wire N__93289;
    wire N__93288;
    wire N__93287;
    wire N__93286;
    wire N__93285;
    wire N__93284;
    wire N__93283;
    wire N__93282;
    wire N__93281;
    wire N__93280;
    wire N__93279;
    wire N__93278;
    wire N__93277;
    wire N__93276;
    wire N__93275;
    wire N__93274;
    wire N__93273;
    wire N__93272;
    wire N__93271;
    wire N__93270;
    wire N__93269;
    wire N__93268;
    wire N__93267;
    wire N__93266;
    wire N__93265;
    wire N__93264;
    wire N__93263;
    wire N__93262;
    wire N__93261;
    wire N__93260;
    wire N__93259;
    wire N__93258;
    wire N__93257;
    wire N__93256;
    wire N__93255;
    wire N__93254;
    wire N__93253;
    wire N__93252;
    wire N__93251;
    wire N__93250;
    wire N__93249;
    wire N__93248;
    wire N__93247;
    wire N__93246;
    wire N__93245;
    wire N__93244;
    wire N__93243;
    wire N__93242;
    wire N__93241;
    wire N__93240;
    wire N__93239;
    wire N__93238;
    wire N__93237;
    wire N__93236;
    wire N__93235;
    wire N__93234;
    wire N__93233;
    wire N__93232;
    wire N__93231;
    wire N__93230;
    wire N__93229;
    wire N__93228;
    wire N__93227;
    wire N__93226;
    wire N__93225;
    wire N__93224;
    wire N__93223;
    wire N__93222;
    wire N__93221;
    wire N__93220;
    wire N__93219;
    wire N__92746;
    wire N__92743;
    wire N__92740;
    wire N__92737;
    wire N__92734;
    wire N__92731;
    wire N__92728;
    wire N__92725;
    wire N__92722;
    wire N__92719;
    wire N__92716;
    wire N__92713;
    wire N__92710;
    wire N__92707;
    wire N__92704;
    wire N__92701;
    wire N__92698;
    wire N__92695;
    wire N__92694;
    wire N__92691;
    wire N__92688;
    wire N__92685;
    wire N__92682;
    wire N__92677;
    wire N__92676;
    wire N__92675;
    wire N__92674;
    wire N__92673;
    wire N__92672;
    wire N__92669;
    wire N__92668;
    wire N__92667;
    wire N__92666;
    wire N__92665;
    wire N__92664;
    wire N__92663;
    wire N__92662;
    wire N__92661;
    wire N__92660;
    wire N__92659;
    wire N__92658;
    wire N__92657;
    wire N__92656;
    wire N__92655;
    wire N__92654;
    wire N__92653;
    wire N__92652;
    wire N__92651;
    wire N__92650;
    wire N__92649;
    wire N__92648;
    wire N__92647;
    wire N__92646;
    wire N__92637;
    wire N__92636;
    wire N__92635;
    wire N__92634;
    wire N__92633;
    wire N__92630;
    wire N__92629;
    wire N__92628;
    wire N__92627;
    wire N__92626;
    wire N__92625;
    wire N__92624;
    wire N__92623;
    wire N__92622;
    wire N__92621;
    wire N__92620;
    wire N__92619;
    wire N__92618;
    wire N__92617;
    wire N__92616;
    wire N__92613;
    wire N__92612;
    wire N__92611;
    wire N__92610;
    wire N__92609;
    wire N__92606;
    wire N__92605;
    wire N__92600;
    wire N__92599;
    wire N__92598;
    wire N__92597;
    wire N__92596;
    wire N__92595;
    wire N__92594;
    wire N__92593;
    wire N__92590;
    wire N__92589;
    wire N__92588;
    wire N__92587;
    wire N__92586;
    wire N__92585;
    wire N__92584;
    wire N__92583;
    wire N__92582;
    wire N__92581;
    wire N__92580;
    wire N__92577;
    wire N__92568;
    wire N__92567;
    wire N__92566;
    wire N__92565;
    wire N__92564;
    wire N__92563;
    wire N__92562;
    wire N__92561;
    wire N__92560;
    wire N__92557;
    wire N__92556;
    wire N__92555;
    wire N__92546;
    wire N__92545;
    wire N__92542;
    wire N__92541;
    wire N__92540;
    wire N__92531;
    wire N__92522;
    wire N__92521;
    wire N__92520;
    wire N__92519;
    wire N__92518;
    wire N__92517;
    wire N__92514;
    wire N__92511;
    wire N__92504;
    wire N__92499;
    wire N__92496;
    wire N__92495;
    wire N__92494;
    wire N__92493;
    wire N__92492;
    wire N__92491;
    wire N__92482;
    wire N__92477;
    wire N__92470;
    wire N__92465;
    wire N__92462;
    wire N__92459;
    wire N__92450;
    wire N__92449;
    wire N__92448;
    wire N__92447;
    wire N__92446;
    wire N__92445;
    wire N__92444;
    wire N__92443;
    wire N__92442;
    wire N__92441;
    wire N__92436;
    wire N__92433;
    wire N__92432;
    wire N__92431;
    wire N__92430;
    wire N__92427;
    wire N__92426;
    wire N__92425;
    wire N__92424;
    wire N__92421;
    wire N__92420;
    wire N__92419;
    wire N__92416;
    wire N__92415;
    wire N__92414;
    wire N__92413;
    wire N__92410;
    wire N__92409;
    wire N__92408;
    wire N__92407;
    wire N__92402;
    wire N__92401;
    wire N__92400;
    wire N__92399;
    wire N__92398;
    wire N__92393;
    wire N__92390;
    wire N__92389;
    wire N__92388;
    wire N__92387;
    wire N__92386;
    wire N__92385;
    wire N__92384;
    wire N__92381;
    wire N__92380;
    wire N__92377;
    wire N__92374;
    wire N__92373;
    wire N__92372;
    wire N__92367;
    wire N__92364;
    wire N__92361;
    wire N__92358;
    wire N__92353;
    wire N__92352;
    wire N__92351;
    wire N__92350;
    wire N__92347;
    wire N__92344;
    wire N__92341;
    wire N__92334;
    wire N__92329;
    wire N__92322;
    wire N__92321;
    wire N__92320;
    wire N__92319;
    wire N__92318;
    wire N__92317;
    wire N__92316;
    wire N__92313;
    wire N__92310;
    wire N__92307;
    wire N__92304;
    wire N__92299;
    wire N__92294;
    wire N__92289;
    wire N__92288;
    wire N__92287;
    wire N__92286;
    wire N__92285;
    wire N__92284;
    wire N__92283;
    wire N__92282;
    wire N__92281;
    wire N__92276;
    wire N__92273;
    wire N__92272;
    wire N__92271;
    wire N__92270;
    wire N__92269;
    wire N__92268;
    wire N__92263;
    wire N__92260;
    wire N__92257;
    wire N__92252;
    wire N__92249;
    wire N__92246;
    wire N__92243;
    wire N__92240;
    wire N__92237;
    wire N__92228;
    wire N__92223;
    wire N__92220;
    wire N__92217;
    wire N__92216;
    wire N__92215;
    wire N__92214;
    wire N__92213;
    wire N__92212;
    wire N__92211;
    wire N__92210;
    wire N__92209;
    wire N__92206;
    wire N__92197;
    wire N__92192;
    wire N__92191;
    wire N__92188;
    wire N__92185;
    wire N__92180;
    wire N__92177;
    wire N__92176;
    wire N__92175;
    wire N__92174;
    wire N__92173;
    wire N__92172;
    wire N__92171;
    wire N__92170;
    wire N__92169;
    wire N__92166;
    wire N__92159;
    wire N__92152;
    wire N__92143;
    wire N__92142;
    wire N__92141;
    wire N__92140;
    wire N__92139;
    wire N__92136;
    wire N__92135;
    wire N__92132;
    wire N__92131;
    wire N__92130;
    wire N__92129;
    wire N__92124;
    wire N__92121;
    wire N__92116;
    wire N__92115;
    wire N__92114;
    wire N__92113;
    wire N__92112;
    wire N__92111;
    wire N__92110;
    wire N__92109;
    wire N__92108;
    wire N__92107;
    wire N__92106;
    wire N__92105;
    wire N__92104;
    wire N__92101;
    wire N__92098;
    wire N__92097;
    wire N__92092;
    wire N__92083;
    wire N__92078;
    wire N__92073;
    wire N__92070;
    wire N__92063;
    wire N__92062;
    wire N__92057;
    wire N__92052;
    wire N__92049;
    wire N__92042;
    wire N__92041;
    wire N__92040;
    wire N__92039;
    wire N__92032;
    wire N__92031;
    wire N__92030;
    wire N__92029;
    wire N__92028;
    wire N__92027;
    wire N__92022;
    wire N__92019;
    wire N__92016;
    wire N__92011;
    wire N__92010;
    wire N__92009;
    wire N__92008;
    wire N__92007;
    wire N__92006;
    wire N__92005;
    wire N__92004;
    wire N__92003;
    wire N__91996;
    wire N__91995;
    wire N__91994;
    wire N__91993;
    wire N__91992;
    wire N__91991;
    wire N__91990;
    wire N__91989;
    wire N__91988;
    wire N__91987;
    wire N__91986;
    wire N__91985;
    wire N__91982;
    wire N__91977;
    wire N__91972;
    wire N__91967;
    wire N__91956;
    wire N__91949;
    wire N__91948;
    wire N__91947;
    wire N__91942;
    wire N__91939;
    wire N__91936;
    wire N__91931;
    wire N__91928;
    wire N__91927;
    wire N__91926;
    wire N__91917;
    wire N__91912;
    wire N__91907;
    wire N__91896;
    wire N__91887;
    wire N__91886;
    wire N__91885;
    wire N__91884;
    wire N__91883;
    wire N__91880;
    wire N__91879;
    wire N__91878;
    wire N__91873;
    wire N__91872;
    wire N__91871;
    wire N__91870;
    wire N__91869;
    wire N__91868;
    wire N__91865;
    wire N__91864;
    wire N__91863;
    wire N__91862;
    wire N__91861;
    wire N__91854;
    wire N__91851;
    wire N__91844;
    wire N__91837;
    wire N__91836;
    wire N__91835;
    wire N__91834;
    wire N__91833;
    wire N__91828;
    wire N__91821;
    wire N__91820;
    wire N__91817;
    wire N__91816;
    wire N__91815;
    wire N__91814;
    wire N__91813;
    wire N__91812;
    wire N__91811;
    wire N__91810;
    wire N__91809;
    wire N__91808;
    wire N__91803;
    wire N__91798;
    wire N__91797;
    wire N__91796;
    wire N__91787;
    wire N__91786;
    wire N__91785;
    wire N__91784;
    wire N__91781;
    wire N__91776;
    wire N__91775;
    wire N__91772;
    wire N__91769;
    wire N__91768;
    wire N__91767;
    wire N__91766;
    wire N__91765;
    wire N__91764;
    wire N__91763;
    wire N__91760;
    wire N__91753;
    wire N__91748;
    wire N__91747;
    wire N__91746;
    wire N__91745;
    wire N__91744;
    wire N__91743;
    wire N__91740;
    wire N__91739;
    wire N__91738;
    wire N__91737;
    wire N__91736;
    wire N__91735;
    wire N__91734;
    wire N__91733;
    wire N__91732;
    wire N__91731;
    wire N__91730;
    wire N__91723;
    wire N__91720;
    wire N__91717;
    wire N__91712;
    wire N__91707;
    wire N__91700;
    wire N__91699;
    wire N__91694;
    wire N__91689;
    wire N__91684;
    wire N__91681;
    wire N__91680;
    wire N__91679;
    wire N__91670;
    wire N__91663;
    wire N__91662;
    wire N__91661;
    wire N__91658;
    wire N__91655;
    wire N__91650;
    wire N__91647;
    wire N__91644;
    wire N__91643;
    wire N__91642;
    wire N__91633;
    wire N__91630;
    wire N__91625;
    wire N__91614;
    wire N__91611;
    wire N__91606;
    wire N__91603;
    wire N__91602;
    wire N__91601;
    wire N__91600;
    wire N__91597;
    wire N__91594;
    wire N__91591;
    wire N__91590;
    wire N__91589;
    wire N__91588;
    wire N__91587;
    wire N__91584;
    wire N__91575;
    wire N__91574;
    wire N__91573;
    wire N__91572;
    wire N__91571;
    wire N__91570;
    wire N__91569;
    wire N__91568;
    wire N__91567;
    wire N__91564;
    wire N__91553;
    wire N__91548;
    wire N__91537;
    wire N__91532;
    wire N__91521;
    wire N__91518;
    wire N__91511;
    wire N__91506;
    wire N__91503;
    wire N__91502;
    wire N__91499;
    wire N__91492;
    wire N__91483;
    wire N__91480;
    wire N__91479;
    wire N__91478;
    wire N__91477;
    wire N__91474;
    wire N__91471;
    wire N__91462;
    wire N__91453;
    wire N__91450;
    wire N__91447;
    wire N__91440;
    wire N__91435;
    wire N__91432;
    wire N__91427;
    wire N__91422;
    wire N__91419;
    wire N__91418;
    wire N__91417;
    wire N__91416;
    wire N__91411;
    wire N__91406;
    wire N__91405;
    wire N__91404;
    wire N__91403;
    wire N__91400;
    wire N__91397;
    wire N__91394;
    wire N__91391;
    wire N__91386;
    wire N__91381;
    wire N__91378;
    wire N__91369;
    wire N__91368;
    wire N__91367;
    wire N__91366;
    wire N__91365;
    wire N__91364;
    wire N__91363;
    wire N__91362;
    wire N__91357;
    wire N__91356;
    wire N__91355;
    wire N__91354;
    wire N__91353;
    wire N__91352;
    wire N__91351;
    wire N__91350;
    wire N__91349;
    wire N__91348;
    wire N__91347;
    wire N__91340;
    wire N__91331;
    wire N__91330;
    wire N__91329;
    wire N__91328;
    wire N__91327;
    wire N__91326;
    wire N__91325;
    wire N__91322;
    wire N__91319;
    wire N__91316;
    wire N__91309;
    wire N__91302;
    wire N__91299;
    wire N__91296;
    wire N__91295;
    wire N__91294;
    wire N__91293;
    wire N__91292;
    wire N__91291;
    wire N__91290;
    wire N__91289;
    wire N__91288;
    wire N__91285;
    wire N__91284;
    wire N__91283;
    wire N__91282;
    wire N__91275;
    wire N__91268;
    wire N__91265;
    wire N__91256;
    wire N__91251;
    wire N__91246;
    wire N__91243;
    wire N__91242;
    wire N__91241;
    wire N__91240;
    wire N__91239;
    wire N__91238;
    wire N__91237;
    wire N__91236;
    wire N__91235;
    wire N__91234;
    wire N__91231;
    wire N__91230;
    wire N__91229;
    wire N__91228;
    wire N__91227;
    wire N__91226;
    wire N__91225;
    wire N__91224;
    wire N__91223;
    wire N__91222;
    wire N__91221;
    wire N__91214;
    wire N__91209;
    wire N__91204;
    wire N__91195;
    wire N__91188;
    wire N__91185;
    wire N__91180;
    wire N__91175;
    wire N__91164;
    wire N__91161;
    wire N__91158;
    wire N__91155;
    wire N__91146;
    wire N__91139;
    wire N__91132;
    wire N__91127;
    wire N__91118;
    wire N__91115;
    wire N__91112;
    wire N__91111;
    wire N__91110;
    wire N__91103;
    wire N__91096;
    wire N__91093;
    wire N__91084;
    wire N__91075;
    wire N__91072;
    wire N__91069;
    wire N__91064;
    wire N__91057;
    wire N__91052;
    wire N__91047;
    wire N__91044;
    wire N__91039;
    wire N__91034;
    wire N__91027;
    wire N__91024;
    wire N__91019;
    wire N__91012;
    wire N__91007;
    wire N__91004;
    wire N__91001;
    wire N__90998;
    wire N__90991;
    wire N__90982;
    wire N__90979;
    wire N__90978;
    wire N__90977;
    wire N__90976;
    wire N__90975;
    wire N__90974;
    wire N__90973;
    wire N__90968;
    wire N__90963;
    wire N__90960;
    wire N__90953;
    wire N__90946;
    wire N__90937;
    wire N__90930;
    wire N__90919;
    wire N__90910;
    wire N__90895;
    wire N__90892;
    wire N__90885;
    wire N__90882;
    wire N__90879;
    wire N__90878;
    wire N__90873;
    wire N__90872;
    wire N__90871;
    wire N__90870;
    wire N__90869;
    wire N__90860;
    wire N__90859;
    wire N__90858;
    wire N__90857;
    wire N__90856;
    wire N__90855;
    wire N__90854;
    wire N__90853;
    wire N__90850;
    wire N__90841;
    wire N__90836;
    wire N__90833;
    wire N__90830;
    wire N__90825;
    wire N__90816;
    wire N__90811;
    wire N__90800;
    wire N__90791;
    wire N__90788;
    wire N__90783;
    wire N__90776;
    wire N__90759;
    wire N__90756;
    wire N__90741;
    wire N__90728;
    wire N__90723;
    wire N__90718;
    wire N__90713;
    wire N__90712;
    wire N__90711;
    wire N__90710;
    wire N__90709;
    wire N__90708;
    wire N__90707;
    wire N__90706;
    wire N__90705;
    wire N__90696;
    wire N__90685;
    wire N__90676;
    wire N__90671;
    wire N__90668;
    wire N__90663;
    wire N__90658;
    wire N__90655;
    wire N__90652;
    wire N__90649;
    wire N__90646;
    wire N__90641;
    wire N__90636;
    wire N__90635;
    wire N__90634;
    wire N__90627;
    wire N__90624;
    wire N__90619;
    wire N__90616;
    wire N__90611;
    wire N__90608;
    wire N__90603;
    wire N__90600;
    wire N__90595;
    wire N__90588;
    wire N__90583;
    wire N__90576;
    wire N__90567;
    wire N__90564;
    wire N__90561;
    wire N__90554;
    wire N__90547;
    wire N__90534;
    wire N__90529;
    wire N__90528;
    wire N__90527;
    wire N__90522;
    wire N__90517;
    wire N__90510;
    wire N__90503;
    wire N__90494;
    wire N__90489;
    wire N__90482;
    wire N__90477;
    wire N__90460;
    wire N__90457;
    wire N__90454;
    wire N__90451;
    wire N__90448;
    wire N__90445;
    wire N__90442;
    wire N__90439;
    wire N__90436;
    wire N__90435;
    wire N__90432;
    wire N__90429;
    wire N__90426;
    wire N__90423;
    wire N__90418;
    wire N__90415;
    wire N__90412;
    wire N__90409;
    wire N__90406;
    wire N__90403;
    wire N__90400;
    wire N__90399;
    wire N__90398;
    wire N__90395;
    wire N__90392;
    wire N__90391;
    wire N__90390;
    wire N__90389;
    wire N__90388;
    wire N__90387;
    wire N__90386;
    wire N__90385;
    wire N__90382;
    wire N__90379;
    wire N__90370;
    wire N__90369;
    wire N__90366;
    wire N__90363;
    wire N__90362;
    wire N__90359;
    wire N__90356;
    wire N__90355;
    wire N__90354;
    wire N__90353;
    wire N__90352;
    wire N__90351;
    wire N__90350;
    wire N__90349;
    wire N__90348;
    wire N__90347;
    wire N__90344;
    wire N__90343;
    wire N__90342;
    wire N__90341;
    wire N__90340;
    wire N__90339;
    wire N__90336;
    wire N__90333;
    wire N__90330;
    wire N__90325;
    wire N__90322;
    wire N__90319;
    wire N__90312;
    wire N__90309;
    wire N__90306;
    wire N__90303;
    wire N__90302;
    wire N__90301;
    wire N__90300;
    wire N__90297;
    wire N__90294;
    wire N__90291;
    wire N__90290;
    wire N__90287;
    wire N__90284;
    wire N__90279;
    wire N__90276;
    wire N__90273;
    wire N__90270;
    wire N__90267;
    wire N__90262;
    wire N__90257;
    wire N__90254;
    wire N__90253;
    wire N__90252;
    wire N__90251;
    wire N__90250;
    wire N__90245;
    wire N__90242;
    wire N__90239;
    wire N__90236;
    wire N__90233;
    wire N__90232;
    wire N__90231;
    wire N__90230;
    wire N__90229;
    wire N__90226;
    wire N__90223;
    wire N__90222;
    wire N__90221;
    wire N__90216;
    wire N__90213;
    wire N__90212;
    wire N__90211;
    wire N__90210;
    wire N__90207;
    wire N__90202;
    wire N__90199;
    wire N__90196;
    wire N__90193;
    wire N__90186;
    wire N__90183;
    wire N__90174;
    wire N__90171;
    wire N__90164;
    wire N__90161;
    wire N__90158;
    wire N__90155;
    wire N__90152;
    wire N__90149;
    wire N__90144;
    wire N__90143;
    wire N__90142;
    wire N__90141;
    wire N__90138;
    wire N__90135;
    wire N__90134;
    wire N__90131;
    wire N__90122;
    wire N__90119;
    wire N__90116;
    wire N__90109;
    wire N__90102;
    wire N__90101;
    wire N__90096;
    wire N__90093;
    wire N__90090;
    wire N__90085;
    wire N__90084;
    wire N__90083;
    wire N__90082;
    wire N__90081;
    wire N__90080;
    wire N__90077;
    wire N__90074;
    wire N__90067;
    wire N__90066;
    wire N__90065;
    wire N__90062;
    wire N__90059;
    wire N__90056;
    wire N__90055;
    wire N__90054;
    wire N__90053;
    wire N__90048;
    wire N__90039;
    wire N__90036;
    wire N__90035;
    wire N__90034;
    wire N__90029;
    wire N__90026;
    wire N__90023;
    wire N__90022;
    wire N__90019;
    wire N__90018;
    wire N__90009;
    wire N__90006;
    wire N__90001;
    wire N__89996;
    wire N__89993;
    wire N__89988;
    wire N__89985;
    wire N__89982;
    wire N__89979;
    wire N__89978;
    wire N__89975;
    wire N__89970;
    wire N__89965;
    wire N__89964;
    wire N__89957;
    wire N__89954;
    wire N__89953;
    wire N__89950;
    wire N__89947;
    wire N__89946;
    wire N__89945;
    wire N__89944;
    wire N__89943;
    wire N__89942;
    wire N__89939;
    wire N__89932;
    wire N__89921;
    wire N__89918;
    wire N__89915;
    wire N__89910;
    wire N__89907;
    wire N__89906;
    wire N__89905;
    wire N__89900;
    wire N__89897;
    wire N__89892;
    wire N__89883;
    wire N__89882;
    wire N__89881;
    wire N__89880;
    wire N__89877;
    wire N__89876;
    wire N__89873;
    wire N__89868;
    wire N__89865;
    wire N__89862;
    wire N__89857;
    wire N__89854;
    wire N__89851;
    wire N__89850;
    wire N__89845;
    wire N__89840;
    wire N__89833;
    wire N__89830;
    wire N__89827;
    wire N__89826;
    wire N__89825;
    wire N__89822;
    wire N__89817;
    wire N__89808;
    wire N__89805;
    wire N__89794;
    wire N__89789;
    wire N__89776;
    wire N__89773;
    wire N__89770;
    wire N__89767;
    wire N__89764;
    wire N__89761;
    wire N__89758;
    wire N__89755;
    wire N__89752;
    wire N__89749;
    wire N__89748;
    wire N__89745;
    wire N__89742;
    wire N__89737;
    wire N__89734;
    wire N__89733;
    wire N__89730;
    wire N__89727;
    wire N__89722;
    wire N__89719;
    wire N__89716;
    wire N__89715;
    wire N__89712;
    wire N__89709;
    wire N__89704;
    wire N__89701;
    wire N__89698;
    wire N__89695;
    wire N__89694;
    wire N__89691;
    wire N__89688;
    wire N__89685;
    wire N__89682;
    wire N__89677;
    wire N__89674;
    wire N__89671;
    wire N__89670;
    wire N__89667;
    wire N__89664;
    wire N__89663;
    wire N__89662;
    wire N__89661;
    wire N__89658;
    wire N__89655;
    wire N__89652;
    wire N__89651;
    wire N__89650;
    wire N__89649;
    wire N__89646;
    wire N__89643;
    wire N__89642;
    wire N__89639;
    wire N__89636;
    wire N__89633;
    wire N__89630;
    wire N__89627;
    wire N__89626;
    wire N__89625;
    wire N__89624;
    wire N__89621;
    wire N__89616;
    wire N__89613;
    wire N__89612;
    wire N__89611;
    wire N__89610;
    wire N__89609;
    wire N__89604;
    wire N__89601;
    wire N__89596;
    wire N__89589;
    wire N__89586;
    wire N__89581;
    wire N__89578;
    wire N__89573;
    wire N__89570;
    wire N__89551;
    wire N__89548;
    wire N__89545;
    wire N__89542;
    wire N__89541;
    wire N__89538;
    wire N__89535;
    wire N__89530;
    wire N__89529;
    wire N__89528;
    wire N__89527;
    wire N__89526;
    wire N__89523;
    wire N__89522;
    wire N__89521;
    wire N__89520;
    wire N__89519;
    wire N__89518;
    wire N__89517;
    wire N__89516;
    wire N__89515;
    wire N__89514;
    wire N__89511;
    wire N__89508;
    wire N__89505;
    wire N__89504;
    wire N__89501;
    wire N__89494;
    wire N__89493;
    wire N__89492;
    wire N__89491;
    wire N__89490;
    wire N__89489;
    wire N__89488;
    wire N__89487;
    wire N__89484;
    wire N__89483;
    wire N__89482;
    wire N__89479;
    wire N__89476;
    wire N__89475;
    wire N__89474;
    wire N__89473;
    wire N__89472;
    wire N__89469;
    wire N__89468;
    wire N__89465;
    wire N__89464;
    wire N__89463;
    wire N__89462;
    wire N__89461;
    wire N__89460;
    wire N__89459;
    wire N__89458;
    wire N__89457;
    wire N__89456;
    wire N__89455;
    wire N__89454;
    wire N__89453;
    wire N__89452;
    wire N__89451;
    wire N__89448;
    wire N__89445;
    wire N__89440;
    wire N__89439;
    wire N__89438;
    wire N__89437;
    wire N__89436;
    wire N__89435;
    wire N__89434;
    wire N__89431;
    wire N__89428;
    wire N__89423;
    wire N__89412;
    wire N__89401;
    wire N__89400;
    wire N__89399;
    wire N__89398;
    wire N__89395;
    wire N__89390;
    wire N__89389;
    wire N__89388;
    wire N__89385;
    wire N__89382;
    wire N__89379;
    wire N__89374;
    wire N__89367;
    wire N__89362;
    wire N__89357;
    wire N__89354;
    wire N__89351;
    wire N__89346;
    wire N__89343;
    wire N__89336;
    wire N__89333;
    wire N__89330;
    wire N__89327;
    wire N__89326;
    wire N__89325;
    wire N__89322;
    wire N__89317;
    wire N__89310;
    wire N__89307;
    wire N__89304;
    wire N__89303;
    wire N__89302;
    wire N__89301;
    wire N__89300;
    wire N__89299;
    wire N__89296;
    wire N__89293;
    wire N__89290;
    wire N__89283;
    wire N__89278;
    wire N__89277;
    wire N__89276;
    wire N__89275;
    wire N__89272;
    wire N__89269;
    wire N__89254;
    wire N__89241;
    wire N__89238;
    wire N__89235;
    wire N__89230;
    wire N__89227;
    wire N__89222;
    wire N__89217;
    wire N__89206;
    wire N__89199;
    wire N__89194;
    wire N__89191;
    wire N__89186;
    wire N__89179;
    wire N__89176;
    wire N__89171;
    wire N__89162;
    wire N__89155;
    wire N__89150;
    wire N__89143;
    wire N__89140;
    wire N__89137;
    wire N__89128;
    wire N__89125;
    wire N__89124;
    wire N__89123;
    wire N__89122;
    wire N__89119;
    wire N__89116;
    wire N__89115;
    wire N__89114;
    wire N__89111;
    wire N__89108;
    wire N__89105;
    wire N__89104;
    wire N__89103;
    wire N__89102;
    wire N__89099;
    wire N__89096;
    wire N__89093;
    wire N__89090;
    wire N__89087;
    wire N__89084;
    wire N__89081;
    wire N__89078;
    wire N__89075;
    wire N__89074;
    wire N__89073;
    wire N__89072;
    wire N__89069;
    wire N__89066;
    wire N__89063;
    wire N__89058;
    wire N__89049;
    wire N__89046;
    wire N__89043;
    wire N__89040;
    wire N__89039;
    wire N__89038;
    wire N__89035;
    wire N__89032;
    wire N__89029;
    wire N__89024;
    wire N__89017;
    wire N__89012;
    wire N__89011;
    wire N__89010;
    wire N__89005;
    wire N__89002;
    wire N__88995;
    wire N__88990;
    wire N__88981;
    wire N__88978;
    wire N__88977;
    wire N__88972;
    wire N__88969;
    wire N__88966;
    wire N__88963;
    wire N__88960;
    wire N__88957;
    wire N__88954;
    wire N__88951;
    wire N__88948;
    wire N__88947;
    wire N__88944;
    wire N__88939;
    wire N__88936;
    wire N__88935;
    wire N__88932;
    wire N__88927;
    wire N__88924;
    wire N__88923;
    wire N__88920;
    wire N__88915;
    wire N__88912;
    wire N__88911;
    wire N__88908;
    wire N__88907;
    wire N__88906;
    wire N__88905;
    wire N__88902;
    wire N__88901;
    wire N__88900;
    wire N__88899;
    wire N__88898;
    wire N__88891;
    wire N__88888;
    wire N__88887;
    wire N__88886;
    wire N__88885;
    wire N__88884;
    wire N__88883;
    wire N__88882;
    wire N__88881;
    wire N__88880;
    wire N__88879;
    wire N__88878;
    wire N__88877;
    wire N__88872;
    wire N__88869;
    wire N__88864;
    wire N__88861;
    wire N__88858;
    wire N__88857;
    wire N__88856;
    wire N__88855;
    wire N__88854;
    wire N__88853;
    wire N__88852;
    wire N__88851;
    wire N__88850;
    wire N__88849;
    wire N__88846;
    wire N__88845;
    wire N__88844;
    wire N__88843;
    wire N__88842;
    wire N__88841;
    wire N__88838;
    wire N__88837;
    wire N__88836;
    wire N__88835;
    wire N__88834;
    wire N__88829;
    wire N__88822;
    wire N__88821;
    wire N__88820;
    wire N__88819;
    wire N__88818;
    wire N__88815;
    wire N__88814;
    wire N__88813;
    wire N__88812;
    wire N__88811;
    wire N__88810;
    wire N__88809;
    wire N__88808;
    wire N__88805;
    wire N__88804;
    wire N__88803;
    wire N__88802;
    wire N__88799;
    wire N__88796;
    wire N__88793;
    wire N__88788;
    wire N__88783;
    wire N__88780;
    wire N__88779;
    wire N__88778;
    wire N__88777;
    wire N__88776;
    wire N__88775;
    wire N__88774;
    wire N__88773;
    wire N__88772;
    wire N__88771;
    wire N__88770;
    wire N__88761;
    wire N__88760;
    wire N__88759;
    wire N__88758;
    wire N__88757;
    wire N__88756;
    wire N__88755;
    wire N__88754;
    wire N__88753;
    wire N__88750;
    wire N__88749;
    wire N__88748;
    wire N__88745;
    wire N__88744;
    wire N__88743;
    wire N__88742;
    wire N__88739;
    wire N__88738;
    wire N__88737;
    wire N__88734;
    wire N__88729;
    wire N__88728;
    wire N__88727;
    wire N__88726;
    wire N__88721;
    wire N__88716;
    wire N__88711;
    wire N__88708;
    wire N__88705;
    wire N__88702;
    wire N__88701;
    wire N__88700;
    wire N__88699;
    wire N__88698;
    wire N__88693;
    wire N__88688;
    wire N__88681;
    wire N__88676;
    wire N__88675;
    wire N__88674;
    wire N__88671;
    wire N__88670;
    wire N__88669;
    wire N__88666;
    wire N__88661;
    wire N__88656;
    wire N__88653;
    wire N__88650;
    wire N__88647;
    wire N__88644;
    wire N__88641;
    wire N__88632;
    wire N__88625;
    wire N__88620;
    wire N__88619;
    wire N__88618;
    wire N__88617;
    wire N__88614;
    wire N__88613;
    wire N__88612;
    wire N__88611;
    wire N__88610;
    wire N__88609;
    wire N__88608;
    wire N__88607;
    wire N__88606;
    wire N__88605;
    wire N__88604;
    wire N__88603;
    wire N__88602;
    wire N__88599;
    wire N__88598;
    wire N__88597;
    wire N__88596;
    wire N__88595;
    wire N__88592;
    wire N__88591;
    wire N__88590;
    wire N__88589;
    wire N__88588;
    wire N__88587;
    wire N__88586;
    wire N__88585;
    wire N__88584;
    wire N__88583;
    wire N__88582;
    wire N__88581;
    wire N__88576;
    wire N__88575;
    wire N__88572;
    wire N__88569;
    wire N__88560;
    wire N__88555;
    wire N__88550;
    wire N__88547;
    wire N__88546;
    wire N__88545;
    wire N__88542;
    wire N__88541;
    wire N__88540;
    wire N__88539;
    wire N__88538;
    wire N__88537;
    wire N__88536;
    wire N__88535;
    wire N__88534;
    wire N__88531;
    wire N__88526;
    wire N__88523;
    wire N__88518;
    wire N__88515;
    wire N__88514;
    wire N__88513;
    wire N__88512;
    wire N__88511;
    wire N__88510;
    wire N__88509;
    wire N__88504;
    wire N__88497;
    wire N__88486;
    wire N__88483;
    wire N__88476;
    wire N__88475;
    wire N__88474;
    wire N__88473;
    wire N__88470;
    wire N__88465;
    wire N__88460;
    wire N__88455;
    wire N__88452;
    wire N__88449;
    wire N__88448;
    wire N__88447;
    wire N__88446;
    wire N__88445;
    wire N__88444;
    wire N__88443;
    wire N__88442;
    wire N__88439;
    wire N__88436;
    wire N__88433;
    wire N__88428;
    wire N__88423;
    wire N__88412;
    wire N__88409;
    wire N__88408;
    wire N__88405;
    wire N__88402;
    wire N__88395;
    wire N__88392;
    wire N__88385;
    wire N__88378;
    wire N__88375;
    wire N__88374;
    wire N__88373;
    wire N__88372;
    wire N__88371;
    wire N__88366;
    wire N__88363;
    wire N__88360;
    wire N__88355;
    wire N__88354;
    wire N__88351;
    wire N__88348;
    wire N__88343;
    wire N__88342;
    wire N__88341;
    wire N__88338;
    wire N__88337;
    wire N__88336;
    wire N__88335;
    wire N__88334;
    wire N__88333;
    wire N__88332;
    wire N__88331;
    wire N__88330;
    wire N__88327;
    wire N__88326;
    wire N__88325;
    wire N__88322;
    wire N__88321;
    wire N__88320;
    wire N__88319;
    wire N__88318;
    wire N__88311;
    wire N__88304;
    wire N__88303;
    wire N__88302;
    wire N__88301;
    wire N__88300;
    wire N__88297;
    wire N__88294;
    wire N__88287;
    wire N__88282;
    wire N__88279;
    wire N__88276;
    wire N__88273;
    wire N__88268;
    wire N__88265;
    wire N__88264;
    wire N__88263;
    wire N__88262;
    wire N__88261;
    wire N__88258;
    wire N__88255;
    wire N__88254;
    wire N__88253;
    wire N__88248;
    wire N__88247;
    wire N__88246;
    wire N__88245;
    wire N__88244;
    wire N__88243;
    wire N__88242;
    wire N__88241;
    wire N__88240;
    wire N__88239;
    wire N__88238;
    wire N__88235;
    wire N__88234;
    wire N__88233;
    wire N__88232;
    wire N__88229;
    wire N__88228;
    wire N__88219;
    wire N__88216;
    wire N__88213;
    wire N__88208;
    wire N__88205;
    wire N__88200;
    wire N__88195;
    wire N__88188;
    wire N__88185;
    wire N__88180;
    wire N__88177;
    wire N__88166;
    wire N__88163;
    wire N__88160;
    wire N__88157;
    wire N__88152;
    wire N__88149;
    wire N__88148;
    wire N__88143;
    wire N__88134;
    wire N__88129;
    wire N__88126;
    wire N__88125;
    wire N__88122;
    wire N__88109;
    wire N__88104;
    wire N__88101;
    wire N__88098;
    wire N__88097;
    wire N__88096;
    wire N__88095;
    wire N__88086;
    wire N__88083;
    wire N__88076;
    wire N__88071;
    wire N__88070;
    wire N__88069;
    wire N__88066;
    wire N__88063;
    wire N__88060;
    wire N__88055;
    wire N__88054;
    wire N__88053;
    wire N__88052;
    wire N__88051;
    wire N__88050;
    wire N__88047;
    wire N__88046;
    wire N__88045;
    wire N__88044;
    wire N__88043;
    wire N__88042;
    wire N__88041;
    wire N__88040;
    wire N__88037;
    wire N__88036;
    wire N__88033;
    wire N__88032;
    wire N__88031;
    wire N__88030;
    wire N__88029;
    wire N__88024;
    wire N__88019;
    wire N__88016;
    wire N__88009;
    wire N__88008;
    wire N__88007;
    wire N__88006;
    wire N__88005;
    wire N__88004;
    wire N__88003;
    wire N__88002;
    wire N__88001;
    wire N__88000;
    wire N__87999;
    wire N__87998;
    wire N__87997;
    wire N__87996;
    wire N__87993;
    wire N__87988;
    wire N__87985;
    wire N__87978;
    wire N__87977;
    wire N__87974;
    wire N__87971;
    wire N__87968;
    wire N__87961;
    wire N__87954;
    wire N__87951;
    wire N__87944;
    wire N__87941;
    wire N__87936;
    wire N__87933;
    wire N__87930;
    wire N__87925;
    wire N__87920;
    wire N__87915;
    wire N__87914;
    wire N__87911;
    wire N__87904;
    wire N__87903;
    wire N__87902;
    wire N__87897;
    wire N__87892;
    wire N__87887;
    wire N__87886;
    wire N__87883;
    wire N__87880;
    wire N__87871;
    wire N__87862;
    wire N__87847;
    wire N__87844;
    wire N__87841;
    wire N__87836;
    wire N__87833;
    wire N__87830;
    wire N__87823;
    wire N__87820;
    wire N__87815;
    wire N__87810;
    wire N__87805;
    wire N__87800;
    wire N__87797;
    wire N__87794;
    wire N__87793;
    wire N__87792;
    wire N__87791;
    wire N__87784;
    wire N__87781;
    wire N__87776;
    wire N__87771;
    wire N__87768;
    wire N__87763;
    wire N__87760;
    wire N__87757;
    wire N__87756;
    wire N__87755;
    wire N__87754;
    wire N__87753;
    wire N__87752;
    wire N__87751;
    wire N__87742;
    wire N__87737;
    wire N__87736;
    wire N__87735;
    wire N__87734;
    wire N__87733;
    wire N__87730;
    wire N__87727;
    wire N__87726;
    wire N__87723;
    wire N__87718;
    wire N__87717;
    wire N__87716;
    wire N__87715;
    wire N__87714;
    wire N__87713;
    wire N__87712;
    wire N__87709;
    wire N__87702;
    wire N__87699;
    wire N__87694;
    wire N__87689;
    wire N__87684;
    wire N__87679;
    wire N__87678;
    wire N__87677;
    wire N__87676;
    wire N__87667;
    wire N__87666;
    wire N__87665;
    wire N__87664;
    wire N__87663;
    wire N__87662;
    wire N__87661;
    wire N__87658;
    wire N__87651;
    wire N__87650;
    wire N__87649;
    wire N__87648;
    wire N__87647;
    wire N__87646;
    wire N__87643;
    wire N__87634;
    wire N__87627;
    wire N__87620;
    wire N__87615;
    wire N__87610;
    wire N__87607;
    wire N__87604;
    wire N__87601;
    wire N__87596;
    wire N__87595;
    wire N__87594;
    wire N__87591;
    wire N__87586;
    wire N__87583;
    wire N__87582;
    wire N__87581;
    wire N__87580;
    wire N__87579;
    wire N__87578;
    wire N__87577;
    wire N__87576;
    wire N__87569;
    wire N__87562;
    wire N__87553;
    wire N__87544;
    wire N__87537;
    wire N__87534;
    wire N__87531;
    wire N__87530;
    wire N__87529;
    wire N__87528;
    wire N__87527;
    wire N__87524;
    wire N__87521;
    wire N__87512;
    wire N__87507;
    wire N__87502;
    wire N__87497;
    wire N__87492;
    wire N__87489;
    wire N__87486;
    wire N__87481;
    wire N__87476;
    wire N__87473;
    wire N__87472;
    wire N__87469;
    wire N__87468;
    wire N__87467;
    wire N__87466;
    wire N__87465;
    wire N__87460;
    wire N__87457;
    wire N__87452;
    wire N__87447;
    wire N__87446;
    wire N__87445;
    wire N__87444;
    wire N__87441;
    wire N__87436;
    wire N__87433;
    wire N__87432;
    wire N__87431;
    wire N__87430;
    wire N__87429;
    wire N__87428;
    wire N__87427;
    wire N__87426;
    wire N__87425;
    wire N__87424;
    wire N__87423;
    wire N__87422;
    wire N__87421;
    wire N__87412;
    wire N__87407;
    wire N__87404;
    wire N__87397;
    wire N__87396;
    wire N__87395;
    wire N__87394;
    wire N__87393;
    wire N__87392;
    wire N__87389;
    wire N__87384;
    wire N__87379;
    wire N__87374;
    wire N__87369;
    wire N__87362;
    wire N__87357;
    wire N__87356;
    wire N__87355;
    wire N__87354;
    wire N__87351;
    wire N__87344;
    wire N__87337;
    wire N__87336;
    wire N__87335;
    wire N__87334;
    wire N__87327;
    wire N__87322;
    wire N__87315;
    wire N__87306;
    wire N__87303;
    wire N__87302;
    wire N__87301;
    wire N__87300;
    wire N__87299;
    wire N__87298;
    wire N__87297;
    wire N__87296;
    wire N__87291;
    wire N__87276;
    wire N__87269;
    wire N__87266;
    wire N__87263;
    wire N__87260;
    wire N__87259;
    wire N__87246;
    wire N__87243;
    wire N__87238;
    wire N__87235;
    wire N__87230;
    wire N__87227;
    wire N__87224;
    wire N__87223;
    wire N__87218;
    wire N__87217;
    wire N__87216;
    wire N__87211;
    wire N__87206;
    wire N__87199;
    wire N__87194;
    wire N__87189;
    wire N__87186;
    wire N__87179;
    wire N__87178;
    wire N__87177;
    wire N__87176;
    wire N__87175;
    wire N__87170;
    wire N__87165;
    wire N__87158;
    wire N__87149;
    wire N__87144;
    wire N__87139;
    wire N__87136;
    wire N__87131;
    wire N__87120;
    wire N__87117;
    wire N__87114;
    wire N__87111;
    wire N__87108;
    wire N__87103;
    wire N__87098;
    wire N__87095;
    wire N__87092;
    wire N__87089;
    wire N__87082;
    wire N__87077;
    wire N__87070;
    wire N__87067;
    wire N__87064;
    wire N__87063;
    wire N__87056;
    wire N__87053;
    wire N__87048;
    wire N__87045;
    wire N__87042;
    wire N__87039;
    wire N__87032;
    wire N__87027;
    wire N__87024;
    wire N__87021;
    wire N__87016;
    wire N__87015;
    wire N__87008;
    wire N__87001;
    wire N__86998;
    wire N__86993;
    wire N__86990;
    wire N__86989;
    wire N__86988;
    wire N__86985;
    wire N__86984;
    wire N__86983;
    wire N__86982;
    wire N__86979;
    wire N__86974;
    wire N__86965;
    wire N__86956;
    wire N__86953;
    wire N__86950;
    wire N__86945;
    wire N__86942;
    wire N__86929;
    wire N__86926;
    wire N__86923;
    wire N__86922;
    wire N__86921;
    wire N__86920;
    wire N__86919;
    wire N__86916;
    wire N__86909;
    wire N__86898;
    wire N__86893;
    wire N__86890;
    wire N__86879;
    wire N__86872;
    wire N__86867;
    wire N__86866;
    wire N__86863;
    wire N__86862;
    wire N__86861;
    wire N__86860;
    wire N__86859;
    wire N__86858;
    wire N__86855;
    wire N__86846;
    wire N__86841;
    wire N__86832;
    wire N__86827;
    wire N__86822;
    wire N__86811;
    wire N__86804;
    wire N__86801;
    wire N__86798;
    wire N__86795;
    wire N__86792;
    wire N__86785;
    wire N__86758;
    wire N__86755;
    wire N__86752;
    wire N__86749;
    wire N__86746;
    wire N__86743;
    wire N__86740;
    wire N__86737;
    wire N__86736;
    wire N__86733;
    wire N__86730;
    wire N__86727;
    wire N__86724;
    wire N__86719;
    wire N__86716;
    wire N__86713;
    wire N__86710;
    wire N__86709;
    wire N__86706;
    wire N__86703;
    wire N__86698;
    wire N__86695;
    wire N__86692;
    wire N__86689;
    wire N__86688;
    wire N__86685;
    wire N__86682;
    wire N__86679;
    wire N__86676;
    wire N__86671;
    wire N__86668;
    wire N__86665;
    wire N__86664;
    wire N__86663;
    wire N__86662;
    wire N__86661;
    wire N__86660;
    wire N__86659;
    wire N__86658;
    wire N__86657;
    wire N__86656;
    wire N__86655;
    wire N__86652;
    wire N__86649;
    wire N__86646;
    wire N__86645;
    wire N__86642;
    wire N__86639;
    wire N__86636;
    wire N__86633;
    wire N__86630;
    wire N__86627;
    wire N__86624;
    wire N__86621;
    wire N__86618;
    wire N__86615;
    wire N__86612;
    wire N__86607;
    wire N__86600;
    wire N__86591;
    wire N__86590;
    wire N__86589;
    wire N__86588;
    wire N__86587;
    wire N__86586;
    wire N__86585;
    wire N__86584;
    wire N__86583;
    wire N__86582;
    wire N__86579;
    wire N__86576;
    wire N__86575;
    wire N__86574;
    wire N__86573;
    wire N__86572;
    wire N__86571;
    wire N__86568;
    wire N__86565;
    wire N__86560;
    wire N__86559;
    wire N__86556;
    wire N__86555;
    wire N__86554;
    wire N__86553;
    wire N__86552;
    wire N__86551;
    wire N__86550;
    wire N__86549;
    wire N__86546;
    wire N__86545;
    wire N__86544;
    wire N__86543;
    wire N__86542;
    wire N__86541;
    wire N__86540;
    wire N__86539;
    wire N__86536;
    wire N__86533;
    wire N__86532;
    wire N__86531;
    wire N__86530;
    wire N__86529;
    wire N__86528;
    wire N__86525;
    wire N__86522;
    wire N__86521;
    wire N__86518;
    wire N__86517;
    wire N__86514;
    wire N__86513;
    wire N__86510;
    wire N__86509;
    wire N__86508;
    wire N__86507;
    wire N__86506;
    wire N__86501;
    wire N__86500;
    wire N__86497;
    wire N__86496;
    wire N__86493;
    wire N__86492;
    wire N__86489;
    wire N__86488;
    wire N__86485;
    wire N__86484;
    wire N__86481;
    wire N__86478;
    wire N__86473;
    wire N__86470;
    wire N__86467;
    wire N__86460;
    wire N__86449;
    wire N__86442;
    wire N__86431;
    wire N__86430;
    wire N__86429;
    wire N__86428;
    wire N__86427;
    wire N__86426;
    wire N__86425;
    wire N__86416;
    wire N__86409;
    wire N__86394;
    wire N__86391;
    wire N__86390;
    wire N__86389;
    wire N__86386;
    wire N__86385;
    wire N__86382;
    wire N__86381;
    wire N__86378;
    wire N__86377;
    wire N__86376;
    wire N__86375;
    wire N__86374;
    wire N__86373;
    wire N__86372;
    wire N__86371;
    wire N__86370;
    wire N__86369;
    wire N__86368;
    wire N__86367;
    wire N__86366;
    wire N__86365;
    wire N__86364;
    wire N__86363;
    wire N__86362;
    wire N__86361;
    wire N__86360;
    wire N__86357;
    wire N__86350;
    wire N__86335;
    wire N__86318;
    wire N__86317;
    wire N__86314;
    wire N__86313;
    wire N__86310;
    wire N__86309;
    wire N__86306;
    wire N__86305;
    wire N__86302;
    wire N__86299;
    wire N__86296;
    wire N__86295;
    wire N__86288;
    wire N__86283;
    wire N__86270;
    wire N__86267;
    wire N__86264;
    wire N__86261;
    wire N__86258;
    wire N__86255;
    wire N__86254;
    wire N__86251;
    wire N__86248;
    wire N__86245;
    wire N__86242;
    wire N__86239;
    wire N__86236;
    wire N__86233;
    wire N__86230;
    wire N__86227;
    wire N__86224;
    wire N__86223;
    wire N__86220;
    wire N__86219;
    wire N__86216;
    wire N__86215;
    wire N__86214;
    wire N__86211;
    wire N__86208;
    wire N__86203;
    wire N__86200;
    wire N__86183;
    wire N__86180;
    wire N__86175;
    wire N__86172;
    wire N__86167;
    wire N__86160;
    wire N__86149;
    wire N__86140;
    wire N__86131;
    wire N__86116;
    wire N__86113;
    wire N__86102;
    wire N__86089;
    wire N__86086;
    wire N__86077;
    wire N__86074;
    wire N__86071;
    wire N__86068;
    wire N__86067;
    wire N__86064;
    wire N__86061;
    wire N__86056;
    wire N__86055;
    wire N__86054;
    wire N__86051;
    wire N__86048;
    wire N__86045;
    wire N__86044;
    wire N__86043;
    wire N__86040;
    wire N__86039;
    wire N__86038;
    wire N__86037;
    wire N__86032;
    wire N__86029;
    wire N__86026;
    wire N__86023;
    wire N__86020;
    wire N__86017;
    wire N__86014;
    wire N__86011;
    wire N__86002;
    wire N__85997;
    wire N__85992;
    wire N__85989;
    wire N__85984;
    wire N__85983;
    wire N__85982;
    wire N__85981;
    wire N__85978;
    wire N__85975;
    wire N__85972;
    wire N__85969;
    wire N__85966;
    wire N__85961;
    wire N__85958;
    wire N__85955;
    wire N__85952;
    wire N__85949;
    wire N__85942;
    wire N__85939;
    wire N__85936;
    wire N__85935;
    wire N__85932;
    wire N__85929;
    wire N__85924;
    wire N__85921;
    wire N__85918;
    wire N__85917;
    wire N__85914;
    wire N__85911;
    wire N__85906;
    wire N__85903;
    wire N__85900;
    wire N__85897;
    wire N__85894;
    wire N__85893;
    wire N__85890;
    wire N__85887;
    wire N__85882;
    wire N__85879;
    wire N__85876;
    wire N__85873;
    wire N__85872;
    wire N__85869;
    wire N__85866;
    wire N__85861;
    wire N__85858;
    wire N__85857;
    wire N__85856;
    wire N__85855;
    wire N__85854;
    wire N__85853;
    wire N__85852;
    wire N__85851;
    wire N__85850;
    wire N__85849;
    wire N__85848;
    wire N__85847;
    wire N__85846;
    wire N__85845;
    wire N__85844;
    wire N__85843;
    wire N__85842;
    wire N__85839;
    wire N__85834;
    wire N__85831;
    wire N__85828;
    wire N__85827;
    wire N__85826;
    wire N__85825;
    wire N__85824;
    wire N__85823;
    wire N__85822;
    wire N__85821;
    wire N__85820;
    wire N__85819;
    wire N__85818;
    wire N__85817;
    wire N__85816;
    wire N__85815;
    wire N__85814;
    wire N__85813;
    wire N__85812;
    wire N__85811;
    wire N__85810;
    wire N__85809;
    wire N__85808;
    wire N__85807;
    wire N__85806;
    wire N__85805;
    wire N__85804;
    wire N__85797;
    wire N__85788;
    wire N__85785;
    wire N__85778;
    wire N__85775;
    wire N__85766;
    wire N__85761;
    wire N__85758;
    wire N__85755;
    wire N__85754;
    wire N__85749;
    wire N__85748;
    wire N__85745;
    wire N__85742;
    wire N__85739;
    wire N__85736;
    wire N__85735;
    wire N__85734;
    wire N__85729;
    wire N__85724;
    wire N__85723;
    wire N__85722;
    wire N__85721;
    wire N__85718;
    wire N__85711;
    wire N__85708;
    wire N__85705;
    wire N__85696;
    wire N__85693;
    wire N__85688;
    wire N__85679;
    wire N__85676;
    wire N__85673;
    wire N__85670;
    wire N__85667;
    wire N__85664;
    wire N__85663;
    wire N__85662;
    wire N__85661;
    wire N__85660;
    wire N__85659;
    wire N__85658;
    wire N__85657;
    wire N__85656;
    wire N__85655;
    wire N__85654;
    wire N__85653;
    wire N__85652;
    wire N__85649;
    wire N__85644;
    wire N__85641;
    wire N__85636;
    wire N__85635;
    wire N__85634;
    wire N__85633;
    wire N__85632;
    wire N__85631;
    wire N__85630;
    wire N__85629;
    wire N__85628;
    wire N__85627;
    wire N__85626;
    wire N__85625;
    wire N__85624;
    wire N__85623;
    wire N__85622;
    wire N__85621;
    wire N__85618;
    wire N__85615;
    wire N__85610;
    wire N__85607;
    wire N__85600;
    wire N__85597;
    wire N__85594;
    wire N__85577;
    wire N__85572;
    wire N__85569;
    wire N__85568;
    wire N__85567;
    wire N__85566;
    wire N__85565;
    wire N__85564;
    wire N__85563;
    wire N__85560;
    wire N__85557;
    wire N__85552;
    wire N__85541;
    wire N__85540;
    wire N__85537;
    wire N__85534;
    wire N__85529;
    wire N__85524;
    wire N__85523;
    wire N__85522;
    wire N__85521;
    wire N__85516;
    wire N__85515;
    wire N__85512;
    wire N__85505;
    wire N__85504;
    wire N__85503;
    wire N__85502;
    wire N__85499;
    wire N__85496;
    wire N__85493;
    wire N__85488;
    wire N__85485;
    wire N__85482;
    wire N__85481;
    wire N__85480;
    wire N__85473;
    wire N__85470;
    wire N__85457;
    wire N__85456;
    wire N__85453;
    wire N__85450;
    wire N__85441;
    wire N__85440;
    wire N__85439;
    wire N__85438;
    wire N__85437;
    wire N__85432;
    wire N__85431;
    wire N__85426;
    wire N__85423;
    wire N__85414;
    wire N__85407;
    wire N__85406;
    wire N__85403;
    wire N__85400;
    wire N__85395;
    wire N__85392;
    wire N__85391;
    wire N__85390;
    wire N__85389;
    wire N__85388;
    wire N__85387;
    wire N__85382;
    wire N__85381;
    wire N__85378;
    wire N__85375;
    wire N__85370;
    wire N__85365;
    wire N__85360;
    wire N__85353;
    wire N__85352;
    wire N__85349;
    wire N__85348;
    wire N__85345;
    wire N__85344;
    wire N__85343;
    wire N__85338;
    wire N__85335;
    wire N__85330;
    wire N__85329;
    wire N__85326;
    wire N__85325;
    wire N__85324;
    wire N__85323;
    wire N__85322;
    wire N__85319;
    wire N__85316;
    wire N__85311;
    wire N__85306;
    wire N__85303;
    wire N__85302;
    wire N__85297;
    wire N__85292;
    wire N__85287;
    wire N__85284;
    wire N__85281;
    wire N__85280;
    wire N__85279;
    wire N__85276;
    wire N__85273;
    wire N__85270;
    wire N__85269;
    wire N__85266;
    wire N__85263;
    wire N__85262;
    wire N__85261;
    wire N__85254;
    wire N__85251;
    wire N__85248;
    wire N__85245;
    wire N__85242;
    wire N__85241;
    wire N__85238;
    wire N__85235;
    wire N__85232;
    wire N__85231;
    wire N__85230;
    wire N__85229;
    wire N__85228;
    wire N__85227;
    wire N__85226;
    wire N__85219;
    wire N__85214;
    wire N__85211;
    wire N__85206;
    wire N__85203;
    wire N__85202;
    wire N__85201;
    wire N__85196;
    wire N__85189;
    wire N__85186;
    wire N__85181;
    wire N__85174;
    wire N__85171;
    wire N__85170;
    wire N__85169;
    wire N__85168;
    wire N__85167;
    wire N__85166;
    wire N__85165;
    wire N__85164;
    wire N__85161;
    wire N__85156;
    wire N__85151;
    wire N__85146;
    wire N__85141;
    wire N__85134;
    wire N__85129;
    wire N__85126;
    wire N__85119;
    wire N__85116;
    wire N__85111;
    wire N__85110;
    wire N__85103;
    wire N__85102;
    wire N__85101;
    wire N__85090;
    wire N__85085;
    wire N__85082;
    wire N__85079;
    wire N__85076;
    wire N__85075;
    wire N__85068;
    wire N__85065;
    wire N__85056;
    wire N__85053;
    wire N__85052;
    wire N__85051;
    wire N__85050;
    wire N__85047;
    wire N__85044;
    wire N__85035;
    wire N__85032;
    wire N__85027;
    wire N__85022;
    wire N__85019;
    wire N__85016;
    wire N__85013;
    wire N__85010;
    wire N__85007;
    wire N__85006;
    wire N__85005;
    wire N__85002;
    wire N__84999;
    wire N__84996;
    wire N__84991;
    wire N__84988;
    wire N__84981;
    wire N__84976;
    wire N__84973;
    wire N__84968;
    wire N__84967;
    wire N__84966;
    wire N__84965;
    wire N__84962;
    wire N__84959;
    wire N__84956;
    wire N__84941;
    wire N__84938;
    wire N__84935;
    wire N__84934;
    wire N__84929;
    wire N__84924;
    wire N__84921;
    wire N__84912;
    wire N__84909;
    wire N__84908;
    wire N__84905;
    wire N__84902;
    wire N__84899;
    wire N__84896;
    wire N__84889;
    wire N__84886;
    wire N__84883;
    wire N__84872;
    wire N__84867;
    wire N__84864;
    wire N__84847;
    wire N__84844;
    wire N__84841;
    wire N__84838;
    wire N__84837;
    wire N__84834;
    wire N__84831;
    wire N__84828;
    wire N__84825;
    wire N__84820;
    wire N__84817;
    wire N__84814;
    wire N__84813;
    wire N__84810;
    wire N__84807;
    wire N__84804;
    wire N__84801;
    wire N__84796;
    wire N__84793;
    wire N__84790;
    wire N__84787;
    wire N__84784;
    wire N__84781;
    wire N__84778;
    wire N__84775;
    wire N__84774;
    wire N__84771;
    wire N__84768;
    wire N__84763;
    wire N__84760;
    wire N__84759;
    wire N__84756;
    wire N__84753;
    wire N__84748;
    wire N__84745;
    wire N__84742;
    wire N__84739;
    wire N__84736;
    wire N__84733;
    wire N__84732;
    wire N__84729;
    wire N__84726;
    wire N__84721;
    wire N__84718;
    wire N__84715;
    wire N__84712;
    wire N__84709;
    wire N__84706;
    wire N__84705;
    wire N__84702;
    wire N__84699;
    wire N__84698;
    wire N__84697;
    wire N__84696;
    wire N__84695;
    wire N__84694;
    wire N__84691;
    wire N__84688;
    wire N__84683;
    wire N__84676;
    wire N__84675;
    wire N__84674;
    wire N__84673;
    wire N__84672;
    wire N__84671;
    wire N__84670;
    wire N__84669;
    wire N__84668;
    wire N__84667;
    wire N__84664;
    wire N__84657;
    wire N__84650;
    wire N__84645;
    wire N__84642;
    wire N__84637;
    wire N__84634;
    wire N__84619;
    wire N__84618;
    wire N__84615;
    wire N__84612;
    wire N__84607;
    wire N__84604;
    wire N__84601;
    wire N__84598;
    wire N__84597;
    wire N__84594;
    wire N__84591;
    wire N__84586;
    wire N__84583;
    wire N__84582;
    wire N__84579;
    wire N__84576;
    wire N__84573;
    wire N__84568;
    wire N__84565;
    wire N__84562;
    wire N__84559;
    wire N__84558;
    wire N__84555;
    wire N__84552;
    wire N__84547;
    wire N__84544;
    wire N__84543;
    wire N__84540;
    wire N__84537;
    wire N__84532;
    wire N__84529;
    wire N__84526;
    wire N__84523;
    wire N__84520;
    wire N__84517;
    wire N__84514;
    wire N__84511;
    wire N__84508;
    wire N__84505;
    wire N__84502;
    wire N__84501;
    wire N__84498;
    wire N__84495;
    wire N__84490;
    wire N__84487;
    wire N__84484;
    wire N__84481;
    wire N__84480;
    wire N__84477;
    wire N__84474;
    wire N__84469;
    wire N__84466;
    wire N__84463;
    wire N__84460;
    wire N__84457;
    wire N__84454;
    wire N__84453;
    wire N__84450;
    wire N__84447;
    wire N__84444;
    wire N__84441;
    wire N__84438;
    wire N__84435;
    wire N__84430;
    wire N__84427;
    wire N__84424;
    wire N__84421;
    wire N__84418;
    wire N__84415;
    wire N__84412;
    wire N__84409;
    wire N__84406;
    wire N__84405;
    wire N__84402;
    wire N__84399;
    wire N__84394;
    wire N__84391;
    wire N__84390;
    wire N__84387;
    wire N__84384;
    wire N__84379;
    wire N__84376;
    wire N__84373;
    wire N__84372;
    wire N__84369;
    wire N__84366;
    wire N__84363;
    wire N__84360;
    wire N__84355;
    wire N__84352;
    wire N__84349;
    wire N__84346;
    wire N__84343;
    wire N__84340;
    wire N__84339;
    wire N__84336;
    wire N__84333;
    wire N__84330;
    wire N__84327;
    wire N__84322;
    wire N__84319;
    wire N__84316;
    wire N__84313;
    wire N__84310;
    wire N__84307;
    wire N__84304;
    wire N__84301;
    wire N__84298;
    wire N__84297;
    wire N__84294;
    wire N__84291;
    wire N__84286;
    wire N__84283;
    wire N__84280;
    wire N__84277;
    wire N__84274;
    wire N__84271;
    wire N__84268;
    wire N__84265;
    wire N__84264;
    wire N__84261;
    wire N__84258;
    wire N__84253;
    wire N__84250;
    wire N__84247;
    wire N__84244;
    wire N__84243;
    wire N__84240;
    wire N__84237;
    wire N__84232;
    wire N__84229;
    wire N__84228;
    wire N__84225;
    wire N__84222;
    wire N__84219;
    wire N__84216;
    wire N__84211;
    wire N__84208;
    wire N__84205;
    wire N__84204;
    wire N__84201;
    wire N__84198;
    wire N__84193;
    wire N__84190;
    wire N__84189;
    wire N__84186;
    wire N__84183;
    wire N__84178;
    wire N__84175;
    wire N__84172;
    wire N__84169;
    wire N__84168;
    wire N__84165;
    wire N__84162;
    wire N__84159;
    wire N__84154;
    wire N__84151;
    wire N__84148;
    wire N__84145;
    wire N__84142;
    wire N__84141;
    wire N__84138;
    wire N__84135;
    wire N__84130;
    wire N__84127;
    wire N__84124;
    wire N__84121;
    wire N__84118;
    wire N__84115;
    wire N__84114;
    wire N__84113;
    wire N__84112;
    wire N__84111;
    wire N__84102;
    wire N__84099;
    wire N__84096;
    wire N__84095;
    wire N__84094;
    wire N__84093;
    wire N__84090;
    wire N__84089;
    wire N__84088;
    wire N__84087;
    wire N__84086;
    wire N__84083;
    wire N__84076;
    wire N__84075;
    wire N__84074;
    wire N__84073;
    wire N__84072;
    wire N__84071;
    wire N__84070;
    wire N__84067;
    wire N__84058;
    wire N__84053;
    wire N__84044;
    wire N__84039;
    wire N__84028;
    wire N__84027;
    wire N__84026;
    wire N__84023;
    wire N__84022;
    wire N__84019;
    wire N__84018;
    wire N__84017;
    wire N__84016;
    wire N__84005;
    wire N__84004;
    wire N__84003;
    wire N__84002;
    wire N__83999;
    wire N__83998;
    wire N__83997;
    wire N__83996;
    wire N__83995;
    wire N__83992;
    wire N__83991;
    wire N__83988;
    wire N__83985;
    wire N__83974;
    wire N__83967;
    wire N__83966;
    wire N__83965;
    wire N__83964;
    wire N__83961;
    wire N__83960;
    wire N__83959;
    wire N__83950;
    wire N__83947;
    wire N__83938;
    wire N__83935;
    wire N__83926;
    wire N__83923;
    wire N__83920;
    wire N__83917;
    wire N__83914;
    wire N__83913;
    wire N__83910;
    wire N__83909;
    wire N__83908;
    wire N__83907;
    wire N__83906;
    wire N__83905;
    wire N__83904;
    wire N__83901;
    wire N__83898;
    wire N__83885;
    wire N__83878;
    wire N__83875;
    wire N__83872;
    wire N__83869;
    wire N__83866;
    wire N__83863;
    wire N__83860;
    wire N__83857;
    wire N__83854;
    wire N__83851;
    wire N__83848;
    wire N__83847;
    wire N__83844;
    wire N__83841;
    wire N__83838;
    wire N__83835;
    wire N__83830;
    wire N__83827;
    wire N__83824;
    wire N__83821;
    wire N__83818;
    wire N__83815;
    wire N__83812;
    wire N__83811;
    wire N__83808;
    wire N__83805;
    wire N__83802;
    wire N__83799;
    wire N__83794;
    wire N__83791;
    wire N__83788;
    wire N__83785;
    wire N__83784;
    wire N__83779;
    wire N__83776;
    wire N__83773;
    wire N__83770;
    wire N__83767;
    wire N__83764;
    wire N__83761;
    wire N__83758;
    wire N__83757;
    wire N__83754;
    wire N__83751;
    wire N__83746;
    wire N__83743;
    wire N__83740;
    wire N__83737;
    wire N__83734;
    wire N__83733;
    wire N__83730;
    wire N__83727;
    wire N__83724;
    wire N__83721;
    wire N__83716;
    wire N__83713;
    wire N__83710;
    wire N__83707;
    wire N__83704;
    wire N__83701;
    wire N__83698;
    wire N__83695;
    wire N__83692;
    wire N__83689;
    wire N__83686;
    wire N__83683;
    wire N__83680;
    wire N__83677;
    wire N__83674;
    wire N__83673;
    wire N__83672;
    wire N__83671;
    wire N__83670;
    wire N__83667;
    wire N__83664;
    wire N__83661;
    wire N__83658;
    wire N__83657;
    wire N__83654;
    wire N__83653;
    wire N__83652;
    wire N__83651;
    wire N__83648;
    wire N__83643;
    wire N__83634;
    wire N__83631;
    wire N__83628;
    wire N__83617;
    wire N__83614;
    wire N__83613;
    wire N__83610;
    wire N__83607;
    wire N__83606;
    wire N__83605;
    wire N__83604;
    wire N__83603;
    wire N__83602;
    wire N__83601;
    wire N__83600;
    wire N__83599;
    wire N__83598;
    wire N__83593;
    wire N__83590;
    wire N__83575;
    wire N__83572;
    wire N__83563;
    wire N__83562;
    wire N__83561;
    wire N__83560;
    wire N__83557;
    wire N__83556;
    wire N__83555;
    wire N__83546;
    wire N__83541;
    wire N__83536;
    wire N__83533;
    wire N__83532;
    wire N__83527;
    wire N__83524;
    wire N__83521;
    wire N__83518;
    wire N__83517;
    wire N__83516;
    wire N__83515;
    wire N__83514;
    wire N__83511;
    wire N__83506;
    wire N__83503;
    wire N__83500;
    wire N__83491;
    wire N__83490;
    wire N__83485;
    wire N__83484;
    wire N__83481;
    wire N__83478;
    wire N__83477;
    wire N__83476;
    wire N__83473;
    wire N__83468;
    wire N__83465;
    wire N__83458;
    wire N__83457;
    wire N__83456;
    wire N__83455;
    wire N__83450;
    wire N__83449;
    wire N__83448;
    wire N__83447;
    wire N__83446;
    wire N__83441;
    wire N__83438;
    wire N__83429;
    wire N__83428;
    wire N__83425;
    wire N__83420;
    wire N__83417;
    wire N__83412;
    wire N__83409;
    wire N__83404;
    wire N__83401;
    wire N__83398;
    wire N__83395;
    wire N__83392;
    wire N__83389;
    wire N__83388;
    wire N__83387;
    wire N__83386;
    wire N__83385;
    wire N__83384;
    wire N__83383;
    wire N__83382;
    wire N__83381;
    wire N__83380;
    wire N__83379;
    wire N__83378;
    wire N__83377;
    wire N__83376;
    wire N__83375;
    wire N__83374;
    wire N__83371;
    wire N__83362;
    wire N__83361;
    wire N__83358;
    wire N__83357;
    wire N__83354;
    wire N__83345;
    wire N__83344;
    wire N__83343;
    wire N__83342;
    wire N__83341;
    wire N__83340;
    wire N__83339;
    wire N__83336;
    wire N__83335;
    wire N__83332;
    wire N__83329;
    wire N__83328;
    wire N__83325;
    wire N__83322;
    wire N__83317;
    wire N__83314;
    wire N__83313;
    wire N__83312;
    wire N__83311;
    wire N__83308;
    wire N__83305;
    wire N__83302;
    wire N__83299;
    wire N__83298;
    wire N__83295;
    wire N__83292;
    wire N__83291;
    wire N__83290;
    wire N__83287;
    wire N__83284;
    wire N__83281;
    wire N__83278;
    wire N__83275;
    wire N__83272;
    wire N__83267;
    wire N__83264;
    wire N__83261;
    wire N__83258;
    wire N__83255;
    wire N__83252;
    wire N__83247;
    wire N__83244;
    wire N__83241;
    wire N__83234;
    wire N__83231;
    wire N__83228;
    wire N__83225;
    wire N__83222;
    wire N__83219;
    wire N__83216;
    wire N__83209;
    wire N__83206;
    wire N__83201;
    wire N__83198;
    wire N__83191;
    wire N__83180;
    wire N__83177;
    wire N__83174;
    wire N__83171;
    wire N__83158;
    wire N__83153;
    wire N__83150;
    wire N__83137;
    wire N__83136;
    wire N__83131;
    wire N__83128;
    wire N__83125;
    wire N__83122;
    wire N__83121;
    wire N__83118;
    wire N__83115;
    wire N__83112;
    wire N__83109;
    wire N__83104;
    wire N__83103;
    wire N__83100;
    wire N__83097;
    wire N__83094;
    wire N__83089;
    wire N__83086;
    wire N__83083;
    wire N__83080;
    wire N__83077;
    wire N__83076;
    wire N__83073;
    wire N__83070;
    wire N__83065;
    wire N__83062;
    wire N__83061;
    wire N__83058;
    wire N__83055;
    wire N__83050;
    wire N__83047;
    wire N__83044;
    wire N__83041;
    wire N__83038;
    wire N__83035;
    wire N__83032;
    wire N__83029;
    wire N__83026;
    wire N__83023;
    wire N__83020;
    wire N__83017;
    wire N__83014;
    wire N__83011;
    wire N__83008;
    wire N__83007;
    wire N__83004;
    wire N__83001;
    wire N__82996;
    wire N__82993;
    wire N__82990;
    wire N__82987;
    wire N__82986;
    wire N__82983;
    wire N__82980;
    wire N__82975;
    wire N__82972;
    wire N__82969;
    wire N__82966;
    wire N__82963;
    wire N__82960;
    wire N__82957;
    wire N__82954;
    wire N__82953;
    wire N__82952;
    wire N__82951;
    wire N__82950;
    wire N__82949;
    wire N__82946;
    wire N__82941;
    wire N__82940;
    wire N__82939;
    wire N__82936;
    wire N__82935;
    wire N__82934;
    wire N__82931;
    wire N__82928;
    wire N__82927;
    wire N__82926;
    wire N__82925;
    wire N__82922;
    wire N__82921;
    wire N__82920;
    wire N__82919;
    wire N__82916;
    wire N__82911;
    wire N__82910;
    wire N__82909;
    wire N__82908;
    wire N__82905;
    wire N__82904;
    wire N__82899;
    wire N__82898;
    wire N__82897;
    wire N__82894;
    wire N__82891;
    wire N__82888;
    wire N__82887;
    wire N__82886;
    wire N__82885;
    wire N__82882;
    wire N__82879;
    wire N__82876;
    wire N__82873;
    wire N__82872;
    wire N__82871;
    wire N__82870;
    wire N__82869;
    wire N__82864;
    wire N__82859;
    wire N__82856;
    wire N__82853;
    wire N__82850;
    wire N__82847;
    wire N__82844;
    wire N__82841;
    wire N__82838;
    wire N__82835;
    wire N__82832;
    wire N__82827;
    wire N__82824;
    wire N__82821;
    wire N__82818;
    wire N__82817;
    wire N__82812;
    wire N__82807;
    wire N__82798;
    wire N__82795;
    wire N__82788;
    wire N__82785;
    wire N__82780;
    wire N__82777;
    wire N__82774;
    wire N__82771;
    wire N__82760;
    wire N__82757;
    wire N__82756;
    wire N__82753;
    wire N__82750;
    wire N__82747;
    wire N__82744;
    wire N__82739;
    wire N__82736;
    wire N__82725;
    wire N__82722;
    wire N__82705;
    wire N__82704;
    wire N__82701;
    wire N__82698;
    wire N__82693;
    wire N__82690;
    wire N__82687;
    wire N__82686;
    wire N__82683;
    wire N__82680;
    wire N__82675;
    wire N__82672;
    wire N__82669;
    wire N__82666;
    wire N__82663;
    wire N__82660;
    wire N__82657;
    wire N__82654;
    wire N__82651;
    wire N__82648;
    wire N__82645;
    wire N__82642;
    wire N__82639;
    wire N__82636;
    wire N__82633;
    wire N__82630;
    wire N__82627;
    wire N__82624;
    wire N__82621;
    wire N__82618;
    wire N__82615;
    wire N__82612;
    wire N__82609;
    wire N__82606;
    wire N__82603;
    wire N__82600;
    wire N__82597;
    wire N__82596;
    wire N__82593;
    wire N__82590;
    wire N__82585;
    wire N__82582;
    wire N__82579;
    wire N__82576;
    wire N__82573;
    wire N__82570;
    wire N__82567;
    wire N__82564;
    wire N__82561;
    wire N__82558;
    wire N__82555;
    wire N__82552;
    wire N__82549;
    wire N__82546;
    wire N__82543;
    wire N__82540;
    wire N__82537;
    wire N__82534;
    wire N__82531;
    wire N__82528;
    wire N__82525;
    wire N__82522;
    wire N__82519;
    wire N__82516;
    wire N__82513;
    wire N__82510;
    wire N__82507;
    wire N__82504;
    wire N__82501;
    wire N__82498;
    wire N__82495;
    wire N__82492;
    wire N__82489;
    wire N__82486;
    wire N__82483;
    wire N__82480;
    wire N__82477;
    wire N__82474;
    wire N__82471;
    wire N__82468;
    wire N__82465;
    wire N__82462;
    wire N__82459;
    wire N__82456;
    wire N__82453;
    wire N__82450;
    wire N__82447;
    wire N__82444;
    wire N__82441;
    wire N__82438;
    wire N__82435;
    wire N__82432;
    wire N__82429;
    wire N__82426;
    wire N__82425;
    wire N__82424;
    wire N__82421;
    wire N__82420;
    wire N__82417;
    wire N__82414;
    wire N__82413;
    wire N__82412;
    wire N__82411;
    wire N__82406;
    wire N__82399;
    wire N__82398;
    wire N__82397;
    wire N__82394;
    wire N__82391;
    wire N__82390;
    wire N__82389;
    wire N__82386;
    wire N__82383;
    wire N__82378;
    wire N__82369;
    wire N__82368;
    wire N__82367;
    wire N__82366;
    wire N__82365;
    wire N__82364;
    wire N__82361;
    wire N__82358;
    wire N__82355;
    wire N__82352;
    wire N__82345;
    wire N__82342;
    wire N__82339;
    wire N__82324;
    wire N__82323;
    wire N__82322;
    wire N__82321;
    wire N__82320;
    wire N__82319;
    wire N__82318;
    wire N__82317;
    wire N__82316;
    wire N__82315;
    wire N__82314;
    wire N__82313;
    wire N__82312;
    wire N__82311;
    wire N__82310;
    wire N__82307;
    wire N__82304;
    wire N__82301;
    wire N__82298;
    wire N__82297;
    wire N__82294;
    wire N__82293;
    wire N__82292;
    wire N__82291;
    wire N__82276;
    wire N__82269;
    wire N__82260;
    wire N__82253;
    wire N__82248;
    wire N__82247;
    wire N__82246;
    wire N__82245;
    wire N__82244;
    wire N__82243;
    wire N__82242;
    wire N__82241;
    wire N__82240;
    wire N__82239;
    wire N__82238;
    wire N__82237;
    wire N__82234;
    wire N__82227;
    wire N__82224;
    wire N__82219;
    wire N__82214;
    wire N__82213;
    wire N__82210;
    wire N__82207;
    wire N__82206;
    wire N__82203;
    wire N__82200;
    wire N__82197;
    wire N__82196;
    wire N__82195;
    wire N__82194;
    wire N__82193;
    wire N__82192;
    wire N__82191;
    wire N__82190;
    wire N__82189;
    wire N__82188;
    wire N__82187;
    wire N__82186;
    wire N__82185;
    wire N__82184;
    wire N__82181;
    wire N__82178;
    wire N__82177;
    wire N__82176;
    wire N__82175;
    wire N__82174;
    wire N__82171;
    wire N__82162;
    wire N__82155;
    wire N__82146;
    wire N__82131;
    wire N__82118;
    wire N__82115;
    wire N__82104;
    wire N__82087;
    wire N__82086;
    wire N__82085;
    wire N__82084;
    wire N__82083;
    wire N__82082;
    wire N__82081;
    wire N__82066;
    wire N__82063;
    wire N__82062;
    wire N__82061;
    wire N__82060;
    wire N__82059;
    wire N__82058;
    wire N__82057;
    wire N__82056;
    wire N__82055;
    wire N__82052;
    wire N__82049;
    wire N__82042;
    wire N__82033;
    wire N__82032;
    wire N__82031;
    wire N__82028;
    wire N__82023;
    wire N__82020;
    wire N__82015;
    wire N__82006;
    wire N__82003;
    wire N__82002;
    wire N__82001;
    wire N__82000;
    wire N__81999;
    wire N__81998;
    wire N__81997;
    wire N__81982;
    wire N__81981;
    wire N__81980;
    wire N__81979;
    wire N__81978;
    wire N__81977;
    wire N__81976;
    wire N__81973;
    wire N__81966;
    wire N__81963;
    wire N__81958;
    wire N__81955;
    wire N__81952;
    wire N__81947;
    wire N__81940;
    wire N__81937;
    wire N__81934;
    wire N__81931;
    wire N__81928;
    wire N__81925;
    wire N__81922;
    wire N__81919;
    wire N__81916;
    wire N__81913;
    wire N__81912;
    wire N__81911;
    wire N__81910;
    wire N__81909;
    wire N__81908;
    wire N__81905;
    wire N__81896;
    wire N__81893;
    wire N__81892;
    wire N__81891;
    wire N__81890;
    wire N__81889;
    wire N__81888;
    wire N__81887;
    wire N__81886;
    wire N__81885;
    wire N__81884;
    wire N__81883;
    wire N__81882;
    wire N__81881;
    wire N__81876;
    wire N__81867;
    wire N__81860;
    wire N__81847;
    wire N__81838;
    wire N__81837;
    wire N__81834;
    wire N__81833;
    wire N__81830;
    wire N__81823;
    wire N__81820;
    wire N__81817;
    wire N__81814;
    wire N__81811;
    wire N__81808;
    wire N__81805;
    wire N__81802;
    wire N__81799;
    wire N__81796;
    wire N__81793;
    wire N__81790;
    wire N__81789;
    wire N__81784;
    wire N__81781;
    wire N__81778;
    wire N__81777;
    wire N__81776;
    wire N__81775;
    wire N__81774;
    wire N__81773;
    wire N__81764;
    wire N__81761;
    wire N__81760;
    wire N__81757;
    wire N__81756;
    wire N__81755;
    wire N__81754;
    wire N__81751;
    wire N__81746;
    wire N__81743;
    wire N__81740;
    wire N__81739;
    wire N__81738;
    wire N__81735;
    wire N__81732;
    wire N__81727;
    wire N__81722;
    wire N__81713;
    wire N__81710;
    wire N__81707;
    wire N__81704;
    wire N__81697;
    wire N__81694;
    wire N__81691;
    wire N__81688;
    wire N__81685;
    wire N__81682;
    wire N__81679;
    wire N__81678;
    wire N__81677;
    wire N__81676;
    wire N__81675;
    wire N__81674;
    wire N__81673;
    wire N__81672;
    wire N__81667;
    wire N__81660;
    wire N__81653;
    wire N__81650;
    wire N__81647;
    wire N__81644;
    wire N__81641;
    wire N__81636;
    wire N__81631;
    wire N__81630;
    wire N__81629;
    wire N__81622;
    wire N__81619;
    wire N__81618;
    wire N__81615;
    wire N__81612;
    wire N__81609;
    wire N__81606;
    wire N__81601;
    wire N__81598;
    wire N__81595;
    wire N__81592;
    wire N__81589;
    wire N__81586;
    wire N__81583;
    wire N__81580;
    wire N__81577;
    wire N__81574;
    wire N__81571;
    wire N__81568;
    wire N__81565;
    wire N__81562;
    wire N__81559;
    wire N__81556;
    wire N__81553;
    wire N__81550;
    wire N__81547;
    wire N__81544;
    wire N__81541;
    wire N__81538;
    wire N__81535;
    wire N__81532;
    wire N__81529;
    wire N__81526;
    wire N__81523;
    wire N__81520;
    wire N__81517;
    wire N__81514;
    wire N__81513;
    wire N__81512;
    wire N__81511;
    wire N__81510;
    wire N__81507;
    wire N__81504;
    wire N__81499;
    wire N__81496;
    wire N__81495;
    wire N__81492;
    wire N__81489;
    wire N__81486;
    wire N__81483;
    wire N__81482;
    wire N__81481;
    wire N__81480;
    wire N__81479;
    wire N__81478;
    wire N__81475;
    wire N__81474;
    wire N__81473;
    wire N__81472;
    wire N__81471;
    wire N__81470;
    wire N__81469;
    wire N__81468;
    wire N__81467;
    wire N__81466;
    wire N__81457;
    wire N__81454;
    wire N__81451;
    wire N__81450;
    wire N__81449;
    wire N__81448;
    wire N__81443;
    wire N__81442;
    wire N__81441;
    wire N__81440;
    wire N__81439;
    wire N__81438;
    wire N__81437;
    wire N__81434;
    wire N__81433;
    wire N__81430;
    wire N__81425;
    wire N__81422;
    wire N__81417;
    wire N__81416;
    wire N__81413;
    wire N__81410;
    wire N__81405;
    wire N__81400;
    wire N__81399;
    wire N__81396;
    wire N__81393;
    wire N__81388;
    wire N__81385;
    wire N__81382;
    wire N__81377;
    wire N__81374;
    wire N__81369;
    wire N__81366;
    wire N__81363;
    wire N__81358;
    wire N__81355;
    wire N__81352;
    wire N__81349;
    wire N__81348;
    wire N__81343;
    wire N__81340;
    wire N__81337;
    wire N__81334;
    wire N__81329;
    wire N__81326;
    wire N__81321;
    wire N__81314;
    wire N__81309;
    wire N__81306;
    wire N__81305;
    wire N__81302;
    wire N__81297;
    wire N__81294;
    wire N__81293;
    wire N__81290;
    wire N__81289;
    wire N__81288;
    wire N__81283;
    wire N__81280;
    wire N__81277;
    wire N__81274;
    wire N__81273;
    wire N__81270;
    wire N__81265;
    wire N__81262;
    wire N__81259;
    wire N__81252;
    wire N__81249;
    wire N__81246;
    wire N__81245;
    wire N__81240;
    wire N__81239;
    wire N__81234;
    wire N__81233;
    wire N__81230;
    wire N__81227;
    wire N__81224;
    wire N__81219;
    wire N__81214;
    wire N__81211;
    wire N__81208;
    wire N__81205;
    wire N__81202;
    wire N__81199;
    wire N__81196;
    wire N__81195;
    wire N__81192;
    wire N__81191;
    wire N__81188;
    wire N__81187;
    wire N__81186;
    wire N__81179;
    wire N__81174;
    wire N__81169;
    wire N__81164;
    wire N__81159;
    wire N__81156;
    wire N__81153;
    wire N__81146;
    wire N__81143;
    wire N__81140;
    wire N__81135;
    wire N__81132;
    wire N__81127;
    wire N__81122;
    wire N__81119;
    wire N__81106;
    wire N__81103;
    wire N__81100;
    wire N__81099;
    wire N__81094;
    wire N__81093;
    wire N__81092;
    wire N__81091;
    wire N__81088;
    wire N__81087;
    wire N__81086;
    wire N__81083;
    wire N__81078;
    wire N__81075;
    wire N__81070;
    wire N__81067;
    wire N__81064;
    wire N__81063;
    wire N__81062;
    wire N__81057;
    wire N__81056;
    wire N__81055;
    wire N__81054;
    wire N__81053;
    wire N__81052;
    wire N__81051;
    wire N__81050;
    wire N__81049;
    wire N__81046;
    wire N__81043;
    wire N__81038;
    wire N__81037;
    wire N__81034;
    wire N__81017;
    wire N__81016;
    wire N__81015;
    wire N__81012;
    wire N__81007;
    wire N__81004;
    wire N__80999;
    wire N__80994;
    wire N__80993;
    wire N__80992;
    wire N__80989;
    wire N__80986;
    wire N__80983;
    wire N__80980;
    wire N__80977;
    wire N__80972;
    wire N__80969;
    wire N__80966;
    wire N__80963;
    wire N__80958;
    wire N__80955;
    wire N__80954;
    wire N__80953;
    wire N__80952;
    wire N__80951;
    wire N__80950;
    wire N__80949;
    wire N__80946;
    wire N__80941;
    wire N__80938;
    wire N__80935;
    wire N__80932;
    wire N__80927;
    wire N__80920;
    wire N__80905;
    wire N__80902;
    wire N__80899;
    wire N__80896;
    wire N__80893;
    wire N__80890;
    wire N__80887;
    wire N__80884;
    wire N__80881;
    wire N__80880;
    wire N__80877;
    wire N__80876;
    wire N__80873;
    wire N__80872;
    wire N__80871;
    wire N__80868;
    wire N__80867;
    wire N__80866;
    wire N__80863;
    wire N__80862;
    wire N__80861;
    wire N__80858;
    wire N__80855;
    wire N__80854;
    wire N__80851;
    wire N__80848;
    wire N__80845;
    wire N__80842;
    wire N__80839;
    wire N__80836;
    wire N__80835;
    wire N__80832;
    wire N__80831;
    wire N__80830;
    wire N__80829;
    wire N__80828;
    wire N__80827;
    wire N__80826;
    wire N__80823;
    wire N__80820;
    wire N__80817;
    wire N__80816;
    wire N__80813;
    wire N__80810;
    wire N__80807;
    wire N__80804;
    wire N__80799;
    wire N__80796;
    wire N__80793;
    wire N__80790;
    wire N__80779;
    wire N__80774;
    wire N__80771;
    wire N__80768;
    wire N__80765;
    wire N__80762;
    wire N__80759;
    wire N__80756;
    wire N__80753;
    wire N__80750;
    wire N__80743;
    wire N__80736;
    wire N__80735;
    wire N__80734;
    wire N__80733;
    wire N__80732;
    wire N__80731;
    wire N__80730;
    wire N__80729;
    wire N__80728;
    wire N__80725;
    wire N__80720;
    wire N__80717;
    wire N__80714;
    wire N__80707;
    wire N__80698;
    wire N__80693;
    wire N__80690;
    wire N__80687;
    wire N__80668;
    wire N__80665;
    wire N__80662;
    wire N__80661;
    wire N__80658;
    wire N__80655;
    wire N__80650;
    wire N__80649;
    wire N__80646;
    wire N__80643;
    wire N__80638;
    wire N__80637;
    wire N__80634;
    wire N__80631;
    wire N__80628;
    wire N__80623;
    wire N__80620;
    wire N__80619;
    wire N__80616;
    wire N__80611;
    wire N__80608;
    wire N__80607;
    wire N__80606;
    wire N__80605;
    wire N__80604;
    wire N__80603;
    wire N__80602;
    wire N__80601;
    wire N__80600;
    wire N__80599;
    wire N__80598;
    wire N__80595;
    wire N__80594;
    wire N__80591;
    wire N__80586;
    wire N__80583;
    wire N__80582;
    wire N__80581;
    wire N__80578;
    wire N__80577;
    wire N__80576;
    wire N__80575;
    wire N__80572;
    wire N__80571;
    wire N__80570;
    wire N__80569;
    wire N__80566;
    wire N__80563;
    wire N__80560;
    wire N__80557;
    wire N__80556;
    wire N__80555;
    wire N__80554;
    wire N__80551;
    wire N__80548;
    wire N__80547;
    wire N__80544;
    wire N__80539;
    wire N__80534;
    wire N__80531;
    wire N__80528;
    wire N__80527;
    wire N__80526;
    wire N__80525;
    wire N__80522;
    wire N__80519;
    wire N__80516;
    wire N__80513;
    wire N__80512;
    wire N__80509;
    wire N__80508;
    wire N__80507;
    wire N__80504;
    wire N__80499;
    wire N__80494;
    wire N__80491;
    wire N__80486;
    wire N__80483;
    wire N__80480;
    wire N__80477;
    wire N__80472;
    wire N__80471;
    wire N__80464;
    wire N__80457;
    wire N__80454;
    wire N__80451;
    wire N__80446;
    wire N__80445;
    wire N__80440;
    wire N__80437;
    wire N__80434;
    wire N__80431;
    wire N__80426;
    wire N__80417;
    wire N__80412;
    wire N__80409;
    wire N__80406;
    wire N__80403;
    wire N__80398;
    wire N__80395;
    wire N__80392;
    wire N__80389;
    wire N__80382;
    wire N__80377;
    wire N__80374;
    wire N__80365;
    wire N__80362;
    wire N__80347;
    wire N__80346;
    wire N__80343;
    wire N__80338;
    wire N__80335;
    wire N__80334;
    wire N__80331;
    wire N__80326;
    wire N__80323;
    wire N__80322;
    wire N__80321;
    wire N__80320;
    wire N__80319;
    wire N__80318;
    wire N__80317;
    wire N__80314;
    wire N__80313;
    wire N__80312;
    wire N__80311;
    wire N__80310;
    wire N__80303;
    wire N__80302;
    wire N__80301;
    wire N__80300;
    wire N__80299;
    wire N__80298;
    wire N__80297;
    wire N__80294;
    wire N__80293;
    wire N__80290;
    wire N__80289;
    wire N__80288;
    wire N__80287;
    wire N__80284;
    wire N__80283;
    wire N__80280;
    wire N__80277;
    wire N__80274;
    wire N__80269;
    wire N__80268;
    wire N__80267;
    wire N__80266;
    wire N__80263;
    wire N__80260;
    wire N__80255;
    wire N__80252;
    wire N__80249;
    wire N__80248;
    wire N__80245;
    wire N__80242;
    wire N__80239;
    wire N__80236;
    wire N__80233;
    wire N__80232;
    wire N__80227;
    wire N__80224;
    wire N__80221;
    wire N__80216;
    wire N__80215;
    wire N__80210;
    wire N__80207;
    wire N__80202;
    wire N__80201;
    wire N__80198;
    wire N__80195;
    wire N__80192;
    wire N__80189;
    wire N__80186;
    wire N__80183;
    wire N__80176;
    wire N__80171;
    wire N__80168;
    wire N__80167;
    wire N__80166;
    wire N__80165;
    wire N__80162;
    wire N__80157;
    wire N__80154;
    wire N__80151;
    wire N__80148;
    wire N__80145;
    wire N__80142;
    wire N__80139;
    wire N__80134;
    wire N__80131;
    wire N__80124;
    wire N__80121;
    wire N__80116;
    wire N__80113;
    wire N__80108;
    wire N__80105;
    wire N__80102;
    wire N__80097;
    wire N__80090;
    wire N__80087;
    wire N__80084;
    wire N__80079;
    wire N__80074;
    wire N__80071;
    wire N__80068;
    wire N__80061;
    wire N__80056;
    wire N__80041;
    wire N__80038;
    wire N__80035;
    wire N__80032;
    wire N__80029;
    wire N__80026;
    wire N__80023;
    wire N__80020;
    wire N__80017;
    wire N__80014;
    wire N__80011;
    wire N__80008;
    wire N__80007;
    wire N__80004;
    wire N__79999;
    wire N__79996;
    wire N__79995;
    wire N__79994;
    wire N__79991;
    wire N__79990;
    wire N__79989;
    wire N__79986;
    wire N__79983;
    wire N__79982;
    wire N__79981;
    wire N__79978;
    wire N__79975;
    wire N__79974;
    wire N__79971;
    wire N__79970;
    wire N__79969;
    wire N__79968;
    wire N__79967;
    wire N__79964;
    wire N__79961;
    wire N__79958;
    wire N__79955;
    wire N__79950;
    wire N__79947;
    wire N__79946;
    wire N__79943;
    wire N__79940;
    wire N__79937;
    wire N__79936;
    wire N__79935;
    wire N__79932;
    wire N__79929;
    wire N__79926;
    wire N__79923;
    wire N__79920;
    wire N__79917;
    wire N__79912;
    wire N__79911;
    wire N__79908;
    wire N__79905;
    wire N__79900;
    wire N__79897;
    wire N__79894;
    wire N__79891;
    wire N__79888;
    wire N__79885;
    wire N__79882;
    wire N__79879;
    wire N__79874;
    wire N__79871;
    wire N__79866;
    wire N__79855;
    wire N__79852;
    wire N__79845;
    wire N__79834;
    wire N__79833;
    wire N__79828;
    wire N__79825;
    wire N__79822;
    wire N__79821;
    wire N__79818;
    wire N__79813;
    wire N__79810;
    wire N__79809;
    wire N__79806;
    wire N__79801;
    wire N__79798;
    wire N__79797;
    wire N__79796;
    wire N__79795;
    wire N__79794;
    wire N__79793;
    wire N__79792;
    wire N__79789;
    wire N__79788;
    wire N__79787;
    wire N__79786;
    wire N__79785;
    wire N__79780;
    wire N__79777;
    wire N__79772;
    wire N__79771;
    wire N__79770;
    wire N__79767;
    wire N__79764;
    wire N__79761;
    wire N__79760;
    wire N__79759;
    wire N__79756;
    wire N__79755;
    wire N__79754;
    wire N__79751;
    wire N__79750;
    wire N__79747;
    wire N__79746;
    wire N__79745;
    wire N__79744;
    wire N__79743;
    wire N__79742;
    wire N__79741;
    wire N__79740;
    wire N__79739;
    wire N__79736;
    wire N__79733;
    wire N__79730;
    wire N__79725;
    wire N__79720;
    wire N__79717;
    wire N__79714;
    wire N__79711;
    wire N__79708;
    wire N__79703;
    wire N__79702;
    wire N__79699;
    wire N__79696;
    wire N__79693;
    wire N__79690;
    wire N__79687;
    wire N__79684;
    wire N__79681;
    wire N__79678;
    wire N__79675;
    wire N__79670;
    wire N__79665;
    wire N__79662;
    wire N__79661;
    wire N__79660;
    wire N__79659;
    wire N__79658;
    wire N__79655;
    wire N__79652;
    wire N__79649;
    wire N__79646;
    wire N__79643;
    wire N__79638;
    wire N__79637;
    wire N__79634;
    wire N__79631;
    wire N__79628;
    wire N__79625;
    wire N__79622;
    wire N__79619;
    wire N__79616;
    wire N__79613;
    wire N__79608;
    wire N__79605;
    wire N__79602;
    wire N__79599;
    wire N__79596;
    wire N__79593;
    wire N__79590;
    wire N__79587;
    wire N__79584;
    wire N__79579;
    wire N__79576;
    wire N__79571;
    wire N__79568;
    wire N__79565;
    wire N__79560;
    wire N__79557;
    wire N__79554;
    wire N__79549;
    wire N__79542;
    wire N__79535;
    wire N__79520;
    wire N__79515;
    wire N__79510;
    wire N__79503;
    wire N__79498;
    wire N__79489;
    wire N__79488;
    wire N__79485;
    wire N__79482;
    wire N__79477;
    wire N__79474;
    wire N__79473;
    wire N__79470;
    wire N__79467;
    wire N__79464;
    wire N__79461;
    wire N__79456;
    wire N__79453;
    wire N__79450;
    wire N__79447;
    wire N__79444;
    wire N__79441;
    wire N__79440;
    wire N__79437;
    wire N__79432;
    wire N__79429;
    wire N__79428;
    wire N__79425;
    wire N__79422;
    wire N__79419;
    wire N__79414;
    wire N__79413;
    wire N__79410;
    wire N__79405;
    wire N__79402;
    wire N__79401;
    wire N__79398;
    wire N__79395;
    wire N__79392;
    wire N__79387;
    wire N__79384;
    wire N__79381;
    wire N__79378;
    wire N__79375;
    wire N__79372;
    wire N__79371;
    wire N__79368;
    wire N__79365;
    wire N__79362;
    wire N__79357;
    wire N__79354;
    wire N__79351;
    wire N__79348;
    wire N__79345;
    wire N__79342;
    wire N__79339;
    wire N__79336;
    wire N__79333;
    wire N__79330;
    wire N__79329;
    wire N__79326;
    wire N__79323;
    wire N__79318;
    wire N__79317;
    wire N__79314;
    wire N__79309;
    wire N__79306;
    wire N__79303;
    wire N__79300;
    wire N__79297;
    wire N__79294;
    wire N__79291;
    wire N__79288;
    wire N__79285;
    wire N__79282;
    wire N__79279;
    wire N__79276;
    wire N__79273;
    wire N__79270;
    wire N__79267;
    wire N__79264;
    wire N__79261;
    wire N__79258;
    wire N__79255;
    wire N__79252;
    wire N__79249;
    wire N__79246;
    wire N__79243;
    wire N__79240;
    wire N__79237;
    wire N__79234;
    wire N__79231;
    wire N__79228;
    wire N__79225;
    wire N__79222;
    wire N__79219;
    wire N__79216;
    wire N__79213;
    wire N__79210;
    wire N__79207;
    wire N__79206;
    wire N__79203;
    wire N__79200;
    wire N__79197;
    wire N__79194;
    wire N__79189;
    wire N__79186;
    wire N__79183;
    wire N__79182;
    wire N__79179;
    wire N__79176;
    wire N__79173;
    wire N__79170;
    wire N__79165;
    wire N__79162;
    wire N__79159;
    wire N__79156;
    wire N__79153;
    wire N__79152;
    wire N__79149;
    wire N__79146;
    wire N__79141;
    wire N__79138;
    wire N__79135;
    wire N__79134;
    wire N__79131;
    wire N__79128;
    wire N__79123;
    wire N__79122;
    wire N__79119;
    wire N__79116;
    wire N__79111;
    wire N__79108;
    wire N__79107;
    wire N__79104;
    wire N__79101;
    wire N__79098;
    wire N__79095;
    wire N__79090;
    wire N__79087;
    wire N__79086;
    wire N__79083;
    wire N__79080;
    wire N__79075;
    wire N__79072;
    wire N__79069;
    wire N__79066;
    wire N__79063;
    wire N__79062;
    wire N__79059;
    wire N__79056;
    wire N__79051;
    wire N__79048;
    wire N__79045;
    wire N__79044;
    wire N__79041;
    wire N__79038;
    wire N__79035;
    wire N__79032;
    wire N__79027;
    wire N__79026;
    wire N__79025;
    wire N__79024;
    wire N__79021;
    wire N__79018;
    wire N__79015;
    wire N__79014;
    wire N__79011;
    wire N__79010;
    wire N__79009;
    wire N__79008;
    wire N__79005;
    wire N__79000;
    wire N__78997;
    wire N__78994;
    wire N__78989;
    wire N__78988;
    wire N__78985;
    wire N__78984;
    wire N__78981;
    wire N__78978;
    wire N__78973;
    wire N__78970;
    wire N__78967;
    wire N__78964;
    wire N__78963;
    wire N__78962;
    wire N__78961;
    wire N__78960;
    wire N__78957;
    wire N__78956;
    wire N__78951;
    wire N__78942;
    wire N__78937;
    wire N__78934;
    wire N__78931;
    wire N__78928;
    wire N__78925;
    wire N__78910;
    wire N__78907;
    wire N__78904;
    wire N__78901;
    wire N__78898;
    wire N__78895;
    wire N__78892;
    wire N__78891;
    wire N__78888;
    wire N__78885;
    wire N__78882;
    wire N__78879;
    wire N__78874;
    wire N__78873;
    wire N__78870;
    wire N__78867;
    wire N__78862;
    wire N__78859;
    wire N__78856;
    wire N__78853;
    wire N__78850;
    wire N__78849;
    wire N__78846;
    wire N__78843;
    wire N__78840;
    wire N__78837;
    wire N__78832;
    wire N__78829;
    wire N__78826;
    wire N__78823;
    wire N__78820;
    wire N__78817;
    wire N__78814;
    wire N__78811;
    wire N__78810;
    wire N__78807;
    wire N__78804;
    wire N__78799;
    wire N__78798;
    wire N__78797;
    wire N__78796;
    wire N__78795;
    wire N__78794;
    wire N__78793;
    wire N__78792;
    wire N__78791;
    wire N__78788;
    wire N__78781;
    wire N__78778;
    wire N__78775;
    wire N__78774;
    wire N__78773;
    wire N__78772;
    wire N__78771;
    wire N__78770;
    wire N__78769;
    wire N__78768;
    wire N__78761;
    wire N__78758;
    wire N__78753;
    wire N__78750;
    wire N__78747;
    wire N__78734;
    wire N__78733;
    wire N__78732;
    wire N__78731;
    wire N__78728;
    wire N__78725;
    wire N__78716;
    wire N__78713;
    wire N__78710;
    wire N__78709;
    wire N__78706;
    wire N__78705;
    wire N__78704;
    wire N__78701;
    wire N__78696;
    wire N__78693;
    wire N__78690;
    wire N__78683;
    wire N__78680;
    wire N__78667;
    wire N__78664;
    wire N__78661;
    wire N__78658;
    wire N__78657;
    wire N__78656;
    wire N__78655;
    wire N__78654;
    wire N__78651;
    wire N__78648;
    wire N__78645;
    wire N__78642;
    wire N__78639;
    wire N__78636;
    wire N__78635;
    wire N__78630;
    wire N__78625;
    wire N__78622;
    wire N__78619;
    wire N__78616;
    wire N__78613;
    wire N__78608;
    wire N__78601;
    wire N__78598;
    wire N__78595;
    wire N__78592;
    wire N__78589;
    wire N__78586;
    wire N__78583;
    wire N__78580;
    wire N__78577;
    wire N__78574;
    wire N__78571;
    wire N__78568;
    wire N__78565;
    wire N__78562;
    wire N__78559;
    wire N__78556;
    wire N__78553;
    wire N__78550;
    wire N__78547;
    wire N__78544;
    wire N__78543;
    wire N__78538;
    wire N__78535;
    wire N__78532;
    wire N__78531;
    wire N__78528;
    wire N__78525;
    wire N__78520;
    wire N__78519;
    wire N__78516;
    wire N__78513;
    wire N__78508;
    wire N__78505;
    wire N__78504;
    wire N__78501;
    wire N__78498;
    wire N__78493;
    wire N__78490;
    wire N__78487;
    wire N__78484;
    wire N__78481;
    wire N__78480;
    wire N__78477;
    wire N__78474;
    wire N__78469;
    wire N__78466;
    wire N__78465;
    wire N__78462;
    wire N__78459;
    wire N__78454;
    wire N__78453;
    wire N__78452;
    wire N__78451;
    wire N__78450;
    wire N__78449;
    wire N__78448;
    wire N__78447;
    wire N__78436;
    wire N__78435;
    wire N__78428;
    wire N__78427;
    wire N__78426;
    wire N__78425;
    wire N__78424;
    wire N__78421;
    wire N__78418;
    wire N__78415;
    wire N__78414;
    wire N__78413;
    wire N__78408;
    wire N__78403;
    wire N__78398;
    wire N__78395;
    wire N__78390;
    wire N__78389;
    wire N__78388;
    wire N__78387;
    wire N__78382;
    wire N__78379;
    wire N__78374;
    wire N__78369;
    wire N__78366;
    wire N__78365;
    wire N__78362;
    wire N__78357;
    wire N__78354;
    wire N__78351;
    wire N__78348;
    wire N__78337;
    wire N__78336;
    wire N__78335;
    wire N__78334;
    wire N__78333;
    wire N__78332;
    wire N__78331;
    wire N__78328;
    wire N__78325;
    wire N__78322;
    wire N__78319;
    wire N__78318;
    wire N__78315;
    wire N__78312;
    wire N__78309;
    wire N__78300;
    wire N__78297;
    wire N__78290;
    wire N__78287;
    wire N__78284;
    wire N__78281;
    wire N__78276;
    wire N__78271;
    wire N__78270;
    wire N__78267;
    wire N__78264;
    wire N__78259;
    wire N__78256;
    wire N__78253;
    wire N__78250;
    wire N__78247;
    wire N__78244;
    wire N__78241;
    wire N__78238;
    wire N__78235;
    wire N__78232;
    wire N__78229;
    wire N__78226;
    wire N__78223;
    wire N__78220;
    wire N__78217;
    wire N__78214;
    wire N__78211;
    wire N__78208;
    wire N__78205;
    wire N__78202;
    wire N__78199;
    wire N__78196;
    wire N__78193;
    wire N__78190;
    wire N__78187;
    wire N__78184;
    wire N__78181;
    wire N__78178;
    wire N__78175;
    wire N__78172;
    wire N__78169;
    wire N__78168;
    wire N__78165;
    wire N__78162;
    wire N__78157;
    wire N__78154;
    wire N__78153;
    wire N__78150;
    wire N__78147;
    wire N__78142;
    wire N__78139;
    wire N__78136;
    wire N__78133;
    wire N__78130;
    wire N__78129;
    wire N__78128;
    wire N__78127;
    wire N__78126;
    wire N__78123;
    wire N__78120;
    wire N__78115;
    wire N__78112;
    wire N__78103;
    wire N__78100;
    wire N__78097;
    wire N__78096;
    wire N__78095;
    wire N__78094;
    wire N__78091;
    wire N__78084;
    wire N__78079;
    wire N__78076;
    wire N__78073;
    wire N__78070;
    wire N__78069;
    wire N__78068;
    wire N__78065;
    wire N__78060;
    wire N__78055;
    wire N__78054;
    wire N__78051;
    wire N__78048;
    wire N__78047;
    wire N__78046;
    wire N__78041;
    wire N__78038;
    wire N__78035;
    wire N__78034;
    wire N__78033;
    wire N__78032;
    wire N__78027;
    wire N__78024;
    wire N__78021;
    wire N__78016;
    wire N__78013;
    wire N__78010;
    wire N__78005;
    wire N__77998;
    wire N__77995;
    wire N__77992;
    wire N__77989;
    wire N__77986;
    wire N__77983;
    wire N__77980;
    wire N__77977;
    wire N__77974;
    wire N__77973;
    wire N__77970;
    wire N__77969;
    wire N__77968;
    wire N__77965;
    wire N__77964;
    wire N__77961;
    wire N__77958;
    wire N__77957;
    wire N__77956;
    wire N__77955;
    wire N__77952;
    wire N__77951;
    wire N__77950;
    wire N__77947;
    wire N__77944;
    wire N__77943;
    wire N__77938;
    wire N__77937;
    wire N__77936;
    wire N__77935;
    wire N__77934;
    wire N__77931;
    wire N__77930;
    wire N__77927;
    wire N__77924;
    wire N__77923;
    wire N__77920;
    wire N__77917;
    wire N__77914;
    wire N__77911;
    wire N__77908;
    wire N__77905;
    wire N__77904;
    wire N__77901;
    wire N__77898;
    wire N__77897;
    wire N__77894;
    wire N__77893;
    wire N__77892;
    wire N__77891;
    wire N__77890;
    wire N__77889;
    wire N__77886;
    wire N__77883;
    wire N__77880;
    wire N__77877;
    wire N__77872;
    wire N__77869;
    wire N__77862;
    wire N__77857;
    wire N__77854;
    wire N__77851;
    wire N__77850;
    wire N__77845;
    wire N__77842;
    wire N__77841;
    wire N__77840;
    wire N__77837;
    wire N__77834;
    wire N__77833;
    wire N__77832;
    wire N__77827;
    wire N__77822;
    wire N__77819;
    wire N__77812;
    wire N__77809;
    wire N__77806;
    wire N__77801;
    wire N__77796;
    wire N__77793;
    wire N__77790;
    wire N__77787;
    wire N__77784;
    wire N__77783;
    wire N__77780;
    wire N__77777;
    wire N__77774;
    wire N__77771;
    wire N__77768;
    wire N__77765;
    wire N__77762;
    wire N__77759;
    wire N__77758;
    wire N__77753;
    wire N__77750;
    wire N__77745;
    wire N__77744;
    wire N__77741;
    wire N__77736;
    wire N__77733;
    wire N__77730;
    wire N__77721;
    wire N__77716;
    wire N__77711;
    wire N__77708;
    wire N__77703;
    wire N__77700;
    wire N__77697;
    wire N__77692;
    wire N__77689;
    wire N__77686;
    wire N__77679;
    wire N__77672;
    wire N__77667;
    wire N__77656;
    wire N__77653;
    wire N__77652;
    wire N__77649;
    wire N__77646;
    wire N__77643;
    wire N__77640;
    wire N__77635;
    wire N__77632;
    wire N__77629;
    wire N__77628;
    wire N__77625;
    wire N__77622;
    wire N__77617;
    wire N__77614;
    wire N__77611;
    wire N__77608;
    wire N__77607;
    wire N__77604;
    wire N__77601;
    wire N__77596;
    wire N__77593;
    wire N__77590;
    wire N__77587;
    wire N__77584;
    wire N__77581;
    wire N__77578;
    wire N__77575;
    wire N__77572;
    wire N__77569;
    wire N__77566;
    wire N__77563;
    wire N__77562;
    wire N__77559;
    wire N__77556;
    wire N__77551;
    wire N__77548;
    wire N__77545;
    wire N__77542;
    wire N__77539;
    wire N__77538;
    wire N__77535;
    wire N__77532;
    wire N__77527;
    wire N__77524;
    wire N__77523;
    wire N__77520;
    wire N__77517;
    wire N__77512;
    wire N__77509;
    wire N__77506;
    wire N__77503;
    wire N__77502;
    wire N__77499;
    wire N__77494;
    wire N__77491;
    wire N__77490;
    wire N__77487;
    wire N__77482;
    wire N__77479;
    wire N__77476;
    wire N__77475;
    wire N__77474;
    wire N__77473;
    wire N__77472;
    wire N__77471;
    wire N__77468;
    wire N__77467;
    wire N__77466;
    wire N__77465;
    wire N__77464;
    wire N__77459;
    wire N__77458;
    wire N__77457;
    wire N__77456;
    wire N__77455;
    wire N__77452;
    wire N__77451;
    wire N__77450;
    wire N__77449;
    wire N__77444;
    wire N__77443;
    wire N__77442;
    wire N__77441;
    wire N__77440;
    wire N__77439;
    wire N__77438;
    wire N__77435;
    wire N__77432;
    wire N__77429;
    wire N__77426;
    wire N__77423;
    wire N__77420;
    wire N__77419;
    wire N__77418;
    wire N__77417;
    wire N__77416;
    wire N__77413;
    wire N__77410;
    wire N__77405;
    wire N__77402;
    wire N__77395;
    wire N__77392;
    wire N__77391;
    wire N__77390;
    wire N__77389;
    wire N__77388;
    wire N__77387;
    wire N__77384;
    wire N__77379;
    wire N__77372;
    wire N__77367;
    wire N__77364;
    wire N__77361;
    wire N__77356;
    wire N__77353;
    wire N__77350;
    wire N__77345;
    wire N__77338;
    wire N__77335;
    wire N__77330;
    wire N__77327;
    wire N__77324;
    wire N__77317;
    wire N__77312;
    wire N__77309;
    wire N__77306;
    wire N__77299;
    wire N__77286;
    wire N__77269;
    wire N__77266;
    wire N__77265;
    wire N__77262;
    wire N__77259;
    wire N__77256;
    wire N__77253;
    wire N__77248;
    wire N__77247;
    wire N__77246;
    wire N__77245;
    wire N__77244;
    wire N__77241;
    wire N__77240;
    wire N__77237;
    wire N__77236;
    wire N__77233;
    wire N__77232;
    wire N__77231;
    wire N__77230;
    wire N__77229;
    wire N__77226;
    wire N__77223;
    wire N__77220;
    wire N__77217;
    wire N__77214;
    wire N__77211;
    wire N__77210;
    wire N__77209;
    wire N__77206;
    wire N__77203;
    wire N__77202;
    wire N__77199;
    wire N__77196;
    wire N__77193;
    wire N__77192;
    wire N__77187;
    wire N__77184;
    wire N__77181;
    wire N__77178;
    wire N__77175;
    wire N__77172;
    wire N__77169;
    wire N__77166;
    wire N__77163;
    wire N__77160;
    wire N__77157;
    wire N__77154;
    wire N__77151;
    wire N__77148;
    wire N__77145;
    wire N__77140;
    wire N__77135;
    wire N__77132;
    wire N__77129;
    wire N__77122;
    wire N__77119;
    wire N__77116;
    wire N__77113;
    wire N__77110;
    wire N__77101;
    wire N__77096;
    wire N__77087;
    wire N__77080;
    wire N__77079;
    wire N__77074;
    wire N__77071;
    wire N__77068;
    wire N__77067;
    wire N__77064;
    wire N__77061;
    wire N__77056;
    wire N__77055;
    wire N__77050;
    wire N__77047;
    wire N__77046;
    wire N__77045;
    wire N__77042;
    wire N__77041;
    wire N__77040;
    wire N__77039;
    wire N__77038;
    wire N__77037;
    wire N__77036;
    wire N__77035;
    wire N__77032;
    wire N__77029;
    wire N__77026;
    wire N__77023;
    wire N__77022;
    wire N__77021;
    wire N__77020;
    wire N__77019;
    wire N__77016;
    wire N__77015;
    wire N__77014;
    wire N__77013;
    wire N__77010;
    wire N__77007;
    wire N__77004;
    wire N__77003;
    wire N__77000;
    wire N__76997;
    wire N__76992;
    wire N__76987;
    wire N__76986;
    wire N__76985;
    wire N__76980;
    wire N__76977;
    wire N__76976;
    wire N__76975;
    wire N__76972;
    wire N__76969;
    wire N__76966;
    wire N__76961;
    wire N__76958;
    wire N__76955;
    wire N__76952;
    wire N__76949;
    wire N__76946;
    wire N__76945;
    wire N__76944;
    wire N__76943;
    wire N__76940;
    wire N__76937;
    wire N__76934;
    wire N__76931;
    wire N__76928;
    wire N__76927;
    wire N__76922;
    wire N__76919;
    wire N__76918;
    wire N__76917;
    wire N__76916;
    wire N__76915;
    wire N__76912;
    wire N__76911;
    wire N__76908;
    wire N__76903;
    wire N__76900;
    wire N__76891;
    wire N__76888;
    wire N__76881;
    wire N__76878;
    wire N__76871;
    wire N__76868;
    wire N__76865;
    wire N__76862;
    wire N__76859;
    wire N__76854;
    wire N__76851;
    wire N__76848;
    wire N__76845;
    wire N__76842;
    wire N__76841;
    wire N__76836;
    wire N__76833;
    wire N__76830;
    wire N__76825;
    wire N__76816;
    wire N__76813;
    wire N__76806;
    wire N__76803;
    wire N__76798;
    wire N__76795;
    wire N__76788;
    wire N__76783;
    wire N__76778;
    wire N__76771;
    wire N__76762;
    wire N__76761;
    wire N__76760;
    wire N__76759;
    wire N__76758;
    wire N__76755;
    wire N__76754;
    wire N__76753;
    wire N__76752;
    wire N__76751;
    wire N__76746;
    wire N__76745;
    wire N__76744;
    wire N__76743;
    wire N__76740;
    wire N__76737;
    wire N__76736;
    wire N__76735;
    wire N__76734;
    wire N__76733;
    wire N__76726;
    wire N__76723;
    wire N__76722;
    wire N__76721;
    wire N__76720;
    wire N__76717;
    wire N__76716;
    wire N__76715;
    wire N__76714;
    wire N__76713;
    wire N__76712;
    wire N__76711;
    wire N__76710;
    wire N__76709;
    wire N__76708;
    wire N__76707;
    wire N__76706;
    wire N__76705;
    wire N__76704;
    wire N__76703;
    wire N__76702;
    wire N__76699;
    wire N__76696;
    wire N__76695;
    wire N__76692;
    wire N__76691;
    wire N__76690;
    wire N__76687;
    wire N__76682;
    wire N__76673;
    wire N__76670;
    wire N__76661;
    wire N__76658;
    wire N__76647;
    wire N__76640;
    wire N__76639;
    wire N__76638;
    wire N__76637;
    wire N__76636;
    wire N__76635;
    wire N__76630;
    wire N__76623;
    wire N__76622;
    wire N__76621;
    wire N__76620;
    wire N__76619;
    wire N__76618;
    wire N__76617;
    wire N__76616;
    wire N__76615;
    wire N__76614;
    wire N__76613;
    wire N__76612;
    wire N__76611;
    wire N__76610;
    wire N__76607;
    wire N__76606;
    wire N__76605;
    wire N__76604;
    wire N__76603;
    wire N__76602;
    wire N__76601;
    wire N__76600;
    wire N__76597;
    wire N__76592;
    wire N__76589;
    wire N__76588;
    wire N__76585;
    wire N__76580;
    wire N__76575;
    wire N__76568;
    wire N__76565;
    wire N__76560;
    wire N__76557;
    wire N__76552;
    wire N__76547;
    wire N__76544;
    wire N__76541;
    wire N__76538;
    wire N__76535;
    wire N__76532;
    wire N__76525;
    wire N__76514;
    wire N__76513;
    wire N__76510;
    wire N__76507;
    wire N__76504;
    wire N__76499;
    wire N__76488;
    wire N__76483;
    wire N__76480;
    wire N__76477;
    wire N__76474;
    wire N__76463;
    wire N__76456;
    wire N__76453;
    wire N__76448;
    wire N__76439;
    wire N__76436;
    wire N__76431;
    wire N__76428;
    wire N__76421;
    wire N__76418;
    wire N__76415;
    wire N__76410;
    wire N__76405;
    wire N__76402;
    wire N__76399;
    wire N__76390;
    wire N__76387;
    wire N__76382;
    wire N__76369;
    wire N__76368;
    wire N__76365;
    wire N__76362;
    wire N__76359;
    wire N__76354;
    wire N__76353;
    wire N__76352;
    wire N__76351;
    wire N__76350;
    wire N__76347;
    wire N__76346;
    wire N__76345;
    wire N__76344;
    wire N__76341;
    wire N__76338;
    wire N__76337;
    wire N__76336;
    wire N__76335;
    wire N__76334;
    wire N__76333;
    wire N__76332;
    wire N__76331;
    wire N__76326;
    wire N__76325;
    wire N__76324;
    wire N__76323;
    wire N__76320;
    wire N__76317;
    wire N__76314;
    wire N__76313;
    wire N__76312;
    wire N__76309;
    wire N__76308;
    wire N__76307;
    wire N__76306;
    wire N__76301;
    wire N__76298;
    wire N__76295;
    wire N__76292;
    wire N__76287;
    wire N__76284;
    wire N__76283;
    wire N__76280;
    wire N__76277;
    wire N__76274;
    wire N__76269;
    wire N__76268;
    wire N__76261;
    wire N__76256;
    wire N__76255;
    wire N__76252;
    wire N__76249;
    wire N__76244;
    wire N__76241;
    wire N__76238;
    wire N__76237;
    wire N__76236;
    wire N__76235;
    wire N__76232;
    wire N__76229;
    wire N__76226;
    wire N__76223;
    wire N__76220;
    wire N__76217;
    wire N__76212;
    wire N__76211;
    wire N__76208;
    wire N__76205;
    wire N__76202;
    wire N__76199;
    wire N__76196;
    wire N__76195;
    wire N__76192;
    wire N__76189;
    wire N__76186;
    wire N__76181;
    wire N__76178;
    wire N__76175;
    wire N__76172;
    wire N__76167;
    wire N__76162;
    wire N__76159;
    wire N__76156;
    wire N__76153;
    wire N__76150;
    wire N__76145;
    wire N__76138;
    wire N__76135;
    wire N__76134;
    wire N__76119;
    wire N__76112;
    wire N__76105;
    wire N__76098;
    wire N__76095;
    wire N__76084;
    wire N__76083;
    wire N__76080;
    wire N__76077;
    wire N__76072;
    wire N__76069;
    wire N__76066;
    wire N__76063;
    wire N__76060;
    wire N__76057;
    wire N__76056;
    wire N__76053;
    wire N__76050;
    wire N__76047;
    wire N__76044;
    wire N__76039;
    wire N__76036;
    wire N__76033;
    wire N__76030;
    wire N__76029;
    wire N__76026;
    wire N__76021;
    wire N__76018;
    wire N__76017;
    wire N__76014;
    wire N__76011;
    wire N__76006;
    wire N__76003;
    wire N__76000;
    wire N__75999;
    wire N__75998;
    wire N__75995;
    wire N__75992;
    wire N__75989;
    wire N__75988;
    wire N__75987;
    wire N__75986;
    wire N__75983;
    wire N__75980;
    wire N__75977;
    wire N__75976;
    wire N__75975;
    wire N__75974;
    wire N__75973;
    wire N__75972;
    wire N__75971;
    wire N__75968;
    wire N__75967;
    wire N__75966;
    wire N__75965;
    wire N__75964;
    wire N__75963;
    wire N__75962;
    wire N__75961;
    wire N__75960;
    wire N__75959;
    wire N__75958;
    wire N__75957;
    wire N__75956;
    wire N__75955;
    wire N__75954;
    wire N__75951;
    wire N__75948;
    wire N__75943;
    wire N__75942;
    wire N__75941;
    wire N__75940;
    wire N__75939;
    wire N__75938;
    wire N__75937;
    wire N__75936;
    wire N__75935;
    wire N__75934;
    wire N__75933;
    wire N__75932;
    wire N__75931;
    wire N__75930;
    wire N__75929;
    wire N__75928;
    wire N__75927;
    wire N__75926;
    wire N__75925;
    wire N__75924;
    wire N__75923;
    wire N__75922;
    wire N__75921;
    wire N__75920;
    wire N__75919;
    wire N__75916;
    wire N__75911;
    wire N__75906;
    wire N__75905;
    wire N__75904;
    wire N__75903;
    wire N__75898;
    wire N__75897;
    wire N__75896;
    wire N__75893;
    wire N__75888;
    wire N__75885;
    wire N__75876;
    wire N__75875;
    wire N__75872;
    wire N__75869;
    wire N__75866;
    wire N__75865;
    wire N__75864;
    wire N__75859;
    wire N__75856;
    wire N__75853;
    wire N__75846;
    wire N__75841;
    wire N__75836;
    wire N__75827;
    wire N__75822;
    wire N__75821;
    wire N__75820;
    wire N__75819;
    wire N__75816;
    wire N__75807;
    wire N__75806;
    wire N__75805;
    wire N__75804;
    wire N__75791;
    wire N__75786;
    wire N__75783;
    wire N__75778;
    wire N__75775;
    wire N__75768;
    wire N__75765;
    wire N__75762;
    wire N__75759;
    wire N__75750;
    wire N__75739;
    wire N__75736;
    wire N__75733;
    wire N__75722;
    wire N__75717;
    wire N__75714;
    wire N__75711;
    wire N__75708;
    wire N__75705;
    wire N__75702;
    wire N__75699;
    wire N__75694;
    wire N__75689;
    wire N__75686;
    wire N__75681;
    wire N__75674;
    wire N__75667;
    wire N__75660;
    wire N__75657;
    wire N__75652;
    wire N__75645;
    wire N__75638;
    wire N__75635;
    wire N__75632;
    wire N__75623;
    wire N__75610;
    wire N__75607;
    wire N__75606;
    wire N__75603;
    wire N__75600;
    wire N__75597;
    wire N__75594;
    wire N__75589;
    wire N__75588;
    wire N__75585;
    wire N__75584;
    wire N__75581;
    wire N__75580;
    wire N__75579;
    wire N__75578;
    wire N__75577;
    wire N__75576;
    wire N__75573;
    wire N__75572;
    wire N__75569;
    wire N__75568;
    wire N__75567;
    wire N__75566;
    wire N__75563;
    wire N__75560;
    wire N__75559;
    wire N__75558;
    wire N__75555;
    wire N__75552;
    wire N__75549;
    wire N__75546;
    wire N__75543;
    wire N__75540;
    wire N__75537;
    wire N__75534;
    wire N__75531;
    wire N__75528;
    wire N__75523;
    wire N__75520;
    wire N__75517;
    wire N__75514;
    wire N__75513;
    wire N__75510;
    wire N__75507;
    wire N__75504;
    wire N__75499;
    wire N__75494;
    wire N__75491;
    wire N__75488;
    wire N__75483;
    wire N__75480;
    wire N__75477;
    wire N__75474;
    wire N__75473;
    wire N__75470;
    wire N__75467;
    wire N__75464;
    wire N__75461;
    wire N__75456;
    wire N__75449;
    wire N__75444;
    wire N__75441;
    wire N__75424;
    wire N__75421;
    wire N__75420;
    wire N__75417;
    wire N__75414;
    wire N__75409;
    wire N__75408;
    wire N__75405;
    wire N__75402;
    wire N__75397;
    wire N__75394;
    wire N__75391;
    wire N__75388;
    wire N__75387;
    wire N__75384;
    wire N__75381;
    wire N__75376;
    wire N__75375;
    wire N__75372;
    wire N__75369;
    wire N__75366;
    wire N__75361;
    wire N__75358;
    wire N__75355;
    wire N__75352;
    wire N__75349;
    wire N__75348;
    wire N__75345;
    wire N__75342;
    wire N__75337;
    wire N__75334;
    wire N__75331;
    wire N__75330;
    wire N__75327;
    wire N__75324;
    wire N__75321;
    wire N__75316;
    wire N__75315;
    wire N__75312;
    wire N__75307;
    wire N__75304;
    wire N__75303;
    wire N__75300;
    wire N__75295;
    wire N__75292;
    wire N__75291;
    wire N__75288;
    wire N__75285;
    wire N__75282;
    wire N__75277;
    wire N__75276;
    wire N__75273;
    wire N__75270;
    wire N__75267;
    wire N__75262;
    wire N__75261;
    wire N__75256;
    wire N__75253;
    wire N__75250;
    wire N__75249;
    wire N__75246;
    wire N__75243;
    wire N__75240;
    wire N__75235;
    wire N__75232;
    wire N__75229;
    wire N__75226;
    wire N__75223;
    wire N__75222;
    wire N__75219;
    wire N__75216;
    wire N__75213;
    wire N__75210;
    wire N__75205;
    wire N__75202;
    wire N__75201;
    wire N__75198;
    wire N__75195;
    wire N__75190;
    wire N__75189;
    wire N__75186;
    wire N__75183;
    wire N__75178;
    wire N__75175;
    wire N__75172;
    wire N__75169;
    wire N__75168;
    wire N__75165;
    wire N__75162;
    wire N__75159;
    wire N__75156;
    wire N__75151;
    wire N__75148;
    wire N__75145;
    wire N__75142;
    wire N__75141;
    wire N__75138;
    wire N__75135;
    wire N__75132;
    wire N__75129;
    wire N__75124;
    wire N__75121;
    wire N__75118;
    wire N__75117;
    wire N__75114;
    wire N__75111;
    wire N__75108;
    wire N__75105;
    wire N__75100;
    wire N__75097;
    wire N__75094;
    wire N__75091;
    wire N__75088;
    wire N__75085;
    wire N__75082;
    wire N__75079;
    wire N__75076;
    wire N__75075;
    wire N__75070;
    wire N__75067;
    wire N__75066;
    wire N__75065;
    wire N__75064;
    wire N__75061;
    wire N__75058;
    wire N__75055;
    wire N__75052;
    wire N__75051;
    wire N__75050;
    wire N__75049;
    wire N__75048;
    wire N__75045;
    wire N__75042;
    wire N__75041;
    wire N__75040;
    wire N__75039;
    wire N__75036;
    wire N__75033;
    wire N__75030;
    wire N__75027;
    wire N__75024;
    wire N__75021;
    wire N__75020;
    wire N__75019;
    wire N__75016;
    wire N__75013;
    wire N__75012;
    wire N__75009;
    wire N__75006;
    wire N__75003;
    wire N__75002;
    wire N__74999;
    wire N__74992;
    wire N__74989;
    wire N__74986;
    wire N__74983;
    wire N__74980;
    wire N__74975;
    wire N__74972;
    wire N__74965;
    wire N__74962;
    wire N__74961;
    wire N__74958;
    wire N__74955;
    wire N__74952;
    wire N__74945;
    wire N__74936;
    wire N__74933;
    wire N__74920;
    wire N__74917;
    wire N__74914;
    wire N__74911;
    wire N__74908;
    wire N__74905;
    wire N__74902;
    wire N__74899;
    wire N__74898;
    wire N__74895;
    wire N__74894;
    wire N__74893;
    wire N__74892;
    wire N__74891;
    wire N__74888;
    wire N__74885;
    wire N__74876;
    wire N__74875;
    wire N__74874;
    wire N__74873;
    wire N__74870;
    wire N__74865;
    wire N__74862;
    wire N__74857;
    wire N__74848;
    wire N__74845;
    wire N__74842;
    wire N__74841;
    wire N__74838;
    wire N__74835;
    wire N__74830;
    wire N__74827;
    wire N__74826;
    wire N__74823;
    wire N__74820;
    wire N__74815;
    wire N__74812;
    wire N__74809;
    wire N__74806;
    wire N__74803;
    wire N__74802;
    wire N__74799;
    wire N__74796;
    wire N__74791;
    wire N__74788;
    wire N__74785;
    wire N__74784;
    wire N__74781;
    wire N__74778;
    wire N__74775;
    wire N__74770;
    wire N__74769;
    wire N__74766;
    wire N__74765;
    wire N__74764;
    wire N__74763;
    wire N__74762;
    wire N__74761;
    wire N__74758;
    wire N__74757;
    wire N__74754;
    wire N__74753;
    wire N__74750;
    wire N__74749;
    wire N__74746;
    wire N__74745;
    wire N__74742;
    wire N__74741;
    wire N__74738;
    wire N__74735;
    wire N__74732;
    wire N__74729;
    wire N__74726;
    wire N__74723;
    wire N__74720;
    wire N__74717;
    wire N__74714;
    wire N__74711;
    wire N__74708;
    wire N__74705;
    wire N__74704;
    wire N__74703;
    wire N__74700;
    wire N__74697;
    wire N__74692;
    wire N__74689;
    wire N__74686;
    wire N__74681;
    wire N__74680;
    wire N__74679;
    wire N__74674;
    wire N__74669;
    wire N__74666;
    wire N__74663;
    wire N__74660;
    wire N__74655;
    wire N__74648;
    wire N__74643;
    wire N__74634;
    wire N__74623;
    wire N__74622;
    wire N__74617;
    wire N__74614;
    wire N__74611;
    wire N__74608;
    wire N__74607;
    wire N__74604;
    wire N__74601;
    wire N__74596;
    wire N__74593;
    wire N__74590;
    wire N__74587;
    wire N__74586;
    wire N__74583;
    wire N__74580;
    wire N__74575;
    wire N__74572;
    wire N__74571;
    wire N__74568;
    wire N__74565;
    wire N__74560;
    wire N__74557;
    wire N__74556;
    wire N__74551;
    wire N__74550;
    wire N__74549;
    wire N__74548;
    wire N__74547;
    wire N__74546;
    wire N__74545;
    wire N__74544;
    wire N__74543;
    wire N__74542;
    wire N__74541;
    wire N__74540;
    wire N__74539;
    wire N__74538;
    wire N__74537;
    wire N__74536;
    wire N__74535;
    wire N__74534;
    wire N__74533;
    wire N__74532;
    wire N__74531;
    wire N__74530;
    wire N__74529;
    wire N__74528;
    wire N__74525;
    wire N__74510;
    wire N__74507;
    wire N__74506;
    wire N__74505;
    wire N__74504;
    wire N__74503;
    wire N__74498;
    wire N__74481;
    wire N__74472;
    wire N__74471;
    wire N__74468;
    wire N__74467;
    wire N__74466;
    wire N__74461;
    wire N__74458;
    wire N__74449;
    wire N__74442;
    wire N__74433;
    wire N__74432;
    wire N__74431;
    wire N__74430;
    wire N__74429;
    wire N__74428;
    wire N__74427;
    wire N__74426;
    wire N__74421;
    wire N__74418;
    wire N__74413;
    wire N__74408;
    wire N__74401;
    wire N__74396;
    wire N__74383;
    wire N__74380;
    wire N__74379;
    wire N__74378;
    wire N__74377;
    wire N__74376;
    wire N__74373;
    wire N__74368;
    wire N__74363;
    wire N__74356;
    wire N__74353;
    wire N__74350;
    wire N__74349;
    wire N__74348;
    wire N__74343;
    wire N__74340;
    wire N__74335;
    wire N__74332;
    wire N__74329;
    wire N__74328;
    wire N__74327;
    wire N__74326;
    wire N__74325;
    wire N__74322;
    wire N__74321;
    wire N__74316;
    wire N__74315;
    wire N__74312;
    wire N__74311;
    wire N__74308;
    wire N__74305;
    wire N__74302;
    wire N__74299;
    wire N__74296;
    wire N__74293;
    wire N__74288;
    wire N__74275;
    wire N__74274;
    wire N__74269;
    wire N__74268;
    wire N__74265;
    wire N__74262;
    wire N__74261;
    wire N__74260;
    wire N__74259;
    wire N__74258;
    wire N__74257;
    wire N__74256;
    wire N__74255;
    wire N__74252;
    wire N__74249;
    wire N__74246;
    wire N__74241;
    wire N__74238;
    wire N__74235;
    wire N__74232;
    wire N__74229;
    wire N__74212;
    wire N__74209;
    wire N__74206;
    wire N__74205;
    wire N__74202;
    wire N__74199;
    wire N__74198;
    wire N__74197;
    wire N__74196;
    wire N__74193;
    wire N__74186;
    wire N__74183;
    wire N__74176;
    wire N__74173;
    wire N__74172;
    wire N__74169;
    wire N__74166;
    wire N__74161;
    wire N__74158;
    wire N__74155;
    wire N__74152;
    wire N__74151;
    wire N__74148;
    wire N__74145;
    wire N__74140;
    wire N__74137;
    wire N__74134;
    wire N__74133;
    wire N__74130;
    wire N__74127;
    wire N__74124;
    wire N__74121;
    wire N__74116;
    wire N__74113;
    wire N__74110;
    wire N__74109;
    wire N__74106;
    wire N__74103;
    wire N__74100;
    wire N__74097;
    wire N__74092;
    wire N__74089;
    wire N__74086;
    wire N__74085;
    wire N__74082;
    wire N__74079;
    wire N__74076;
    wire N__74073;
    wire N__74068;
    wire N__74065;
    wire N__74062;
    wire N__74059;
    wire N__74056;
    wire N__74053;
    wire N__74050;
    wire N__74047;
    wire N__74044;
    wire N__74041;
    wire N__74038;
    wire N__74035;
    wire N__74032;
    wire N__74031;
    wire N__74028;
    wire N__74025;
    wire N__74024;
    wire N__74021;
    wire N__74016;
    wire N__74015;
    wire N__74014;
    wire N__74011;
    wire N__74008;
    wire N__74005;
    wire N__74002;
    wire N__73993;
    wire N__73992;
    wire N__73991;
    wire N__73988;
    wire N__73987;
    wire N__73986;
    wire N__73983;
    wire N__73982;
    wire N__73977;
    wire N__73976;
    wire N__73975;
    wire N__73972;
    wire N__73971;
    wire N__73970;
    wire N__73965;
    wire N__73962;
    wire N__73959;
    wire N__73954;
    wire N__73951;
    wire N__73950;
    wire N__73947;
    wire N__73946;
    wire N__73945;
    wire N__73944;
    wire N__73943;
    wire N__73940;
    wire N__73937;
    wire N__73934;
    wire N__73927;
    wire N__73924;
    wire N__73911;
    wire N__73900;
    wire N__73897;
    wire N__73896;
    wire N__73895;
    wire N__73892;
    wire N__73889;
    wire N__73886;
    wire N__73885;
    wire N__73882;
    wire N__73879;
    wire N__73874;
    wire N__73873;
    wire N__73870;
    wire N__73865;
    wire N__73862;
    wire N__73855;
    wire N__73854;
    wire N__73851;
    wire N__73848;
    wire N__73843;
    wire N__73840;
    wire N__73839;
    wire N__73836;
    wire N__73833;
    wire N__73828;
    wire N__73825;
    wire N__73822;
    wire N__73821;
    wire N__73816;
    wire N__73813;
    wire N__73810;
    wire N__73807;
    wire N__73806;
    wire N__73801;
    wire N__73798;
    wire N__73795;
    wire N__73792;
    wire N__73789;
    wire N__73786;
    wire N__73785;
    wire N__73780;
    wire N__73777;
    wire N__73774;
    wire N__73771;
    wire N__73768;
    wire N__73767;
    wire N__73764;
    wire N__73761;
    wire N__73756;
    wire N__73755;
    wire N__73754;
    wire N__73751;
    wire N__73748;
    wire N__73747;
    wire N__73746;
    wire N__73743;
    wire N__73740;
    wire N__73737;
    wire N__73734;
    wire N__73731;
    wire N__73728;
    wire N__73719;
    wire N__73718;
    wire N__73713;
    wire N__73712;
    wire N__73711;
    wire N__73710;
    wire N__73709;
    wire N__73708;
    wire N__73705;
    wire N__73704;
    wire N__73701;
    wire N__73698;
    wire N__73695;
    wire N__73692;
    wire N__73691;
    wire N__73690;
    wire N__73689;
    wire N__73686;
    wire N__73685;
    wire N__73682;
    wire N__73681;
    wire N__73678;
    wire N__73675;
    wire N__73670;
    wire N__73665;
    wire N__73662;
    wire N__73657;
    wire N__73656;
    wire N__73653;
    wire N__73650;
    wire N__73647;
    wire N__73644;
    wire N__73639;
    wire N__73636;
    wire N__73633;
    wire N__73630;
    wire N__73627;
    wire N__73624;
    wire N__73621;
    wire N__73618;
    wire N__73613;
    wire N__73610;
    wire N__73605;
    wire N__73600;
    wire N__73597;
    wire N__73592;
    wire N__73589;
    wire N__73586;
    wire N__73581;
    wire N__73576;
    wire N__73567;
    wire N__73564;
    wire N__73561;
    wire N__73560;
    wire N__73559;
    wire N__73558;
    wire N__73557;
    wire N__73556;
    wire N__73553;
    wire N__73548;
    wire N__73545;
    wire N__73542;
    wire N__73539;
    wire N__73538;
    wire N__73537;
    wire N__73536;
    wire N__73533;
    wire N__73530;
    wire N__73527;
    wire N__73524;
    wire N__73521;
    wire N__73518;
    wire N__73513;
    wire N__73510;
    wire N__73507;
    wire N__73502;
    wire N__73499;
    wire N__73494;
    wire N__73483;
    wire N__73482;
    wire N__73481;
    wire N__73478;
    wire N__73477;
    wire N__73476;
    wire N__73475;
    wire N__73474;
    wire N__73473;
    wire N__73470;
    wire N__73469;
    wire N__73468;
    wire N__73467;
    wire N__73466;
    wire N__73465;
    wire N__73464;
    wire N__73463;
    wire N__73462;
    wire N__73461;
    wire N__73460;
    wire N__73459;
    wire N__73458;
    wire N__73457;
    wire N__73456;
    wire N__73453;
    wire N__73450;
    wire N__73447;
    wire N__73444;
    wire N__73441;
    wire N__73440;
    wire N__73437;
    wire N__73436;
    wire N__73433;
    wire N__73430;
    wire N__73429;
    wire N__73428;
    wire N__73427;
    wire N__73426;
    wire N__73425;
    wire N__73424;
    wire N__73423;
    wire N__73422;
    wire N__73421;
    wire N__73420;
    wire N__73419;
    wire N__73418;
    wire N__73417;
    wire N__73416;
    wire N__73415;
    wire N__73414;
    wire N__73413;
    wire N__73402;
    wire N__73399;
    wire N__73396;
    wire N__73385;
    wire N__73382;
    wire N__73381;
    wire N__73380;
    wire N__73379;
    wire N__73374;
    wire N__73373;
    wire N__73372;
    wire N__73369;
    wire N__73366;
    wire N__73363;
    wire N__73352;
    wire N__73349;
    wire N__73344;
    wire N__73339;
    wire N__73322;
    wire N__73313;
    wire N__73310;
    wire N__73307;
    wire N__73304;
    wire N__73303;
    wire N__73302;
    wire N__73301;
    wire N__73300;
    wire N__73299;
    wire N__73298;
    wire N__73297;
    wire N__73296;
    wire N__73295;
    wire N__73294;
    wire N__73293;
    wire N__73286;
    wire N__73279;
    wire N__73276;
    wire N__73273;
    wire N__73270;
    wire N__73267;
    wire N__73264;
    wire N__73261;
    wire N__73258;
    wire N__73245;
    wire N__73240;
    wire N__73237;
    wire N__73226;
    wire N__73223;
    wire N__73220;
    wire N__73213;
    wire N__73204;
    wire N__73203;
    wire N__73202;
    wire N__73201;
    wire N__73200;
    wire N__73199;
    wire N__73198;
    wire N__73197;
    wire N__73196;
    wire N__73193;
    wire N__73190;
    wire N__73187;
    wire N__73184;
    wire N__73179;
    wire N__73172;
    wire N__73165;
    wire N__73162;
    wire N__73145;
    wire N__73142;
    wire N__73139;
    wire N__73136;
    wire N__73131;
    wire N__73128;
    wire N__73121;
    wire N__73108;
    wire N__73105;
    wire N__73102;
    wire N__73099;
    wire N__73096;
    wire N__73093;
    wire N__73090;
    wire N__73087;
    wire N__73084;
    wire N__73081;
    wire N__73078;
    wire N__73075;
    wire N__73072;
    wire N__73069;
    wire N__73066;
    wire N__73063;
    wire N__73060;
    wire N__73057;
    wire N__73054;
    wire N__73053;
    wire N__73052;
    wire N__73051;
    wire N__73050;
    wire N__73047;
    wire N__73046;
    wire N__73043;
    wire N__73040;
    wire N__73037;
    wire N__73034;
    wire N__73033;
    wire N__73032;
    wire N__73029;
    wire N__73026;
    wire N__73025;
    wire N__73022;
    wire N__73019;
    wire N__73018;
    wire N__73017;
    wire N__73014;
    wire N__73013;
    wire N__73010;
    wire N__73007;
    wire N__73004;
    wire N__73001;
    wire N__72998;
    wire N__72995;
    wire N__72994;
    wire N__72993;
    wire N__72988;
    wire N__72985;
    wire N__72982;
    wire N__72981;
    wire N__72978;
    wire N__72975;
    wire N__72970;
    wire N__72967;
    wire N__72960;
    wire N__72957;
    wire N__72954;
    wire N__72951;
    wire N__72948;
    wire N__72945;
    wire N__72942;
    wire N__72941;
    wire N__72936;
    wire N__72931;
    wire N__72928;
    wire N__72923;
    wire N__72914;
    wire N__72911;
    wire N__72898;
    wire N__72895;
    wire N__72892;
    wire N__72889;
    wire N__72888;
    wire N__72885;
    wire N__72882;
    wire N__72877;
    wire N__72874;
    wire N__72871;
    wire N__72868;
    wire N__72865;
    wire N__72862;
    wire N__72859;
    wire N__72856;
    wire N__72853;
    wire N__72850;
    wire N__72847;
    wire N__72844;
    wire N__72841;
    wire N__72838;
    wire N__72835;
    wire N__72832;
    wire N__72829;
    wire N__72826;
    wire N__72823;
    wire N__72820;
    wire N__72817;
    wire N__72814;
    wire N__72811;
    wire N__72808;
    wire N__72805;
    wire N__72802;
    wire N__72799;
    wire N__72796;
    wire N__72793;
    wire N__72790;
    wire N__72787;
    wire N__72784;
    wire N__72781;
    wire N__72778;
    wire N__72775;
    wire N__72772;
    wire N__72769;
    wire N__72766;
    wire N__72763;
    wire N__72760;
    wire N__72757;
    wire N__72754;
    wire N__72751;
    wire N__72748;
    wire N__72745;
    wire N__72742;
    wire N__72739;
    wire N__72738;
    wire N__72733;
    wire N__72730;
    wire N__72729;
    wire N__72728;
    wire N__72725;
    wire N__72724;
    wire N__72721;
    wire N__72720;
    wire N__72717;
    wire N__72716;
    wire N__72713;
    wire N__72712;
    wire N__72711;
    wire N__72710;
    wire N__72709;
    wire N__72706;
    wire N__72703;
    wire N__72702;
    wire N__72701;
    wire N__72700;
    wire N__72697;
    wire N__72694;
    wire N__72691;
    wire N__72688;
    wire N__72687;
    wire N__72684;
    wire N__72681;
    wire N__72678;
    wire N__72675;
    wire N__72672;
    wire N__72669;
    wire N__72668;
    wire N__72667;
    wire N__72664;
    wire N__72661;
    wire N__72658;
    wire N__72653;
    wire N__72648;
    wire N__72645;
    wire N__72640;
    wire N__72637;
    wire N__72632;
    wire N__72629;
    wire N__72624;
    wire N__72621;
    wire N__72618;
    wire N__72615;
    wire N__72610;
    wire N__72605;
    wire N__72598;
    wire N__72583;
    wire N__72580;
    wire N__72579;
    wire N__72576;
    wire N__72573;
    wire N__72568;
    wire N__72567;
    wire N__72566;
    wire N__72565;
    wire N__72564;
    wire N__72561;
    wire N__72560;
    wire N__72555;
    wire N__72552;
    wire N__72551;
    wire N__72550;
    wire N__72547;
    wire N__72544;
    wire N__72541;
    wire N__72540;
    wire N__72539;
    wire N__72536;
    wire N__72535;
    wire N__72532;
    wire N__72529;
    wire N__72526;
    wire N__72523;
    wire N__72520;
    wire N__72517;
    wire N__72516;
    wire N__72515;
    wire N__72514;
    wire N__72511;
    wire N__72508;
    wire N__72505;
    wire N__72502;
    wire N__72501;
    wire N__72498;
    wire N__72495;
    wire N__72492;
    wire N__72491;
    wire N__72488;
    wire N__72485;
    wire N__72482;
    wire N__72479;
    wire N__72476;
    wire N__72473;
    wire N__72470;
    wire N__72467;
    wire N__72464;
    wire N__72461;
    wire N__72458;
    wire N__72455;
    wire N__72452;
    wire N__72449;
    wire N__72446;
    wire N__72443;
    wire N__72436;
    wire N__72431;
    wire N__72426;
    wire N__72419;
    wire N__72410;
    wire N__72397;
    wire N__72394;
    wire N__72393;
    wire N__72390;
    wire N__72387;
    wire N__72382;
    wire N__72381;
    wire N__72376;
    wire N__72373;
    wire N__72370;
    wire N__72367;
    wire N__72366;
    wire N__72363;
    wire N__72360;
    wire N__72355;
    wire N__72352;
    wire N__72351;
    wire N__72348;
    wire N__72345;
    wire N__72342;
    wire N__72339;
    wire N__72334;
    wire N__72333;
    wire N__72330;
    wire N__72327;
    wire N__72324;
    wire N__72319;
    wire N__72316;
    wire N__72315;
    wire N__72310;
    wire N__72307;
    wire N__72304;
    wire N__72301;
    wire N__72300;
    wire N__72297;
    wire N__72294;
    wire N__72289;
    wire N__72286;
    wire N__72285;
    wire N__72282;
    wire N__72279;
    wire N__72274;
    wire N__72271;
    wire N__72268;
    wire N__72265;
    wire N__72264;
    wire N__72263;
    wire N__72262;
    wire N__72261;
    wire N__72258;
    wire N__72257;
    wire N__72254;
    wire N__72251;
    wire N__72248;
    wire N__72247;
    wire N__72246;
    wire N__72245;
    wire N__72244;
    wire N__72243;
    wire N__72240;
    wire N__72237;
    wire N__72234;
    wire N__72233;
    wire N__72230;
    wire N__72229;
    wire N__72228;
    wire N__72225;
    wire N__72222;
    wire N__72219;
    wire N__72214;
    wire N__72211;
    wire N__72208;
    wire N__72207;
    wire N__72204;
    wire N__72203;
    wire N__72200;
    wire N__72197;
    wire N__72194;
    wire N__72191;
    wire N__72188;
    wire N__72185;
    wire N__72182;
    wire N__72177;
    wire N__72172;
    wire N__72169;
    wire N__72166;
    wire N__72163;
    wire N__72160;
    wire N__72155;
    wire N__72148;
    wire N__72145;
    wire N__72136;
    wire N__72133;
    wire N__72128;
    wire N__72115;
    wire N__72114;
    wire N__72113;
    wire N__72112;
    wire N__72111;
    wire N__72110;
    wire N__72109;
    wire N__72106;
    wire N__72105;
    wire N__72102;
    wire N__72101;
    wire N__72100;
    wire N__72097;
    wire N__72094;
    wire N__72093;
    wire N__72092;
    wire N__72089;
    wire N__72086;
    wire N__72085;
    wire N__72082;
    wire N__72079;
    wire N__72076;
    wire N__72075;
    wire N__72072;
    wire N__72069;
    wire N__72066;
    wire N__72065;
    wire N__72062;
    wire N__72059;
    wire N__72056;
    wire N__72053;
    wire N__72050;
    wire N__72047;
    wire N__72044;
    wire N__72041;
    wire N__72038;
    wire N__72035;
    wire N__72032;
    wire N__72029;
    wire N__72026;
    wire N__72023;
    wire N__72020;
    wire N__72019;
    wire N__72016;
    wire N__72013;
    wire N__72010;
    wire N__72007;
    wire N__72004;
    wire N__71999;
    wire N__71996;
    wire N__71989;
    wire N__71980;
    wire N__71977;
    wire N__71974;
    wire N__71969;
    wire N__71966;
    wire N__71961;
    wire N__71952;
    wire N__71941;
    wire N__71938;
    wire N__71937;
    wire N__71934;
    wire N__71931;
    wire N__71926;
    wire N__71923;
    wire N__71920;
    wire N__71919;
    wire N__71916;
    wire N__71913;
    wire N__71908;
    wire N__71905;
    wire N__71904;
    wire N__71903;
    wire N__71902;
    wire N__71899;
    wire N__71896;
    wire N__71893;
    wire N__71892;
    wire N__71889;
    wire N__71888;
    wire N__71887;
    wire N__71886;
    wire N__71885;
    wire N__71884;
    wire N__71879;
    wire N__71878;
    wire N__71875;
    wire N__71872;
    wire N__71869;
    wire N__71866;
    wire N__71865;
    wire N__71864;
    wire N__71863;
    wire N__71860;
    wire N__71857;
    wire N__71854;
    wire N__71851;
    wire N__71850;
    wire N__71847;
    wire N__71844;
    wire N__71839;
    wire N__71836;
    wire N__71833;
    wire N__71830;
    wire N__71827;
    wire N__71824;
    wire N__71821;
    wire N__71818;
    wire N__71813;
    wire N__71810;
    wire N__71809;
    wire N__71806;
    wire N__71803;
    wire N__71796;
    wire N__71789;
    wire N__71780;
    wire N__71777;
    wire N__71764;
    wire N__71763;
    wire N__71762;
    wire N__71759;
    wire N__71756;
    wire N__71755;
    wire N__71752;
    wire N__71749;
    wire N__71746;
    wire N__71743;
    wire N__71742;
    wire N__71741;
    wire N__71740;
    wire N__71739;
    wire N__71738;
    wire N__71737;
    wire N__71736;
    wire N__71733;
    wire N__71730;
    wire N__71727;
    wire N__71724;
    wire N__71721;
    wire N__71718;
    wire N__71715;
    wire N__71712;
    wire N__71711;
    wire N__71710;
    wire N__71707;
    wire N__71704;
    wire N__71703;
    wire N__71700;
    wire N__71699;
    wire N__71696;
    wire N__71689;
    wire N__71686;
    wire N__71679;
    wire N__71676;
    wire N__71673;
    wire N__71670;
    wire N__71667;
    wire N__71664;
    wire N__71661;
    wire N__71658;
    wire N__71657;
    wire N__71654;
    wire N__71643;
    wire N__71636;
    wire N__71631;
    wire N__71628;
    wire N__71617;
    wire N__71614;
    wire N__71613;
    wire N__71610;
    wire N__71607;
    wire N__71602;
    wire N__71601;
    wire N__71600;
    wire N__71599;
    wire N__71598;
    wire N__71597;
    wire N__71596;
    wire N__71591;
    wire N__71588;
    wire N__71587;
    wire N__71586;
    wire N__71581;
    wire N__71578;
    wire N__71575;
    wire N__71570;
    wire N__71569;
    wire N__71568;
    wire N__71565;
    wire N__71562;
    wire N__71561;
    wire N__71560;
    wire N__71559;
    wire N__71558;
    wire N__71557;
    wire N__71556;
    wire N__71555;
    wire N__71554;
    wire N__71553;
    wire N__71552;
    wire N__71551;
    wire N__71546;
    wire N__71545;
    wire N__71544;
    wire N__71543;
    wire N__71542;
    wire N__71541;
    wire N__71540;
    wire N__71535;
    wire N__71532;
    wire N__71529;
    wire N__71528;
    wire N__71527;
    wire N__71526;
    wire N__71525;
    wire N__71524;
    wire N__71523;
    wire N__71522;
    wire N__71521;
    wire N__71520;
    wire N__71519;
    wire N__71518;
    wire N__71517;
    wire N__71512;
    wire N__71507;
    wire N__71504;
    wire N__71499;
    wire N__71498;
    wire N__71495;
    wire N__71494;
    wire N__71493;
    wire N__71492;
    wire N__71487;
    wire N__71480;
    wire N__71477;
    wire N__71472;
    wire N__71471;
    wire N__71470;
    wire N__71463;
    wire N__71462;
    wire N__71461;
    wire N__71458;
    wire N__71457;
    wire N__71456;
    wire N__71455;
    wire N__71450;
    wire N__71447;
    wire N__71444;
    wire N__71437;
    wire N__71432;
    wire N__71425;
    wire N__71418;
    wire N__71409;
    wire N__71406;
    wire N__71405;
    wire N__71404;
    wire N__71401;
    wire N__71400;
    wire N__71399;
    wire N__71398;
    wire N__71395;
    wire N__71390;
    wire N__71387;
    wire N__71384;
    wire N__71379;
    wire N__71376;
    wire N__71373;
    wire N__71370;
    wire N__71365;
    wire N__71362;
    wire N__71359;
    wire N__71358;
    wire N__71357;
    wire N__71354;
    wire N__71353;
    wire N__71350;
    wire N__71347;
    wire N__71332;
    wire N__71331;
    wire N__71330;
    wire N__71329;
    wire N__71326;
    wire N__71325;
    wire N__71322;
    wire N__71319;
    wire N__71316;
    wire N__71309;
    wire N__71304;
    wire N__71299;
    wire N__71296;
    wire N__71295;
    wire N__71290;
    wire N__71285;
    wire N__71280;
    wire N__71277;
    wire N__71274;
    wire N__71271;
    wire N__71268;
    wire N__71261;
    wire N__71258;
    wire N__71255;
    wire N__71252;
    wire N__71249;
    wire N__71246;
    wire N__71239;
    wire N__71230;
    wire N__71227;
    wire N__71220;
    wire N__71215;
    wire N__71212;
    wire N__71207;
    wire N__71198;
    wire N__71191;
    wire N__71186;
    wire N__71173;
    wire N__71170;
    wire N__71169;
    wire N__71166;
    wire N__71163;
    wire N__71158;
    wire N__71157;
    wire N__71154;
    wire N__71151;
    wire N__71146;
    wire N__71143;
    wire N__71142;
    wire N__71139;
    wire N__71136;
    wire N__71133;
    wire N__71130;
    wire N__71125;
    wire N__71122;
    wire N__71121;
    wire N__71116;
    wire N__71113;
    wire N__71110;
    wire N__71109;
    wire N__71106;
    wire N__71103;
    wire N__71100;
    wire N__71097;
    wire N__71092;
    wire N__71091;
    wire N__71088;
    wire N__71083;
    wire N__71080;
    wire N__71077;
    wire N__71074;
    wire N__71071;
    wire N__71068;
    wire N__71065;
    wire N__71062;
    wire N__71061;
    wire N__71058;
    wire N__71055;
    wire N__71052;
    wire N__71047;
    wire N__71046;
    wire N__71043;
    wire N__71040;
    wire N__71037;
    wire N__71032;
    wire N__71029;
    wire N__71026;
    wire N__71023;
    wire N__71022;
    wire N__71019;
    wire N__71016;
    wire N__71011;
    wire N__71008;
    wire N__71007;
    wire N__71006;
    wire N__71005;
    wire N__71000;
    wire N__70999;
    wire N__70998;
    wire N__70995;
    wire N__70992;
    wire N__70991;
    wire N__70990;
    wire N__70989;
    wire N__70988;
    wire N__70987;
    wire N__70986;
    wire N__70983;
    wire N__70978;
    wire N__70977;
    wire N__70976;
    wire N__70975;
    wire N__70974;
    wire N__70969;
    wire N__70966;
    wire N__70965;
    wire N__70964;
    wire N__70961;
    wire N__70956;
    wire N__70951;
    wire N__70950;
    wire N__70949;
    wire N__70948;
    wire N__70945;
    wire N__70942;
    wire N__70939;
    wire N__70938;
    wire N__70937;
    wire N__70932;
    wire N__70929;
    wire N__70928;
    wire N__70925;
    wire N__70922;
    wire N__70919;
    wire N__70916;
    wire N__70915;
    wire N__70912;
    wire N__70909;
    wire N__70906;
    wire N__70903;
    wire N__70898;
    wire N__70897;
    wire N__70896;
    wire N__70889;
    wire N__70886;
    wire N__70883;
    wire N__70882;
    wire N__70879;
    wire N__70876;
    wire N__70873;
    wire N__70864;
    wire N__70861;
    wire N__70860;
    wire N__70857;
    wire N__70852;
    wire N__70847;
    wire N__70844;
    wire N__70841;
    wire N__70838;
    wire N__70833;
    wire N__70830;
    wire N__70827;
    wire N__70822;
    wire N__70817;
    wire N__70814;
    wire N__70813;
    wire N__70812;
    wire N__70807;
    wire N__70804;
    wire N__70799;
    wire N__70792;
    wire N__70783;
    wire N__70778;
    wire N__70765;
    wire N__70764;
    wire N__70761;
    wire N__70756;
    wire N__70753;
    wire N__70752;
    wire N__70749;
    wire N__70744;
    wire N__70741;
    wire N__70740;
    wire N__70737;
    wire N__70732;
    wire N__70729;
    wire N__70728;
    wire N__70725;
    wire N__70722;
    wire N__70721;
    wire N__70720;
    wire N__70719;
    wire N__70718;
    wire N__70717;
    wire N__70716;
    wire N__70715;
    wire N__70714;
    wire N__70713;
    wire N__70708;
    wire N__70707;
    wire N__70706;
    wire N__70705;
    wire N__70702;
    wire N__70699;
    wire N__70696;
    wire N__70693;
    wire N__70692;
    wire N__70689;
    wire N__70686;
    wire N__70683;
    wire N__70682;
    wire N__70681;
    wire N__70680;
    wire N__70677;
    wire N__70676;
    wire N__70675;
    wire N__70672;
    wire N__70669;
    wire N__70664;
    wire N__70663;
    wire N__70662;
    wire N__70661;
    wire N__70658;
    wire N__70655;
    wire N__70652;
    wire N__70649;
    wire N__70646;
    wire N__70643;
    wire N__70640;
    wire N__70637;
    wire N__70634;
    wire N__70633;
    wire N__70632;
    wire N__70631;
    wire N__70626;
    wire N__70623;
    wire N__70620;
    wire N__70615;
    wire N__70608;
    wire N__70605;
    wire N__70602;
    wire N__70599;
    wire N__70596;
    wire N__70591;
    wire N__70586;
    wire N__70585;
    wire N__70582;
    wire N__70579;
    wire N__70576;
    wire N__70573;
    wire N__70572;
    wire N__70571;
    wire N__70570;
    wire N__70569;
    wire N__70566;
    wire N__70565;
    wire N__70560;
    wire N__70557;
    wire N__70552;
    wire N__70549;
    wire N__70546;
    wire N__70543;
    wire N__70540;
    wire N__70531;
    wire N__70528;
    wire N__70523;
    wire N__70518;
    wire N__70513;
    wire N__70508;
    wire N__70505;
    wire N__70502;
    wire N__70497;
    wire N__70490;
    wire N__70483;
    wire N__70476;
    wire N__70473;
    wire N__70456;
    wire N__70455;
    wire N__70452;
    wire N__70449;
    wire N__70446;
    wire N__70443;
    wire N__70438;
    wire N__70435;
    wire N__70434;
    wire N__70429;
    wire N__70426;
    wire N__70423;
    wire N__70422;
    wire N__70417;
    wire N__70414;
    wire N__70411;
    wire N__70408;
    wire N__70405;
    wire N__70404;
    wire N__70401;
    wire N__70398;
    wire N__70393;
    wire N__70392;
    wire N__70391;
    wire N__70388;
    wire N__70387;
    wire N__70386;
    wire N__70385;
    wire N__70384;
    wire N__70383;
    wire N__70380;
    wire N__70379;
    wire N__70378;
    wire N__70375;
    wire N__70374;
    wire N__70373;
    wire N__70370;
    wire N__70367;
    wire N__70364;
    wire N__70361;
    wire N__70358;
    wire N__70355;
    wire N__70352;
    wire N__70349;
    wire N__70346;
    wire N__70343;
    wire N__70340;
    wire N__70337;
    wire N__70336;
    wire N__70333;
    wire N__70330;
    wire N__70327;
    wire N__70324;
    wire N__70321;
    wire N__70318;
    wire N__70317;
    wire N__70314;
    wire N__70311;
    wire N__70308;
    wire N__70305;
    wire N__70302;
    wire N__70299;
    wire N__70296;
    wire N__70295;
    wire N__70294;
    wire N__70289;
    wire N__70286;
    wire N__70283;
    wire N__70280;
    wire N__70277;
    wire N__70274;
    wire N__70271;
    wire N__70268;
    wire N__70265;
    wire N__70262;
    wire N__70257;
    wire N__70254;
    wire N__70251;
    wire N__70248;
    wire N__70245;
    wire N__70240;
    wire N__70235;
    wire N__70232;
    wire N__70225;
    wire N__70220;
    wire N__70213;
    wire N__70198;
    wire N__70195;
    wire N__70194;
    wire N__70191;
    wire N__70188;
    wire N__70183;
    wire N__70180;
    wire N__70177;
    wire N__70174;
    wire N__70171;
    wire N__70168;
    wire N__70165;
    wire N__70164;
    wire N__70161;
    wire N__70158;
    wire N__70153;
    wire N__70152;
    wire N__70149;
    wire N__70146;
    wire N__70141;
    wire N__70140;
    wire N__70139;
    wire N__70138;
    wire N__70137;
    wire N__70134;
    wire N__70133;
    wire N__70132;
    wire N__70129;
    wire N__70126;
    wire N__70123;
    wire N__70122;
    wire N__70121;
    wire N__70120;
    wire N__70117;
    wire N__70114;
    wire N__70113;
    wire N__70110;
    wire N__70109;
    wire N__70106;
    wire N__70103;
    wire N__70102;
    wire N__70101;
    wire N__70100;
    wire N__70097;
    wire N__70094;
    wire N__70091;
    wire N__70086;
    wire N__70083;
    wire N__70080;
    wire N__70079;
    wire N__70076;
    wire N__70073;
    wire N__70070;
    wire N__70067;
    wire N__70064;
    wire N__70061;
    wire N__70058;
    wire N__70055;
    wire N__70052;
    wire N__70049;
    wire N__70044;
    wire N__70039;
    wire N__70036;
    wire N__70033;
    wire N__70030;
    wire N__70025;
    wire N__70022;
    wire N__70013;
    wire N__70006;
    wire N__69991;
    wire N__69988;
    wire N__69985;
    wire N__69982;
    wire N__69981;
    wire N__69978;
    wire N__69975;
    wire N__69972;
    wire N__69969;
    wire N__69964;
    wire N__69961;
    wire N__69958;
    wire N__69955;
    wire N__69952;
    wire N__69951;
    wire N__69948;
    wire N__69945;
    wire N__69942;
    wire N__69939;
    wire N__69938;
    wire N__69935;
    wire N__69932;
    wire N__69929;
    wire N__69922;
    wire N__69919;
    wire N__69918;
    wire N__69915;
    wire N__69912;
    wire N__69909;
    wire N__69906;
    wire N__69903;
    wire N__69898;
    wire N__69895;
    wire N__69892;
    wire N__69891;
    wire N__69890;
    wire N__69889;
    wire N__69884;
    wire N__69879;
    wire N__69874;
    wire N__69873;
    wire N__69872;
    wire N__69865;
    wire N__69862;
    wire N__69859;
    wire N__69856;
    wire N__69853;
    wire N__69850;
    wire N__69847;
    wire N__69846;
    wire N__69843;
    wire N__69840;
    wire N__69837;
    wire N__69834;
    wire N__69829;
    wire N__69826;
    wire N__69823;
    wire N__69822;
    wire N__69819;
    wire N__69816;
    wire N__69811;
    wire N__69808;
    wire N__69807;
    wire N__69804;
    wire N__69801;
    wire N__69796;
    wire N__69793;
    wire N__69790;
    wire N__69787;
    wire N__69784;
    wire N__69781;
    wire N__69778;
    wire N__69775;
    wire N__69774;
    wire N__69773;
    wire N__69772;
    wire N__69769;
    wire N__69766;
    wire N__69763;
    wire N__69760;
    wire N__69753;
    wire N__69750;
    wire N__69749;
    wire N__69744;
    wire N__69741;
    wire N__69736;
    wire N__69735;
    wire N__69732;
    wire N__69729;
    wire N__69726;
    wire N__69723;
    wire N__69718;
    wire N__69715;
    wire N__69712;
    wire N__69709;
    wire N__69706;
    wire N__69705;
    wire N__69704;
    wire N__69703;
    wire N__69702;
    wire N__69701;
    wire N__69696;
    wire N__69687;
    wire N__69682;
    wire N__69679;
    wire N__69676;
    wire N__69673;
    wire N__69670;
    wire N__69667;
    wire N__69664;
    wire N__69663;
    wire N__69660;
    wire N__69657;
    wire N__69652;
    wire N__69649;
    wire N__69648;
    wire N__69645;
    wire N__69642;
    wire N__69637;
    wire N__69634;
    wire N__69631;
    wire N__69630;
    wire N__69625;
    wire N__69622;
    wire N__69621;
    wire N__69620;
    wire N__69619;
    wire N__69618;
    wire N__69617;
    wire N__69616;
    wire N__69615;
    wire N__69614;
    wire N__69613;
    wire N__69612;
    wire N__69611;
    wire N__69606;
    wire N__69605;
    wire N__69604;
    wire N__69601;
    wire N__69586;
    wire N__69585;
    wire N__69582;
    wire N__69579;
    wire N__69576;
    wire N__69569;
    wire N__69566;
    wire N__69563;
    wire N__69558;
    wire N__69547;
    wire N__69546;
    wire N__69545;
    wire N__69544;
    wire N__69543;
    wire N__69540;
    wire N__69533;
    wire N__69530;
    wire N__69523;
    wire N__69522;
    wire N__69517;
    wire N__69514;
    wire N__69511;
    wire N__69510;
    wire N__69507;
    wire N__69504;
    wire N__69499;
    wire N__69498;
    wire N__69495;
    wire N__69492;
    wire N__69487;
    wire N__69486;
    wire N__69483;
    wire N__69480;
    wire N__69477;
    wire N__69474;
    wire N__69469;
    wire N__69468;
    wire N__69467;
    wire N__69466;
    wire N__69465;
    wire N__69462;
    wire N__69453;
    wire N__69448;
    wire N__69445;
    wire N__69444;
    wire N__69443;
    wire N__69440;
    wire N__69437;
    wire N__69434;
    wire N__69433;
    wire N__69430;
    wire N__69427;
    wire N__69424;
    wire N__69421;
    wire N__69412;
    wire N__69409;
    wire N__69408;
    wire N__69407;
    wire N__69406;
    wire N__69405;
    wire N__69404;
    wire N__69403;
    wire N__69402;
    wire N__69401;
    wire N__69400;
    wire N__69397;
    wire N__69386;
    wire N__69383;
    wire N__69380;
    wire N__69379;
    wire N__69378;
    wire N__69377;
    wire N__69376;
    wire N__69375;
    wire N__69370;
    wire N__69369;
    wire N__69368;
    wire N__69367;
    wire N__69366;
    wire N__69363;
    wire N__69356;
    wire N__69353;
    wire N__69344;
    wire N__69341;
    wire N__69332;
    wire N__69319;
    wire N__69316;
    wire N__69313;
    wire N__69312;
    wire N__69309;
    wire N__69306;
    wire N__69301;
    wire N__69298;
    wire N__69297;
    wire N__69294;
    wire N__69291;
    wire N__69286;
    wire N__69283;
    wire N__69282;
    wire N__69279;
    wire N__69276;
    wire N__69271;
    wire N__69270;
    wire N__69269;
    wire N__69266;
    wire N__69265;
    wire N__69262;
    wire N__69259;
    wire N__69256;
    wire N__69255;
    wire N__69248;
    wire N__69245;
    wire N__69242;
    wire N__69235;
    wire N__69232;
    wire N__69229;
    wire N__69228;
    wire N__69225;
    wire N__69222;
    wire N__69217;
    wire N__69214;
    wire N__69213;
    wire N__69210;
    wire N__69207;
    wire N__69204;
    wire N__69199;
    wire N__69198;
    wire N__69195;
    wire N__69192;
    wire N__69187;
    wire N__69184;
    wire N__69181;
    wire N__69178;
    wire N__69175;
    wire N__69172;
    wire N__69171;
    wire N__69170;
    wire N__69169;
    wire N__69168;
    wire N__69165;
    wire N__69162;
    wire N__69159;
    wire N__69156;
    wire N__69155;
    wire N__69154;
    wire N__69153;
    wire N__69152;
    wire N__69149;
    wire N__69146;
    wire N__69139;
    wire N__69136;
    wire N__69131;
    wire N__69128;
    wire N__69125;
    wire N__69120;
    wire N__69113;
    wire N__69106;
    wire N__69103;
    wire N__69100;
    wire N__69097;
    wire N__69096;
    wire N__69093;
    wire N__69092;
    wire N__69089;
    wire N__69086;
    wire N__69083;
    wire N__69080;
    wire N__69073;
    wire N__69070;
    wire N__69067;
    wire N__69064;
    wire N__69061;
    wire N__69060;
    wire N__69059;
    wire N__69056;
    wire N__69051;
    wire N__69046;
    wire N__69043;
    wire N__69040;
    wire N__69039;
    wire N__69038;
    wire N__69037;
    wire N__69036;
    wire N__69033;
    wire N__69024;
    wire N__69019;
    wire N__69016;
    wire N__69015;
    wire N__69014;
    wire N__69013;
    wire N__69012;
    wire N__69011;
    wire N__69010;
    wire N__69009;
    wire N__68992;
    wire N__68991;
    wire N__68990;
    wire N__68989;
    wire N__68988;
    wire N__68987;
    wire N__68986;
    wire N__68985;
    wire N__68982;
    wire N__68981;
    wire N__68966;
    wire N__68965;
    wire N__68964;
    wire N__68963;
    wire N__68960;
    wire N__68957;
    wire N__68954;
    wire N__68947;
    wire N__68938;
    wire N__68935;
    wire N__68932;
    wire N__68931;
    wire N__68928;
    wire N__68925;
    wire N__68922;
    wire N__68919;
    wire N__68914;
    wire N__68913;
    wire N__68912;
    wire N__68911;
    wire N__68910;
    wire N__68909;
    wire N__68908;
    wire N__68907;
    wire N__68906;
    wire N__68905;
    wire N__68904;
    wire N__68903;
    wire N__68902;
    wire N__68901;
    wire N__68884;
    wire N__68879;
    wire N__68870;
    wire N__68869;
    wire N__68868;
    wire N__68867;
    wire N__68866;
    wire N__68865;
    wire N__68864;
    wire N__68863;
    wire N__68860;
    wire N__68855;
    wire N__68846;
    wire N__68839;
    wire N__68830;
    wire N__68829;
    wire N__68826;
    wire N__68823;
    wire N__68820;
    wire N__68817;
    wire N__68814;
    wire N__68811;
    wire N__68808;
    wire N__68805;
    wire N__68802;
    wire N__68799;
    wire N__68796;
    wire N__68791;
    wire N__68788;
    wire N__68785;
    wire N__68782;
    wire N__68779;
    wire N__68776;
    wire N__68775;
    wire N__68772;
    wire N__68769;
    wire N__68766;
    wire N__68763;
    wire N__68758;
    wire N__68757;
    wire N__68754;
    wire N__68751;
    wire N__68748;
    wire N__68745;
    wire N__68740;
    wire N__68739;
    wire N__68736;
    wire N__68733;
    wire N__68728;
    wire N__68725;
    wire N__68724;
    wire N__68721;
    wire N__68718;
    wire N__68713;
    wire N__68710;
    wire N__68707;
    wire N__68704;
    wire N__68701;
    wire N__68698;
    wire N__68697;
    wire N__68692;
    wire N__68691;
    wire N__68688;
    wire N__68685;
    wire N__68680;
    wire N__68679;
    wire N__68676;
    wire N__68673;
    wire N__68672;
    wire N__68667;
    wire N__68664;
    wire N__68659;
    wire N__68656;
    wire N__68655;
    wire N__68654;
    wire N__68649;
    wire N__68646;
    wire N__68643;
    wire N__68640;
    wire N__68635;
    wire N__68632;
    wire N__68629;
    wire N__68626;
    wire N__68623;
    wire N__68622;
    wire N__68619;
    wire N__68616;
    wire N__68611;
    wire N__68608;
    wire N__68605;
    wire N__68604;
    wire N__68603;
    wire N__68602;
    wire N__68601;
    wire N__68600;
    wire N__68599;
    wire N__68598;
    wire N__68595;
    wire N__68592;
    wire N__68581;
    wire N__68580;
    wire N__68579;
    wire N__68576;
    wire N__68575;
    wire N__68572;
    wire N__68567;
    wire N__68558;
    wire N__68555;
    wire N__68552;
    wire N__68549;
    wire N__68542;
    wire N__68539;
    wire N__68538;
    wire N__68535;
    wire N__68532;
    wire N__68529;
    wire N__68528;
    wire N__68527;
    wire N__68524;
    wire N__68521;
    wire N__68516;
    wire N__68513;
    wire N__68506;
    wire N__68503;
    wire N__68500;
    wire N__68497;
    wire N__68496;
    wire N__68493;
    wire N__68490;
    wire N__68485;
    wire N__68482;
    wire N__68481;
    wire N__68478;
    wire N__68475;
    wire N__68472;
    wire N__68469;
    wire N__68466;
    wire N__68463;
    wire N__68460;
    wire N__68457;
    wire N__68454;
    wire N__68451;
    wire N__68448;
    wire N__68445;
    wire N__68440;
    wire N__68437;
    wire N__68434;
    wire N__68433;
    wire N__68430;
    wire N__68427;
    wire N__68422;
    wire N__68419;
    wire N__68416;
    wire N__68413;
    wire N__68410;
    wire N__68407;
    wire N__68406;
    wire N__68403;
    wire N__68400;
    wire N__68395;
    wire N__68392;
    wire N__68389;
    wire N__68386;
    wire N__68383;
    wire N__68380;
    wire N__68377;
    wire N__68374;
    wire N__68371;
    wire N__68368;
    wire N__68367;
    wire N__68364;
    wire N__68361;
    wire N__68356;
    wire N__68355;
    wire N__68352;
    wire N__68349;
    wire N__68344;
    wire N__68341;
    wire N__68338;
    wire N__68337;
    wire N__68334;
    wire N__68331;
    wire N__68326;
    wire N__68323;
    wire N__68322;
    wire N__68319;
    wire N__68316;
    wire N__68311;
    wire N__68310;
    wire N__68307;
    wire N__68302;
    wire N__68299;
    wire N__68298;
    wire N__68297;
    wire N__68296;
    wire N__68295;
    wire N__68294;
    wire N__68293;
    wire N__68292;
    wire N__68289;
    wire N__68288;
    wire N__68285;
    wire N__68282;
    wire N__68279;
    wire N__68278;
    wire N__68275;
    wire N__68274;
    wire N__68269;
    wire N__68266;
    wire N__68265;
    wire N__68262;
    wire N__68259;
    wire N__68256;
    wire N__68253;
    wire N__68250;
    wire N__68247;
    wire N__68246;
    wire N__68245;
    wire N__68244;
    wire N__68241;
    wire N__68238;
    wire N__68237;
    wire N__68232;
    wire N__68229;
    wire N__68226;
    wire N__68223;
    wire N__68220;
    wire N__68217;
    wire N__68212;
    wire N__68207;
    wire N__68204;
    wire N__68201;
    wire N__68198;
    wire N__68195;
    wire N__68190;
    wire N__68185;
    wire N__68178;
    wire N__68173;
    wire N__68168;
    wire N__68165;
    wire N__68156;
    wire N__68149;
    wire N__68146;
    wire N__68145;
    wire N__68142;
    wire N__68139;
    wire N__68134;
    wire N__68133;
    wire N__68130;
    wire N__68125;
    wire N__68122;
    wire N__68121;
    wire N__68118;
    wire N__68115;
    wire N__68110;
    wire N__68109;
    wire N__68106;
    wire N__68103;
    wire N__68098;
    wire N__68095;
    wire N__68092;
    wire N__68089;
    wire N__68088;
    wire N__68087;
    wire N__68086;
    wire N__68085;
    wire N__68082;
    wire N__68079;
    wire N__68078;
    wire N__68077;
    wire N__68076;
    wire N__68075;
    wire N__68072;
    wire N__68071;
    wire N__68068;
    wire N__68065;
    wire N__68060;
    wire N__68057;
    wire N__68054;
    wire N__68051;
    wire N__68050;
    wire N__68049;
    wire N__68046;
    wire N__68045;
    wire N__68042;
    wire N__68039;
    wire N__68038;
    wire N__68035;
    wire N__68034;
    wire N__68031;
    wire N__68026;
    wire N__68023;
    wire N__68020;
    wire N__68015;
    wire N__68012;
    wire N__68009;
    wire N__68004;
    wire N__68001;
    wire N__68000;
    wire N__67997;
    wire N__67994;
    wire N__67991;
    wire N__67988;
    wire N__67985;
    wire N__67980;
    wire N__67977;
    wire N__67974;
    wire N__67969;
    wire N__67966;
    wire N__67961;
    wire N__67952;
    wire N__67947;
    wire N__67940;
    wire N__67933;
    wire N__67930;
    wire N__67927;
    wire N__67924;
    wire N__67921;
    wire N__67918;
    wire N__67915;
    wire N__67912;
    wire N__67909;
    wire N__67906;
    wire N__67903;
    wire N__67900;
    wire N__67897;
    wire N__67894;
    wire N__67891;
    wire N__67888;
    wire N__67887;
    wire N__67884;
    wire N__67883;
    wire N__67880;
    wire N__67879;
    wire N__67876;
    wire N__67875;
    wire N__67874;
    wire N__67873;
    wire N__67870;
    wire N__67869;
    wire N__67868;
    wire N__67865;
    wire N__67864;
    wire N__67861;
    wire N__67858;
    wire N__67855;
    wire N__67854;
    wire N__67851;
    wire N__67848;
    wire N__67847;
    wire N__67846;
    wire N__67843;
    wire N__67840;
    wire N__67837;
    wire N__67834;
    wire N__67831;
    wire N__67828;
    wire N__67823;
    wire N__67820;
    wire N__67815;
    wire N__67812;
    wire N__67809;
    wire N__67804;
    wire N__67801;
    wire N__67800;
    wire N__67799;
    wire N__67798;
    wire N__67795;
    wire N__67792;
    wire N__67789;
    wire N__67786;
    wire N__67783;
    wire N__67776;
    wire N__67771;
    wire N__67768;
    wire N__67765;
    wire N__67762;
    wire N__67741;
    wire N__67740;
    wire N__67737;
    wire N__67732;
    wire N__67729;
    wire N__67728;
    wire N__67725;
    wire N__67720;
    wire N__67717;
    wire N__67716;
    wire N__67715;
    wire N__67714;
    wire N__67711;
    wire N__67708;
    wire N__67707;
    wire N__67704;
    wire N__67701;
    wire N__67700;
    wire N__67697;
    wire N__67696;
    wire N__67693;
    wire N__67690;
    wire N__67687;
    wire N__67684;
    wire N__67681;
    wire N__67678;
    wire N__67675;
    wire N__67674;
    wire N__67673;
    wire N__67672;
    wire N__67671;
    wire N__67670;
    wire N__67669;
    wire N__67668;
    wire N__67667;
    wire N__67664;
    wire N__67661;
    wire N__67658;
    wire N__67653;
    wire N__67650;
    wire N__67647;
    wire N__67644;
    wire N__67641;
    wire N__67638;
    wire N__67633;
    wire N__67630;
    wire N__67627;
    wire N__67624;
    wire N__67623;
    wire N__67618;
    wire N__67613;
    wire N__67608;
    wire N__67603;
    wire N__67594;
    wire N__67591;
    wire N__67588;
    wire N__67573;
    wire N__67572;
    wire N__67569;
    wire N__67566;
    wire N__67561;
    wire N__67558;
    wire N__67557;
    wire N__67554;
    wire N__67551;
    wire N__67546;
    wire N__67543;
    wire N__67542;
    wire N__67537;
    wire N__67534;
    wire N__67531;
    wire N__67528;
    wire N__67525;
    wire N__67524;
    wire N__67521;
    wire N__67518;
    wire N__67513;
    wire N__67512;
    wire N__67511;
    wire N__67510;
    wire N__67509;
    wire N__67506;
    wire N__67505;
    wire N__67504;
    wire N__67503;
    wire N__67500;
    wire N__67499;
    wire N__67496;
    wire N__67493;
    wire N__67492;
    wire N__67491;
    wire N__67490;
    wire N__67487;
    wire N__67486;
    wire N__67483;
    wire N__67480;
    wire N__67477;
    wire N__67474;
    wire N__67471;
    wire N__67468;
    wire N__67467;
    wire N__67464;
    wire N__67461;
    wire N__67460;
    wire N__67455;
    wire N__67452;
    wire N__67449;
    wire N__67446;
    wire N__67441;
    wire N__67438;
    wire N__67435;
    wire N__67430;
    wire N__67427;
    wire N__67422;
    wire N__67421;
    wire N__67418;
    wire N__67415;
    wire N__67412;
    wire N__67409;
    wire N__67404;
    wire N__67401;
    wire N__67398;
    wire N__67395;
    wire N__67390;
    wire N__67387;
    wire N__67384;
    wire N__67381;
    wire N__67372;
    wire N__67365;
    wire N__67354;
    wire N__67353;
    wire N__67348;
    wire N__67345;
    wire N__67344;
    wire N__67341;
    wire N__67340;
    wire N__67339;
    wire N__67338;
    wire N__67337;
    wire N__67336;
    wire N__67333;
    wire N__67330;
    wire N__67327;
    wire N__67326;
    wire N__67323;
    wire N__67322;
    wire N__67319;
    wire N__67316;
    wire N__67313;
    wire N__67312;
    wire N__67311;
    wire N__67308;
    wire N__67305;
    wire N__67302;
    wire N__67301;
    wire N__67298;
    wire N__67295;
    wire N__67292;
    wire N__67285;
    wire N__67282;
    wire N__67279;
    wire N__67278;
    wire N__67275;
    wire N__67270;
    wire N__67267;
    wire N__67266;
    wire N__67263;
    wire N__67260;
    wire N__67257;
    wire N__67250;
    wire N__67247;
    wire N__67240;
    wire N__67237;
    wire N__67236;
    wire N__67235;
    wire N__67232;
    wire N__67227;
    wire N__67224;
    wire N__67217;
    wire N__67214;
    wire N__67211;
    wire N__67198;
    wire N__67197;
    wire N__67196;
    wire N__67195;
    wire N__67194;
    wire N__67193;
    wire N__67192;
    wire N__67189;
    wire N__67188;
    wire N__67187;
    wire N__67184;
    wire N__67179;
    wire N__67176;
    wire N__67173;
    wire N__67170;
    wire N__67167;
    wire N__67164;
    wire N__67163;
    wire N__67160;
    wire N__67157;
    wire N__67156;
    wire N__67155;
    wire N__67154;
    wire N__67153;
    wire N__67150;
    wire N__67147;
    wire N__67142;
    wire N__67137;
    wire N__67134;
    wire N__67133;
    wire N__67130;
    wire N__67127;
    wire N__67124;
    wire N__67121;
    wire N__67118;
    wire N__67115;
    wire N__67110;
    wire N__67107;
    wire N__67102;
    wire N__67099;
    wire N__67098;
    wire N__67095;
    wire N__67090;
    wire N__67087;
    wire N__67082;
    wire N__67073;
    wire N__67070;
    wire N__67057;
    wire N__67056;
    wire N__67053;
    wire N__67050;
    wire N__67045;
    wire N__67042;
    wire N__67039;
    wire N__67036;
    wire N__67033;
    wire N__67032;
    wire N__67029;
    wire N__67026;
    wire N__67021;
    wire N__67018;
    wire N__67015;
    wire N__67012;
    wire N__67009;
    wire N__67006;
    wire N__67003;
    wire N__67000;
    wire N__66997;
    wire N__66996;
    wire N__66995;
    wire N__66992;
    wire N__66989;
    wire N__66986;
    wire N__66985;
    wire N__66984;
    wire N__66981;
    wire N__66980;
    wire N__66979;
    wire N__66978;
    wire N__66975;
    wire N__66974;
    wire N__66973;
    wire N__66972;
    wire N__66971;
    wire N__66968;
    wire N__66965;
    wire N__66962;
    wire N__66961;
    wire N__66960;
    wire N__66959;
    wire N__66956;
    wire N__66953;
    wire N__66948;
    wire N__66945;
    wire N__66942;
    wire N__66939;
    wire N__66934;
    wire N__66931;
    wire N__66928;
    wire N__66925;
    wire N__66922;
    wire N__66919;
    wire N__66916;
    wire N__66915;
    wire N__66910;
    wire N__66907;
    wire N__66904;
    wire N__66901;
    wire N__66898;
    wire N__66895;
    wire N__66890;
    wire N__66887;
    wire N__66882;
    wire N__66879;
    wire N__66876;
    wire N__66871;
    wire N__66864;
    wire N__66861;
    wire N__66854;
    wire N__66849;
    wire N__66838;
    wire N__66837;
    wire N__66832;
    wire N__66829;
    wire N__66828;
    wire N__66827;
    wire N__66826;
    wire N__66825;
    wire N__66822;
    wire N__66819;
    wire N__66818;
    wire N__66817;
    wire N__66816;
    wire N__66813;
    wire N__66812;
    wire N__66809;
    wire N__66808;
    wire N__66805;
    wire N__66804;
    wire N__66803;
    wire N__66802;
    wire N__66799;
    wire N__66796;
    wire N__66793;
    wire N__66790;
    wire N__66787;
    wire N__66784;
    wire N__66781;
    wire N__66778;
    wire N__66775;
    wire N__66772;
    wire N__66769;
    wire N__66766;
    wire N__66763;
    wire N__66762;
    wire N__66761;
    wire N__66758;
    wire N__66755;
    wire N__66750;
    wire N__66747;
    wire N__66742;
    wire N__66739;
    wire N__66736;
    wire N__66733;
    wire N__66730;
    wire N__66727;
    wire N__66724;
    wire N__66721;
    wire N__66718;
    wire N__66717;
    wire N__66710;
    wire N__66705;
    wire N__66700;
    wire N__66691;
    wire N__66688;
    wire N__66685;
    wire N__66682;
    wire N__66667;
    wire N__66666;
    wire N__66661;
    wire N__66658;
    wire N__66655;
    wire N__66652;
    wire N__66649;
    wire N__66648;
    wire N__66645;
    wire N__66642;
    wire N__66637;
    wire N__66636;
    wire N__66633;
    wire N__66630;
    wire N__66625;
    wire N__66622;
    wire N__66619;
    wire N__66616;
    wire N__66615;
    wire N__66612;
    wire N__66609;
    wire N__66604;
    wire N__66603;
    wire N__66598;
    wire N__66595;
    wire N__66592;
    wire N__66589;
    wire N__66588;
    wire N__66587;
    wire N__66586;
    wire N__66583;
    wire N__66582;
    wire N__66581;
    wire N__66580;
    wire N__66579;
    wire N__66578;
    wire N__66577;
    wire N__66574;
    wire N__66573;
    wire N__66570;
    wire N__66567;
    wire N__66566;
    wire N__66563;
    wire N__66560;
    wire N__66557;
    wire N__66554;
    wire N__66551;
    wire N__66548;
    wire N__66545;
    wire N__66542;
    wire N__66539;
    wire N__66534;
    wire N__66531;
    wire N__66530;
    wire N__66529;
    wire N__66526;
    wire N__66523;
    wire N__66520;
    wire N__66517;
    wire N__66514;
    wire N__66511;
    wire N__66508;
    wire N__66505;
    wire N__66502;
    wire N__66497;
    wire N__66494;
    wire N__66491;
    wire N__66490;
    wire N__66489;
    wire N__66486;
    wire N__66483;
    wire N__66480;
    wire N__66477;
    wire N__66474;
    wire N__66469;
    wire N__66462;
    wire N__66457;
    wire N__66454;
    wire N__66451;
    wire N__66430;
    wire N__66429;
    wire N__66426;
    wire N__66425;
    wire N__66424;
    wire N__66423;
    wire N__66422;
    wire N__66421;
    wire N__66420;
    wire N__66417;
    wire N__66416;
    wire N__66415;
    wire N__66414;
    wire N__66413;
    wire N__66412;
    wire N__66409;
    wire N__66406;
    wire N__66403;
    wire N__66402;
    wire N__66399;
    wire N__66396;
    wire N__66391;
    wire N__66388;
    wire N__66387;
    wire N__66384;
    wire N__66381;
    wire N__66376;
    wire N__66373;
    wire N__66370;
    wire N__66367;
    wire N__66364;
    wire N__66361;
    wire N__66358;
    wire N__66355;
    wire N__66352;
    wire N__66349;
    wire N__66348;
    wire N__66345;
    wire N__66342;
    wire N__66339;
    wire N__66336;
    wire N__66333;
    wire N__66328;
    wire N__66325;
    wire N__66320;
    wire N__66313;
    wire N__66310;
    wire N__66307;
    wire N__66304;
    wire N__66301;
    wire N__66298;
    wire N__66287;
    wire N__66274;
    wire N__66271;
    wire N__66270;
    wire N__66269;
    wire N__66268;
    wire N__66267;
    wire N__66266;
    wire N__66263;
    wire N__66260;
    wire N__66259;
    wire N__66256;
    wire N__66255;
    wire N__66252;
    wire N__66251;
    wire N__66250;
    wire N__66247;
    wire N__66244;
    wire N__66239;
    wire N__66236;
    wire N__66233;
    wire N__66230;
    wire N__66227;
    wire N__66224;
    wire N__66221;
    wire N__66220;
    wire N__66219;
    wire N__66218;
    wire N__66215;
    wire N__66212;
    wire N__66209;
    wire N__66206;
    wire N__66203;
    wire N__66200;
    wire N__66197;
    wire N__66194;
    wire N__66191;
    wire N__66184;
    wire N__66183;
    wire N__66182;
    wire N__66181;
    wire N__66178;
    wire N__66175;
    wire N__66172;
    wire N__66169;
    wire N__66164;
    wire N__66155;
    wire N__66152;
    wire N__66147;
    wire N__66130;
    wire N__66127;
    wire N__66126;
    wire N__66123;
    wire N__66120;
    wire N__66117;
    wire N__66114;
    wire N__66109;
    wire N__66106;
    wire N__66103;
    wire N__66100;
    wire N__66097;
    wire N__66094;
    wire N__66091;
    wire N__66088;
    wire N__66087;
    wire N__66082;
    wire N__66079;
    wire N__66076;
    wire N__66073;
    wire N__66072;
    wire N__66069;
    wire N__66066;
    wire N__66061;
    wire N__66058;
    wire N__66057;
    wire N__66054;
    wire N__66051;
    wire N__66046;
    wire N__66045;
    wire N__66042;
    wire N__66039;
    wire N__66036;
    wire N__66033;
    wire N__66028;
    wire N__66027;
    wire N__66026;
    wire N__66023;
    wire N__66022;
    wire N__66021;
    wire N__66018;
    wire N__66017;
    wire N__66016;
    wire N__66015;
    wire N__66012;
    wire N__66009;
    wire N__66008;
    wire N__66007;
    wire N__66006;
    wire N__66005;
    wire N__66004;
    wire N__66003;
    wire N__66000;
    wire N__65997;
    wire N__65994;
    wire N__65993;
    wire N__65990;
    wire N__65985;
    wire N__65980;
    wire N__65979;
    wire N__65976;
    wire N__65973;
    wire N__65970;
    wire N__65967;
    wire N__65964;
    wire N__65961;
    wire N__65954;
    wire N__65951;
    wire N__65948;
    wire N__65943;
    wire N__65940;
    wire N__65935;
    wire N__65932;
    wire N__65927;
    wire N__65922;
    wire N__65915;
    wire N__65902;
    wire N__65901;
    wire N__65898;
    wire N__65897;
    wire N__65896;
    wire N__65893;
    wire N__65892;
    wire N__65889;
    wire N__65888;
    wire N__65887;
    wire N__65884;
    wire N__65881;
    wire N__65880;
    wire N__65879;
    wire N__65878;
    wire N__65877;
    wire N__65876;
    wire N__65873;
    wire N__65870;
    wire N__65867;
    wire N__65864;
    wire N__65861;
    wire N__65860;
    wire N__65855;
    wire N__65852;
    wire N__65849;
    wire N__65846;
    wire N__65843;
    wire N__65840;
    wire N__65839;
    wire N__65836;
    wire N__65833;
    wire N__65830;
    wire N__65825;
    wire N__65822;
    wire N__65815;
    wire N__65808;
    wire N__65805;
    wire N__65804;
    wire N__65803;
    wire N__65798;
    wire N__65793;
    wire N__65790;
    wire N__65783;
    wire N__65780;
    wire N__65777;
    wire N__65764;
    wire N__65761;
    wire N__65758;
    wire N__65755;
    wire N__65752;
    wire N__65749;
    wire N__65746;
    wire N__65743;
    wire N__65740;
    wire N__65737;
    wire N__65734;
    wire N__65731;
    wire N__65728;
    wire N__65725;
    wire N__65722;
    wire N__65719;
    wire N__65716;
    wire N__65713;
    wire N__65710;
    wire N__65707;
    wire N__65704;
    wire N__65703;
    wire N__65698;
    wire N__65695;
    wire N__65692;
    wire N__65689;
    wire N__65688;
    wire N__65687;
    wire N__65686;
    wire N__65685;
    wire N__65682;
    wire N__65679;
    wire N__65678;
    wire N__65677;
    wire N__65676;
    wire N__65673;
    wire N__65670;
    wire N__65669;
    wire N__65666;
    wire N__65665;
    wire N__65664;
    wire N__65659;
    wire N__65654;
    wire N__65651;
    wire N__65650;
    wire N__65647;
    wire N__65644;
    wire N__65641;
    wire N__65640;
    wire N__65637;
    wire N__65634;
    wire N__65631;
    wire N__65628;
    wire N__65625;
    wire N__65622;
    wire N__65619;
    wire N__65618;
    wire N__65615;
    wire N__65612;
    wire N__65609;
    wire N__65606;
    wire N__65605;
    wire N__65604;
    wire N__65601;
    wire N__65596;
    wire N__65587;
    wire N__65584;
    wire N__65575;
    wire N__65572;
    wire N__65569;
    wire N__65554;
    wire N__65553;
    wire N__65548;
    wire N__65545;
    wire N__65544;
    wire N__65539;
    wire N__65536;
    wire N__65533;
    wire N__65532;
    wire N__65529;
    wire N__65526;
    wire N__65523;
    wire N__65520;
    wire N__65515;
    wire N__65512;
    wire N__65509;
    wire N__65508;
    wire N__65505;
    wire N__65502;
    wire N__65499;
    wire N__65496;
    wire N__65493;
    wire N__65490;
    wire N__65485;
    wire N__65482;
    wire N__65479;
    wire N__65476;
    wire N__65475;
    wire N__65472;
    wire N__65469;
    wire N__65464;
    wire N__65461;
    wire N__65458;
    wire N__65457;
    wire N__65454;
    wire N__65451;
    wire N__65448;
    wire N__65445;
    wire N__65442;
    wire N__65439;
    wire N__65434;
    wire N__65431;
    wire N__65428;
    wire N__65425;
    wire N__65424;
    wire N__65421;
    wire N__65418;
    wire N__65413;
    wire N__65412;
    wire N__65409;
    wire N__65406;
    wire N__65403;
    wire N__65400;
    wire N__65397;
    wire N__65394;
    wire N__65391;
    wire N__65388;
    wire N__65385;
    wire N__65380;
    wire N__65377;
    wire N__65374;
    wire N__65373;
    wire N__65370;
    wire N__65367;
    wire N__65362;
    wire N__65359;
    wire N__65358;
    wire N__65355;
    wire N__65352;
    wire N__65349;
    wire N__65346;
    wire N__65343;
    wire N__65340;
    wire N__65335;
    wire N__65332;
    wire N__65329;
    wire N__65328;
    wire N__65325;
    wire N__65322;
    wire N__65317;
    wire N__65314;
    wire N__65313;
    wire N__65310;
    wire N__65307;
    wire N__65304;
    wire N__65301;
    wire N__65298;
    wire N__65295;
    wire N__65292;
    wire N__65287;
    wire N__65284;
    wire N__65283;
    wire N__65278;
    wire N__65275;
    wire N__65272;
    wire N__65269;
    wire N__65266;
    wire N__65263;
    wire N__65260;
    wire N__65259;
    wire N__65258;
    wire N__65251;
    wire N__65248;
    wire N__65247;
    wire N__65246;
    wire N__65243;
    wire N__65240;
    wire N__65237;
    wire N__65230;
    wire N__65227;
    wire N__65226;
    wire N__65225;
    wire N__65224;
    wire N__65223;
    wire N__65222;
    wire N__65221;
    wire N__65220;
    wire N__65217;
    wire N__65210;
    wire N__65207;
    wire N__65202;
    wire N__65199;
    wire N__65196;
    wire N__65191;
    wire N__65186;
    wire N__65183;
    wire N__65180;
    wire N__65177;
    wire N__65174;
    wire N__65171;
    wire N__65168;
    wire N__65161;
    wire N__65160;
    wire N__65159;
    wire N__65158;
    wire N__65157;
    wire N__65156;
    wire N__65155;
    wire N__65154;
    wire N__65151;
    wire N__65148;
    wire N__65141;
    wire N__65134;
    wire N__65131;
    wire N__65124;
    wire N__65121;
    wire N__65118;
    wire N__65113;
    wire N__65110;
    wire N__65109;
    wire N__65108;
    wire N__65105;
    wire N__65100;
    wire N__65095;
    wire N__65092;
    wire N__65089;
    wire N__65088;
    wire N__65085;
    wire N__65082;
    wire N__65077;
    wire N__65074;
    wire N__65073;
    wire N__65070;
    wire N__65067;
    wire N__65064;
    wire N__65061;
    wire N__65056;
    wire N__65053;
    wire N__65050;
    wire N__65047;
    wire N__65044;
    wire N__65043;
    wire N__65040;
    wire N__65037;
    wire N__65034;
    wire N__65031;
    wire N__65026;
    wire N__65023;
    wire N__65020;
    wire N__65019;
    wire N__65016;
    wire N__65013;
    wire N__65008;
    wire N__65005;
    wire N__65002;
    wire N__64999;
    wire N__64996;
    wire N__64993;
    wire N__64990;
    wire N__64989;
    wire N__64986;
    wire N__64983;
    wire N__64980;
    wire N__64977;
    wire N__64972;
    wire N__64969;
    wire N__64968;
    wire N__64965;
    wire N__64962;
    wire N__64957;
    wire N__64954;
    wire N__64951;
    wire N__64948;
    wire N__64945;
    wire N__64942;
    wire N__64941;
    wire N__64940;
    wire N__64937;
    wire N__64932;
    wire N__64927;
    wire N__64924;
    wire N__64921;
    wire N__64920;
    wire N__64917;
    wire N__64914;
    wire N__64909;
    wire N__64906;
    wire N__64905;
    wire N__64902;
    wire N__64899;
    wire N__64894;
    wire N__64893;
    wire N__64888;
    wire N__64885;
    wire N__64884;
    wire N__64883;
    wire N__64878;
    wire N__64875;
    wire N__64870;
    wire N__64869;
    wire N__64866;
    wire N__64865;
    wire N__64864;
    wire N__64861;
    wire N__64860;
    wire N__64851;
    wire N__64848;
    wire N__64843;
    wire N__64840;
    wire N__64839;
    wire N__64836;
    wire N__64833;
    wire N__64830;
    wire N__64825;
    wire N__64822;
    wire N__64821;
    wire N__64818;
    wire N__64815;
    wire N__64812;
    wire N__64807;
    wire N__64804;
    wire N__64801;
    wire N__64798;
    wire N__64797;
    wire N__64794;
    wire N__64791;
    wire N__64786;
    wire N__64783;
    wire N__64780;
    wire N__64779;
    wire N__64776;
    wire N__64773;
    wire N__64768;
    wire N__64767;
    wire N__64764;
    wire N__64761;
    wire N__64756;
    wire N__64755;
    wire N__64752;
    wire N__64749;
    wire N__64746;
    wire N__64741;
    wire N__64740;
    wire N__64739;
    wire N__64732;
    wire N__64729;
    wire N__64728;
    wire N__64725;
    wire N__64720;
    wire N__64717;
    wire N__64714;
    wire N__64713;
    wire N__64710;
    wire N__64709;
    wire N__64702;
    wire N__64699;
    wire N__64698;
    wire N__64695;
    wire N__64692;
    wire N__64687;
    wire N__64684;
    wire N__64681;
    wire N__64678;
    wire N__64675;
    wire N__64674;
    wire N__64671;
    wire N__64668;
    wire N__64663;
    wire N__64660;
    wire N__64657;
    wire N__64656;
    wire N__64653;
    wire N__64650;
    wire N__64647;
    wire N__64644;
    wire N__64639;
    wire N__64636;
    wire N__64633;
    wire N__64630;
    wire N__64629;
    wire N__64626;
    wire N__64623;
    wire N__64620;
    wire N__64615;
    wire N__64614;
    wire N__64611;
    wire N__64608;
    wire N__64605;
    wire N__64602;
    wire N__64599;
    wire N__64594;
    wire N__64591;
    wire N__64588;
    wire N__64587;
    wire N__64584;
    wire N__64581;
    wire N__64578;
    wire N__64573;
    wire N__64570;
    wire N__64567;
    wire N__64564;
    wire N__64561;
    wire N__64558;
    wire N__64557;
    wire N__64554;
    wire N__64551;
    wire N__64548;
    wire N__64543;
    wire N__64542;
    wire N__64539;
    wire N__64536;
    wire N__64533;
    wire N__64530;
    wire N__64527;
    wire N__64522;
    wire N__64519;
    wire N__64518;
    wire N__64517;
    wire N__64516;
    wire N__64511;
    wire N__64508;
    wire N__64505;
    wire N__64498;
    wire N__64495;
    wire N__64492;
    wire N__64489;
    wire N__64486;
    wire N__64483;
    wire N__64482;
    wire N__64481;
    wire N__64474;
    wire N__64473;
    wire N__64470;
    wire N__64467;
    wire N__64462;
    wire N__64461;
    wire N__64460;
    wire N__64457;
    wire N__64456;
    wire N__64449;
    wire N__64446;
    wire N__64441;
    wire N__64440;
    wire N__64439;
    wire N__64436;
    wire N__64431;
    wire N__64426;
    wire N__64423;
    wire N__64420;
    wire N__64419;
    wire N__64418;
    wire N__64417;
    wire N__64416;
    wire N__64415;
    wire N__64404;
    wire N__64401;
    wire N__64396;
    wire N__64395;
    wire N__64392;
    wire N__64389;
    wire N__64386;
    wire N__64381;
    wire N__64378;
    wire N__64375;
    wire N__64372;
    wire N__64369;
    wire N__64368;
    wire N__64367;
    wire N__64364;
    wire N__64363;
    wire N__64362;
    wire N__64361;
    wire N__64360;
    wire N__64359;
    wire N__64358;
    wire N__64355;
    wire N__64354;
    wire N__64353;
    wire N__64350;
    wire N__64349;
    wire N__64346;
    wire N__64345;
    wire N__64344;
    wire N__64341;
    wire N__64330;
    wire N__64325;
    wire N__64322;
    wire N__64317;
    wire N__64314;
    wire N__64313;
    wire N__64308;
    wire N__64303;
    wire N__64300;
    wire N__64297;
    wire N__64294;
    wire N__64293;
    wire N__64292;
    wire N__64291;
    wire N__64288;
    wire N__64285;
    wire N__64280;
    wire N__64275;
    wire N__64272;
    wire N__64265;
    wire N__64260;
    wire N__64257;
    wire N__64254;
    wire N__64243;
    wire N__64242;
    wire N__64239;
    wire N__64234;
    wire N__64231;
    wire N__64228;
    wire N__64225;
    wire N__64222;
    wire N__64219;
    wire N__64216;
    wire N__64215;
    wire N__64212;
    wire N__64207;
    wire N__64204;
    wire N__64203;
    wire N__64200;
    wire N__64197;
    wire N__64194;
    wire N__64191;
    wire N__64186;
    wire N__64185;
    wire N__64182;
    wire N__64177;
    wire N__64174;
    wire N__64173;
    wire N__64170;
    wire N__64165;
    wire N__64162;
    wire N__64159;
    wire N__64156;
    wire N__64153;
    wire N__64150;
    wire N__64149;
    wire N__64146;
    wire N__64145;
    wire N__64144;
    wire N__64143;
    wire N__64142;
    wire N__64141;
    wire N__64138;
    wire N__64135;
    wire N__64130;
    wire N__64129;
    wire N__64126;
    wire N__64121;
    wire N__64118;
    wire N__64113;
    wire N__64110;
    wire N__64109;
    wire N__64108;
    wire N__64105;
    wire N__64098;
    wire N__64091;
    wire N__64086;
    wire N__64081;
    wire N__64080;
    wire N__64077;
    wire N__64076;
    wire N__64073;
    wire N__64072;
    wire N__64071;
    wire N__64070;
    wire N__64069;
    wire N__64068;
    wire N__64065;
    wire N__64062;
    wire N__64057;
    wire N__64054;
    wire N__64049;
    wire N__64046;
    wire N__64043;
    wire N__64034;
    wire N__64027;
    wire N__64024;
    wire N__64021;
    wire N__64018;
    wire N__64015;
    wire N__64012;
    wire N__64011;
    wire N__64010;
    wire N__64009;
    wire N__64008;
    wire N__64007;
    wire N__64006;
    wire N__64005;
    wire N__64002;
    wire N__63999;
    wire N__63998;
    wire N__63995;
    wire N__63992;
    wire N__63989;
    wire N__63986;
    wire N__63985;
    wire N__63984;
    wire N__63981;
    wire N__63980;
    wire N__63977;
    wire N__63974;
    wire N__63971;
    wire N__63968;
    wire N__63965;
    wire N__63962;
    wire N__63959;
    wire N__63956;
    wire N__63955;
    wire N__63954;
    wire N__63953;
    wire N__63952;
    wire N__63949;
    wire N__63946;
    wire N__63943;
    wire N__63940;
    wire N__63937;
    wire N__63934;
    wire N__63931;
    wire N__63928;
    wire N__63925;
    wire N__63922;
    wire N__63917;
    wire N__63912;
    wire N__63909;
    wire N__63906;
    wire N__63901;
    wire N__63898;
    wire N__63895;
    wire N__63890;
    wire N__63887;
    wire N__63878;
    wire N__63859;
    wire N__63856;
    wire N__63855;
    wire N__63852;
    wire N__63849;
    wire N__63846;
    wire N__63841;
    wire N__63840;
    wire N__63837;
    wire N__63832;
    wire N__63829;
    wire N__63826;
    wire N__63823;
    wire N__63820;
    wire N__63817;
    wire N__63816;
    wire N__63811;
    wire N__63808;
    wire N__63807;
    wire N__63804;
    wire N__63801;
    wire N__63798;
    wire N__63793;
    wire N__63790;
    wire N__63787;
    wire N__63786;
    wire N__63783;
    wire N__63780;
    wire N__63775;
    wire N__63772;
    wire N__63769;
    wire N__63766;
    wire N__63765;
    wire N__63762;
    wire N__63759;
    wire N__63754;
    wire N__63751;
    wire N__63750;
    wire N__63747;
    wire N__63744;
    wire N__63741;
    wire N__63738;
    wire N__63733;
    wire N__63730;
    wire N__63729;
    wire N__63728;
    wire N__63727;
    wire N__63724;
    wire N__63721;
    wire N__63718;
    wire N__63717;
    wire N__63714;
    wire N__63713;
    wire N__63712;
    wire N__63711;
    wire N__63708;
    wire N__63705;
    wire N__63702;
    wire N__63699;
    wire N__63696;
    wire N__63693;
    wire N__63690;
    wire N__63689;
    wire N__63686;
    wire N__63685;
    wire N__63684;
    wire N__63681;
    wire N__63678;
    wire N__63677;
    wire N__63676;
    wire N__63673;
    wire N__63670;
    wire N__63667;
    wire N__63664;
    wire N__63661;
    wire N__63658;
    wire N__63655;
    wire N__63650;
    wire N__63649;
    wire N__63648;
    wire N__63643;
    wire N__63640;
    wire N__63637;
    wire N__63636;
    wire N__63631;
    wire N__63624;
    wire N__63621;
    wire N__63616;
    wire N__63613;
    wire N__63610;
    wire N__63603;
    wire N__63600;
    wire N__63583;
    wire N__63580;
    wire N__63579;
    wire N__63576;
    wire N__63573;
    wire N__63568;
    wire N__63565;
    wire N__63562;
    wire N__63561;
    wire N__63558;
    wire N__63555;
    wire N__63552;
    wire N__63549;
    wire N__63544;
    wire N__63543;
    wire N__63542;
    wire N__63541;
    wire N__63540;
    wire N__63539;
    wire N__63538;
    wire N__63537;
    wire N__63536;
    wire N__63535;
    wire N__63534;
    wire N__63533;
    wire N__63532;
    wire N__63531;
    wire N__63530;
    wire N__63529;
    wire N__63528;
    wire N__63527;
    wire N__63526;
    wire N__63525;
    wire N__63522;
    wire N__63513;
    wire N__63510;
    wire N__63509;
    wire N__63506;
    wire N__63505;
    wire N__63504;
    wire N__63503;
    wire N__63500;
    wire N__63497;
    wire N__63494;
    wire N__63493;
    wire N__63492;
    wire N__63491;
    wire N__63490;
    wire N__63487;
    wire N__63486;
    wire N__63485;
    wire N__63482;
    wire N__63477;
    wire N__63474;
    wire N__63473;
    wire N__63472;
    wire N__63471;
    wire N__63466;
    wire N__63463;
    wire N__63458;
    wire N__63455;
    wire N__63450;
    wire N__63449;
    wire N__63448;
    wire N__63447;
    wire N__63446;
    wire N__63445;
    wire N__63442;
    wire N__63441;
    wire N__63440;
    wire N__63439;
    wire N__63438;
    wire N__63437;
    wire N__63436;
    wire N__63433;
    wire N__63430;
    wire N__63425;
    wire N__63422;
    wire N__63417;
    wire N__63410;
    wire N__63407;
    wire N__63404;
    wire N__63399;
    wire N__63398;
    wire N__63393;
    wire N__63386;
    wire N__63383;
    wire N__63382;
    wire N__63381;
    wire N__63380;
    wire N__63379;
    wire N__63378;
    wire N__63377;
    wire N__63366;
    wire N__63363;
    wire N__63354;
    wire N__63353;
    wire N__63350;
    wire N__63347;
    wire N__63344;
    wire N__63343;
    wire N__63342;
    wire N__63341;
    wire N__63340;
    wire N__63339;
    wire N__63338;
    wire N__63333;
    wire N__63328;
    wire N__63325;
    wire N__63322;
    wire N__63313;
    wire N__63312;
    wire N__63311;
    wire N__63308;
    wire N__63303;
    wire N__63300;
    wire N__63297;
    wire N__63294;
    wire N__63291;
    wire N__63288;
    wire N__63283;
    wire N__63280;
    wire N__63277;
    wire N__63276;
    wire N__63273;
    wire N__63268;
    wire N__63265;
    wire N__63262;
    wire N__63259;
    wire N__63258;
    wire N__63247;
    wire N__63242;
    wire N__63239;
    wire N__63234;
    wire N__63231;
    wire N__63230;
    wire N__63227;
    wire N__63224;
    wire N__63221;
    wire N__63218;
    wire N__63215;
    wire N__63212;
    wire N__63209;
    wire N__63204;
    wire N__63199;
    wire N__63196;
    wire N__63189;
    wire N__63182;
    wire N__63177;
    wire N__63174;
    wire N__63169;
    wire N__63164;
    wire N__63163;
    wire N__63160;
    wire N__63157;
    wire N__63154;
    wire N__63151;
    wire N__63148;
    wire N__63135;
    wire N__63126;
    wire N__63119;
    wire N__63116;
    wire N__63103;
    wire N__63100;
    wire N__63097;
    wire N__63092;
    wire N__63085;
    wire N__63082;
    wire N__63079;
    wire N__63076;
    wire N__63075;
    wire N__63072;
    wire N__63069;
    wire N__63064;
    wire N__63061;
    wire N__63060;
    wire N__63057;
    wire N__63054;
    wire N__63049;
    wire N__63046;
    wire N__63043;
    wire N__63042;
    wire N__63039;
    wire N__63036;
    wire N__63033;
    wire N__63028;
    wire N__63025;
    wire N__63022;
    wire N__63019;
    wire N__63018;
    wire N__63015;
    wire N__63012;
    wire N__63007;
    wire N__63006;
    wire N__63005;
    wire N__63002;
    wire N__63001;
    wire N__62998;
    wire N__62997;
    wire N__62996;
    wire N__62993;
    wire N__62990;
    wire N__62989;
    wire N__62988;
    wire N__62987;
    wire N__62986;
    wire N__62985;
    wire N__62984;
    wire N__62983;
    wire N__62980;
    wire N__62979;
    wire N__62978;
    wire N__62975;
    wire N__62972;
    wire N__62969;
    wire N__62966;
    wire N__62963;
    wire N__62962;
    wire N__62959;
    wire N__62956;
    wire N__62953;
    wire N__62950;
    wire N__62947;
    wire N__62944;
    wire N__62941;
    wire N__62938;
    wire N__62935;
    wire N__62932;
    wire N__62927;
    wire N__62920;
    wire N__62917;
    wire N__62914;
    wire N__62905;
    wire N__62900;
    wire N__62897;
    wire N__62890;
    wire N__62887;
    wire N__62872;
    wire N__62871;
    wire N__62866;
    wire N__62863;
    wire N__62862;
    wire N__62861;
    wire N__62860;
    wire N__62859;
    wire N__62858;
    wire N__62857;
    wire N__62856;
    wire N__62855;
    wire N__62854;
    wire N__62853;
    wire N__62852;
    wire N__62849;
    wire N__62846;
    wire N__62845;
    wire N__62844;
    wire N__62843;
    wire N__62842;
    wire N__62839;
    wire N__62836;
    wire N__62835;
    wire N__62834;
    wire N__62833;
    wire N__62824;
    wire N__62823;
    wire N__62822;
    wire N__62821;
    wire N__62818;
    wire N__62817;
    wire N__62814;
    wire N__62813;
    wire N__62812;
    wire N__62811;
    wire N__62810;
    wire N__62809;
    wire N__62808;
    wire N__62807;
    wire N__62804;
    wire N__62803;
    wire N__62802;
    wire N__62801;
    wire N__62800;
    wire N__62799;
    wire N__62798;
    wire N__62797;
    wire N__62796;
    wire N__62793;
    wire N__62792;
    wire N__62791;
    wire N__62790;
    wire N__62783;
    wire N__62782;
    wire N__62781;
    wire N__62780;
    wire N__62779;
    wire N__62778;
    wire N__62777;
    wire N__62770;
    wire N__62765;
    wire N__62758;
    wire N__62755;
    wire N__62750;
    wire N__62747;
    wire N__62744;
    wire N__62741;
    wire N__62734;
    wire N__62725;
    wire N__62724;
    wire N__62723;
    wire N__62720;
    wire N__62719;
    wire N__62718;
    wire N__62717;
    wire N__62716;
    wire N__62713;
    wire N__62710;
    wire N__62707;
    wire N__62704;
    wire N__62699;
    wire N__62694;
    wire N__62691;
    wire N__62690;
    wire N__62689;
    wire N__62688;
    wire N__62685;
    wire N__62680;
    wire N__62679;
    wire N__62678;
    wire N__62677;
    wire N__62676;
    wire N__62673;
    wire N__62670;
    wire N__62665;
    wire N__62656;
    wire N__62641;
    wire N__62636;
    wire N__62635;
    wire N__62634;
    wire N__62633;
    wire N__62630;
    wire N__62625;
    wire N__62618;
    wire N__62613;
    wire N__62612;
    wire N__62607;
    wire N__62596;
    wire N__62593;
    wire N__62590;
    wire N__62587;
    wire N__62582;
    wire N__62579;
    wire N__62576;
    wire N__62573;
    wire N__62570;
    wire N__62557;
    wire N__62550;
    wire N__62547;
    wire N__62542;
    wire N__62539;
    wire N__62536;
    wire N__62531;
    wire N__62522;
    wire N__62517;
    wire N__62510;
    wire N__62507;
    wire N__62504;
    wire N__62501;
    wire N__62498;
    wire N__62491;
    wire N__62486;
    wire N__62481;
    wire N__62470;
    wire N__62467;
    wire N__62464;
    wire N__62463;
    wire N__62460;
    wire N__62457;
    wire N__62454;
    wire N__62451;
    wire N__62446;
    wire N__62445;
    wire N__62444;
    wire N__62439;
    wire N__62436;
    wire N__62431;
    wire N__62430;
    wire N__62429;
    wire N__62426;
    wire N__62425;
    wire N__62424;
    wire N__62423;
    wire N__62422;
    wire N__62421;
    wire N__62420;
    wire N__62419;
    wire N__62416;
    wire N__62415;
    wire N__62414;
    wire N__62413;
    wire N__62412;
    wire N__62411;
    wire N__62408;
    wire N__62407;
    wire N__62404;
    wire N__62401;
    wire N__62400;
    wire N__62395;
    wire N__62388;
    wire N__62385;
    wire N__62384;
    wire N__62383;
    wire N__62380;
    wire N__62379;
    wire N__62378;
    wire N__62377;
    wire N__62376;
    wire N__62375;
    wire N__62374;
    wire N__62373;
    wire N__62372;
    wire N__62371;
    wire N__62368;
    wire N__62367;
    wire N__62364;
    wire N__62361;
    wire N__62360;
    wire N__62359;
    wire N__62358;
    wire N__62357;
    wire N__62356;
    wire N__62355;
    wire N__62354;
    wire N__62353;
    wire N__62352;
    wire N__62351;
    wire N__62350;
    wire N__62349;
    wire N__62346;
    wire N__62341;
    wire N__62338;
    wire N__62333;
    wire N__62332;
    wire N__62331;
    wire N__62330;
    wire N__62329;
    wire N__62326;
    wire N__62321;
    wire N__62318;
    wire N__62317;
    wire N__62316;
    wire N__62315;
    wire N__62312;
    wire N__62309;
    wire N__62306;
    wire N__62297;
    wire N__62292;
    wire N__62285;
    wire N__62282;
    wire N__62279;
    wire N__62274;
    wire N__62273;
    wire N__62270;
    wire N__62269;
    wire N__62268;
    wire N__62263;
    wire N__62256;
    wire N__62255;
    wire N__62254;
    wire N__62253;
    wire N__62252;
    wire N__62251;
    wire N__62248;
    wire N__62245;
    wire N__62244;
    wire N__62243;
    wire N__62240;
    wire N__62237;
    wire N__62232;
    wire N__62229;
    wire N__62222;
    wire N__62219;
    wire N__62218;
    wire N__62217;
    wire N__62216;
    wire N__62213;
    wire N__62208;
    wire N__62205;
    wire N__62202;
    wire N__62199;
    wire N__62198;
    wire N__62195;
    wire N__62192;
    wire N__62189;
    wire N__62186;
    wire N__62179;
    wire N__62168;
    wire N__62159;
    wire N__62154;
    wire N__62149;
    wire N__62142;
    wire N__62137;
    wire N__62132;
    wire N__62125;
    wire N__62118;
    wire N__62111;
    wire N__62108;
    wire N__62103;
    wire N__62098;
    wire N__62095;
    wire N__62084;
    wire N__62081;
    wire N__62078;
    wire N__62075;
    wire N__62068;
    wire N__62061;
    wire N__62052;
    wire N__62045;
    wire N__62032;
    wire N__62029;
    wire N__62026;
    wire N__62023;
    wire N__62020;
    wire N__62019;
    wire N__62016;
    wire N__62013;
    wire N__62008;
    wire N__62005;
    wire N__62002;
    wire N__62001;
    wire N__61998;
    wire N__61995;
    wire N__61990;
    wire N__61987;
    wire N__61986;
    wire N__61981;
    wire N__61978;
    wire N__61975;
    wire N__61972;
    wire N__61969;
    wire N__61966;
    wire N__61963;
    wire N__61960;
    wire N__61957;
    wire N__61954;
    wire N__61951;
    wire N__61948;
    wire N__61945;
    wire N__61942;
    wire N__61939;
    wire N__61936;
    wire N__61935;
    wire N__61932;
    wire N__61929;
    wire N__61924;
    wire N__61921;
    wire N__61918;
    wire N__61915;
    wire N__61912;
    wire N__61909;
    wire N__61906;
    wire N__61905;
    wire N__61902;
    wire N__61899;
    wire N__61894;
    wire N__61893;
    wire N__61892;
    wire N__61891;
    wire N__61890;
    wire N__61889;
    wire N__61886;
    wire N__61885;
    wire N__61882;
    wire N__61881;
    wire N__61880;
    wire N__61879;
    wire N__61878;
    wire N__61875;
    wire N__61872;
    wire N__61867;
    wire N__61864;
    wire N__61861;
    wire N__61858;
    wire N__61855;
    wire N__61852;
    wire N__61849;
    wire N__61846;
    wire N__61839;
    wire N__61836;
    wire N__61831;
    wire N__61830;
    wire N__61829;
    wire N__61828;
    wire N__61827;
    wire N__61824;
    wire N__61821;
    wire N__61818;
    wire N__61815;
    wire N__61810;
    wire N__61807;
    wire N__61804;
    wire N__61801;
    wire N__61798;
    wire N__61795;
    wire N__61792;
    wire N__61783;
    wire N__61780;
    wire N__61765;
    wire N__61764;
    wire N__61759;
    wire N__61756;
    wire N__61753;
    wire N__61750;
    wire N__61747;
    wire N__61746;
    wire N__61743;
    wire N__61740;
    wire N__61735;
    wire N__61732;
    wire N__61729;
    wire N__61728;
    wire N__61725;
    wire N__61722;
    wire N__61717;
    wire N__61716;
    wire N__61713;
    wire N__61710;
    wire N__61705;
    wire N__61702;
    wire N__61699;
    wire N__61696;
    wire N__61695;
    wire N__61692;
    wire N__61689;
    wire N__61684;
    wire N__61681;
    wire N__61680;
    wire N__61677;
    wire N__61674;
    wire N__61669;
    wire N__61666;
    wire N__61665;
    wire N__61662;
    wire N__61659;
    wire N__61654;
    wire N__61651;
    wire N__61648;
    wire N__61647;
    wire N__61644;
    wire N__61641;
    wire N__61638;
    wire N__61635;
    wire N__61630;
    wire N__61627;
    wire N__61624;
    wire N__61621;
    wire N__61618;
    wire N__61617;
    wire N__61614;
    wire N__61611;
    wire N__61606;
    wire N__61603;
    wire N__61600;
    wire N__61597;
    wire N__61594;
    wire N__61591;
    wire N__61588;
    wire N__61585;
    wire N__61582;
    wire N__61579;
    wire N__61576;
    wire N__61573;
    wire N__61570;
    wire N__61567;
    wire N__61564;
    wire N__61561;
    wire N__61558;
    wire N__61555;
    wire N__61552;
    wire N__61549;
    wire N__61546;
    wire N__61543;
    wire N__61540;
    wire N__61537;
    wire N__61534;
    wire N__61531;
    wire N__61528;
    wire N__61525;
    wire N__61522;
    wire N__61519;
    wire N__61516;
    wire N__61513;
    wire N__61512;
    wire N__61509;
    wire N__61506;
    wire N__61501;
    wire N__61498;
    wire N__61495;
    wire N__61494;
    wire N__61491;
    wire N__61488;
    wire N__61483;
    wire N__61480;
    wire N__61477;
    wire N__61474;
    wire N__61473;
    wire N__61470;
    wire N__61467;
    wire N__61462;
    wire N__61461;
    wire N__61456;
    wire N__61453;
    wire N__61450;
    wire N__61449;
    wire N__61446;
    wire N__61443;
    wire N__61440;
    wire N__61437;
    wire N__61432;
    wire N__61429;
    wire N__61428;
    wire N__61425;
    wire N__61422;
    wire N__61419;
    wire N__61416;
    wire N__61411;
    wire N__61408;
    wire N__61405;
    wire N__61404;
    wire N__61403;
    wire N__61400;
    wire N__61399;
    wire N__61398;
    wire N__61397;
    wire N__61396;
    wire N__61395;
    wire N__61390;
    wire N__61389;
    wire N__61388;
    wire N__61387;
    wire N__61386;
    wire N__61385;
    wire N__61384;
    wire N__61379;
    wire N__61374;
    wire N__61373;
    wire N__61372;
    wire N__61367;
    wire N__61364;
    wire N__61359;
    wire N__61350;
    wire N__61349;
    wire N__61348;
    wire N__61347;
    wire N__61346;
    wire N__61345;
    wire N__61344;
    wire N__61343;
    wire N__61342;
    wire N__61341;
    wire N__61340;
    wire N__61337;
    wire N__61334;
    wire N__61333;
    wire N__61332;
    wire N__61329;
    wire N__61326;
    wire N__61317;
    wire N__61308;
    wire N__61307;
    wire N__61306;
    wire N__61305;
    wire N__61304;
    wire N__61301;
    wire N__61296;
    wire N__61295;
    wire N__61292;
    wire N__61291;
    wire N__61290;
    wire N__61289;
    wire N__61288;
    wire N__61287;
    wire N__61286;
    wire N__61283;
    wire N__61282;
    wire N__61281;
    wire N__61280;
    wire N__61277;
    wire N__61272;
    wire N__61269;
    wire N__61268;
    wire N__61265;
    wire N__61264;
    wire N__61263;
    wire N__61262;
    wire N__61259;
    wire N__61252;
    wire N__61251;
    wire N__61250;
    wire N__61249;
    wire N__61248;
    wire N__61247;
    wire N__61246;
    wire N__61241;
    wire N__61240;
    wire N__61239;
    wire N__61234;
    wire N__61231;
    wire N__61228;
    wire N__61225;
    wire N__61222;
    wire N__61221;
    wire N__61220;
    wire N__61217;
    wire N__61214;
    wire N__61211;
    wire N__61208;
    wire N__61203;
    wire N__61194;
    wire N__61187;
    wire N__61184;
    wire N__61179;
    wire N__61174;
    wire N__61169;
    wire N__61166;
    wire N__61161;
    wire N__61158;
    wire N__61155;
    wire N__61152;
    wire N__61149;
    wire N__61144;
    wire N__61137;
    wire N__61134;
    wire N__61131;
    wire N__61128;
    wire N__61125;
    wire N__61116;
    wire N__61113;
    wire N__61112;
    wire N__61111;
    wire N__61110;
    wire N__61109;
    wire N__61108;
    wire N__61107;
    wire N__61100;
    wire N__61091;
    wire N__61088;
    wire N__61085;
    wire N__61080;
    wire N__61077;
    wire N__61072;
    wire N__61069;
    wire N__61064;
    wire N__61057;
    wire N__61056;
    wire N__61055;
    wire N__61042;
    wire N__61035;
    wire N__61030;
    wire N__61027;
    wire N__61024;
    wire N__61021;
    wire N__61018;
    wire N__61015;
    wire N__61010;
    wire N__61005;
    wire N__61002;
    wire N__60999;
    wire N__60996;
    wire N__60989;
    wire N__60984;
    wire N__60979;
    wire N__60972;
    wire N__60967;
    wire N__60964;
    wire N__60961;
    wire N__60958;
    wire N__60955;
    wire N__60952;
    wire N__60949;
    wire N__60946;
    wire N__60943;
    wire N__60940;
    wire N__60937;
    wire N__60934;
    wire N__60931;
    wire N__60928;
    wire N__60925;
    wire N__60922;
    wire N__60919;
    wire N__60916;
    wire N__60913;
    wire N__60910;
    wire N__60907;
    wire N__60904;
    wire N__60901;
    wire N__60898;
    wire N__60895;
    wire N__60892;
    wire N__60889;
    wire N__60888;
    wire N__60887;
    wire N__60886;
    wire N__60885;
    wire N__60874;
    wire N__60871;
    wire N__60870;
    wire N__60869;
    wire N__60862;
    wire N__60859;
    wire N__60858;
    wire N__60857;
    wire N__60856;
    wire N__60853;
    wire N__60848;
    wire N__60843;
    wire N__60838;
    wire N__60835;
    wire N__60834;
    wire N__60833;
    wire N__60826;
    wire N__60823;
    wire N__60820;
    wire N__60819;
    wire N__60818;
    wire N__60817;
    wire N__60814;
    wire N__60813;
    wire N__60812;
    wire N__60799;
    wire N__60796;
    wire N__60795;
    wire N__60794;
    wire N__60793;
    wire N__60788;
    wire N__60787;
    wire N__60782;
    wire N__60781;
    wire N__60780;
    wire N__60777;
    wire N__60774;
    wire N__60771;
    wire N__60770;
    wire N__60769;
    wire N__60768;
    wire N__60767;
    wire N__60764;
    wire N__60761;
    wire N__60754;
    wire N__60751;
    wire N__60742;
    wire N__60733;
    wire N__60730;
    wire N__60727;
    wire N__60726;
    wire N__60725;
    wire N__60724;
    wire N__60723;
    wire N__60722;
    wire N__60721;
    wire N__60718;
    wire N__60713;
    wire N__60710;
    wire N__60707;
    wire N__60702;
    wire N__60701;
    wire N__60700;
    wire N__60699;
    wire N__60698;
    wire N__60697;
    wire N__60694;
    wire N__60691;
    wire N__60684;
    wire N__60675;
    wire N__60672;
    wire N__60661;
    wire N__60660;
    wire N__60657;
    wire N__60654;
    wire N__60649;
    wire N__60646;
    wire N__60643;
    wire N__60640;
    wire N__60637;
    wire N__60634;
    wire N__60631;
    wire N__60628;
    wire N__60625;
    wire N__60622;
    wire N__60619;
    wire N__60616;
    wire N__60613;
    wire N__60610;
    wire N__60607;
    wire N__60604;
    wire N__60601;
    wire N__60598;
    wire N__60595;
    wire N__60592;
    wire N__60589;
    wire N__60586;
    wire N__60583;
    wire N__60580;
    wire N__60579;
    wire N__60576;
    wire N__60573;
    wire N__60568;
    wire N__60567;
    wire N__60564;
    wire N__60561;
    wire N__60556;
    wire N__60553;
    wire N__60550;
    wire N__60549;
    wire N__60548;
    wire N__60543;
    wire N__60540;
    wire N__60535;
    wire N__60534;
    wire N__60533;
    wire N__60528;
    wire N__60525;
    wire N__60520;
    wire N__60517;
    wire N__60516;
    wire N__60515;
    wire N__60510;
    wire N__60507;
    wire N__60502;
    wire N__60501;
    wire N__60500;
    wire N__60495;
    wire N__60492;
    wire N__60487;
    wire N__60486;
    wire N__60481;
    wire N__60478;
    wire N__60475;
    wire N__60474;
    wire N__60473;
    wire N__60468;
    wire N__60465;
    wire N__60460;
    wire N__60457;
    wire N__60454;
    wire N__60451;
    wire N__60448;
    wire N__60445;
    wire N__60442;
    wire N__60439;
    wire N__60436;
    wire N__60435;
    wire N__60432;
    wire N__60429;
    wire N__60424;
    wire N__60421;
    wire N__60418;
    wire N__60415;
    wire N__60414;
    wire N__60411;
    wire N__60408;
    wire N__60407;
    wire N__60404;
    wire N__60401;
    wire N__60398;
    wire N__60395;
    wire N__60392;
    wire N__60385;
    wire N__60384;
    wire N__60379;
    wire N__60378;
    wire N__60377;
    wire N__60374;
    wire N__60369;
    wire N__60366;
    wire N__60363;
    wire N__60358;
    wire N__60357;
    wire N__60356;
    wire N__60353;
    wire N__60352;
    wire N__60351;
    wire N__60350;
    wire N__60349;
    wire N__60346;
    wire N__60345;
    wire N__60344;
    wire N__60343;
    wire N__60340;
    wire N__60337;
    wire N__60334;
    wire N__60331;
    wire N__60318;
    wire N__60307;
    wire N__60304;
    wire N__60301;
    wire N__60300;
    wire N__60299;
    wire N__60298;
    wire N__60297;
    wire N__60296;
    wire N__60295;
    wire N__60290;
    wire N__60279;
    wire N__60274;
    wire N__60271;
    wire N__60270;
    wire N__60267;
    wire N__60264;
    wire N__60259;
    wire N__60256;
    wire N__60255;
    wire N__60252;
    wire N__60249;
    wire N__60244;
    wire N__60243;
    wire N__60240;
    wire N__60237;
    wire N__60232;
    wire N__60229;
    wire N__60226;
    wire N__60225;
    wire N__60224;
    wire N__60223;
    wire N__60222;
    wire N__60221;
    wire N__60218;
    wire N__60215;
    wire N__60206;
    wire N__60199;
    wire N__60196;
    wire N__60193;
    wire N__60190;
    wire N__60187;
    wire N__60184;
    wire N__60181;
    wire N__60178;
    wire N__60175;
    wire N__60174;
    wire N__60169;
    wire N__60168;
    wire N__60165;
    wire N__60162;
    wire N__60159;
    wire N__60156;
    wire N__60151;
    wire N__60148;
    wire N__60147;
    wire N__60144;
    wire N__60141;
    wire N__60136;
    wire N__60133;
    wire N__60132;
    wire N__60129;
    wire N__60126;
    wire N__60121;
    wire N__60118;
    wire N__60115;
    wire N__60112;
    wire N__60109;
    wire N__60106;
    wire N__60105;
    wire N__60104;
    wire N__60103;
    wire N__60102;
    wire N__60101;
    wire N__60090;
    wire N__60087;
    wire N__60082;
    wire N__60081;
    wire N__60076;
    wire N__60073;
    wire N__60072;
    wire N__60071;
    wire N__60070;
    wire N__60069;
    wire N__60068;
    wire N__60065;
    wire N__60062;
    wire N__60057;
    wire N__60052;
    wire N__60043;
    wire N__60042;
    wire N__60041;
    wire N__60040;
    wire N__60039;
    wire N__60038;
    wire N__60037;
    wire N__60026;
    wire N__60021;
    wire N__60016;
    wire N__60013;
    wire N__60010;
    wire N__60007;
    wire N__60004;
    wire N__60001;
    wire N__59998;
    wire N__59997;
    wire N__59994;
    wire N__59991;
    wire N__59986;
    wire N__59983;
    wire N__59980;
    wire N__59977;
    wire N__59976;
    wire N__59973;
    wire N__59970;
    wire N__59965;
    wire N__59962;
    wire N__59959;
    wire N__59956;
    wire N__59953;
    wire N__59952;
    wire N__59949;
    wire N__59946;
    wire N__59941;
    wire N__59938;
    wire N__59935;
    wire N__59932;
    wire N__59929;
    wire N__59926;
    wire N__59925;
    wire N__59922;
    wire N__59919;
    wire N__59914;
    wire N__59911;
    wire N__59908;
    wire N__59907;
    wire N__59904;
    wire N__59901;
    wire N__59896;
    wire N__59893;
    wire N__59890;
    wire N__59887;
    wire N__59886;
    wire N__59883;
    wire N__59880;
    wire N__59875;
    wire N__59872;
    wire N__59869;
    wire N__59868;
    wire N__59865;
    wire N__59862;
    wire N__59857;
    wire N__59854;
    wire N__59851;
    wire N__59848;
    wire N__59845;
    wire N__59842;
    wire N__59839;
    wire N__59836;
    wire N__59835;
    wire N__59832;
    wire N__59829;
    wire N__59824;
    wire N__59821;
    wire N__59818;
    wire N__59815;
    wire N__59812;
    wire N__59809;
    wire N__59806;
    wire N__59805;
    wire N__59802;
    wire N__59799;
    wire N__59796;
    wire N__59793;
    wire N__59788;
    wire N__59785;
    wire N__59784;
    wire N__59781;
    wire N__59776;
    wire N__59773;
    wire N__59772;
    wire N__59769;
    wire N__59764;
    wire N__59761;
    wire N__59760;
    wire N__59757;
    wire N__59754;
    wire N__59749;
    wire N__59746;
    wire N__59745;
    wire N__59740;
    wire N__59737;
    wire N__59734;
    wire N__59731;
    wire N__59728;
    wire N__59727;
    wire N__59724;
    wire N__59721;
    wire N__59716;
    wire N__59713;
    wire N__59712;
    wire N__59709;
    wire N__59706;
    wire N__59701;
    wire N__59698;
    wire N__59695;
    wire N__59694;
    wire N__59691;
    wire N__59688;
    wire N__59683;
    wire N__59680;
    wire N__59679;
    wire N__59674;
    wire N__59671;
    wire N__59670;
    wire N__59665;
    wire N__59662;
    wire N__59659;
    wire N__59658;
    wire N__59657;
    wire N__59654;
    wire N__59653;
    wire N__59652;
    wire N__59651;
    wire N__59648;
    wire N__59645;
    wire N__59644;
    wire N__59641;
    wire N__59638;
    wire N__59635;
    wire N__59634;
    wire N__59633;
    wire N__59632;
    wire N__59629;
    wire N__59626;
    wire N__59623;
    wire N__59620;
    wire N__59615;
    wire N__59612;
    wire N__59611;
    wire N__59608;
    wire N__59605;
    wire N__59602;
    wire N__59601;
    wire N__59600;
    wire N__59597;
    wire N__59594;
    wire N__59589;
    wire N__59586;
    wire N__59583;
    wire N__59580;
    wire N__59577;
    wire N__59572;
    wire N__59569;
    wire N__59566;
    wire N__59565;
    wire N__59564;
    wire N__59561;
    wire N__59554;
    wire N__59549;
    wire N__59546;
    wire N__59541;
    wire N__59538;
    wire N__59535;
    wire N__59532;
    wire N__59515;
    wire N__59514;
    wire N__59509;
    wire N__59506;
    wire N__59503;
    wire N__59500;
    wire N__59497;
    wire N__59494;
    wire N__59491;
    wire N__59488;
    wire N__59485;
    wire N__59482;
    wire N__59479;
    wire N__59478;
    wire N__59475;
    wire N__59472;
    wire N__59467;
    wire N__59464;
    wire N__59461;
    wire N__59460;
    wire N__59457;
    wire N__59454;
    wire N__59449;
    wire N__59448;
    wire N__59443;
    wire N__59440;
    wire N__59437;
    wire N__59434;
    wire N__59431;
    wire N__59428;
    wire N__59425;
    wire N__59422;
    wire N__59419;
    wire N__59418;
    wire N__59413;
    wire N__59410;
    wire N__59407;
    wire N__59406;
    wire N__59403;
    wire N__59400;
    wire N__59395;
    wire N__59392;
    wire N__59389;
    wire N__59386;
    wire N__59385;
    wire N__59382;
    wire N__59379;
    wire N__59374;
    wire N__59371;
    wire N__59370;
    wire N__59367;
    wire N__59362;
    wire N__59359;
    wire N__59358;
    wire N__59355;
    wire N__59350;
    wire N__59347;
    wire N__59346;
    wire N__59343;
    wire N__59338;
    wire N__59335;
    wire N__59332;
    wire N__59329;
    wire N__59328;
    wire N__59325;
    wire N__59322;
    wire N__59319;
    wire N__59316;
    wire N__59311;
    wire N__59308;
    wire N__59307;
    wire N__59304;
    wire N__59301;
    wire N__59296;
    wire N__59293;
    wire N__59290;
    wire N__59287;
    wire N__59284;
    wire N__59283;
    wire N__59282;
    wire N__59281;
    wire N__59280;
    wire N__59279;
    wire N__59276;
    wire N__59275;
    wire N__59274;
    wire N__59273;
    wire N__59272;
    wire N__59269;
    wire N__59264;
    wire N__59261;
    wire N__59258;
    wire N__59255;
    wire N__59252;
    wire N__59249;
    wire N__59248;
    wire N__59247;
    wire N__59244;
    wire N__59243;
    wire N__59240;
    wire N__59239;
    wire N__59236;
    wire N__59233;
    wire N__59230;
    wire N__59227;
    wire N__59222;
    wire N__59219;
    wire N__59216;
    wire N__59213;
    wire N__59210;
    wire N__59207;
    wire N__59206;
    wire N__59203;
    wire N__59200;
    wire N__59199;
    wire N__59196;
    wire N__59191;
    wire N__59184;
    wire N__59179;
    wire N__59174;
    wire N__59171;
    wire N__59166;
    wire N__59163;
    wire N__59146;
    wire N__59143;
    wire N__59142;
    wire N__59139;
    wire N__59136;
    wire N__59131;
    wire N__59128;
    wire N__59125;
    wire N__59122;
    wire N__59121;
    wire N__59118;
    wire N__59115;
    wire N__59110;
    wire N__59107;
    wire N__59104;
    wire N__59101;
    wire N__59098;
    wire N__59097;
    wire N__59094;
    wire N__59091;
    wire N__59086;
    wire N__59083;
    wire N__59082;
    wire N__59079;
    wire N__59074;
    wire N__59071;
    wire N__59070;
    wire N__59067;
    wire N__59062;
    wire N__59059;
    wire N__59058;
    wire N__59055;
    wire N__59052;
    wire N__59049;
    wire N__59044;
    wire N__59041;
    wire N__59038;
    wire N__59035;
    wire N__59032;
    wire N__59029;
    wire N__59026;
    wire N__59025;
    wire N__59020;
    wire N__59017;
    wire N__59016;
    wire N__59013;
    wire N__59010;
    wire N__59005;
    wire N__59002;
    wire N__58999;
    wire N__58996;
    wire N__58993;
    wire N__58992;
    wire N__58989;
    wire N__58986;
    wire N__58983;
    wire N__58980;
    wire N__58975;
    wire N__58974;
    wire N__58971;
    wire N__58968;
    wire N__58965;
    wire N__58960;
    wire N__58957;
    wire N__58954;
    wire N__58951;
    wire N__58948;
    wire N__58945;
    wire N__58944;
    wire N__58939;
    wire N__58936;
    wire N__58933;
    wire N__58932;
    wire N__58929;
    wire N__58926;
    wire N__58921;
    wire N__58918;
    wire N__58915;
    wire N__58914;
    wire N__58911;
    wire N__58908;
    wire N__58903;
    wire N__58902;
    wire N__58899;
    wire N__58896;
    wire N__58893;
    wire N__58888;
    wire N__58885;
    wire N__58882;
    wire N__58879;
    wire N__58876;
    wire N__58873;
    wire N__58872;
    wire N__58869;
    wire N__58866;
    wire N__58861;
    wire N__58860;
    wire N__58857;
    wire N__58852;
    wire N__58849;
    wire N__58846;
    wire N__58843;
    wire N__58840;
    wire N__58837;
    wire N__58834;
    wire N__58831;
    wire N__58828;
    wire N__58825;
    wire N__58822;
    wire N__58819;
    wire N__58816;
    wire N__58813;
    wire N__58810;
    wire N__58807;
    wire N__58806;
    wire N__58801;
    wire N__58798;
    wire N__58797;
    wire N__58794;
    wire N__58789;
    wire N__58786;
    wire N__58783;
    wire N__58780;
    wire N__58779;
    wire N__58776;
    wire N__58773;
    wire N__58768;
    wire N__58765;
    wire N__58762;
    wire N__58759;
    wire N__58756;
    wire N__58753;
    wire N__58752;
    wire N__58749;
    wire N__58746;
    wire N__58741;
    wire N__58738;
    wire N__58735;
    wire N__58732;
    wire N__58729;
    wire N__58726;
    wire N__58723;
    wire N__58720;
    wire N__58717;
    wire N__58714;
    wire N__58713;
    wire N__58710;
    wire N__58707;
    wire N__58704;
    wire N__58701;
    wire N__58696;
    wire N__58693;
    wire N__58690;
    wire N__58687;
    wire N__58684;
    wire N__58681;
    wire N__58678;
    wire N__58675;
    wire N__58672;
    wire N__58671;
    wire N__58668;
    wire N__58665;
    wire N__58660;
    wire N__58657;
    wire N__58654;
    wire N__58653;
    wire N__58650;
    wire N__58647;
    wire N__58644;
    wire N__58639;
    wire N__58636;
    wire N__58635;
    wire N__58632;
    wire N__58629;
    wire N__58626;
    wire N__58623;
    wire N__58618;
    wire N__58615;
    wire N__58612;
    wire N__58609;
    wire N__58608;
    wire N__58605;
    wire N__58602;
    wire N__58599;
    wire N__58594;
    wire N__58593;
    wire N__58590;
    wire N__58587;
    wire N__58582;
    wire N__58581;
    wire N__58578;
    wire N__58575;
    wire N__58572;
    wire N__58567;
    wire N__58566;
    wire N__58563;
    wire N__58560;
    wire N__58555;
    wire N__58552;
    wire N__58549;
    wire N__58546;
    wire N__58543;
    wire N__58540;
    wire N__58537;
    wire N__58534;
    wire N__58531;
    wire N__58528;
    wire N__58525;
    wire N__58522;
    wire N__58519;
    wire N__58518;
    wire N__58517;
    wire N__58510;
    wire N__58507;
    wire N__58504;
    wire N__58501;
    wire N__58498;
    wire N__58495;
    wire N__58494;
    wire N__58491;
    wire N__58490;
    wire N__58483;
    wire N__58480;
    wire N__58479;
    wire N__58474;
    wire N__58471;
    wire N__58470;
    wire N__58467;
    wire N__58464;
    wire N__58459;
    wire N__58458;
    wire N__58455;
    wire N__58452;
    wire N__58451;
    wire N__58450;
    wire N__58445;
    wire N__58442;
    wire N__58439;
    wire N__58432;
    wire N__58429;
    wire N__58426;
    wire N__58425;
    wire N__58422;
    wire N__58419;
    wire N__58414;
    wire N__58413;
    wire N__58410;
    wire N__58407;
    wire N__58402;
    wire N__58401;
    wire N__58398;
    wire N__58395;
    wire N__58390;
    wire N__58387;
    wire N__58384;
    wire N__58381;
    wire N__58378;
    wire N__58375;
    wire N__58372;
    wire N__58369;
    wire N__58366;
    wire N__58363;
    wire N__58360;
    wire N__58357;
    wire N__58354;
    wire N__58351;
    wire N__58348;
    wire N__58345;
    wire N__58342;
    wire N__58339;
    wire N__58336;
    wire N__58335;
    wire N__58332;
    wire N__58329;
    wire N__58324;
    wire N__58321;
    wire N__58320;
    wire N__58317;
    wire N__58314;
    wire N__58311;
    wire N__58306;
    wire N__58305;
    wire N__58302;
    wire N__58299;
    wire N__58296;
    wire N__58291;
    wire N__58288;
    wire N__58285;
    wire N__58282;
    wire N__58279;
    wire N__58276;
    wire N__58273;
    wire N__58270;
    wire N__58267;
    wire N__58264;
    wire N__58261;
    wire N__58258;
    wire N__58255;
    wire N__58252;
    wire N__58251;
    wire N__58248;
    wire N__58245;
    wire N__58240;
    wire N__58239;
    wire N__58236;
    wire N__58233;
    wire N__58228;
    wire N__58227;
    wire N__58226;
    wire N__58223;
    wire N__58220;
    wire N__58219;
    wire N__58216;
    wire N__58213;
    wire N__58210;
    wire N__58207;
    wire N__58198;
    wire N__58197;
    wire N__58194;
    wire N__58191;
    wire N__58186;
    wire N__58185;
    wire N__58184;
    wire N__58177;
    wire N__58174;
    wire N__58173;
    wire N__58170;
    wire N__58167;
    wire N__58164;
    wire N__58159;
    wire N__58156;
    wire N__58153;
    wire N__58150;
    wire N__58147;
    wire N__58146;
    wire N__58143;
    wire N__58140;
    wire N__58135;
    wire N__58134;
    wire N__58131;
    wire N__58128;
    wire N__58125;
    wire N__58122;
    wire N__58119;
    wire N__58116;
    wire N__58113;
    wire N__58110;
    wire N__58105;
    wire N__58102;
    wire N__58101;
    wire N__58098;
    wire N__58095;
    wire N__58092;
    wire N__58089;
    wire N__58084;
    wire N__58083;
    wire N__58080;
    wire N__58077;
    wire N__58074;
    wire N__58071;
    wire N__58068;
    wire N__58065;
    wire N__58060;
    wire N__58057;
    wire N__58056;
    wire N__58053;
    wire N__58050;
    wire N__58047;
    wire N__58044;
    wire N__58041;
    wire N__58038;
    wire N__58035;
    wire N__58032;
    wire N__58027;
    wire N__58024;
    wire N__58021;
    wire N__58020;
    wire N__58019;
    wire N__58018;
    wire N__58015;
    wire N__58012;
    wire N__58007;
    wire N__58000;
    wire N__57997;
    wire N__57994;
    wire N__57991;
    wire N__57988;
    wire N__57987;
    wire N__57984;
    wire N__57981;
    wire N__57980;
    wire N__57977;
    wire N__57974;
    wire N__57971;
    wire N__57968;
    wire N__57963;
    wire N__57962;
    wire N__57957;
    wire N__57954;
    wire N__57949;
    wire N__57946;
    wire N__57943;
    wire N__57942;
    wire N__57939;
    wire N__57936;
    wire N__57931;
    wire N__57930;
    wire N__57925;
    wire N__57924;
    wire N__57923;
    wire N__57922;
    wire N__57921;
    wire N__57920;
    wire N__57919;
    wire N__57918;
    wire N__57917;
    wire N__57914;
    wire N__57897;
    wire N__57896;
    wire N__57895;
    wire N__57894;
    wire N__57893;
    wire N__57892;
    wire N__57891;
    wire N__57886;
    wire N__57873;
    wire N__57868;
    wire N__57865;
    wire N__57862;
    wire N__57859;
    wire N__57856;
    wire N__57853;
    wire N__57850;
    wire N__57847;
    wire N__57844;
    wire N__57841;
    wire N__57838;
    wire N__57835;
    wire N__57832;
    wire N__57829;
    wire N__57826;
    wire N__57823;
    wire N__57820;
    wire N__57819;
    wire N__57816;
    wire N__57813;
    wire N__57810;
    wire N__57805;
    wire N__57802;
    wire N__57799;
    wire N__57796;
    wire N__57793;
    wire N__57790;
    wire N__57789;
    wire N__57786;
    wire N__57783;
    wire N__57780;
    wire N__57775;
    wire N__57772;
    wire N__57769;
    wire N__57766;
    wire N__57763;
    wire N__57760;
    wire N__57757;
    wire N__57754;
    wire N__57753;
    wire N__57752;
    wire N__57751;
    wire N__57750;
    wire N__57749;
    wire N__57748;
    wire N__57745;
    wire N__57740;
    wire N__57737;
    wire N__57732;
    wire N__57731;
    wire N__57728;
    wire N__57725;
    wire N__57722;
    wire N__57717;
    wire N__57712;
    wire N__57711;
    wire N__57710;
    wire N__57709;
    wire N__57708;
    wire N__57707;
    wire N__57706;
    wire N__57703;
    wire N__57700;
    wire N__57697;
    wire N__57694;
    wire N__57691;
    wire N__57680;
    wire N__57667;
    wire N__57666;
    wire N__57663;
    wire N__57660;
    wire N__57655;
    wire N__57652;
    wire N__57649;
    wire N__57648;
    wire N__57647;
    wire N__57646;
    wire N__57645;
    wire N__57642;
    wire N__57639;
    wire N__57638;
    wire N__57637;
    wire N__57634;
    wire N__57631;
    wire N__57630;
    wire N__57629;
    wire N__57626;
    wire N__57625;
    wire N__57622;
    wire N__57619;
    wire N__57610;
    wire N__57607;
    wire N__57600;
    wire N__57599;
    wire N__57596;
    wire N__57591;
    wire N__57588;
    wire N__57585;
    wire N__57584;
    wire N__57583;
    wire N__57580;
    wire N__57577;
    wire N__57574;
    wire N__57571;
    wire N__57568;
    wire N__57561;
    wire N__57558;
    wire N__57553;
    wire N__57548;
    wire N__57545;
    wire N__57540;
    wire N__57537;
    wire N__57534;
    wire N__57531;
    wire N__57528;
    wire N__57525;
    wire N__57522;
    wire N__57517;
    wire N__57514;
    wire N__57513;
    wire N__57510;
    wire N__57507;
    wire N__57502;
    wire N__57501;
    wire N__57500;
    wire N__57497;
    wire N__57492;
    wire N__57491;
    wire N__57488;
    wire N__57485;
    wire N__57482;
    wire N__57479;
    wire N__57474;
    wire N__57471;
    wire N__57468;
    wire N__57463;
    wire N__57460;
    wire N__57457;
    wire N__57454;
    wire N__57451;
    wire N__57448;
    wire N__57445;
    wire N__57444;
    wire N__57441;
    wire N__57438;
    wire N__57435;
    wire N__57432;
    wire N__57429;
    wire N__57426;
    wire N__57423;
    wire N__57418;
    wire N__57415;
    wire N__57412;
    wire N__57409;
    wire N__57406;
    wire N__57403;
    wire N__57400;
    wire N__57399;
    wire N__57398;
    wire N__57397;
    wire N__57394;
    wire N__57393;
    wire N__57392;
    wire N__57389;
    wire N__57388;
    wire N__57387;
    wire N__57386;
    wire N__57385;
    wire N__57382;
    wire N__57379;
    wire N__57376;
    wire N__57371;
    wire N__57362;
    wire N__57359;
    wire N__57356;
    wire N__57347;
    wire N__57344;
    wire N__57341;
    wire N__57334;
    wire N__57333;
    wire N__57330;
    wire N__57327;
    wire N__57322;
    wire N__57319;
    wire N__57316;
    wire N__57315;
    wire N__57312;
    wire N__57309;
    wire N__57304;
    wire N__57303;
    wire N__57300;
    wire N__57297;
    wire N__57294;
    wire N__57291;
    wire N__57288;
    wire N__57285;
    wire N__57282;
    wire N__57279;
    wire N__57276;
    wire N__57273;
    wire N__57270;
    wire N__57267;
    wire N__57262;
    wire N__57261;
    wire N__57258;
    wire N__57255;
    wire N__57252;
    wire N__57249;
    wire N__57246;
    wire N__57243;
    wire N__57240;
    wire N__57237;
    wire N__57234;
    wire N__57231;
    wire N__57226;
    wire N__57225;
    wire N__57224;
    wire N__57223;
    wire N__57222;
    wire N__57215;
    wire N__57210;
    wire N__57205;
    wire N__57204;
    wire N__57203;
    wire N__57198;
    wire N__57195;
    wire N__57192;
    wire N__57187;
    wire N__57184;
    wire N__57181;
    wire N__57178;
    wire N__57175;
    wire N__57172;
    wire N__57169;
    wire N__57166;
    wire N__57163;
    wire N__57160;
    wire N__57157;
    wire N__57156;
    wire N__57151;
    wire N__57148;
    wire N__57145;
    wire N__57142;
    wire N__57139;
    wire N__57136;
    wire N__57133;
    wire N__57130;
    wire N__57127;
    wire N__57124;
    wire N__57121;
    wire N__57120;
    wire N__57115;
    wire N__57112;
    wire N__57111;
    wire N__57108;
    wire N__57105;
    wire N__57100;
    wire N__57097;
    wire N__57094;
    wire N__57091;
    wire N__57088;
    wire N__57085;
    wire N__57082;
    wire N__57081;
    wire N__57078;
    wire N__57075;
    wire N__57070;
    wire N__57067;
    wire N__57064;
    wire N__57061;
    wire N__57060;
    wire N__57057;
    wire N__57054;
    wire N__57049;
    wire N__57046;
    wire N__57043;
    wire N__57042;
    wire N__57039;
    wire N__57036;
    wire N__57031;
    wire N__57028;
    wire N__57025;
    wire N__57024;
    wire N__57021;
    wire N__57018;
    wire N__57013;
    wire N__57010;
    wire N__57007;
    wire N__57004;
    wire N__57003;
    wire N__57000;
    wire N__56997;
    wire N__56992;
    wire N__56989;
    wire N__56986;
    wire N__56983;
    wire N__56982;
    wire N__56979;
    wire N__56976;
    wire N__56971;
    wire N__56968;
    wire N__56965;
    wire N__56962;
    wire N__56959;
    wire N__56956;
    wire N__56955;
    wire N__56952;
    wire N__56949;
    wire N__56944;
    wire N__56941;
    wire N__56940;
    wire N__56937;
    wire N__56934;
    wire N__56929;
    wire N__56926;
    wire N__56923;
    wire N__56922;
    wire N__56919;
    wire N__56916;
    wire N__56911;
    wire N__56908;
    wire N__56905;
    wire N__56902;
    wire N__56899;
    wire N__56898;
    wire N__56895;
    wire N__56892;
    wire N__56887;
    wire N__56884;
    wire N__56881;
    wire N__56878;
    wire N__56875;
    wire N__56872;
    wire N__56871;
    wire N__56868;
    wire N__56863;
    wire N__56860;
    wire N__56859;
    wire N__56856;
    wire N__56851;
    wire N__56848;
    wire N__56847;
    wire N__56844;
    wire N__56839;
    wire N__56836;
    wire N__56833;
    wire N__56832;
    wire N__56829;
    wire N__56826;
    wire N__56823;
    wire N__56820;
    wire N__56815;
    wire N__56812;
    wire N__56811;
    wire N__56808;
    wire N__56805;
    wire N__56800;
    wire N__56797;
    wire N__56794;
    wire N__56793;
    wire N__56790;
    wire N__56787;
    wire N__56782;
    wire N__56779;
    wire N__56776;
    wire N__56773;
    wire N__56770;
    wire N__56767;
    wire N__56764;
    wire N__56763;
    wire N__56760;
    wire N__56757;
    wire N__56752;
    wire N__56749;
    wire N__56748;
    wire N__56745;
    wire N__56742;
    wire N__56737;
    wire N__56736;
    wire N__56733;
    wire N__56728;
    wire N__56725;
    wire N__56724;
    wire N__56721;
    wire N__56718;
    wire N__56715;
    wire N__56710;
    wire N__56709;
    wire N__56704;
    wire N__56701;
    wire N__56698;
    wire N__56697;
    wire N__56694;
    wire N__56691;
    wire N__56686;
    wire N__56683;
    wire N__56680;
    wire N__56679;
    wire N__56676;
    wire N__56673;
    wire N__56668;
    wire N__56667;
    wire N__56662;
    wire N__56659;
    wire N__56656;
    wire N__56653;
    wire N__56652;
    wire N__56647;
    wire N__56644;
    wire N__56643;
    wire N__56640;
    wire N__56637;
    wire N__56632;
    wire N__56629;
    wire N__56626;
    wire N__56625;
    wire N__56624;
    wire N__56621;
    wire N__56620;
    wire N__56619;
    wire N__56616;
    wire N__56615;
    wire N__56614;
    wire N__56613;
    wire N__56610;
    wire N__56607;
    wire N__56606;
    wire N__56605;
    wire N__56604;
    wire N__56603;
    wire N__56600;
    wire N__56599;
    wire N__56596;
    wire N__56595;
    wire N__56594;
    wire N__56593;
    wire N__56592;
    wire N__56589;
    wire N__56586;
    wire N__56583;
    wire N__56580;
    wire N__56575;
    wire N__56572;
    wire N__56571;
    wire N__56570;
    wire N__56569;
    wire N__56568;
    wire N__56567;
    wire N__56566;
    wire N__56565;
    wire N__56558;
    wire N__56557;
    wire N__56556;
    wire N__56555;
    wire N__56550;
    wire N__56549;
    wire N__56548;
    wire N__56547;
    wire N__56546;
    wire N__56543;
    wire N__56538;
    wire N__56535;
    wire N__56532;
    wire N__56527;
    wire N__56524;
    wire N__56521;
    wire N__56520;
    wire N__56519;
    wire N__56518;
    wire N__56517;
    wire N__56516;
    wire N__56515;
    wire N__56514;
    wire N__56513;
    wire N__56512;
    wire N__56511;
    wire N__56510;
    wire N__56509;
    wire N__56508;
    wire N__56507;
    wire N__56504;
    wire N__56499;
    wire N__56494;
    wire N__56491;
    wire N__56490;
    wire N__56489;
    wire N__56488;
    wire N__56483;
    wire N__56480;
    wire N__56477;
    wire N__56476;
    wire N__56475;
    wire N__56474;
    wire N__56473;
    wire N__56466;
    wire N__56463;
    wire N__56460;
    wire N__56459;
    wire N__56458;
    wire N__56457;
    wire N__56450;
    wire N__56443;
    wire N__56438;
    wire N__56433;
    wire N__56430;
    wire N__56421;
    wire N__56416;
    wire N__56415;
    wire N__56410;
    wire N__56409;
    wire N__56408;
    wire N__56403;
    wire N__56400;
    wire N__56395;
    wire N__56388;
    wire N__56383;
    wire N__56378;
    wire N__56375;
    wire N__56370;
    wire N__56367;
    wire N__56364;
    wire N__56359;
    wire N__56354;
    wire N__56353;
    wire N__56352;
    wire N__56343;
    wire N__56340;
    wire N__56333;
    wire N__56332;
    wire N__56331;
    wire N__56330;
    wire N__56329;
    wire N__56322;
    wire N__56319;
    wire N__56316;
    wire N__56313;
    wire N__56310;
    wire N__56301;
    wire N__56298;
    wire N__56295;
    wire N__56290;
    wire N__56281;
    wire N__56278;
    wire N__56275;
    wire N__56268;
    wire N__56263;
    wire N__56258;
    wire N__56255;
    wire N__56250;
    wire N__56243;
    wire N__56234;
    wire N__56227;
    wire N__56212;
    wire N__56209;
    wire N__56206;
    wire N__56203;
    wire N__56202;
    wire N__56199;
    wire N__56196;
    wire N__56191;
    wire N__56188;
    wire N__56187;
    wire N__56184;
    wire N__56181;
    wire N__56178;
    wire N__56175;
    wire N__56170;
    wire N__56167;
    wire N__56164;
    wire N__56161;
    wire N__56160;
    wire N__56155;
    wire N__56152;
    wire N__56149;
    wire N__56146;
    wire N__56143;
    wire N__56140;
    wire N__56139;
    wire N__56136;
    wire N__56133;
    wire N__56128;
    wire N__56127;
    wire N__56122;
    wire N__56119;
    wire N__56116;
    wire N__56113;
    wire N__56110;
    wire N__56109;
    wire N__56106;
    wire N__56103;
    wire N__56098;
    wire N__56095;
    wire N__56092;
    wire N__56089;
    wire N__56086;
    wire N__56085;
    wire N__56082;
    wire N__56079;
    wire N__56074;
    wire N__56073;
    wire N__56068;
    wire N__56065;
    wire N__56062;
    wire N__56061;
    wire N__56058;
    wire N__56055;
    wire N__56050;
    wire N__56047;
    wire N__56046;
    wire N__56043;
    wire N__56040;
    wire N__56035;
    wire N__56034;
    wire N__56029;
    wire N__56026;
    wire N__56023;
    wire N__56020;
    wire N__56017;
    wire N__56014;
    wire N__56011;
    wire N__56008;
    wire N__56005;
    wire N__56002;
    wire N__55999;
    wire N__55996;
    wire N__55993;
    wire N__55990;
    wire N__55987;
    wire N__55984;
    wire N__55981;
    wire N__55980;
    wire N__55977;
    wire N__55974;
    wire N__55969;
    wire N__55966;
    wire N__55963;
    wire N__55962;
    wire N__55959;
    wire N__55956;
    wire N__55951;
    wire N__55948;
    wire N__55947;
    wire N__55944;
    wire N__55941;
    wire N__55938;
    wire N__55935;
    wire N__55930;
    wire N__55927;
    wire N__55926;
    wire N__55923;
    wire N__55920;
    wire N__55917;
    wire N__55914;
    wire N__55909;
    wire N__55906;
    wire N__55903;
    wire N__55900;
    wire N__55899;
    wire N__55896;
    wire N__55893;
    wire N__55890;
    wire N__55887;
    wire N__55882;
    wire N__55879;
    wire N__55876;
    wire N__55873;
    wire N__55870;
    wire N__55867;
    wire N__55864;
    wire N__55861;
    wire N__55858;
    wire N__55855;
    wire N__55852;
    wire N__55849;
    wire N__55846;
    wire N__55843;
    wire N__55842;
    wire N__55839;
    wire N__55836;
    wire N__55831;
    wire N__55828;
    wire N__55827;
    wire N__55824;
    wire N__55821;
    wire N__55816;
    wire N__55813;
    wire N__55810;
    wire N__55807;
    wire N__55804;
    wire N__55801;
    wire N__55800;
    wire N__55797;
    wire N__55794;
    wire N__55789;
    wire N__55786;
    wire N__55785;
    wire N__55782;
    wire N__55779;
    wire N__55774;
    wire N__55771;
    wire N__55768;
    wire N__55767;
    wire N__55766;
    wire N__55765;
    wire N__55764;
    wire N__55763;
    wire N__55760;
    wire N__55757;
    wire N__55756;
    wire N__55753;
    wire N__55752;
    wire N__55749;
    wire N__55748;
    wire N__55745;
    wire N__55744;
    wire N__55741;
    wire N__55740;
    wire N__55737;
    wire N__55734;
    wire N__55717;
    wire N__55714;
    wire N__55705;
    wire N__55702;
    wire N__55701;
    wire N__55698;
    wire N__55695;
    wire N__55692;
    wire N__55687;
    wire N__55684;
    wire N__55681;
    wire N__55678;
    wire N__55675;
    wire N__55672;
    wire N__55669;
    wire N__55666;
    wire N__55663;
    wire N__55660;
    wire N__55657;
    wire N__55654;
    wire N__55651;
    wire N__55648;
    wire N__55645;
    wire N__55644;
    wire N__55639;
    wire N__55636;
    wire N__55633;
    wire N__55632;
    wire N__55629;
    wire N__55626;
    wire N__55621;
    wire N__55618;
    wire N__55615;
    wire N__55614;
    wire N__55613;
    wire N__55612;
    wire N__55609;
    wire N__55608;
    wire N__55607;
    wire N__55604;
    wire N__55603;
    wire N__55600;
    wire N__55599;
    wire N__55596;
    wire N__55591;
    wire N__55590;
    wire N__55589;
    wire N__55588;
    wire N__55587;
    wire N__55586;
    wire N__55585;
    wire N__55584;
    wire N__55583;
    wire N__55582;
    wire N__55581;
    wire N__55580;
    wire N__55579;
    wire N__55578;
    wire N__55577;
    wire N__55574;
    wire N__55571;
    wire N__55562;
    wire N__55559;
    wire N__55554;
    wire N__55551;
    wire N__55544;
    wire N__55533;
    wire N__55526;
    wire N__55507;
    wire N__55504;
    wire N__55501;
    wire N__55498;
    wire N__55497;
    wire N__55494;
    wire N__55493;
    wire N__55490;
    wire N__55489;
    wire N__55488;
    wire N__55487;
    wire N__55484;
    wire N__55483;
    wire N__55482;
    wire N__55481;
    wire N__55480;
    wire N__55479;
    wire N__55478;
    wire N__55467;
    wire N__55466;
    wire N__55465;
    wire N__55464;
    wire N__55463;
    wire N__55462;
    wire N__55461;
    wire N__55460;
    wire N__55459;
    wire N__55456;
    wire N__55447;
    wire N__55446;
    wire N__55443;
    wire N__55440;
    wire N__55439;
    wire N__55438;
    wire N__55437;
    wire N__55436;
    wire N__55435;
    wire N__55434;
    wire N__55433;
    wire N__55432;
    wire N__55431;
    wire N__55430;
    wire N__55427;
    wire N__55420;
    wire N__55417;
    wire N__55408;
    wire N__55403;
    wire N__55400;
    wire N__55397;
    wire N__55392;
    wire N__55383;
    wire N__55372;
    wire N__55351;
    wire N__55348;
    wire N__55345;
    wire N__55342;
    wire N__55341;
    wire N__55338;
    wire N__55335;
    wire N__55330;
    wire N__55327;
    wire N__55324;
    wire N__55323;
    wire N__55320;
    wire N__55317;
    wire N__55312;
    wire N__55309;
    wire N__55306;
    wire N__55305;
    wire N__55302;
    wire N__55299;
    wire N__55294;
    wire N__55291;
    wire N__55288;
    wire N__55285;
    wire N__55284;
    wire N__55281;
    wire N__55278;
    wire N__55273;
    wire N__55270;
    wire N__55269;
    wire N__55266;
    wire N__55265;
    wire N__55262;
    wire N__55261;
    wire N__55260;
    wire N__55259;
    wire N__55258;
    wire N__55257;
    wire N__55256;
    wire N__55255;
    wire N__55254;
    wire N__55253;
    wire N__55252;
    wire N__55251;
    wire N__55244;
    wire N__55239;
    wire N__55236;
    wire N__55235;
    wire N__55234;
    wire N__55233;
    wire N__55232;
    wire N__55231;
    wire N__55230;
    wire N__55219;
    wire N__55218;
    wire N__55215;
    wire N__55214;
    wire N__55211;
    wire N__55210;
    wire N__55207;
    wire N__55204;
    wire N__55201;
    wire N__55192;
    wire N__55189;
    wire N__55186;
    wire N__55185;
    wire N__55184;
    wire N__55183;
    wire N__55180;
    wire N__55179;
    wire N__55178;
    wire N__55177;
    wire N__55176;
    wire N__55173;
    wire N__55170;
    wire N__55161;
    wire N__55152;
    wire N__55145;
    wire N__55138;
    wire N__55129;
    wire N__55114;
    wire N__55111;
    wire N__55108;
    wire N__55105;
    wire N__55102;
    wire N__55099;
    wire N__55096;
    wire N__55093;
    wire N__55090;
    wire N__55087;
    wire N__55084;
    wire N__55081;
    wire N__55078;
    wire N__55075;
    wire N__55074;
    wire N__55073;
    wire N__55072;
    wire N__55071;
    wire N__55070;
    wire N__55069;
    wire N__55068;
    wire N__55067;
    wire N__55066;
    wire N__55065;
    wire N__55064;
    wire N__55063;
    wire N__55062;
    wire N__55061;
    wire N__55060;
    wire N__55059;
    wire N__55052;
    wire N__55051;
    wire N__55050;
    wire N__55049;
    wire N__55048;
    wire N__55047;
    wire N__55038;
    wire N__55029;
    wire N__55016;
    wire N__55015;
    wire N__55014;
    wire N__55013;
    wire N__55012;
    wire N__55011;
    wire N__55010;
    wire N__55009;
    wire N__55008;
    wire N__55005;
    wire N__54998;
    wire N__54993;
    wire N__54986;
    wire N__54977;
    wire N__54968;
    wire N__54955;
    wire N__54952;
    wire N__54951;
    wire N__54950;
    wire N__54949;
    wire N__54946;
    wire N__54945;
    wire N__54942;
    wire N__54937;
    wire N__54934;
    wire N__54929;
    wire N__54928;
    wire N__54927;
    wire N__54926;
    wire N__54923;
    wire N__54920;
    wire N__54917;
    wire N__54914;
    wire N__54909;
    wire N__54898;
    wire N__54895;
    wire N__54892;
    wire N__54889;
    wire N__54886;
    wire N__54885;
    wire N__54882;
    wire N__54879;
    wire N__54874;
    wire N__54871;
    wire N__54870;
    wire N__54869;
    wire N__54868;
    wire N__54865;
    wire N__54862;
    wire N__54857;
    wire N__54850;
    wire N__54847;
    wire N__54846;
    wire N__54845;
    wire N__54844;
    wire N__54841;
    wire N__54838;
    wire N__54835;
    wire N__54832;
    wire N__54823;
    wire N__54820;
    wire N__54817;
    wire N__54816;
    wire N__54815;
    wire N__54814;
    wire N__54811;
    wire N__54808;
    wire N__54803;
    wire N__54796;
    wire N__54793;
    wire N__54792;
    wire N__54791;
    wire N__54790;
    wire N__54787;
    wire N__54784;
    wire N__54781;
    wire N__54778;
    wire N__54769;
    wire N__54766;
    wire N__54763;
    wire N__54760;
    wire N__54757;
    wire N__54756;
    wire N__54753;
    wire N__54752;
    wire N__54749;
    wire N__54742;
    wire N__54739;
    wire N__54736;
    wire N__54733;
    wire N__54730;
    wire N__54729;
    wire N__54726;
    wire N__54723;
    wire N__54718;
    wire N__54717;
    wire N__54714;
    wire N__54709;
    wire N__54706;
    wire N__54705;
    wire N__54702;
    wire N__54699;
    wire N__54694;
    wire N__54691;
    wire N__54690;
    wire N__54685;
    wire N__54682;
    wire N__54679;
    wire N__54678;
    wire N__54675;
    wire N__54672;
    wire N__54667;
    wire N__54664;
    wire N__54661;
    wire N__54658;
    wire N__54655;
    wire N__54652;
    wire N__54649;
    wire N__54646;
    wire N__54643;
    wire N__54640;
    wire N__54637;
    wire N__54634;
    wire N__54631;
    wire N__54628;
    wire N__54625;
    wire N__54622;
    wire N__54621;
    wire N__54618;
    wire N__54615;
    wire N__54610;
    wire N__54607;
    wire N__54604;
    wire N__54601;
    wire N__54598;
    wire N__54597;
    wire N__54594;
    wire N__54591;
    wire N__54588;
    wire N__54583;
    wire N__54580;
    wire N__54577;
    wire N__54576;
    wire N__54573;
    wire N__54570;
    wire N__54567;
    wire N__54564;
    wire N__54561;
    wire N__54556;
    wire N__54553;
    wire N__54550;
    wire N__54547;
    wire N__54544;
    wire N__54541;
    wire N__54538;
    wire N__54535;
    wire N__54532;
    wire N__54529;
    wire N__54526;
    wire N__54523;
    wire N__54520;
    wire N__54517;
    wire N__54514;
    wire N__54513;
    wire N__54510;
    wire N__54507;
    wire N__54504;
    wire N__54501;
    wire N__54496;
    wire N__54493;
    wire N__54492;
    wire N__54489;
    wire N__54486;
    wire N__54483;
    wire N__54482;
    wire N__54479;
    wire N__54476;
    wire N__54473;
    wire N__54470;
    wire N__54467;
    wire N__54462;
    wire N__54457;
    wire N__54454;
    wire N__54451;
    wire N__54448;
    wire N__54445;
    wire N__54442;
    wire N__54441;
    wire N__54438;
    wire N__54435;
    wire N__54432;
    wire N__54427;
    wire N__54424;
    wire N__54421;
    wire N__54420;
    wire N__54417;
    wire N__54414;
    wire N__54411;
    wire N__54408;
    wire N__54405;
    wire N__54400;
    wire N__54397;
    wire N__54394;
    wire N__54393;
    wire N__54388;
    wire N__54385;
    wire N__54384;
    wire N__54379;
    wire N__54376;
    wire N__54375;
    wire N__54372;
    wire N__54367;
    wire N__54364;
    wire N__54363;
    wire N__54358;
    wire N__54355;
    wire N__54352;
    wire N__54351;
    wire N__54350;
    wire N__54349;
    wire N__54348;
    wire N__54345;
    wire N__54340;
    wire N__54335;
    wire N__54328;
    wire N__54327;
    wire N__54326;
    wire N__54325;
    wire N__54324;
    wire N__54323;
    wire N__54322;
    wire N__54319;
    wire N__54314;
    wire N__54305;
    wire N__54298;
    wire N__54295;
    wire N__54292;
    wire N__54291;
    wire N__54288;
    wire N__54285;
    wire N__54282;
    wire N__54279;
    wire N__54274;
    wire N__54271;
    wire N__54270;
    wire N__54267;
    wire N__54264;
    wire N__54259;
    wire N__54256;
    wire N__54253;
    wire N__54252;
    wire N__54249;
    wire N__54246;
    wire N__54243;
    wire N__54240;
    wire N__54235;
    wire N__54232;
    wire N__54229;
    wire N__54228;
    wire N__54225;
    wire N__54220;
    wire N__54217;
    wire N__54214;
    wire N__54213;
    wire N__54208;
    wire N__54205;
    wire N__54204;
    wire N__54201;
    wire N__54198;
    wire N__54195;
    wire N__54190;
    wire N__54187;
    wire N__54186;
    wire N__54183;
    wire N__54180;
    wire N__54175;
    wire N__54172;
    wire N__54169;
    wire N__54166;
    wire N__54163;
    wire N__54160;
    wire N__54157;
    wire N__54156;
    wire N__54153;
    wire N__54150;
    wire N__54145;
    wire N__54142;
    wire N__54139;
    wire N__54136;
    wire N__54133;
    wire N__54130;
    wire N__54127;
    wire N__54126;
    wire N__54121;
    wire N__54118;
    wire N__54117;
    wire N__54112;
    wire N__54109;
    wire N__54108;
    wire N__54105;
    wire N__54102;
    wire N__54099;
    wire N__54098;
    wire N__54095;
    wire N__54094;
    wire N__54093;
    wire N__54090;
    wire N__54087;
    wire N__54086;
    wire N__54083;
    wire N__54082;
    wire N__54081;
    wire N__54080;
    wire N__54077;
    wire N__54074;
    wire N__54073;
    wire N__54072;
    wire N__54069;
    wire N__54066;
    wire N__54065;
    wire N__54064;
    wire N__54063;
    wire N__54060;
    wire N__54057;
    wire N__54054;
    wire N__54051;
    wire N__54048;
    wire N__54045;
    wire N__54042;
    wire N__54041;
    wire N__54038;
    wire N__54035;
    wire N__54030;
    wire N__54029;
    wire N__54026;
    wire N__54021;
    wire N__54018;
    wire N__54015;
    wire N__54012;
    wire N__54007;
    wire N__54004;
    wire N__54001;
    wire N__53998;
    wire N__53995;
    wire N__53990;
    wire N__53987;
    wire N__53984;
    wire N__53979;
    wire N__53976;
    wire N__53973;
    wire N__53966;
    wire N__53959;
    wire N__53944;
    wire N__53943;
    wire N__53940;
    wire N__53937;
    wire N__53932;
    wire N__53929;
    wire N__53926;
    wire N__53923;
    wire N__53922;
    wire N__53919;
    wire N__53916;
    wire N__53911;
    wire N__53908;
    wire N__53907;
    wire N__53904;
    wire N__53901;
    wire N__53896;
    wire N__53893;
    wire N__53890;
    wire N__53889;
    wire N__53886;
    wire N__53883;
    wire N__53880;
    wire N__53877;
    wire N__53872;
    wire N__53869;
    wire N__53866;
    wire N__53865;
    wire N__53862;
    wire N__53859;
    wire N__53854;
    wire N__53851;
    wire N__53850;
    wire N__53845;
    wire N__53842;
    wire N__53839;
    wire N__53838;
    wire N__53835;
    wire N__53832;
    wire N__53827;
    wire N__53824;
    wire N__53821;
    wire N__53820;
    wire N__53817;
    wire N__53814;
    wire N__53809;
    wire N__53806;
    wire N__53805;
    wire N__53802;
    wire N__53799;
    wire N__53794;
    wire N__53791;
    wire N__53790;
    wire N__53787;
    wire N__53784;
    wire N__53781;
    wire N__53778;
    wire N__53773;
    wire N__53770;
    wire N__53767;
    wire N__53764;
    wire N__53761;
    wire N__53758;
    wire N__53757;
    wire N__53754;
    wire N__53751;
    wire N__53746;
    wire N__53743;
    wire N__53740;
    wire N__53737;
    wire N__53734;
    wire N__53731;
    wire N__53730;
    wire N__53725;
    wire N__53722;
    wire N__53719;
    wire N__53716;
    wire N__53713;
    wire N__53712;
    wire N__53709;
    wire N__53706;
    wire N__53701;
    wire N__53700;
    wire N__53697;
    wire N__53694;
    wire N__53689;
    wire N__53686;
    wire N__53683;
    wire N__53680;
    wire N__53679;
    wire N__53676;
    wire N__53673;
    wire N__53668;
    wire N__53667;
    wire N__53662;
    wire N__53659;
    wire N__53656;
    wire N__53655;
    wire N__53650;
    wire N__53647;
    wire N__53644;
    wire N__53641;
    wire N__53640;
    wire N__53637;
    wire N__53634;
    wire N__53629;
    wire N__53626;
    wire N__53623;
    wire N__53620;
    wire N__53617;
    wire N__53616;
    wire N__53611;
    wire N__53608;
    wire N__53607;
    wire N__53604;
    wire N__53601;
    wire N__53596;
    wire N__53593;
    wire N__53590;
    wire N__53589;
    wire N__53586;
    wire N__53583;
    wire N__53578;
    wire N__53575;
    wire N__53572;
    wire N__53571;
    wire N__53568;
    wire N__53565;
    wire N__53560;
    wire N__53557;
    wire N__53556;
    wire N__53553;
    wire N__53550;
    wire N__53545;
    wire N__53542;
    wire N__53539;
    wire N__53536;
    wire N__53533;
    wire N__53530;
    wire N__53527;
    wire N__53524;
    wire N__53521;
    wire N__53518;
    wire N__53515;
    wire N__53512;
    wire N__53509;
    wire N__53506;
    wire N__53503;
    wire N__53500;
    wire N__53497;
    wire N__53494;
    wire N__53491;
    wire N__53488;
    wire N__53485;
    wire N__53482;
    wire N__53479;
    wire N__53476;
    wire N__53473;
    wire N__53470;
    wire N__53467;
    wire N__53466;
    wire N__53463;
    wire N__53460;
    wire N__53455;
    wire N__53452;
    wire N__53449;
    wire N__53448;
    wire N__53445;
    wire N__53442;
    wire N__53437;
    wire N__53434;
    wire N__53433;
    wire N__53428;
    wire N__53425;
    wire N__53422;
    wire N__53419;
    wire N__53416;
    wire N__53415;
    wire N__53412;
    wire N__53409;
    wire N__53406;
    wire N__53403;
    wire N__53398;
    wire N__53395;
    wire N__53392;
    wire N__53391;
    wire N__53388;
    wire N__53383;
    wire N__53380;
    wire N__53379;
    wire N__53376;
    wire N__53373;
    wire N__53368;
    wire N__53365;
    wire N__53362;
    wire N__53359;
    wire N__53358;
    wire N__53355;
    wire N__53352;
    wire N__53347;
    wire N__53346;
    wire N__53343;
    wire N__53340;
    wire N__53337;
    wire N__53332;
    wire N__53331;
    wire N__53328;
    wire N__53325;
    wire N__53322;
    wire N__53317;
    wire N__53314;
    wire N__53311;
    wire N__53308;
    wire N__53305;
    wire N__53302;
    wire N__53299;
    wire N__53296;
    wire N__53293;
    wire N__53290;
    wire N__53287;
    wire N__53284;
    wire N__53281;
    wire N__53278;
    wire N__53275;
    wire N__53272;
    wire N__53271;
    wire N__53268;
    wire N__53265;
    wire N__53260;
    wire N__53259;
    wire N__53256;
    wire N__53253;
    wire N__53248;
    wire N__53247;
    wire N__53242;
    wire N__53239;
    wire N__53236;
    wire N__53233;
    wire N__53230;
    wire N__53229;
    wire N__53226;
    wire N__53223;
    wire N__53218;
    wire N__53215;
    wire N__53212;
    wire N__53209;
    wire N__53208;
    wire N__53205;
    wire N__53202;
    wire N__53197;
    wire N__53194;
    wire N__53191;
    wire N__53190;
    wire N__53185;
    wire N__53182;
    wire N__53179;
    wire N__53176;
    wire N__53173;
    wire N__53172;
    wire N__53169;
    wire N__53164;
    wire N__53161;
    wire N__53158;
    wire N__53155;
    wire N__53154;
    wire N__53151;
    wire N__53148;
    wire N__53145;
    wire N__53142;
    wire N__53137;
    wire N__53134;
    wire N__53133;
    wire N__53130;
    wire N__53127;
    wire N__53124;
    wire N__53121;
    wire N__53116;
    wire N__53115;
    wire N__53110;
    wire N__53107;
    wire N__53104;
    wire N__53101;
    wire N__53100;
    wire N__53097;
    wire N__53094;
    wire N__53089;
    wire N__53086;
    wire N__53083;
    wire N__53082;
    wire N__53079;
    wire N__53076;
    wire N__53073;
    wire N__53070;
    wire N__53065;
    wire N__53062;
    wire N__53059;
    wire N__53056;
    wire N__53053;
    wire N__53050;
    wire N__53047;
    wire N__53044;
    wire N__53041;
    wire N__53038;
    wire N__53035;
    wire N__53032;
    wire N__53031;
    wire N__53028;
    wire N__53025;
    wire N__53022;
    wire N__53019;
    wire N__53016;
    wire N__53013;
    wire N__53008;
    wire N__53005;
    wire N__53002;
    wire N__52999;
    wire N__52996;
    wire N__52993;
    wire N__52990;
    wire N__52987;
    wire N__52984;
    wire N__52981;
    wire N__52978;
    wire N__52977;
    wire N__52974;
    wire N__52971;
    wire N__52966;
    wire N__52963;
    wire N__52960;
    wire N__52957;
    wire N__52956;
    wire N__52951;
    wire N__52948;
    wire N__52945;
    wire N__52942;
    wire N__52939;
    wire N__52938;
    wire N__52935;
    wire N__52932;
    wire N__52927;
    wire N__52924;
    wire N__52921;
    wire N__52918;
    wire N__52915;
    wire N__52912;
    wire N__52909;
    wire N__52906;
    wire N__52903;
    wire N__52900;
    wire N__52897;
    wire N__52894;
    wire N__52891;
    wire N__52888;
    wire N__52885;
    wire N__52882;
    wire N__52879;
    wire N__52876;
    wire N__52873;
    wire N__52870;
    wire N__52867;
    wire N__52864;
    wire N__52863;
    wire N__52860;
    wire N__52857;
    wire N__52854;
    wire N__52853;
    wire N__52852;
    wire N__52847;
    wire N__52844;
    wire N__52841;
    wire N__52834;
    wire N__52831;
    wire N__52828;
    wire N__52825;
    wire N__52822;
    wire N__52819;
    wire N__52818;
    wire N__52817;
    wire N__52814;
    wire N__52809;
    wire N__52804;
    wire N__52801;
    wire N__52798;
    wire N__52797;
    wire N__52796;
    wire N__52795;
    wire N__52794;
    wire N__52793;
    wire N__52790;
    wire N__52783;
    wire N__52780;
    wire N__52777;
    wire N__52768;
    wire N__52765;
    wire N__52762;
    wire N__52759;
    wire N__52756;
    wire N__52753;
    wire N__52750;
    wire N__52747;
    wire N__52744;
    wire N__52743;
    wire N__52742;
    wire N__52739;
    wire N__52736;
    wire N__52733;
    wire N__52726;
    wire N__52723;
    wire N__52720;
    wire N__52717;
    wire N__52714;
    wire N__52711;
    wire N__52708;
    wire N__52705;
    wire N__52704;
    wire N__52701;
    wire N__52698;
    wire N__52697;
    wire N__52696;
    wire N__52693;
    wire N__52690;
    wire N__52685;
    wire N__52678;
    wire N__52675;
    wire N__52672;
    wire N__52669;
    wire N__52668;
    wire N__52663;
    wire N__52662;
    wire N__52659;
    wire N__52656;
    wire N__52651;
    wire N__52648;
    wire N__52645;
    wire N__52644;
    wire N__52641;
    wire N__52638;
    wire N__52633;
    wire N__52630;
    wire N__52627;
    wire N__52624;
    wire N__52621;
    wire N__52618;
    wire N__52615;
    wire N__52612;
    wire N__52609;
    wire N__52606;
    wire N__52603;
    wire N__52600;
    wire N__52597;
    wire N__52594;
    wire N__52591;
    wire N__52588;
    wire N__52585;
    wire N__52582;
    wire N__52579;
    wire N__52578;
    wire N__52575;
    wire N__52574;
    wire N__52573;
    wire N__52572;
    wire N__52571;
    wire N__52568;
    wire N__52563;
    wire N__52562;
    wire N__52561;
    wire N__52560;
    wire N__52559;
    wire N__52558;
    wire N__52557;
    wire N__52556;
    wire N__52553;
    wire N__52546;
    wire N__52543;
    wire N__52540;
    wire N__52527;
    wire N__52522;
    wire N__52515;
    wire N__52512;
    wire N__52509;
    wire N__52506;
    wire N__52503;
    wire N__52498;
    wire N__52495;
    wire N__52492;
    wire N__52489;
    wire N__52486;
    wire N__52483;
    wire N__52480;
    wire N__52477;
    wire N__52474;
    wire N__52471;
    wire N__52468;
    wire N__52465;
    wire N__52462;
    wire N__52459;
    wire N__52456;
    wire N__52453;
    wire N__52450;
    wire N__52447;
    wire N__52446;
    wire N__52443;
    wire N__52442;
    wire N__52439;
    wire N__52436;
    wire N__52435;
    wire N__52434;
    wire N__52431;
    wire N__52428;
    wire N__52425;
    wire N__52422;
    wire N__52419;
    wire N__52416;
    wire N__52413;
    wire N__52406;
    wire N__52399;
    wire N__52396;
    wire N__52393;
    wire N__52390;
    wire N__52389;
    wire N__52388;
    wire N__52387;
    wire N__52386;
    wire N__52385;
    wire N__52382;
    wire N__52379;
    wire N__52370;
    wire N__52363;
    wire N__52360;
    wire N__52357;
    wire N__52354;
    wire N__52351;
    wire N__52348;
    wire N__52345;
    wire N__52342;
    wire N__52339;
    wire N__52336;
    wire N__52333;
    wire N__52330;
    wire N__52327;
    wire N__52324;
    wire N__52321;
    wire N__52318;
    wire N__52315;
    wire N__52312;
    wire N__52309;
    wire N__52306;
    wire N__52303;
    wire N__52300;
    wire N__52299;
    wire N__52296;
    wire N__52291;
    wire N__52288;
    wire N__52287;
    wire N__52284;
    wire N__52281;
    wire N__52276;
    wire N__52273;
    wire N__52270;
    wire N__52267;
    wire N__52264;
    wire N__52261;
    wire N__52258;
    wire N__52255;
    wire N__52252;
    wire N__52249;
    wire N__52246;
    wire N__52243;
    wire N__52240;
    wire N__52237;
    wire N__52234;
    wire N__52231;
    wire N__52228;
    wire N__52225;
    wire N__52222;
    wire N__52219;
    wire N__52216;
    wire N__52213;
    wire N__52210;
    wire N__52207;
    wire N__52204;
    wire N__52201;
    wire N__52198;
    wire N__52195;
    wire N__52192;
    wire N__52189;
    wire N__52186;
    wire N__52183;
    wire N__52180;
    wire N__52179;
    wire N__52176;
    wire N__52171;
    wire N__52168;
    wire N__52165;
    wire N__52162;
    wire N__52159;
    wire N__52158;
    wire N__52155;
    wire N__52150;
    wire N__52147;
    wire N__52144;
    wire N__52143;
    wire N__52140;
    wire N__52137;
    wire N__52132;
    wire N__52129;
    wire N__52126;
    wire N__52123;
    wire N__52122;
    wire N__52119;
    wire N__52116;
    wire N__52113;
    wire N__52110;
    wire N__52105;
    wire N__52104;
    wire N__52099;
    wire N__52096;
    wire N__52093;
    wire N__52092;
    wire N__52087;
    wire N__52084;
    wire N__52081;
    wire N__52078;
    wire N__52075;
    wire N__52072;
    wire N__52069;
    wire N__52066;
    wire N__52063;
    wire N__52060;
    wire N__52057;
    wire N__52054;
    wire N__52051;
    wire N__52048;
    wire N__52045;
    wire N__52042;
    wire N__52039;
    wire N__52036;
    wire N__52033;
    wire N__52030;
    wire N__52027;
    wire N__52024;
    wire N__52023;
    wire N__52020;
    wire N__52017;
    wire N__52012;
    wire N__52009;
    wire N__52006;
    wire N__52005;
    wire N__52002;
    wire N__51999;
    wire N__51994;
    wire N__51993;
    wire N__51988;
    wire N__51985;
    wire N__51982;
    wire N__51979;
    wire N__51976;
    wire N__51975;
    wire N__51972;
    wire N__51969;
    wire N__51964;
    wire N__51963;
    wire N__51960;
    wire N__51957;
    wire N__51952;
    wire N__51951;
    wire N__51948;
    wire N__51945;
    wire N__51940;
    wire N__51937;
    wire N__51936;
    wire N__51933;
    wire N__51930;
    wire N__51925;
    wire N__51922;
    wire N__51919;
    wire N__51918;
    wire N__51915;
    wire N__51912;
    wire N__51909;
    wire N__51906;
    wire N__51901;
    wire N__51898;
    wire N__51897;
    wire N__51894;
    wire N__51891;
    wire N__51886;
    wire N__51885;
    wire N__51882;
    wire N__51879;
    wire N__51874;
    wire N__51871;
    wire N__51868;
    wire N__51865;
    wire N__51862;
    wire N__51859;
    wire N__51858;
    wire N__51855;
    wire N__51852;
    wire N__51847;
    wire N__51844;
    wire N__51841;
    wire N__51838;
    wire N__51837;
    wire N__51834;
    wire N__51831;
    wire N__51826;
    wire N__51825;
    wire N__51822;
    wire N__51819;
    wire N__51814;
    wire N__51811;
    wire N__51810;
    wire N__51807;
    wire N__51804;
    wire N__51799;
    wire N__51796;
    wire N__51793;
    wire N__51792;
    wire N__51789;
    wire N__51786;
    wire N__51781;
    wire N__51778;
    wire N__51775;
    wire N__51772;
    wire N__51769;
    wire N__51766;
    wire N__51763;
    wire N__51760;
    wire N__51759;
    wire N__51756;
    wire N__51753;
    wire N__51748;
    wire N__51745;
    wire N__51744;
    wire N__51741;
    wire N__51738;
    wire N__51735;
    wire N__51730;
    wire N__51729;
    wire N__51726;
    wire N__51723;
    wire N__51720;
    wire N__51717;
    wire N__51714;
    wire N__51711;
    wire N__51706;
    wire N__51705;
    wire N__51702;
    wire N__51699;
    wire N__51696;
    wire N__51691;
    wire N__51688;
    wire N__51685;
    wire N__51684;
    wire N__51681;
    wire N__51678;
    wire N__51673;
    wire N__51670;
    wire N__51669;
    wire N__51666;
    wire N__51663;
    wire N__51658;
    wire N__51655;
    wire N__51654;
    wire N__51649;
    wire N__51646;
    wire N__51645;
    wire N__51642;
    wire N__51639;
    wire N__51634;
    wire N__51633;
    wire N__51628;
    wire N__51625;
    wire N__51622;
    wire N__51619;
    wire N__51616;
    wire N__51613;
    wire N__51610;
    wire N__51609;
    wire N__51606;
    wire N__51603;
    wire N__51598;
    wire N__51595;
    wire N__51592;
    wire N__51589;
    wire N__51586;
    wire N__51583;
    wire N__51582;
    wire N__51579;
    wire N__51576;
    wire N__51571;
    wire N__51568;
    wire N__51565;
    wire N__51562;
    wire N__51559;
    wire N__51556;
    wire N__51553;
    wire N__51550;
    wire N__51547;
    wire N__51546;
    wire N__51543;
    wire N__51540;
    wire N__51535;
    wire N__51532;
    wire N__51529;
    wire N__51526;
    wire N__51525;
    wire N__51522;
    wire N__51517;
    wire N__51514;
    wire N__51511;
    wire N__51508;
    wire N__51505;
    wire N__51502;
    wire N__51499;
    wire N__51496;
    wire N__51493;
    wire N__51490;
    wire N__51489;
    wire N__51486;
    wire N__51483;
    wire N__51478;
    wire N__51477;
    wire N__51474;
    wire N__51469;
    wire N__51466;
    wire N__51465;
    wire N__51462;
    wire N__51459;
    wire N__51456;
    wire N__51453;
    wire N__51448;
    wire N__51445;
    wire N__51442;
    wire N__51441;
    wire N__51438;
    wire N__51435;
    wire N__51432;
    wire N__51429;
    wire N__51424;
    wire N__51421;
    wire N__51418;
    wire N__51415;
    wire N__51414;
    wire N__51411;
    wire N__51408;
    wire N__51403;
    wire N__51400;
    wire N__51397;
    wire N__51394;
    wire N__51391;
    wire N__51388;
    wire N__51385;
    wire N__51382;
    wire N__51379;
    wire N__51376;
    wire N__51373;
    wire N__51370;
    wire N__51369;
    wire N__51366;
    wire N__51363;
    wire N__51358;
    wire N__51355;
    wire N__51352;
    wire N__51349;
    wire N__51346;
    wire N__51343;
    wire N__51340;
    wire N__51337;
    wire N__51334;
    wire N__51331;
    wire N__51328;
    wire N__51325;
    wire N__51322;
    wire N__51319;
    wire N__51316;
    wire N__51315;
    wire N__51312;
    wire N__51309;
    wire N__51304;
    wire N__51301;
    wire N__51298;
    wire N__51295;
    wire N__51292;
    wire N__51289;
    wire N__51286;
    wire N__51283;
    wire N__51280;
    wire N__51277;
    wire N__51274;
    wire N__51271;
    wire N__51268;
    wire N__51265;
    wire N__51262;
    wire N__51259;
    wire N__51256;
    wire N__51253;
    wire N__51250;
    wire N__51247;
    wire N__51244;
    wire N__51241;
    wire N__51238;
    wire N__51235;
    wire N__51232;
    wire N__51229;
    wire N__51226;
    wire N__51223;
    wire N__51220;
    wire N__51217;
    wire N__51214;
    wire N__51213;
    wire N__51210;
    wire N__51207;
    wire N__51202;
    wire N__51199;
    wire N__51196;
    wire N__51193;
    wire N__51190;
    wire N__51187;
    wire N__51184;
    wire N__51181;
    wire N__51178;
    wire N__51177;
    wire N__51172;
    wire N__51169;
    wire N__51166;
    wire N__51163;
    wire N__51160;
    wire N__51157;
    wire N__51154;
    wire N__51151;
    wire N__51148;
    wire N__51145;
    wire N__51142;
    wire N__51139;
    wire N__51136;
    wire N__51133;
    wire N__51130;
    wire N__51129;
    wire N__51126;
    wire N__51123;
    wire N__51122;
    wire N__51119;
    wire N__51116;
    wire N__51113;
    wire N__51110;
    wire N__51107;
    wire N__51104;
    wire N__51097;
    wire N__51094;
    wire N__51091;
    wire N__51088;
    wire N__51085;
    wire N__51082;
    wire N__51079;
    wire N__51076;
    wire N__51073;
    wire N__51070;
    wire N__51067;
    wire N__51064;
    wire N__51063;
    wire N__51060;
    wire N__51057;
    wire N__51052;
    wire N__51051;
    wire N__51048;
    wire N__51045;
    wire N__51040;
    wire N__51037;
    wire N__51036;
    wire N__51033;
    wire N__51030;
    wire N__51025;
    wire N__51024;
    wire N__51021;
    wire N__51018;
    wire N__51013;
    wire N__51012;
    wire N__51009;
    wire N__51006;
    wire N__51001;
    wire N__51000;
    wire N__50999;
    wire N__50998;
    wire N__50991;
    wire N__50988;
    wire N__50983;
    wire N__50982;
    wire N__50981;
    wire N__50980;
    wire N__50973;
    wire N__50970;
    wire N__50965;
    wire N__50964;
    wire N__50963;
    wire N__50960;
    wire N__50959;
    wire N__50956;
    wire N__50951;
    wire N__50948;
    wire N__50941;
    wire N__50940;
    wire N__50937;
    wire N__50936;
    wire N__50935;
    wire N__50928;
    wire N__50925;
    wire N__50920;
    wire N__50917;
    wire N__50914;
    wire N__50911;
    wire N__50908;
    wire N__50905;
    wire N__50902;
    wire N__50899;
    wire N__50896;
    wire N__50893;
    wire N__50890;
    wire N__50887;
    wire N__50884;
    wire N__50881;
    wire N__50878;
    wire N__50875;
    wire N__50872;
    wire N__50869;
    wire N__50866;
    wire N__50863;
    wire N__50860;
    wire N__50857;
    wire N__50854;
    wire N__50851;
    wire N__50848;
    wire N__50845;
    wire N__50842;
    wire N__50839;
    wire N__50836;
    wire N__50833;
    wire N__50830;
    wire N__50827;
    wire N__50824;
    wire N__50821;
    wire N__50818;
    wire N__50815;
    wire N__50814;
    wire N__50811;
    wire N__50808;
    wire N__50805;
    wire N__50802;
    wire N__50799;
    wire N__50796;
    wire N__50791;
    wire N__50790;
    wire N__50787;
    wire N__50784;
    wire N__50781;
    wire N__50780;
    wire N__50777;
    wire N__50774;
    wire N__50771;
    wire N__50768;
    wire N__50763;
    wire N__50758;
    wire N__50755;
    wire N__50754;
    wire N__50751;
    wire N__50750;
    wire N__50747;
    wire N__50742;
    wire N__50741;
    wire N__50738;
    wire N__50735;
    wire N__50732;
    wire N__50729;
    wire N__50724;
    wire N__50719;
    wire N__50716;
    wire N__50713;
    wire N__50710;
    wire N__50709;
    wire N__50706;
    wire N__50703;
    wire N__50698;
    wire N__50695;
    wire N__50694;
    wire N__50691;
    wire N__50688;
    wire N__50685;
    wire N__50682;
    wire N__50677;
    wire N__50674;
    wire N__50671;
    wire N__50668;
    wire N__50665;
    wire N__50662;
    wire N__50659;
    wire N__50656;
    wire N__50655;
    wire N__50650;
    wire N__50649;
    wire N__50646;
    wire N__50643;
    wire N__50638;
    wire N__50637;
    wire N__50636;
    wire N__50633;
    wire N__50628;
    wire N__50625;
    wire N__50624;
    wire N__50621;
    wire N__50618;
    wire N__50615;
    wire N__50612;
    wire N__50607;
    wire N__50602;
    wire N__50599;
    wire N__50596;
    wire N__50593;
    wire N__50590;
    wire N__50587;
    wire N__50584;
    wire N__50581;
    wire N__50580;
    wire N__50577;
    wire N__50574;
    wire N__50571;
    wire N__50568;
    wire N__50565;
    wire N__50562;
    wire N__50559;
    wire N__50556;
    wire N__50551;
    wire N__50548;
    wire N__50547;
    wire N__50546;
    wire N__50545;
    wire N__50536;
    wire N__50533;
    wire N__50532;
    wire N__50529;
    wire N__50526;
    wire N__50523;
    wire N__50518;
    wire N__50517;
    wire N__50512;
    wire N__50509;
    wire N__50508;
    wire N__50503;
    wire N__50500;
    wire N__50497;
    wire N__50494;
    wire N__50491;
    wire N__50488;
    wire N__50485;
    wire N__50482;
    wire N__50479;
    wire N__50476;
    wire N__50473;
    wire N__50470;
    wire N__50467;
    wire N__50464;
    wire N__50461;
    wire N__50458;
    wire N__50455;
    wire N__50452;
    wire N__50449;
    wire N__50448;
    wire N__50443;
    wire N__50440;
    wire N__50437;
    wire N__50436;
    wire N__50433;
    wire N__50430;
    wire N__50425;
    wire N__50422;
    wire N__50419;
    wire N__50416;
    wire N__50413;
    wire N__50410;
    wire N__50407;
    wire N__50404;
    wire N__50401;
    wire N__50398;
    wire N__50395;
    wire N__50392;
    wire N__50389;
    wire N__50386;
    wire N__50383;
    wire N__50380;
    wire N__50377;
    wire N__50374;
    wire N__50371;
    wire N__50368;
    wire N__50365;
    wire N__50362;
    wire N__50359;
    wire N__50356;
    wire N__50353;
    wire N__50350;
    wire N__50347;
    wire N__50344;
    wire N__50341;
    wire N__50338;
    wire N__50335;
    wire N__50332;
    wire N__50329;
    wire N__50326;
    wire N__50323;
    wire N__50320;
    wire N__50317;
    wire N__50314;
    wire N__50311;
    wire N__50308;
    wire N__50305;
    wire N__50302;
    wire N__50299;
    wire N__50296;
    wire N__50293;
    wire N__50290;
    wire N__50287;
    wire N__50284;
    wire N__50281;
    wire N__50278;
    wire N__50275;
    wire N__50272;
    wire N__50269;
    wire N__50266;
    wire N__50263;
    wire N__50260;
    wire N__50257;
    wire N__50254;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50242;
    wire N__50239;
    wire N__50236;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50224;
    wire N__50221;
    wire N__50218;
    wire N__50215;
    wire N__50212;
    wire N__50209;
    wire N__50206;
    wire N__50203;
    wire N__50200;
    wire N__50197;
    wire N__50194;
    wire N__50191;
    wire N__50188;
    wire N__50185;
    wire N__50182;
    wire N__50179;
    wire N__50176;
    wire N__50173;
    wire N__50170;
    wire N__50167;
    wire N__50164;
    wire N__50163;
    wire N__50162;
    wire N__50161;
    wire N__50160;
    wire N__50159;
    wire N__50158;
    wire N__50157;
    wire N__50156;
    wire N__50155;
    wire N__50146;
    wire N__50143;
    wire N__50142;
    wire N__50139;
    wire N__50134;
    wire N__50131;
    wire N__50128;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50114;
    wire N__50111;
    wire N__50104;
    wire N__50095;
    wire N__50092;
    wire N__50091;
    wire N__50090;
    wire N__50085;
    wire N__50084;
    wire N__50081;
    wire N__50078;
    wire N__50075;
    wire N__50072;
    wire N__50069;
    wire N__50064;
    wire N__50059;
    wire N__50056;
    wire N__50055;
    wire N__50054;
    wire N__50053;
    wire N__50050;
    wire N__50047;
    wire N__50044;
    wire N__50043;
    wire N__50042;
    wire N__50041;
    wire N__50040;
    wire N__50039;
    wire N__50038;
    wire N__50037;
    wire N__50036;
    wire N__50035;
    wire N__50034;
    wire N__50033;
    wire N__50030;
    wire N__50029;
    wire N__50028;
    wire N__50027;
    wire N__50026;
    wire N__50025;
    wire N__50024;
    wire N__50021;
    wire N__50018;
    wire N__50011;
    wire N__50002;
    wire N__49993;
    wire N__49986;
    wire N__49983;
    wire N__49978;
    wire N__49975;
    wire N__49972;
    wire N__49969;
    wire N__49958;
    wire N__49953;
    wire N__49950;
    wire N__49947;
    wire N__49942;
    wire N__49941;
    wire N__49938;
    wire N__49935;
    wire N__49932;
    wire N__49929;
    wire N__49926;
    wire N__49921;
    wire N__49912;
    wire N__49911;
    wire N__49908;
    wire N__49905;
    wire N__49902;
    wire N__49899;
    wire N__49896;
    wire N__49893;
    wire N__49888;
    wire N__49885;
    wire N__49884;
    wire N__49883;
    wire N__49882;
    wire N__49879;
    wire N__49878;
    wire N__49877;
    wire N__49876;
    wire N__49871;
    wire N__49860;
    wire N__49859;
    wire N__49858;
    wire N__49857;
    wire N__49856;
    wire N__49851;
    wire N__49850;
    wire N__49847;
    wire N__49846;
    wire N__49845;
    wire N__49842;
    wire N__49841;
    wire N__49840;
    wire N__49839;
    wire N__49838;
    wire N__49837;
    wire N__49832;
    wire N__49831;
    wire N__49828;
    wire N__49817;
    wire N__49816;
    wire N__49815;
    wire N__49812;
    wire N__49811;
    wire N__49810;
    wire N__49809;
    wire N__49808;
    wire N__49807;
    wire N__49806;
    wire N__49805;
    wire N__49804;
    wire N__49801;
    wire N__49800;
    wire N__49799;
    wire N__49798;
    wire N__49797;
    wire N__49796;
    wire N__49795;
    wire N__49794;
    wire N__49793;
    wire N__49792;
    wire N__49789;
    wire N__49786;
    wire N__49785;
    wire N__49784;
    wire N__49783;
    wire N__49782;
    wire N__49779;
    wire N__49776;
    wire N__49773;
    wire N__49768;
    wire N__49765;
    wire N__49750;
    wire N__49743;
    wire N__49736;
    wire N__49733;
    wire N__49724;
    wire N__49709;
    wire N__49706;
    wire N__49703;
    wire N__49702;
    wire N__49701;
    wire N__49694;
    wire N__49689;
    wire N__49680;
    wire N__49679;
    wire N__49676;
    wire N__49671;
    wire N__49668;
    wire N__49665;
    wire N__49662;
    wire N__49657;
    wire N__49654;
    wire N__49649;
    wire N__49636;
    wire N__49633;
    wire N__49632;
    wire N__49631;
    wire N__49626;
    wire N__49623;
    wire N__49620;
    wire N__49619;
    wire N__49616;
    wire N__49613;
    wire N__49610;
    wire N__49607;
    wire N__49600;
    wire N__49597;
    wire N__49596;
    wire N__49595;
    wire N__49594;
    wire N__49593;
    wire N__49592;
    wire N__49591;
    wire N__49590;
    wire N__49589;
    wire N__49586;
    wire N__49583;
    wire N__49582;
    wire N__49581;
    wire N__49580;
    wire N__49579;
    wire N__49576;
    wire N__49573;
    wire N__49572;
    wire N__49571;
    wire N__49570;
    wire N__49569;
    wire N__49568;
    wire N__49565;
    wire N__49562;
    wire N__49559;
    wire N__49556;
    wire N__49555;
    wire N__49554;
    wire N__49553;
    wire N__49550;
    wire N__49549;
    wire N__49548;
    wire N__49547;
    wire N__49546;
    wire N__49545;
    wire N__49544;
    wire N__49543;
    wire N__49542;
    wire N__49541;
    wire N__49540;
    wire N__49539;
    wire N__49538;
    wire N__49537;
    wire N__49528;
    wire N__49527;
    wire N__49524;
    wire N__49523;
    wire N__49520;
    wire N__49519;
    wire N__49516;
    wire N__49513;
    wire N__49512;
    wire N__49511;
    wire N__49510;
    wire N__49509;
    wire N__49506;
    wire N__49503;
    wire N__49502;
    wire N__49501;
    wire N__49500;
    wire N__49493;
    wire N__49488;
    wire N__49485;
    wire N__49482;
    wire N__49481;
    wire N__49480;
    wire N__49479;
    wire N__49478;
    wire N__49477;
    wire N__49476;
    wire N__49467;
    wire N__49456;
    wire N__49449;
    wire N__49448;
    wire N__49447;
    wire N__49446;
    wire N__49435;
    wire N__49432;
    wire N__49423;
    wire N__49420;
    wire N__49415;
    wire N__49408;
    wire N__49407;
    wire N__49394;
    wire N__49389;
    wire N__49384;
    wire N__49371;
    wire N__49366;
    wire N__49363;
    wire N__49356;
    wire N__49349;
    wire N__49342;
    wire N__49341;
    wire N__49338;
    wire N__49333;
    wire N__49330;
    wire N__49323;
    wire N__49318;
    wire N__49315;
    wire N__49312;
    wire N__49297;
    wire N__49296;
    wire N__49293;
    wire N__49290;
    wire N__49287;
    wire N__49284;
    wire N__49279;
    wire N__49276;
    wire N__49275;
    wire N__49274;
    wire N__49271;
    wire N__49270;
    wire N__49265;
    wire N__49262;
    wire N__49259;
    wire N__49256;
    wire N__49253;
    wire N__49246;
    wire N__49243;
    wire N__49240;
    wire N__49239;
    wire N__49238;
    wire N__49235;
    wire N__49230;
    wire N__49225;
    wire N__49222;
    wire N__49219;
    wire N__49216;
    wire N__49213;
    wire N__49210;
    wire N__49207;
    wire N__49204;
    wire N__49201;
    wire N__49198;
    wire N__49195;
    wire N__49192;
    wire N__49189;
    wire N__49186;
    wire N__49183;
    wire N__49180;
    wire N__49177;
    wire N__49174;
    wire N__49171;
    wire N__49168;
    wire N__49165;
    wire N__49162;
    wire N__49161;
    wire N__49158;
    wire N__49155;
    wire N__49150;
    wire N__49149;
    wire N__49148;
    wire N__49141;
    wire N__49140;
    wire N__49139;
    wire N__49138;
    wire N__49135;
    wire N__49128;
    wire N__49127;
    wire N__49126;
    wire N__49125;
    wire N__49124;
    wire N__49123;
    wire N__49122;
    wire N__49121;
    wire N__49120;
    wire N__49119;
    wire N__49118;
    wire N__49117;
    wire N__49112;
    wire N__49095;
    wire N__49090;
    wire N__49087;
    wire N__49084;
    wire N__49081;
    wire N__49072;
    wire N__49069;
    wire N__49068;
    wire N__49065;
    wire N__49062;
    wire N__49059;
    wire N__49054;
    wire N__49051;
    wire N__49048;
    wire N__49047;
    wire N__49044;
    wire N__49041;
    wire N__49036;
    wire N__49035;
    wire N__49034;
    wire N__49031;
    wire N__49030;
    wire N__49029;
    wire N__49028;
    wire N__49021;
    wire N__49020;
    wire N__49017;
    wire N__49016;
    wire N__49013;
    wire N__49010;
    wire N__49007;
    wire N__49006;
    wire N__49003;
    wire N__48998;
    wire N__48995;
    wire N__48992;
    wire N__48989;
    wire N__48986;
    wire N__48983;
    wire N__48982;
    wire N__48979;
    wire N__48976;
    wire N__48971;
    wire N__48966;
    wire N__48963;
    wire N__48958;
    wire N__48949;
    wire N__48946;
    wire N__48945;
    wire N__48942;
    wire N__48939;
    wire N__48938;
    wire N__48935;
    wire N__48932;
    wire N__48929;
    wire N__48924;
    wire N__48919;
    wire N__48916;
    wire N__48913;
    wire N__48910;
    wire N__48909;
    wire N__48906;
    wire N__48903;
    wire N__48898;
    wire N__48897;
    wire N__48896;
    wire N__48895;
    wire N__48894;
    wire N__48893;
    wire N__48892;
    wire N__48891;
    wire N__48886;
    wire N__48883;
    wire N__48882;
    wire N__48881;
    wire N__48880;
    wire N__48879;
    wire N__48878;
    wire N__48877;
    wire N__48876;
    wire N__48875;
    wire N__48874;
    wire N__48873;
    wire N__48872;
    wire N__48871;
    wire N__48870;
    wire N__48869;
    wire N__48868;
    wire N__48867;
    wire N__48866;
    wire N__48865;
    wire N__48862;
    wire N__48859;
    wire N__48856;
    wire N__48855;
    wire N__48854;
    wire N__48853;
    wire N__48852;
    wire N__48851;
    wire N__48850;
    wire N__48847;
    wire N__48846;
    wire N__48843;
    wire N__48842;
    wire N__48837;
    wire N__48832;
    wire N__48823;
    wire N__48814;
    wire N__48813;
    wire N__48812;
    wire N__48811;
    wire N__48810;
    wire N__48799;
    wire N__48796;
    wire N__48791;
    wire N__48788;
    wire N__48777;
    wire N__48770;
    wire N__48769;
    wire N__48768;
    wire N__48767;
    wire N__48766;
    wire N__48765;
    wire N__48764;
    wire N__48763;
    wire N__48762;
    wire N__48761;
    wire N__48760;
    wire N__48759;
    wire N__48756;
    wire N__48755;
    wire N__48752;
    wire N__48751;
    wire N__48748;
    wire N__48745;
    wire N__48744;
    wire N__48735;
    wire N__48734;
    wire N__48733;
    wire N__48732;
    wire N__48731;
    wire N__48726;
    wire N__48725;
    wire N__48722;
    wire N__48719;
    wire N__48712;
    wire N__48711;
    wire N__48710;
    wire N__48709;
    wire N__48708;
    wire N__48705;
    wire N__48700;
    wire N__48697;
    wire N__48694;
    wire N__48693;
    wire N__48692;
    wire N__48685;
    wire N__48676;
    wire N__48673;
    wire N__48670;
    wire N__48667;
    wire N__48664;
    wire N__48661;
    wire N__48658;
    wire N__48655;
    wire N__48652;
    wire N__48649;
    wire N__48648;
    wire N__48645;
    wire N__48638;
    wire N__48635;
    wire N__48632;
    wire N__48629;
    wire N__48626;
    wire N__48621;
    wire N__48616;
    wire N__48613;
    wire N__48610;
    wire N__48603;
    wire N__48600;
    wire N__48597;
    wire N__48594;
    wire N__48589;
    wire N__48584;
    wire N__48579;
    wire N__48568;
    wire N__48565;
    wire N__48558;
    wire N__48553;
    wire N__48542;
    wire N__48539;
    wire N__48536;
    wire N__48521;
    wire N__48518;
    wire N__48513;
    wire N__48502;
    wire N__48499;
    wire N__48496;
    wire N__48493;
    wire N__48490;
    wire N__48489;
    wire N__48486;
    wire N__48483;
    wire N__48478;
    wire N__48475;
    wire N__48472;
    wire N__48469;
    wire N__48466;
    wire N__48463;
    wire N__48462;
    wire N__48459;
    wire N__48456;
    wire N__48451;
    wire N__48448;
    wire N__48447;
    wire N__48444;
    wire N__48441;
    wire N__48436;
    wire N__48433;
    wire N__48430;
    wire N__48429;
    wire N__48426;
    wire N__48423;
    wire N__48418;
    wire N__48417;
    wire N__48414;
    wire N__48409;
    wire N__48406;
    wire N__48403;
    wire N__48402;
    wire N__48399;
    wire N__48396;
    wire N__48391;
    wire N__48388;
    wire N__48385;
    wire N__48382;
    wire N__48379;
    wire N__48376;
    wire N__48373;
    wire N__48372;
    wire N__48369;
    wire N__48366;
    wire N__48361;
    wire N__48358;
    wire N__48357;
    wire N__48354;
    wire N__48351;
    wire N__48346;
    wire N__48345;
    wire N__48342;
    wire N__48339;
    wire N__48334;
    wire N__48331;
    wire N__48328;
    wire N__48325;
    wire N__48322;
    wire N__48319;
    wire N__48316;
    wire N__48313;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48301;
    wire N__48300;
    wire N__48297;
    wire N__48294;
    wire N__48289;
    wire N__48288;
    wire N__48285;
    wire N__48282;
    wire N__48277;
    wire N__48274;
    wire N__48271;
    wire N__48270;
    wire N__48265;
    wire N__48262;
    wire N__48259;
    wire N__48256;
    wire N__48255;
    wire N__48252;
    wire N__48249;
    wire N__48244;
    wire N__48241;
    wire N__48238;
    wire N__48235;
    wire N__48234;
    wire N__48231;
    wire N__48228;
    wire N__48223;
    wire N__48220;
    wire N__48217;
    wire N__48216;
    wire N__48213;
    wire N__48210;
    wire N__48207;
    wire N__48204;
    wire N__48199;
    wire N__48198;
    wire N__48195;
    wire N__48190;
    wire N__48187;
    wire N__48184;
    wire N__48181;
    wire N__48178;
    wire N__48175;
    wire N__48172;
    wire N__48171;
    wire N__48168;
    wire N__48163;
    wire N__48160;
    wire N__48157;
    wire N__48156;
    wire N__48153;
    wire N__48150;
    wire N__48147;
    wire N__48144;
    wire N__48139;
    wire N__48136;
    wire N__48133;
    wire N__48132;
    wire N__48129;
    wire N__48126;
    wire N__48121;
    wire N__48118;
    wire N__48117;
    wire N__48114;
    wire N__48111;
    wire N__48106;
    wire N__48105;
    wire N__48100;
    wire N__48097;
    wire N__48094;
    wire N__48091;
    wire N__48090;
    wire N__48087;
    wire N__48084;
    wire N__48079;
    wire N__48076;
    wire N__48075;
    wire N__48072;
    wire N__48069;
    wire N__48066;
    wire N__48063;
    wire N__48058;
    wire N__48057;
    wire N__48054;
    wire N__48051;
    wire N__48046;
    wire N__48043;
    wire N__48040;
    wire N__48037;
    wire N__48034;
    wire N__48031;
    wire N__48028;
    wire N__48025;
    wire N__48022;
    wire N__48019;
    wire N__48016;
    wire N__48013;
    wire N__48010;
    wire N__48007;
    wire N__48004;
    wire N__48001;
    wire N__48000;
    wire N__47997;
    wire N__47994;
    wire N__47989;
    wire N__47988;
    wire N__47985;
    wire N__47982;
    wire N__47977;
    wire N__47974;
    wire N__47973;
    wire N__47970;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47958;
    wire N__47955;
    wire N__47950;
    wire N__47949;
    wire N__47946;
    wire N__47943;
    wire N__47938;
    wire N__47935;
    wire N__47934;
    wire N__47931;
    wire N__47928;
    wire N__47923;
    wire N__47922;
    wire N__47919;
    wire N__47916;
    wire N__47911;
    wire N__47910;
    wire N__47907;
    wire N__47904;
    wire N__47899;
    wire N__47896;
    wire N__47893;
    wire N__47890;
    wire N__47889;
    wire N__47886;
    wire N__47883;
    wire N__47878;
    wire N__47875;
    wire N__47872;
    wire N__47869;
    wire N__47866;
    wire N__47865;
    wire N__47862;
    wire N__47859;
    wire N__47856;
    wire N__47853;
    wire N__47848;
    wire N__47845;
    wire N__47842;
    wire N__47841;
    wire N__47836;
    wire N__47833;
    wire N__47832;
    wire N__47827;
    wire N__47824;
    wire N__47823;
    wire N__47820;
    wire N__47817;
    wire N__47812;
    wire N__47811;
    wire N__47808;
    wire N__47805;
    wire N__47800;
    wire N__47799;
    wire N__47796;
    wire N__47793;
    wire N__47788;
    wire N__47787;
    wire N__47784;
    wire N__47781;
    wire N__47778;
    wire N__47773;
    wire N__47770;
    wire N__47767;
    wire N__47764;
    wire N__47763;
    wire N__47760;
    wire N__47757;
    wire N__47752;
    wire N__47749;
    wire N__47746;
    wire N__47743;
    wire N__47740;
    wire N__47737;
    wire N__47736;
    wire N__47733;
    wire N__47730;
    wire N__47725;
    wire N__47722;
    wire N__47721;
    wire N__47718;
    wire N__47715;
    wire N__47712;
    wire N__47709;
    wire N__47704;
    wire N__47701;
    wire N__47698;
    wire N__47697;
    wire N__47694;
    wire N__47691;
    wire N__47688;
    wire N__47685;
    wire N__47680;
    wire N__47677;
    wire N__47676;
    wire N__47673;
    wire N__47670;
    wire N__47665;
    wire N__47662;
    wire N__47659;
    wire N__47656;
    wire N__47655;
    wire N__47652;
    wire N__47649;
    wire N__47646;
    wire N__47643;
    wire N__47638;
    wire N__47637;
    wire N__47634;
    wire N__47631;
    wire N__47628;
    wire N__47625;
    wire N__47620;
    wire N__47617;
    wire N__47616;
    wire N__47613;
    wire N__47610;
    wire N__47607;
    wire N__47604;
    wire N__47599;
    wire N__47596;
    wire N__47593;
    wire N__47590;
    wire N__47589;
    wire N__47586;
    wire N__47583;
    wire N__47580;
    wire N__47577;
    wire N__47572;
    wire N__47569;
    wire N__47566;
    wire N__47563;
    wire N__47560;
    wire N__47557;
    wire N__47554;
    wire N__47551;
    wire N__47548;
    wire N__47545;
    wire N__47542;
    wire N__47539;
    wire N__47536;
    wire N__47533;
    wire N__47530;
    wire N__47527;
    wire N__47524;
    wire N__47521;
    wire N__47518;
    wire N__47515;
    wire N__47512;
    wire N__47509;
    wire N__47508;
    wire N__47503;
    wire N__47500;
    wire N__47497;
    wire N__47494;
    wire N__47491;
    wire N__47490;
    wire N__47485;
    wire N__47482;
    wire N__47481;
    wire N__47476;
    wire N__47473;
    wire N__47470;
    wire N__47469;
    wire N__47464;
    wire N__47461;
    wire N__47460;
    wire N__47459;
    wire N__47458;
    wire N__47455;
    wire N__47454;
    wire N__47453;
    wire N__47452;
    wire N__47451;
    wire N__47448;
    wire N__47447;
    wire N__47446;
    wire N__47445;
    wire N__47444;
    wire N__47443;
    wire N__47438;
    wire N__47437;
    wire N__47436;
    wire N__47435;
    wire N__47434;
    wire N__47433;
    wire N__47432;
    wire N__47431;
    wire N__47430;
    wire N__47429;
    wire N__47428;
    wire N__47419;
    wire N__47418;
    wire N__47417;
    wire N__47416;
    wire N__47413;
    wire N__47412;
    wire N__47411;
    wire N__47410;
    wire N__47409;
    wire N__47408;
    wire N__47397;
    wire N__47394;
    wire N__47393;
    wire N__47392;
    wire N__47391;
    wire N__47390;
    wire N__47389;
    wire N__47388;
    wire N__47387;
    wire N__47386;
    wire N__47385;
    wire N__47384;
    wire N__47383;
    wire N__47382;
    wire N__47379;
    wire N__47374;
    wire N__47373;
    wire N__47364;
    wire N__47361;
    wire N__47356;
    wire N__47353;
    wire N__47350;
    wire N__47343;
    wire N__47342;
    wire N__47341;
    wire N__47340;
    wire N__47339;
    wire N__47338;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47326;
    wire N__47321;
    wire N__47318;
    wire N__47317;
    wire N__47316;
    wire N__47315;
    wire N__47314;
    wire N__47313;
    wire N__47312;
    wire N__47311;
    wire N__47310;
    wire N__47297;
    wire N__47296;
    wire N__47293;
    wire N__47290;
    wire N__47279;
    wire N__47274;
    wire N__47271;
    wire N__47268;
    wire N__47257;
    wire N__47252;
    wire N__47247;
    wire N__47244;
    wire N__47241;
    wire N__47230;
    wire N__47223;
    wire N__47214;
    wire N__47213;
    wire N__47210;
    wire N__47207;
    wire N__47204;
    wire N__47199;
    wire N__47196;
    wire N__47193;
    wire N__47184;
    wire N__47181;
    wire N__47180;
    wire N__47177;
    wire N__47174;
    wire N__47169;
    wire N__47166;
    wire N__47163;
    wire N__47158;
    wire N__47157;
    wire N__47156;
    wire N__47155;
    wire N__47152;
    wire N__47143;
    wire N__47140;
    wire N__47137;
    wire N__47134;
    wire N__47127;
    wire N__47122;
    wire N__47119;
    wire N__47116;
    wire N__47113;
    wire N__47110;
    wire N__47107;
    wire N__47104;
    wire N__47101;
    wire N__47096;
    wire N__47093;
    wire N__47080;
    wire N__47073;
    wire N__47070;
    wire N__47067;
    wire N__47062;
    wire N__47059;
    wire N__47056;
    wire N__47053;
    wire N__47052;
    wire N__47049;
    wire N__47046;
    wire N__47041;
    wire N__47040;
    wire N__47039;
    wire N__47038;
    wire N__47035;
    wire N__47032;
    wire N__47031;
    wire N__47030;
    wire N__47027;
    wire N__47026;
    wire N__47025;
    wire N__47024;
    wire N__47023;
    wire N__47022;
    wire N__47021;
    wire N__47020;
    wire N__47017;
    wire N__47016;
    wire N__47015;
    wire N__47014;
    wire N__47013;
    wire N__47012;
    wire N__47011;
    wire N__47010;
    wire N__47009;
    wire N__47006;
    wire N__47005;
    wire N__47004;
    wire N__47001;
    wire N__47000;
    wire N__46999;
    wire N__46998;
    wire N__46997;
    wire N__46996;
    wire N__46995;
    wire N__46994;
    wire N__46991;
    wire N__46990;
    wire N__46989;
    wire N__46988;
    wire N__46987;
    wire N__46986;
    wire N__46985;
    wire N__46984;
    wire N__46977;
    wire N__46976;
    wire N__46975;
    wire N__46974;
    wire N__46973;
    wire N__46966;
    wire N__46965;
    wire N__46964;
    wire N__46963;
    wire N__46962;
    wire N__46957;
    wire N__46952;
    wire N__46949;
    wire N__46942;
    wire N__46939;
    wire N__46936;
    wire N__46935;
    wire N__46930;
    wire N__46929;
    wire N__46926;
    wire N__46921;
    wire N__46918;
    wire N__46915;
    wire N__46910;
    wire N__46903;
    wire N__46902;
    wire N__46901;
    wire N__46900;
    wire N__46899;
    wire N__46896;
    wire N__46891;
    wire N__46888;
    wire N__46885;
    wire N__46876;
    wire N__46873;
    wire N__46864;
    wire N__46861;
    wire N__46860;
    wire N__46859;
    wire N__46858;
    wire N__46857;
    wire N__46856;
    wire N__46855;
    wire N__46854;
    wire N__46847;
    wire N__46844;
    wire N__46839;
    wire N__46836;
    wire N__46831;
    wire N__46828;
    wire N__46825;
    wire N__46822;
    wire N__46819;
    wire N__46806;
    wire N__46803;
    wire N__46798;
    wire N__46795;
    wire N__46792;
    wire N__46789;
    wire N__46782;
    wire N__46779;
    wire N__46776;
    wire N__46775;
    wire N__46774;
    wire N__46773;
    wire N__46772;
    wire N__46769;
    wire N__46762;
    wire N__46759;
    wire N__46756;
    wire N__46751;
    wire N__46742;
    wire N__46733;
    wire N__46732;
    wire N__46731;
    wire N__46722;
    wire N__46719;
    wire N__46710;
    wire N__46707;
    wire N__46704;
    wire N__46701;
    wire N__46696;
    wire N__46693;
    wire N__46690;
    wire N__46679;
    wire N__46676;
    wire N__46673;
    wire N__46670;
    wire N__46663;
    wire N__46650;
    wire N__46643;
    wire N__46640;
    wire N__46637;
    wire N__46634;
    wire N__46627;
    wire N__46624;
    wire N__46621;
    wire N__46620;
    wire N__46617;
    wire N__46614;
    wire N__46609;
    wire N__46606;
    wire N__46603;
    wire N__46600;
    wire N__46599;
    wire N__46596;
    wire N__46593;
    wire N__46588;
    wire N__46587;
    wire N__46586;
    wire N__46585;
    wire N__46584;
    wire N__46583;
    wire N__46582;
    wire N__46581;
    wire N__46580;
    wire N__46579;
    wire N__46576;
    wire N__46573;
    wire N__46570;
    wire N__46569;
    wire N__46568;
    wire N__46567;
    wire N__46566;
    wire N__46565;
    wire N__46562;
    wire N__46555;
    wire N__46554;
    wire N__46553;
    wire N__46552;
    wire N__46549;
    wire N__46548;
    wire N__46545;
    wire N__46542;
    wire N__46541;
    wire N__46540;
    wire N__46539;
    wire N__46538;
    wire N__46537;
    wire N__46534;
    wire N__46531;
    wire N__46526;
    wire N__46521;
    wire N__46516;
    wire N__46513;
    wire N__46510;
    wire N__46509;
    wire N__46508;
    wire N__46501;
    wire N__46498;
    wire N__46497;
    wire N__46494;
    wire N__46493;
    wire N__46492;
    wire N__46491;
    wire N__46488;
    wire N__46487;
    wire N__46484;
    wire N__46483;
    wire N__46482;
    wire N__46473;
    wire N__46472;
    wire N__46471;
    wire N__46470;
    wire N__46469;
    wire N__46468;
    wire N__46465;
    wire N__46464;
    wire N__46463;
    wire N__46462;
    wire N__46457;
    wire N__46456;
    wire N__46455;
    wire N__46454;
    wire N__46453;
    wire N__46452;
    wire N__46451;
    wire N__46448;
    wire N__46443;
    wire N__46438;
    wire N__46433;
    wire N__46430;
    wire N__46427;
    wire N__46416;
    wire N__46413;
    wire N__46410;
    wire N__46409;
    wire N__46408;
    wire N__46407;
    wire N__46406;
    wire N__46403;
    wire N__46398;
    wire N__46397;
    wire N__46396;
    wire N__46395;
    wire N__46394;
    wire N__46391;
    wire N__46388;
    wire N__46387;
    wire N__46386;
    wire N__46385;
    wire N__46384;
    wire N__46381;
    wire N__46380;
    wire N__46373;
    wire N__46370;
    wire N__46363;
    wire N__46360;
    wire N__46357;
    wire N__46350;
    wire N__46349;
    wire N__46348;
    wire N__46347;
    wire N__46344;
    wire N__46341;
    wire N__46336;
    wire N__46327;
    wire N__46320;
    wire N__46317;
    wire N__46312;
    wire N__46309;
    wire N__46308;
    wire N__46303;
    wire N__46300;
    wire N__46293;
    wire N__46290;
    wire N__46287;
    wire N__46278;
    wire N__46275;
    wire N__46272;
    wire N__46269;
    wire N__46264;
    wire N__46261;
    wire N__46256;
    wire N__46253;
    wire N__46248;
    wire N__46245;
    wire N__46236;
    wire N__46229;
    wire N__46226;
    wire N__46211;
    wire N__46198;
    wire N__46191;
    wire N__46188;
    wire N__46183;
    wire N__46180;
    wire N__46177;
    wire N__46168;
    wire N__46167;
    wire N__46164;
    wire N__46161;
    wire N__46156;
    wire N__46153;
    wire N__46152;
    wire N__46149;
    wire N__46146;
    wire N__46141;
    wire N__46138;
    wire N__46135;
    wire N__46132;
    wire N__46129;
    wire N__46126;
    wire N__46123;
    wire N__46120;
    wire N__46117;
    wire N__46116;
    wire N__46113;
    wire N__46110;
    wire N__46105;
    wire N__46102;
    wire N__46099;
    wire N__46098;
    wire N__46095;
    wire N__46092;
    wire N__46091;
    wire N__46088;
    wire N__46083;
    wire N__46078;
    wire N__46075;
    wire N__46072;
    wire N__46069;
    wire N__46066;
    wire N__46063;
    wire N__46060;
    wire N__46057;
    wire N__46054;
    wire N__46053;
    wire N__46050;
    wire N__46047;
    wire N__46042;
    wire N__46041;
    wire N__46036;
    wire N__46033;
    wire N__46030;
    wire N__46027;
    wire N__46026;
    wire N__46023;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46009;
    wire N__46006;
    wire N__46003;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45991;
    wire N__45990;
    wire N__45985;
    wire N__45982;
    wire N__45979;
    wire N__45976;
    wire N__45975;
    wire N__45972;
    wire N__45969;
    wire N__45964;
    wire N__45961;
    wire N__45958;
    wire N__45955;
    wire N__45952;
    wire N__45949;
    wire N__45946;
    wire N__45943;
    wire N__45942;
    wire N__45939;
    wire N__45936;
    wire N__45935;
    wire N__45934;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45919;
    wire N__45910;
    wire N__45909;
    wire N__45904;
    wire N__45901;
    wire N__45898;
    wire N__45897;
    wire N__45892;
    wire N__45889;
    wire N__45886;
    wire N__45885;
    wire N__45880;
    wire N__45877;
    wire N__45876;
    wire N__45871;
    wire N__45868;
    wire N__45865;
    wire N__45864;
    wire N__45861;
    wire N__45858;
    wire N__45853;
    wire N__45852;
    wire N__45847;
    wire N__45844;
    wire N__45841;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45829;
    wire N__45826;
    wire N__45823;
    wire N__45820;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45808;
    wire N__45805;
    wire N__45802;
    wire N__45801;
    wire N__45798;
    wire N__45795;
    wire N__45790;
    wire N__45787;
    wire N__45784;
    wire N__45781;
    wire N__45778;
    wire N__45777;
    wire N__45774;
    wire N__45771;
    wire N__45766;
    wire N__45763;
    wire N__45760;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45748;
    wire N__45745;
    wire N__45744;
    wire N__45741;
    wire N__45736;
    wire N__45733;
    wire N__45730;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45720;
    wire N__45717;
    wire N__45714;
    wire N__45709;
    wire N__45706;
    wire N__45703;
    wire N__45700;
    wire N__45699;
    wire N__45696;
    wire N__45693;
    wire N__45688;
    wire N__45685;
    wire N__45682;
    wire N__45681;
    wire N__45678;
    wire N__45675;
    wire N__45670;
    wire N__45669;
    wire N__45664;
    wire N__45661;
    wire N__45658;
    wire N__45655;
    wire N__45652;
    wire N__45649;
    wire N__45646;
    wire N__45643;
    wire N__45642;
    wire N__45637;
    wire N__45634;
    wire N__45631;
    wire N__45630;
    wire N__45627;
    wire N__45624;
    wire N__45619;
    wire N__45616;
    wire N__45615;
    wire N__45612;
    wire N__45609;
    wire N__45604;
    wire N__45601;
    wire N__45598;
    wire N__45595;
    wire N__45594;
    wire N__45591;
    wire N__45588;
    wire N__45583;
    wire N__45580;
    wire N__45577;
    wire N__45574;
    wire N__45573;
    wire N__45570;
    wire N__45567;
    wire N__45562;
    wire N__45561;
    wire N__45560;
    wire N__45559;
    wire N__45556;
    wire N__45549;
    wire N__45544;
    wire N__45541;
    wire N__45538;
    wire N__45535;
    wire N__45534;
    wire N__45531;
    wire N__45528;
    wire N__45523;
    wire N__45520;
    wire N__45517;
    wire N__45514;
    wire N__45513;
    wire N__45510;
    wire N__45507;
    wire N__45502;
    wire N__45499;
    wire N__45496;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45484;
    wire N__45481;
    wire N__45478;
    wire N__45475;
    wire N__45474;
    wire N__45473;
    wire N__45472;
    wire N__45463;
    wire N__45460;
    wire N__45459;
    wire N__45458;
    wire N__45455;
    wire N__45450;
    wire N__45445;
    wire N__45442;
    wire N__45439;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45424;
    wire N__45421;
    wire N__45420;
    wire N__45417;
    wire N__45414;
    wire N__45409;
    wire N__45408;
    wire N__45407;
    wire N__45406;
    wire N__45397;
    wire N__45394;
    wire N__45391;
    wire N__45388;
    wire N__45385;
    wire N__45384;
    wire N__45381;
    wire N__45378;
    wire N__45373;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45352;
    wire N__45349;
    wire N__45346;
    wire N__45343;
    wire N__45342;
    wire N__45337;
    wire N__45334;
    wire N__45331;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45319;
    wire N__45318;
    wire N__45313;
    wire N__45310;
    wire N__45307;
    wire N__45304;
    wire N__45301;
    wire N__45300;
    wire N__45297;
    wire N__45294;
    wire N__45289;
    wire N__45286;
    wire N__45283;
    wire N__45282;
    wire N__45279;
    wire N__45276;
    wire N__45271;
    wire N__45268;
    wire N__45267;
    wire N__45264;
    wire N__45261;
    wire N__45256;
    wire N__45253;
    wire N__45252;
    wire N__45249;
    wire N__45246;
    wire N__45241;
    wire N__45238;
    wire N__45235;
    wire N__45232;
    wire N__45229;
    wire N__45228;
    wire N__45225;
    wire N__45222;
    wire N__45217;
    wire N__45214;
    wire N__45213;
    wire N__45210;
    wire N__45207;
    wire N__45204;
    wire N__45201;
    wire N__45196;
    wire N__45193;
    wire N__45190;
    wire N__45187;
    wire N__45184;
    wire N__45181;
    wire N__45178;
    wire N__45175;
    wire N__45172;
    wire N__45171;
    wire N__45166;
    wire N__45163;
    wire N__45160;
    wire N__45157;
    wire N__45156;
    wire N__45153;
    wire N__45150;
    wire N__45145;
    wire N__45142;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45130;
    wire N__45127;
    wire N__45124;
    wire N__45121;
    wire N__45120;
    wire N__45117;
    wire N__45114;
    wire N__45109;
    wire N__45106;
    wire N__45103;
    wire N__45102;
    wire N__45099;
    wire N__45096;
    wire N__45091;
    wire N__45088;
    wire N__45085;
    wire N__45082;
    wire N__45081;
    wire N__45078;
    wire N__45075;
    wire N__45072;
    wire N__45069;
    wire N__45064;
    wire N__45061;
    wire N__45060;
    wire N__45057;
    wire N__45054;
    wire N__45049;
    wire N__45046;
    wire N__45043;
    wire N__45040;
    wire N__45037;
    wire N__45034;
    wire N__45031;
    wire N__45028;
    wire N__45025;
    wire N__45022;
    wire N__45019;
    wire N__45016;
    wire N__45013;
    wire N__45012;
    wire N__45007;
    wire N__45004;
    wire N__45003;
    wire N__44998;
    wire N__44995;
    wire N__44992;
    wire N__44991;
    wire N__44988;
    wire N__44985;
    wire N__44982;
    wire N__44979;
    wire N__44974;
    wire N__44971;
    wire N__44968;
    wire N__44965;
    wire N__44964;
    wire N__44959;
    wire N__44956;
    wire N__44955;
    wire N__44952;
    wire N__44949;
    wire N__44944;
    wire N__44943;
    wire N__44938;
    wire N__44935;
    wire N__44934;
    wire N__44931;
    wire N__44928;
    wire N__44923;
    wire N__44920;
    wire N__44917;
    wire N__44916;
    wire N__44913;
    wire N__44910;
    wire N__44907;
    wire N__44904;
    wire N__44901;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44887;
    wire N__44884;
    wire N__44881;
    wire N__44878;
    wire N__44875;
    wire N__44874;
    wire N__44871;
    wire N__44868;
    wire N__44863;
    wire N__44860;
    wire N__44857;
    wire N__44854;
    wire N__44851;
    wire N__44850;
    wire N__44847;
    wire N__44844;
    wire N__44841;
    wire N__44838;
    wire N__44833;
    wire N__44832;
    wire N__44829;
    wire N__44826;
    wire N__44823;
    wire N__44820;
    wire N__44815;
    wire N__44812;
    wire N__44811;
    wire N__44808;
    wire N__44805;
    wire N__44802;
    wire N__44799;
    wire N__44794;
    wire N__44791;
    wire N__44788;
    wire N__44787;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44775;
    wire N__44770;
    wire N__44767;
    wire N__44764;
    wire N__44763;
    wire N__44760;
    wire N__44757;
    wire N__44752;
    wire N__44749;
    wire N__44746;
    wire N__44743;
    wire N__44740;
    wire N__44737;
    wire N__44734;
    wire N__44733;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44721;
    wire N__44716;
    wire N__44713;
    wire N__44712;
    wire N__44709;
    wire N__44706;
    wire N__44701;
    wire N__44698;
    wire N__44695;
    wire N__44692;
    wire N__44689;
    wire N__44686;
    wire N__44683;
    wire N__44680;
    wire N__44677;
    wire N__44674;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44662;
    wire N__44659;
    wire N__44656;
    wire N__44655;
    wire N__44650;
    wire N__44647;
    wire N__44644;
    wire N__44641;
    wire N__44640;
    wire N__44637;
    wire N__44634;
    wire N__44629;
    wire N__44626;
    wire N__44623;
    wire N__44620;
    wire N__44617;
    wire N__44614;
    wire N__44611;
    wire N__44608;
    wire N__44605;
    wire N__44602;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44592;
    wire N__44589;
    wire N__44586;
    wire N__44583;
    wire N__44580;
    wire N__44575;
    wire N__44574;
    wire N__44571;
    wire N__44568;
    wire N__44563;
    wire N__44560;
    wire N__44557;
    wire N__44554;
    wire N__44553;
    wire N__44550;
    wire N__44547;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44533;
    wire N__44532;
    wire N__44529;
    wire N__44526;
    wire N__44521;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44511;
    wire N__44508;
    wire N__44503;
    wire N__44500;
    wire N__44497;
    wire N__44496;
    wire N__44493;
    wire N__44490;
    wire N__44485;
    wire N__44484;
    wire N__44479;
    wire N__44476;
    wire N__44473;
    wire N__44470;
    wire N__44467;
    wire N__44464;
    wire N__44461;
    wire N__44458;
    wire N__44455;
    wire N__44452;
    wire N__44451;
    wire N__44448;
    wire N__44445;
    wire N__44440;
    wire N__44437;
    wire N__44434;
    wire N__44431;
    wire N__44428;
    wire N__44425;
    wire N__44422;
    wire N__44421;
    wire N__44418;
    wire N__44415;
    wire N__44410;
    wire N__44407;
    wire N__44404;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44392;
    wire N__44391;
    wire N__44390;
    wire N__44387;
    wire N__44386;
    wire N__44385;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44368;
    wire N__44359;
    wire N__44356;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44344;
    wire N__44343;
    wire N__44338;
    wire N__44335;
    wire N__44334;
    wire N__44329;
    wire N__44326;
    wire N__44323;
    wire N__44320;
    wire N__44319;
    wire N__44316;
    wire N__44313;
    wire N__44308;
    wire N__44305;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44293;
    wire N__44290;
    wire N__44287;
    wire N__44284;
    wire N__44281;
    wire N__44278;
    wire N__44275;
    wire N__44274;
    wire N__44273;
    wire N__44270;
    wire N__44265;
    wire N__44262;
    wire N__44259;
    wire N__44254;
    wire N__44251;
    wire N__44248;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44236;
    wire N__44233;
    wire N__44230;
    wire N__44227;
    wire N__44224;
    wire N__44221;
    wire N__44218;
    wire N__44215;
    wire N__44212;
    wire N__44209;
    wire N__44208;
    wire N__44205;
    wire N__44204;
    wire N__44201;
    wire N__44198;
    wire N__44195;
    wire N__44188;
    wire N__44185;
    wire N__44182;
    wire N__44179;
    wire N__44176;
    wire N__44173;
    wire N__44170;
    wire N__44167;
    wire N__44164;
    wire N__44161;
    wire N__44158;
    wire N__44155;
    wire N__44152;
    wire N__44151;
    wire N__44148;
    wire N__44145;
    wire N__44140;
    wire N__44137;
    wire N__44134;
    wire N__44131;
    wire N__44128;
    wire N__44125;
    wire N__44124;
    wire N__44119;
    wire N__44116;
    wire N__44113;
    wire N__44112;
    wire N__44107;
    wire N__44104;
    wire N__44101;
    wire N__44100;
    wire N__44095;
    wire N__44092;
    wire N__44089;
    wire N__44086;
    wire N__44083;
    wire N__44080;
    wire N__44077;
    wire N__44074;
    wire N__44071;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44059;
    wire N__44056;
    wire N__44053;
    wire N__44052;
    wire N__44047;
    wire N__44046;
    wire N__44045;
    wire N__44044;
    wire N__44041;
    wire N__44038;
    wire N__44033;
    wire N__44026;
    wire N__44023;
    wire N__44020;
    wire N__44017;
    wire N__44014;
    wire N__44013;
    wire N__44010;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43998;
    wire N__43995;
    wire N__43992;
    wire N__43989;
    wire N__43986;
    wire N__43983;
    wire N__43980;
    wire N__43977;
    wire N__43974;
    wire N__43971;
    wire N__43970;
    wire N__43965;
    wire N__43962;
    wire N__43957;
    wire N__43954;
    wire N__43951;
    wire N__43948;
    wire N__43945;
    wire N__43942;
    wire N__43941;
    wire N__43940;
    wire N__43939;
    wire N__43936;
    wire N__43933;
    wire N__43928;
    wire N__43927;
    wire N__43924;
    wire N__43921;
    wire N__43918;
    wire N__43915;
    wire N__43906;
    wire N__43903;
    wire N__43900;
    wire N__43897;
    wire N__43894;
    wire N__43891;
    wire N__43888;
    wire N__43885;
    wire N__43882;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43870;
    wire N__43869;
    wire N__43868;
    wire N__43861;
    wire N__43858;
    wire N__43855;
    wire N__43852;
    wire N__43849;
    wire N__43846;
    wire N__43843;
    wire N__43842;
    wire N__43837;
    wire N__43836;
    wire N__43833;
    wire N__43830;
    wire N__43825;
    wire N__43824;
    wire N__43819;
    wire N__43816;
    wire N__43813;
    wire N__43810;
    wire N__43809;
    wire N__43808;
    wire N__43807;
    wire N__43798;
    wire N__43795;
    wire N__43792;
    wire N__43791;
    wire N__43788;
    wire N__43785;
    wire N__43782;
    wire N__43779;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43765;
    wire N__43764;
    wire N__43761;
    wire N__43758;
    wire N__43753;
    wire N__43750;
    wire N__43747;
    wire N__43744;
    wire N__43741;
    wire N__43740;
    wire N__43737;
    wire N__43734;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43716;
    wire N__43715;
    wire N__43714;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43700;
    wire N__43693;
    wire N__43690;
    wire N__43689;
    wire N__43686;
    wire N__43685;
    wire N__43682;
    wire N__43679;
    wire N__43674;
    wire N__43673;
    wire N__43672;
    wire N__43667;
    wire N__43662;
    wire N__43657;
    wire N__43654;
    wire N__43651;
    wire N__43650;
    wire N__43649;
    wire N__43648;
    wire N__43645;
    wire N__43642;
    wire N__43637;
    wire N__43630;
    wire N__43627;
    wire N__43626;
    wire N__43625;
    wire N__43622;
    wire N__43617;
    wire N__43612;
    wire N__43611;
    wire N__43610;
    wire N__43609;
    wire N__43604;
    wire N__43599;
    wire N__43596;
    wire N__43591;
    wire N__43588;
    wire N__43587;
    wire N__43586;
    wire N__43585;
    wire N__43582;
    wire N__43575;
    wire N__43570;
    wire N__43567;
    wire N__43564;
    wire N__43563;
    wire N__43562;
    wire N__43555;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43543;
    wire N__43542;
    wire N__43539;
    wire N__43536;
    wire N__43531;
    wire N__43528;
    wire N__43525;
    wire N__43522;
    wire N__43519;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43509;
    wire N__43506;
    wire N__43501;
    wire N__43498;
    wire N__43495;
    wire N__43494;
    wire N__43491;
    wire N__43488;
    wire N__43483;
    wire N__43480;
    wire N__43477;
    wire N__43476;
    wire N__43473;
    wire N__43470;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43453;
    wire N__43452;
    wire N__43449;
    wire N__43446;
    wire N__43441;
    wire N__43438;
    wire N__43435;
    wire N__43434;
    wire N__43431;
    wire N__43428;
    wire N__43423;
    wire N__43420;
    wire N__43417;
    wire N__43414;
    wire N__43411;
    wire N__43408;
    wire N__43407;
    wire N__43404;
    wire N__43401;
    wire N__43396;
    wire N__43395;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43375;
    wire N__43372;
    wire N__43369;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43357;
    wire N__43354;
    wire N__43353;
    wire N__43350;
    wire N__43347;
    wire N__43342;
    wire N__43339;
    wire N__43336;
    wire N__43335;
    wire N__43332;
    wire N__43329;
    wire N__43326;
    wire N__43323;
    wire N__43318;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43305;
    wire N__43302;
    wire N__43299;
    wire N__43294;
    wire N__43291;
    wire N__43288;
    wire N__43287;
    wire N__43284;
    wire N__43281;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43269;
    wire N__43266;
    wire N__43263;
    wire N__43258;
    wire N__43255;
    wire N__43254;
    wire N__43251;
    wire N__43248;
    wire N__43243;
    wire N__43240;
    wire N__43237;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43216;
    wire N__43213;
    wire N__43210;
    wire N__43207;
    wire N__43204;
    wire N__43201;
    wire N__43198;
    wire N__43195;
    wire N__43192;
    wire N__43189;
    wire N__43186;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43174;
    wire N__43171;
    wire N__43170;
    wire N__43167;
    wire N__43164;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43150;
    wire N__43147;
    wire N__43146;
    wire N__43143;
    wire N__43140;
    wire N__43137;
    wire N__43134;
    wire N__43129;
    wire N__43126;
    wire N__43125;
    wire N__43120;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43108;
    wire N__43105;
    wire N__43102;
    wire N__43099;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43087;
    wire N__43084;
    wire N__43081;
    wire N__43078;
    wire N__43075;
    wire N__43072;
    wire N__43069;
    wire N__43068;
    wire N__43063;
    wire N__43060;
    wire N__43059;
    wire N__43054;
    wire N__43051;
    wire N__43050;
    wire N__43047;
    wire N__43042;
    wire N__43039;
    wire N__43038;
    wire N__43035;
    wire N__43032;
    wire N__43029;
    wire N__43026;
    wire N__43021;
    wire N__43018;
    wire N__43015;
    wire N__43012;
    wire N__43011;
    wire N__43008;
    wire N__43005;
    wire N__43000;
    wire N__42997;
    wire N__42996;
    wire N__42991;
    wire N__42988;
    wire N__42985;
    wire N__42984;
    wire N__42981;
    wire N__42978;
    wire N__42973;
    wire N__42970;
    wire N__42967;
    wire N__42964;
    wire N__42961;
    wire N__42960;
    wire N__42955;
    wire N__42952;
    wire N__42951;
    wire N__42946;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42931;
    wire N__42928;
    wire N__42925;
    wire N__42922;
    wire N__42919;
    wire N__42916;
    wire N__42913;
    wire N__42910;
    wire N__42907;
    wire N__42904;
    wire N__42903;
    wire N__42900;
    wire N__42897;
    wire N__42892;
    wire N__42889;
    wire N__42888;
    wire N__42885;
    wire N__42882;
    wire N__42879;
    wire N__42876;
    wire N__42871;
    wire N__42868;
    wire N__42865;
    wire N__42862;
    wire N__42859;
    wire N__42856;
    wire N__42855;
    wire N__42852;
    wire N__42847;
    wire N__42844;
    wire N__42843;
    wire N__42840;
    wire N__42835;
    wire N__42832;
    wire N__42829;
    wire N__42826;
    wire N__42823;
    wire N__42820;
    wire N__42817;
    wire N__42814;
    wire N__42811;
    wire N__42808;
    wire N__42807;
    wire N__42802;
    wire N__42799;
    wire N__42796;
    wire N__42793;
    wire N__42792;
    wire N__42789;
    wire N__42786;
    wire N__42783;
    wire N__42780;
    wire N__42775;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42765;
    wire N__42762;
    wire N__42757;
    wire N__42754;
    wire N__42753;
    wire N__42750;
    wire N__42747;
    wire N__42742;
    wire N__42739;
    wire N__42738;
    wire N__42735;
    wire N__42732;
    wire N__42727;
    wire N__42724;
    wire N__42721;
    wire N__42718;
    wire N__42717;
    wire N__42714;
    wire N__42713;
    wire N__42710;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42694;
    wire N__42691;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42678;
    wire N__42673;
    wire N__42670;
    wire N__42667;
    wire N__42664;
    wire N__42661;
    wire N__42660;
    wire N__42657;
    wire N__42652;
    wire N__42649;
    wire N__42648;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42636;
    wire N__42633;
    wire N__42630;
    wire N__42627;
    wire N__42622;
    wire N__42619;
    wire N__42616;
    wire N__42613;
    wire N__42610;
    wire N__42607;
    wire N__42604;
    wire N__42603;
    wire N__42600;
    wire N__42597;
    wire N__42592;
    wire N__42589;
    wire N__42586;
    wire N__42583;
    wire N__42582;
    wire N__42579;
    wire N__42576;
    wire N__42573;
    wire N__42570;
    wire N__42565;
    wire N__42562;
    wire N__42559;
    wire N__42558;
    wire N__42553;
    wire N__42550;
    wire N__42547;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42535;
    wire N__42532;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42520;
    wire N__42517;
    wire N__42514;
    wire N__42511;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42499;
    wire N__42496;
    wire N__42493;
    wire N__42490;
    wire N__42489;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42477;
    wire N__42474;
    wire N__42471;
    wire N__42466;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42448;
    wire N__42445;
    wire N__42442;
    wire N__42439;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42427;
    wire N__42424;
    wire N__42421;
    wire N__42420;
    wire N__42417;
    wire N__42414;
    wire N__42409;
    wire N__42406;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42394;
    wire N__42391;
    wire N__42388;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42376;
    wire N__42373;
    wire N__42370;
    wire N__42367;
    wire N__42364;
    wire N__42361;
    wire N__42358;
    wire N__42355;
    wire N__42352;
    wire N__42349;
    wire N__42346;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42328;
    wire N__42325;
    wire N__42322;
    wire N__42319;
    wire N__42316;
    wire N__42315;
    wire N__42312;
    wire N__42309;
    wire N__42304;
    wire N__42301;
    wire N__42298;
    wire N__42297;
    wire N__42294;
    wire N__42291;
    wire N__42286;
    wire N__42283;
    wire N__42280;
    wire N__42277;
    wire N__42276;
    wire N__42273;
    wire N__42270;
    wire N__42265;
    wire N__42264;
    wire N__42259;
    wire N__42256;
    wire N__42253;
    wire N__42252;
    wire N__42247;
    wire N__42244;
    wire N__42241;
    wire N__42238;
    wire N__42235;
    wire N__42234;
    wire N__42231;
    wire N__42228;
    wire N__42223;
    wire N__42220;
    wire N__42217;
    wire N__42214;
    wire N__42211;
    wire N__42208;
    wire N__42205;
    wire N__42202;
    wire N__42199;
    wire N__42196;
    wire N__42193;
    wire N__42190;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42180;
    wire N__42177;
    wire N__42172;
    wire N__42169;
    wire N__42166;
    wire N__42165;
    wire N__42162;
    wire N__42159;
    wire N__42154;
    wire N__42153;
    wire N__42148;
    wire N__42145;
    wire N__42142;
    wire N__42139;
    wire N__42136;
    wire N__42133;
    wire N__42130;
    wire N__42127;
    wire N__42124;
    wire N__42123;
    wire N__42118;
    wire N__42115;
    wire N__42114;
    wire N__42113;
    wire N__42112;
    wire N__42111;
    wire N__42110;
    wire N__42107;
    wire N__42096;
    wire N__42091;
    wire N__42088;
    wire N__42085;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42073;
    wire N__42070;
    wire N__42069;
    wire N__42066;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42052;
    wire N__42049;
    wire N__42046;
    wire N__42045;
    wire N__42042;
    wire N__42039;
    wire N__42034;
    wire N__42031;
    wire N__42028;
    wire N__42027;
    wire N__42024;
    wire N__42021;
    wire N__42016;
    wire N__42013;
    wire N__42010;
    wire N__42007;
    wire N__42006;
    wire N__42003;
    wire N__42000;
    wire N__41995;
    wire N__41992;
    wire N__41989;
    wire N__41986;
    wire N__41983;
    wire N__41980;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41968;
    wire N__41967;
    wire N__41966;
    wire N__41965;
    wire N__41964;
    wire N__41963;
    wire N__41952;
    wire N__41949;
    wire N__41944;
    wire N__41941;
    wire N__41940;
    wire N__41937;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41923;
    wire N__41920;
    wire N__41917;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41896;
    wire N__41893;
    wire N__41890;
    wire N__41887;
    wire N__41884;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41872;
    wire N__41871;
    wire N__41866;
    wire N__41863;
    wire N__41860;
    wire N__41857;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41845;
    wire N__41842;
    wire N__41839;
    wire N__41838;
    wire N__41835;
    wire N__41832;
    wire N__41827;
    wire N__41824;
    wire N__41821;
    wire N__41818;
    wire N__41815;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41803;
    wire N__41802;
    wire N__41801;
    wire N__41798;
    wire N__41797;
    wire N__41794;
    wire N__41793;
    wire N__41792;
    wire N__41791;
    wire N__41790;
    wire N__41787;
    wire N__41786;
    wire N__41785;
    wire N__41784;
    wire N__41783;
    wire N__41782;
    wire N__41779;
    wire N__41776;
    wire N__41775;
    wire N__41774;
    wire N__41773;
    wire N__41772;
    wire N__41771;
    wire N__41770;
    wire N__41769;
    wire N__41768;
    wire N__41767;
    wire N__41766;
    wire N__41765;
    wire N__41762;
    wire N__41759;
    wire N__41752;
    wire N__41751;
    wire N__41750;
    wire N__41749;
    wire N__41748;
    wire N__41747;
    wire N__41746;
    wire N__41745;
    wire N__41744;
    wire N__41741;
    wire N__41738;
    wire N__41735;
    wire N__41732;
    wire N__41727;
    wire N__41726;
    wire N__41725;
    wire N__41724;
    wire N__41723;
    wire N__41722;
    wire N__41721;
    wire N__41720;
    wire N__41719;
    wire N__41714;
    wire N__41711;
    wire N__41704;
    wire N__41701;
    wire N__41690;
    wire N__41689;
    wire N__41688;
    wire N__41687;
    wire N__41686;
    wire N__41685;
    wire N__41682;
    wire N__41675;
    wire N__41672;
    wire N__41671;
    wire N__41670;
    wire N__41669;
    wire N__41668;
    wire N__41667;
    wire N__41660;
    wire N__41651;
    wire N__41650;
    wire N__41649;
    wire N__41648;
    wire N__41647;
    wire N__41646;
    wire N__41639;
    wire N__41636;
    wire N__41633;
    wire N__41630;
    wire N__41623;
    wire N__41614;
    wire N__41613;
    wire N__41612;
    wire N__41603;
    wire N__41600;
    wire N__41589;
    wire N__41586;
    wire N__41581;
    wire N__41578;
    wire N__41575;
    wire N__41572;
    wire N__41567;
    wire N__41562;
    wire N__41561;
    wire N__41560;
    wire N__41559;
    wire N__41558;
    wire N__41547;
    wire N__41542;
    wire N__41533;
    wire N__41530;
    wire N__41529;
    wire N__41528;
    wire N__41527;
    wire N__41524;
    wire N__41521;
    wire N__41512;
    wire N__41509;
    wire N__41504;
    wire N__41499;
    wire N__41496;
    wire N__41489;
    wire N__41480;
    wire N__41473;
    wire N__41470;
    wire N__41467;
    wire N__41464;
    wire N__41449;
    wire N__41440;
    wire N__41437;
    wire N__41436;
    wire N__41433;
    wire N__41430;
    wire N__41425;
    wire N__41422;
    wire N__41419;
    wire N__41416;
    wire N__41413;
    wire N__41412;
    wire N__41409;
    wire N__41406;
    wire N__41401;
    wire N__41398;
    wire N__41395;
    wire N__41394;
    wire N__41391;
    wire N__41388;
    wire N__41383;
    wire N__41380;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41367;
    wire N__41362;
    wire N__41361;
    wire N__41356;
    wire N__41353;
    wire N__41350;
    wire N__41349;
    wire N__41346;
    wire N__41343;
    wire N__41338;
    wire N__41337;
    wire N__41334;
    wire N__41331;
    wire N__41326;
    wire N__41323;
    wire N__41322;
    wire N__41319;
    wire N__41316;
    wire N__41311;
    wire N__41310;
    wire N__41307;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41293;
    wire N__41292;
    wire N__41289;
    wire N__41286;
    wire N__41283;
    wire N__41280;
    wire N__41275;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41263;
    wire N__41262;
    wire N__41259;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41245;
    wire N__41244;
    wire N__41239;
    wire N__41236;
    wire N__41233;
    wire N__41230;
    wire N__41229;
    wire N__41226;
    wire N__41223;
    wire N__41218;
    wire N__41215;
    wire N__41212;
    wire N__41209;
    wire N__41206;
    wire N__41203;
    wire N__41200;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41187;
    wire N__41182;
    wire N__41181;
    wire N__41178;
    wire N__41173;
    wire N__41170;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41155;
    wire N__41154;
    wire N__41149;
    wire N__41146;
    wire N__41143;
    wire N__41140;
    wire N__41137;
    wire N__41134;
    wire N__41131;
    wire N__41128;
    wire N__41125;
    wire N__41122;
    wire N__41119;
    wire N__41116;
    wire N__41113;
    wire N__41110;
    wire N__41107;
    wire N__41104;
    wire N__41101;
    wire N__41098;
    wire N__41095;
    wire N__41092;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41080;
    wire N__41077;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41065;
    wire N__41062;
    wire N__41059;
    wire N__41056;
    wire N__41053;
    wire N__41050;
    wire N__41047;
    wire N__41046;
    wire N__41043;
    wire N__41040;
    wire N__41037;
    wire N__41034;
    wire N__41029;
    wire N__41026;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41016;
    wire N__41013;
    wire N__41008;
    wire N__41005;
    wire N__41002;
    wire N__40999;
    wire N__40996;
    wire N__40993;
    wire N__40992;
    wire N__40989;
    wire N__40986;
    wire N__40983;
    wire N__40980;
    wire N__40975;
    wire N__40972;
    wire N__40969;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40957;
    wire N__40954;
    wire N__40951;
    wire N__40948;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40936;
    wire N__40933;
    wire N__40930;
    wire N__40927;
    wire N__40924;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40912;
    wire N__40909;
    wire N__40906;
    wire N__40903;
    wire N__40900;
    wire N__40897;
    wire N__40896;
    wire N__40893;
    wire N__40890;
    wire N__40885;
    wire N__40884;
    wire N__40881;
    wire N__40876;
    wire N__40873;
    wire N__40872;
    wire N__40869;
    wire N__40864;
    wire N__40861;
    wire N__40860;
    wire N__40857;
    wire N__40854;
    wire N__40851;
    wire N__40846;
    wire N__40845;
    wire N__40842;
    wire N__40837;
    wire N__40834;
    wire N__40833;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40819;
    wire N__40818;
    wire N__40815;
    wire N__40812;
    wire N__40809;
    wire N__40804;
    wire N__40803;
    wire N__40800;
    wire N__40797;
    wire N__40794;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40771;
    wire N__40768;
    wire N__40765;
    wire N__40764;
    wire N__40761;
    wire N__40758;
    wire N__40753;
    wire N__40750;
    wire N__40747;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40737;
    wire N__40734;
    wire N__40731;
    wire N__40728;
    wire N__40723;
    wire N__40720;
    wire N__40717;
    wire N__40714;
    wire N__40711;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40701;
    wire N__40698;
    wire N__40695;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40680;
    wire N__40677;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40663;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40626;
    wire N__40623;
    wire N__40620;
    wire N__40615;
    wire N__40614;
    wire N__40609;
    wire N__40606;
    wire N__40605;
    wire N__40600;
    wire N__40597;
    wire N__40596;
    wire N__40591;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40578;
    wire N__40575;
    wire N__40572;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40560;
    wire N__40555;
    wire N__40552;
    wire N__40549;
    wire N__40548;
    wire N__40545;
    wire N__40542;
    wire N__40539;
    wire N__40536;
    wire N__40531;
    wire N__40528;
    wire N__40525;
    wire N__40522;
    wire N__40519;
    wire N__40518;
    wire N__40515;
    wire N__40512;
    wire N__40509;
    wire N__40506;
    wire N__40501;
    wire N__40500;
    wire N__40497;
    wire N__40492;
    wire N__40489;
    wire N__40488;
    wire N__40485;
    wire N__40482;
    wire N__40477;
    wire N__40474;
    wire N__40473;
    wire N__40470;
    wire N__40465;
    wire N__40462;
    wire N__40459;
    wire N__40456;
    wire N__40453;
    wire N__40450;
    wire N__40447;
    wire N__40444;
    wire N__40441;
    wire N__40438;
    wire N__40435;
    wire N__40432;
    wire N__40431;
    wire N__40428;
    wire N__40425;
    wire N__40420;
    wire N__40417;
    wire N__40414;
    wire N__40411;
    wire N__40410;
    wire N__40407;
    wire N__40404;
    wire N__40399;
    wire N__40396;
    wire N__40393;
    wire N__40390;
    wire N__40387;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40375;
    wire N__40372;
    wire N__40369;
    wire N__40368;
    wire N__40363;
    wire N__40360;
    wire N__40359;
    wire N__40354;
    wire N__40351;
    wire N__40350;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40338;
    wire N__40333;
    wire N__40332;
    wire N__40327;
    wire N__40324;
    wire N__40321;
    wire N__40318;
    wire N__40315;
    wire N__40312;
    wire N__40309;
    wire N__40308;
    wire N__40303;
    wire N__40300;
    wire N__40299;
    wire N__40296;
    wire N__40293;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40279;
    wire N__40276;
    wire N__40273;
    wire N__40272;
    wire N__40269;
    wire N__40266;
    wire N__40261;
    wire N__40258;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40246;
    wire N__40243;
    wire N__40242;
    wire N__40239;
    wire N__40236;
    wire N__40231;
    wire N__40228;
    wire N__40225;
    wire N__40222;
    wire N__40221;
    wire N__40218;
    wire N__40215;
    wire N__40210;
    wire N__40209;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40192;
    wire N__40189;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40171;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40159;
    wire N__40156;
    wire N__40155;
    wire N__40152;
    wire N__40149;
    wire N__40144;
    wire N__40143;
    wire N__40140;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40108;
    wire N__40105;
    wire N__40102;
    wire N__40099;
    wire N__40096;
    wire N__40093;
    wire N__40090;
    wire N__40087;
    wire N__40086;
    wire N__40083;
    wire N__40080;
    wire N__40077;
    wire N__40074;
    wire N__40069;
    wire N__40066;
    wire N__40065;
    wire N__40062;
    wire N__40059;
    wire N__40054;
    wire N__40053;
    wire N__40050;
    wire N__40047;
    wire N__40042;
    wire N__40039;
    wire N__40038;
    wire N__40035;
    wire N__40032;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40017;
    wire N__40014;
    wire N__40011;
    wire N__40008;
    wire N__40005;
    wire N__40000;
    wire N__39997;
    wire N__39994;
    wire N__39991;
    wire N__39988;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39976;
    wire N__39973;
    wire N__39970;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39958;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39948;
    wire N__39943;
    wire N__39942;
    wire N__39939;
    wire N__39936;
    wire N__39933;
    wire N__39930;
    wire N__39925;
    wire N__39922;
    wire N__39919;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39901;
    wire N__39898;
    wire N__39895;
    wire N__39894;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39877;
    wire N__39874;
    wire N__39871;
    wire N__39868;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39856;
    wire N__39853;
    wire N__39852;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39840;
    wire N__39835;
    wire N__39832;
    wire N__39831;
    wire N__39828;
    wire N__39825;
    wire N__39822;
    wire N__39819;
    wire N__39814;
    wire N__39811;
    wire N__39808;
    wire N__39805;
    wire N__39804;
    wire N__39801;
    wire N__39798;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39784;
    wire N__39783;
    wire N__39780;
    wire N__39777;
    wire N__39772;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39757;
    wire N__39754;
    wire N__39751;
    wire N__39750;
    wire N__39747;
    wire N__39744;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39729;
    wire N__39726;
    wire N__39723;
    wire N__39718;
    wire N__39715;
    wire N__39714;
    wire N__39711;
    wire N__39708;
    wire N__39705;
    wire N__39702;
    wire N__39697;
    wire N__39694;
    wire N__39691;
    wire N__39688;
    wire N__39685;
    wire N__39684;
    wire N__39681;
    wire N__39678;
    wire N__39673;
    wire N__39670;
    wire N__39669;
    wire N__39666;
    wire N__39663;
    wire N__39658;
    wire N__39655;
    wire N__39654;
    wire N__39651;
    wire N__39648;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39636;
    wire N__39633;
    wire N__39630;
    wire N__39625;
    wire N__39622;
    wire N__39619;
    wire N__39616;
    wire N__39613;
    wire N__39610;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39600;
    wire N__39597;
    wire N__39594;
    wire N__39589;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39576;
    wire N__39573;
    wire N__39568;
    wire N__39567;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39550;
    wire N__39547;
    wire N__39544;
    wire N__39543;
    wire N__39540;
    wire N__39537;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39523;
    wire N__39522;
    wire N__39519;
    wire N__39516;
    wire N__39513;
    wire N__39510;
    wire N__39505;
    wire N__39502;
    wire N__39499;
    wire N__39496;
    wire N__39495;
    wire N__39490;
    wire N__39487;
    wire N__39486;
    wire N__39481;
    wire N__39478;
    wire N__39475;
    wire N__39472;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39451;
    wire N__39448;
    wire N__39445;
    wire N__39442;
    wire N__39439;
    wire N__39436;
    wire N__39433;
    wire N__39430;
    wire N__39427;
    wire N__39424;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39406;
    wire N__39405;
    wire N__39402;
    wire N__39399;
    wire N__39394;
    wire N__39391;
    wire N__39388;
    wire N__39385;
    wire N__39382;
    wire N__39379;
    wire N__39376;
    wire N__39373;
    wire N__39370;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39358;
    wire N__39355;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39342;
    wire N__39339;
    wire N__39336;
    wire N__39331;
    wire N__39330;
    wire N__39327;
    wire N__39324;
    wire N__39319;
    wire N__39318;
    wire N__39315;
    wire N__39312;
    wire N__39307;
    wire N__39304;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39292;
    wire N__39289;
    wire N__39286;
    wire N__39283;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39271;
    wire N__39270;
    wire N__39267;
    wire N__39262;
    wire N__39259;
    wire N__39258;
    wire N__39255;
    wire N__39250;
    wire N__39247;
    wire N__39244;
    wire N__39241;
    wire N__39238;
    wire N__39235;
    wire N__39232;
    wire N__39229;
    wire N__39226;
    wire N__39223;
    wire N__39220;
    wire N__39217;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39204;
    wire N__39199;
    wire N__39196;
    wire N__39193;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39181;
    wire N__39178;
    wire N__39175;
    wire N__39172;
    wire N__39169;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39150;
    wire N__39145;
    wire N__39142;
    wire N__39139;
    wire N__39136;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39084;
    wire N__39081;
    wire N__39078;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39066;
    wire N__39061;
    wire N__39058;
    wire N__39057;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39045;
    wire N__39042;
    wire N__39039;
    wire N__39036;
    wire N__39033;
    wire N__39028;
    wire N__39025;
    wire N__39022;
    wire N__39021;
    wire N__39018;
    wire N__39015;
    wire N__39010;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38989;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38974;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38955;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38941;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38929;
    wire N__38928;
    wire N__38923;
    wire N__38920;
    wire N__38919;
    wire N__38914;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38901;
    wire N__38898;
    wire N__38895;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38883;
    wire N__38880;
    wire N__38877;
    wire N__38872;
    wire N__38869;
    wire N__38866;
    wire N__38863;
    wire N__38860;
    wire N__38857;
    wire N__38854;
    wire N__38851;
    wire N__38848;
    wire N__38845;
    wire N__38844;
    wire N__38841;
    wire N__38838;
    wire N__38833;
    wire N__38830;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38812;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38800;
    wire N__38797;
    wire N__38794;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38782;
    wire N__38779;
    wire N__38778;
    wire N__38775;
    wire N__38772;
    wire N__38769;
    wire N__38766;
    wire N__38761;
    wire N__38758;
    wire N__38755;
    wire N__38752;
    wire N__38749;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38737;
    wire N__38736;
    wire N__38731;
    wire N__38728;
    wire N__38725;
    wire N__38722;
    wire N__38719;
    wire N__38716;
    wire N__38713;
    wire N__38710;
    wire N__38707;
    wire N__38704;
    wire N__38701;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38689;
    wire N__38686;
    wire N__38683;
    wire N__38680;
    wire N__38679;
    wire N__38674;
    wire N__38671;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38653;
    wire N__38650;
    wire N__38647;
    wire N__38644;
    wire N__38641;
    wire N__38638;
    wire N__38635;
    wire N__38632;
    wire N__38629;
    wire N__38626;
    wire N__38623;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38610;
    wire N__38605;
    wire N__38604;
    wire N__38599;
    wire N__38596;
    wire N__38595;
    wire N__38592;
    wire N__38589;
    wire N__38584;
    wire N__38581;
    wire N__38578;
    wire N__38575;
    wire N__38572;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38560;
    wire N__38557;
    wire N__38554;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38542;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38523;
    wire N__38520;
    wire N__38517;
    wire N__38512;
    wire N__38509;
    wire N__38508;
    wire N__38505;
    wire N__38502;
    wire N__38497;
    wire N__38494;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38481;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38458;
    wire N__38455;
    wire N__38452;
    wire N__38451;
    wire N__38448;
    wire N__38445;
    wire N__38440;
    wire N__38437;
    wire N__38434;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38424;
    wire N__38421;
    wire N__38416;
    wire N__38413;
    wire N__38410;
    wire N__38407;
    wire N__38406;
    wire N__38403;
    wire N__38400;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38377;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38365;
    wire N__38362;
    wire N__38359;
    wire N__38356;
    wire N__38353;
    wire N__38350;
    wire N__38349;
    wire N__38344;
    wire N__38341;
    wire N__38340;
    wire N__38335;
    wire N__38332;
    wire N__38329;
    wire N__38326;
    wire N__38325;
    wire N__38322;
    wire N__38319;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38304;
    wire N__38301;
    wire N__38298;
    wire N__38293;
    wire N__38290;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38280;
    wire N__38277;
    wire N__38272;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38260;
    wire N__38257;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38245;
    wire N__38244;
    wire N__38241;
    wire N__38238;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38223;
    wire N__38220;
    wire N__38217;
    wire N__38212;
    wire N__38211;
    wire N__38208;
    wire N__38205;
    wire N__38202;
    wire N__38199;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38187;
    wire N__38184;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38170;
    wire N__38169;
    wire N__38166;
    wire N__38163;
    wire N__38160;
    wire N__38155;
    wire N__38152;
    wire N__38151;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38122;
    wire N__38121;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38109;
    wire N__38106;
    wire N__38103;
    wire N__38098;
    wire N__38097;
    wire N__38094;
    wire N__38091;
    wire N__38086;
    wire N__38085;
    wire N__38082;
    wire N__38079;
    wire N__38076;
    wire N__38073;
    wire N__38068;
    wire N__38065;
    wire N__38062;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38050;
    wire N__38047;
    wire N__38046;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38034;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38020;
    wire N__38019;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38002;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37992;
    wire N__37987;
    wire N__37984;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37971;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37959;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37947;
    wire N__37942;
    wire N__37939;
    wire N__37936;
    wire N__37933;
    wire N__37930;
    wire N__37927;
    wire N__37924;
    wire N__37921;
    wire N__37920;
    wire N__37917;
    wire N__37914;
    wire N__37911;
    wire N__37908;
    wire N__37903;
    wire N__37900;
    wire N__37897;
    wire N__37894;
    wire N__37891;
    wire N__37890;
    wire N__37887;
    wire N__37884;
    wire N__37879;
    wire N__37876;
    wire N__37873;
    wire N__37872;
    wire N__37869;
    wire N__37866;
    wire N__37861;
    wire N__37858;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37846;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37834;
    wire N__37831;
    wire N__37828;
    wire N__37827;
    wire N__37824;
    wire N__37821;
    wire N__37816;
    wire N__37815;
    wire N__37812;
    wire N__37809;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37795;
    wire N__37792;
    wire N__37789;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37771;
    wire N__37768;
    wire N__37765;
    wire N__37762;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37747;
    wire N__37744;
    wire N__37741;
    wire N__37738;
    wire N__37735;
    wire N__37732;
    wire N__37731;
    wire N__37726;
    wire N__37723;
    wire N__37720;
    wire N__37717;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37705;
    wire N__37702;
    wire N__37701;
    wire N__37696;
    wire N__37693;
    wire N__37690;
    wire N__37687;
    wire N__37684;
    wire N__37681;
    wire N__37680;
    wire N__37677;
    wire N__37672;
    wire N__37669;
    wire N__37666;
    wire N__37665;
    wire N__37662;
    wire N__37659;
    wire N__37656;
    wire N__37651;
    wire N__37648;
    wire N__37645;
    wire N__37642;
    wire N__37641;
    wire N__37638;
    wire N__37635;
    wire N__37630;
    wire N__37627;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37615;
    wire N__37612;
    wire N__37609;
    wire N__37608;
    wire N__37603;
    wire N__37600;
    wire N__37599;
    wire N__37594;
    wire N__37591;
    wire N__37590;
    wire N__37585;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37575;
    wire N__37572;
    wire N__37569;
    wire N__37564;
    wire N__37561;
    wire N__37558;
    wire N__37555;
    wire N__37552;
    wire N__37549;
    wire N__37546;
    wire N__37543;
    wire N__37540;
    wire N__37537;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37524;
    wire N__37521;
    wire N__37518;
    wire N__37513;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37501;
    wire N__37500;
    wire N__37497;
    wire N__37494;
    wire N__37489;
    wire N__37486;
    wire N__37483;
    wire N__37480;
    wire N__37477;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37464;
    wire N__37461;
    wire N__37458;
    wire N__37453;
    wire N__37450;
    wire N__37447;
    wire N__37446;
    wire N__37441;
    wire N__37438;
    wire N__37435;
    wire N__37432;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37420;
    wire N__37417;
    wire N__37414;
    wire N__37413;
    wire N__37410;
    wire N__37407;
    wire N__37402;
    wire N__37399;
    wire N__37396;
    wire N__37393;
    wire N__37392;
    wire N__37387;
    wire N__37384;
    wire N__37381;
    wire N__37378;
    wire N__37375;
    wire N__37374;
    wire N__37371;
    wire N__37368;
    wire N__37363;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37351;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37341;
    wire N__37336;
    wire N__37333;
    wire N__37332;
    wire N__37329;
    wire N__37326;
    wire N__37321;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37311;
    wire N__37306;
    wire N__37303;
    wire N__37300;
    wire N__37297;
    wire N__37294;
    wire N__37291;
    wire N__37288;
    wire N__37285;
    wire N__37282;
    wire N__37279;
    wire N__37276;
    wire N__37273;
    wire N__37270;
    wire N__37267;
    wire N__37264;
    wire N__37261;
    wire N__37258;
    wire N__37255;
    wire N__37252;
    wire N__37251;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37236;
    wire N__37233;
    wire N__37230;
    wire N__37225;
    wire N__37222;
    wire N__37219;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37207;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37192;
    wire N__37191;
    wire N__37188;
    wire N__37185;
    wire N__37180;
    wire N__37179;
    wire N__37174;
    wire N__37171;
    wire N__37168;
    wire N__37167;
    wire N__37164;
    wire N__37161;
    wire N__37156;
    wire N__37153;
    wire N__37150;
    wire N__37147;
    wire N__37146;
    wire N__37143;
    wire N__37140;
    wire N__37135;
    wire N__37132;
    wire N__37129;
    wire N__37126;
    wire N__37123;
    wire N__37120;
    wire N__37117;
    wire N__37114;
    wire N__37113;
    wire N__37110;
    wire N__37107;
    wire N__37102;
    wire N__37101;
    wire N__37098;
    wire N__37095;
    wire N__37090;
    wire N__37087;
    wire N__37084;
    wire N__37081;
    wire N__37078;
    wire N__37075;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37063;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37038;
    wire N__37033;
    wire N__37030;
    wire N__37029;
    wire N__37024;
    wire N__37021;
    wire N__37020;
    wire N__37017;
    wire N__37014;
    wire N__37009;
    wire N__37008;
    wire N__37005;
    wire N__37002;
    wire N__36999;
    wire N__36994;
    wire N__36991;
    wire N__36990;
    wire N__36987;
    wire N__36984;
    wire N__36979;
    wire N__36976;
    wire N__36973;
    wire N__36972;
    wire N__36969;
    wire N__36966;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36943;
    wire N__36942;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36930;
    wire N__36925;
    wire N__36922;
    wire N__36919;
    wire N__36918;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36895;
    wire N__36892;
    wire N__36891;
    wire N__36888;
    wire N__36885;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36873;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36849;
    wire N__36846;
    wire N__36843;
    wire N__36838;
    wire N__36837;
    wire N__36834;
    wire N__36831;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36802;
    wire N__36799;
    wire N__36796;
    wire N__36793;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36774;
    wire N__36771;
    wire N__36766;
    wire N__36765;
    wire N__36760;
    wire N__36757;
    wire N__36756;
    wire N__36751;
    wire N__36748;
    wire N__36745;
    wire N__36742;
    wire N__36739;
    wire N__36736;
    wire N__36733;
    wire N__36730;
    wire N__36727;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36715;
    wire N__36712;
    wire N__36709;
    wire N__36708;
    wire N__36705;
    wire N__36702;
    wire N__36699;
    wire N__36696;
    wire N__36691;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36676;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36666;
    wire N__36663;
    wire N__36658;
    wire N__36657;
    wire N__36654;
    wire N__36651;
    wire N__36648;
    wire N__36643;
    wire N__36642;
    wire N__36639;
    wire N__36636;
    wire N__36631;
    wire N__36628;
    wire N__36625;
    wire N__36622;
    wire N__36621;
    wire N__36618;
    wire N__36615;
    wire N__36610;
    wire N__36607;
    wire N__36606;
    wire N__36601;
    wire N__36598;
    wire N__36597;
    wire N__36594;
    wire N__36591;
    wire N__36588;
    wire N__36583;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36573;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36556;
    wire N__36555;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36538;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36528;
    wire N__36523;
    wire N__36520;
    wire N__36517;
    wire N__36514;
    wire N__36511;
    wire N__36508;
    wire N__36505;
    wire N__36504;
    wire N__36501;
    wire N__36498;
    wire N__36495;
    wire N__36490;
    wire N__36487;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36474;
    wire N__36469;
    wire N__36468;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36454;
    wire N__36453;
    wire N__36450;
    wire N__36445;
    wire N__36442;
    wire N__36439;
    wire N__36436;
    wire N__36433;
    wire N__36430;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36418;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36403;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36376;
    wire N__36373;
    wire N__36370;
    wire N__36369;
    wire N__36364;
    wire N__36361;
    wire N__36360;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36348;
    wire N__36345;
    wire N__36340;
    wire N__36337;
    wire N__36336;
    wire N__36333;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36319;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36307;
    wire N__36304;
    wire N__36301;
    wire N__36298;
    wire N__36295;
    wire N__36294;
    wire N__36291;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36274;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36262;
    wire N__36261;
    wire N__36258;
    wire N__36255;
    wire N__36250;
    wire N__36249;
    wire N__36246;
    wire N__36243;
    wire N__36238;
    wire N__36235;
    wire N__36234;
    wire N__36231;
    wire N__36226;
    wire N__36223;
    wire N__36222;
    wire N__36217;
    wire N__36214;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36189;
    wire N__36186;
    wire N__36183;
    wire N__36180;
    wire N__36177;
    wire N__36172;
    wire N__36169;
    wire N__36166;
    wire N__36163;
    wire N__36160;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36127;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36109;
    wire N__36106;
    wire N__36103;
    wire N__36100;
    wire N__36097;
    wire N__36094;
    wire N__36093;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36076;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36066;
    wire N__36063;
    wire N__36060;
    wire N__36055;
    wire N__36054;
    wire N__36051;
    wire N__36048;
    wire N__36045;
    wire N__36040;
    wire N__36037;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36025;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36012;
    wire N__36007;
    wire N__36004;
    wire N__36003;
    wire N__36000;
    wire N__35997;
    wire N__35994;
    wire N__35991;
    wire N__35986;
    wire N__35983;
    wire N__35980;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35962;
    wire N__35959;
    wire N__35956;
    wire N__35953;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35937;
    wire N__35934;
    wire N__35931;
    wire N__35926;
    wire N__35923;
    wire N__35922;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35908;
    wire N__35907;
    wire N__35904;
    wire N__35901;
    wire N__35896;
    wire N__35895;
    wire N__35892;
    wire N__35889;
    wire N__35886;
    wire N__35883;
    wire N__35878;
    wire N__35875;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35851;
    wire N__35848;
    wire N__35845;
    wire N__35842;
    wire N__35839;
    wire N__35836;
    wire N__35835;
    wire N__35832;
    wire N__35829;
    wire N__35824;
    wire N__35823;
    wire N__35820;
    wire N__35815;
    wire N__35812;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35802;
    wire N__35799;
    wire N__35796;
    wire N__35793;
    wire N__35790;
    wire N__35785;
    wire N__35782;
    wire N__35781;
    wire N__35778;
    wire N__35775;
    wire N__35772;
    wire N__35769;
    wire N__35764;
    wire N__35761;
    wire N__35758;
    wire N__35757;
    wire N__35754;
    wire N__35751;
    wire N__35746;
    wire N__35743;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35731;
    wire N__35728;
    wire N__35727;
    wire N__35722;
    wire N__35719;
    wire N__35716;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35706;
    wire N__35703;
    wire N__35700;
    wire N__35697;
    wire N__35694;
    wire N__35689;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35676;
    wire N__35673;
    wire N__35670;
    wire N__35665;
    wire N__35662;
    wire N__35661;
    wire N__35658;
    wire N__35655;
    wire N__35650;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35638;
    wire N__35637;
    wire N__35634;
    wire N__35631;
    wire N__35628;
    wire N__35625;
    wire N__35620;
    wire N__35617;
    wire N__35616;
    wire N__35613;
    wire N__35610;
    wire N__35605;
    wire N__35602;
    wire N__35601;
    wire N__35596;
    wire N__35593;
    wire N__35590;
    wire N__35587;
    wire N__35584;
    wire N__35583;
    wire N__35578;
    wire N__35575;
    wire N__35572;
    wire N__35569;
    wire N__35566;
    wire N__35563;
    wire N__35560;
    wire N__35559;
    wire N__35554;
    wire N__35551;
    wire N__35550;
    wire N__35545;
    wire N__35542;
    wire N__35539;
    wire N__35538;
    wire N__35535;
    wire N__35532;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35512;
    wire N__35509;
    wire N__35506;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35485;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35470;
    wire N__35467;
    wire N__35464;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35454;
    wire N__35451;
    wire N__35448;
    wire N__35445;
    wire N__35442;
    wire N__35437;
    wire N__35434;
    wire N__35431;
    wire N__35428;
    wire N__35425;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35397;
    wire N__35394;
    wire N__35391;
    wire N__35386;
    wire N__35383;
    wire N__35382;
    wire N__35379;
    wire N__35376;
    wire N__35373;
    wire N__35370;
    wire N__35365;
    wire N__35362;
    wire N__35359;
    wire N__35358;
    wire N__35355;
    wire N__35352;
    wire N__35349;
    wire N__35346;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35332;
    wire N__35329;
    wire N__35326;
    wire N__35325;
    wire N__35320;
    wire N__35317;
    wire N__35316;
    wire N__35313;
    wire N__35310;
    wire N__35307;
    wire N__35304;
    wire N__35299;
    wire N__35296;
    wire N__35293;
    wire N__35292;
    wire N__35289;
    wire N__35284;
    wire N__35281;
    wire N__35278;
    wire N__35275;
    wire N__35274;
    wire N__35269;
    wire N__35266;
    wire N__35265;
    wire N__35260;
    wire N__35257;
    wire N__35256;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35242;
    wire N__35239;
    wire N__35238;
    wire N__35235;
    wire N__35230;
    wire N__35227;
    wire N__35226;
    wire N__35223;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35155;
    wire N__35152;
    wire N__35149;
    wire N__35146;
    wire N__35143;
    wire N__35140;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35101;
    wire N__35100;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35085;
    wire N__35082;
    wire N__35077;
    wire N__35074;
    wire N__35073;
    wire N__35068;
    wire N__35065;
    wire N__35064;
    wire N__35061;
    wire N__35058;
    wire N__35055;
    wire N__35050;
    wire N__35047;
    wire N__35046;
    wire N__35043;
    wire N__35040;
    wire N__35037;
    wire N__35034;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35011;
    wire N__35008;
    wire N__35005;
    wire N__35004;
    wire N__34999;
    wire N__34996;
    wire N__34995;
    wire N__34990;
    wire N__34987;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34936;
    wire N__34933;
    wire N__34930;
    wire N__34927;
    wire N__34924;
    wire N__34921;
    wire N__34920;
    wire N__34915;
    wire N__34912;
    wire N__34909;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34893;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34879;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34854;
    wire N__34849;
    wire N__34846;
    wire N__34845;
    wire N__34842;
    wire N__34837;
    wire N__34834;
    wire N__34831;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34819;
    wire N__34818;
    wire N__34815;
    wire N__34812;
    wire N__34807;
    wire N__34806;
    wire N__34801;
    wire N__34798;
    wire N__34797;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34780;
    wire N__34777;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34767;
    wire N__34764;
    wire N__34759;
    wire N__34756;
    wire N__34755;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34743;
    wire N__34738;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34720;
    wire N__34717;
    wire N__34714;
    wire N__34711;
    wire N__34710;
    wire N__34707;
    wire N__34704;
    wire N__34701;
    wire N__34698;
    wire N__34693;
    wire N__34692;
    wire N__34687;
    wire N__34684;
    wire N__34683;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34669;
    wire N__34666;
    wire N__34665;
    wire N__34662;
    wire N__34657;
    wire N__34654;
    wire N__34651;
    wire N__34650;
    wire N__34647;
    wire N__34644;
    wire N__34641;
    wire N__34638;
    wire N__34633;
    wire N__34630;
    wire N__34629;
    wire N__34626;
    wire N__34623;
    wire N__34620;
    wire N__34617;
    wire N__34612;
    wire N__34609;
    wire N__34606;
    wire N__34603;
    wire N__34602;
    wire N__34599;
    wire N__34596;
    wire N__34591;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34579;
    wire N__34576;
    wire N__34573;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34561;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34551;
    wire N__34548;
    wire N__34545;
    wire N__34542;
    wire N__34537;
    wire N__34536;
    wire N__34533;
    wire N__34528;
    wire N__34525;
    wire N__34522;
    wire N__34519;
    wire N__34516;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34506;
    wire N__34501;
    wire N__34498;
    wire N__34495;
    wire N__34492;
    wire N__34491;
    wire N__34488;
    wire N__34485;
    wire N__34480;
    wire N__34479;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34462;
    wire N__34461;
    wire N__34456;
    wire N__34453;
    wire N__34450;
    wire N__34449;
    wire N__34446;
    wire N__34443;
    wire N__34438;
    wire N__34435;
    wire N__34432;
    wire N__34429;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34410;
    wire N__34405;
    wire N__34402;
    wire N__34401;
    wire N__34396;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34384;
    wire N__34381;
    wire N__34378;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34357;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34324;
    wire N__34321;
    wire N__34320;
    wire N__34315;
    wire N__34312;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34296;
    wire N__34291;
    wire N__34288;
    wire N__34287;
    wire N__34284;
    wire N__34281;
    wire N__34276;
    wire N__34273;
    wire N__34272;
    wire N__34269;
    wire N__34266;
    wire N__34263;
    wire N__34260;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34230;
    wire N__34227;
    wire N__34222;
    wire N__34219;
    wire N__34218;
    wire N__34215;
    wire N__34212;
    wire N__34209;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34171;
    wire N__34168;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34156;
    wire N__34155;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34135;
    wire N__34132;
    wire N__34129;
    wire N__34128;
    wire N__34123;
    wire N__34120;
    wire N__34119;
    wire N__34114;
    wire N__34111;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34099;
    wire N__34096;
    wire N__34095;
    wire N__34090;
    wire N__34087;
    wire N__34086;
    wire N__34083;
    wire N__34080;
    wire N__34077;
    wire N__34074;
    wire N__34069;
    wire N__34066;
    wire N__34063;
    wire N__34060;
    wire N__34057;
    wire N__34054;
    wire N__34053;
    wire N__34050;
    wire N__34045;
    wire N__34042;
    wire N__34041;
    wire N__34038;
    wire N__34033;
    wire N__34030;
    wire N__34029;
    wire N__34026;
    wire N__34023;
    wire N__34018;
    wire N__34015;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33970;
    wire N__33969;
    wire N__33966;
    wire N__33963;
    wire N__33960;
    wire N__33957;
    wire N__33952;
    wire N__33949;
    wire N__33946;
    wire N__33945;
    wire N__33942;
    wire N__33939;
    wire N__33934;
    wire N__33931;
    wire N__33928;
    wire N__33925;
    wire N__33922;
    wire N__33921;
    wire N__33918;
    wire N__33915;
    wire N__33910;
    wire N__33907;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33885;
    wire N__33882;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33822;
    wire N__33817;
    wire N__33814;
    wire N__33813;
    wire N__33808;
    wire N__33805;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33769;
    wire N__33768;
    wire N__33763;
    wire N__33760;
    wire N__33759;
    wire N__33756;
    wire N__33751;
    wire N__33748;
    wire N__33747;
    wire N__33742;
    wire N__33739;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33721;
    wire N__33718;
    wire N__33717;
    wire N__33714;
    wire N__33711;
    wire N__33708;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33693;
    wire N__33690;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33672;
    wire N__33669;
    wire N__33666;
    wire N__33661;
    wire N__33660;
    wire N__33657;
    wire N__33654;
    wire N__33649;
    wire N__33648;
    wire N__33645;
    wire N__33640;
    wire N__33637;
    wire N__33636;
    wire N__33631;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33618;
    wire N__33615;
    wire N__33612;
    wire N__33609;
    wire N__33606;
    wire N__33601;
    wire N__33598;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33573;
    wire N__33568;
    wire N__33567;
    wire N__33564;
    wire N__33561;
    wire N__33556;
    wire N__33555;
    wire N__33552;
    wire N__33547;
    wire N__33544;
    wire N__33543;
    wire N__33540;
    wire N__33535;
    wire N__33532;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33514;
    wire N__33513;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33487;
    wire N__33484;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33472;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33442;
    wire N__33439;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33421;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33399;
    wire N__33396;
    wire N__33391;
    wire N__33388;
    wire N__33385;
    wire N__33382;
    wire N__33379;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33360;
    wire N__33355;
    wire N__33352;
    wire N__33351;
    wire N__33348;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33325;
    wire N__33324;
    wire N__33321;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33300;
    wire N__33295;
    wire N__33292;
    wire N__33291;
    wire N__33286;
    wire N__33283;
    wire N__33282;
    wire N__33279;
    wire N__33274;
    wire N__33271;
    wire N__33270;
    wire N__33267;
    wire N__33264;
    wire N__33261;
    wire N__33256;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33244;
    wire N__33241;
    wire N__33240;
    wire N__33237;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33223;
    wire N__33220;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33210;
    wire N__33205;
    wire N__33202;
    wire N__33201;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33126;
    wire N__33123;
    wire N__33118;
    wire N__33115;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33064;
    wire N__33063;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33046;
    wire N__33045;
    wire N__33042;
    wire N__33037;
    wire N__33034;
    wire N__33031;
    wire N__33030;
    wire N__33027;
    wire N__33022;
    wire N__33019;
    wire N__33018;
    wire N__33015;
    wire N__33012;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32973;
    wire N__32970;
    wire N__32965;
    wire N__32962;
    wire N__32961;
    wire N__32958;
    wire N__32953;
    wire N__32950;
    wire N__32949;
    wire N__32946;
    wire N__32941;
    wire N__32938;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire VCCG0;
    wire ICE_SYSCLK_c;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12836 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14273_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12839 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11573_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11543 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13628_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13472_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12956_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13199 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13256 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12842_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12845_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11636_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_10 ;
    wire REG_mem_26_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11545 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13265_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11621 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13298_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13259 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14006 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14009_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11627 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12914 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12917 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14048 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14036_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12129_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12126 ;
    wire REG_mem_13_7;
    wire REG_mem_58_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11524 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12776 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14384_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14387_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12779 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12071_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13688_cascade_ ;
    wire REG_mem_23_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14270 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13328_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12977_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11572 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12866_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12869 ;
    wire REG_mem_55_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_14 ;
    wire REG_mem_48_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12332 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12331 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_10 ;
    wire REG_mem_36_14;
    wire REG_mem_37_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_14 ;
    wire REG_mem_31_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13898_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13901 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11527 ;
    wire REG_mem_16_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12965 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11635 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11548 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13262 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11546 ;
    wire REG_mem_18_10;
    wire REG_mem_19_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14228 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11528 ;
    wire REG_mem_58_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12998_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13001_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_3 ;
    wire REG_mem_26_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12355 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13196 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14264_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11549 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11578 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11579_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13271 ;
    wire REG_mem_36_10;
    wire REG_mem_37_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11584 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13268 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11525 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_10 ;
    wire FIFO_D13_c_13;
    wire FIFO_D14_c_14;
    wire FIFO_D15_c_15;
    wire \usb3_if_inst.usb3_data_in_latched_14 ;
    wire \INVusb3_if_inst.dc32_fifo_data_in_i15C_net ;
    wire REG_mem_31_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12980_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13817_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13226 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11513_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13160_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12185 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13163 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13475 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13331 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11534 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13106_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13109 ;
    wire REG_mem_46_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13046_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13049 ;
    wire REG_mem_44_14;
    wire REG_mem_31_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12272 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13190_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12248 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13193 ;
    wire REG_mem_18_14;
    wire REG_mem_19_14;
    wire REG_mem_49_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12974 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12271 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12191 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_3 ;
    wire REG_mem_31_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14000_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_9 ;
    wire REG_mem_63_14;
    wire REG_mem_6_10;
    wire REG_mem_5_10;
    wire REG_mem_10_10;
    wire REG_mem_11_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14180_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14183 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14096 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13052_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13055 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14336 ;
    wire REG_mem_26_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12012 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11991_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14312_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14003 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14099 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11975_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11976 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11523 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12806 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12809 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13322 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13274_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12339_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12327 ;
    wire REG_mem_63_13;
    wire REG_mem_58_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11830_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13490 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11792_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11791 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13493 ;
    wire REG_mem_36_3;
    wire REG_mem_37_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11531_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11509_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14186 ;
    wire REG_mem_58_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11510 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_12 ;
    wire FIFO_D11_c_11;
    wire FIFO_D12_c_12;
    wire \usb3_if_inst.usb3_data_in_latched_15 ;
    wire \INVusb3_if_inst.dc32_fifo_data_in_i16C_net ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13166_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13169_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12446 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12466 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14330_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11516 ;
    wire REG_mem_50_9;
    wire REG_mem_51_9;
    wire REG_mem_55_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12031 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12032_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12035 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14150_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12034 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12043 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12857_cascade_ ;
    wire REG_mem_42_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12854 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12959 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14300 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11501 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11500_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12467 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13127 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12962 ;
    wire REG_mem_48_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13025 ;
    wire REG_mem_55_10;
    wire REG_mem_49_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11674 ;
    wire REG_mem_13_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13664_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13667 ;
    wire REG_mem_12_14;
    wire REG_mem_14_14;
    wire REG_mem_15_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_13 ;
    wire REG_mem_63_3;
    wire REG_mem_63_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13124 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12464 ;
    wire REG_mem_58_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11675 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_14 ;
    wire REG_mem_12_7;
    wire REG_mem_8_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13184_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12890_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13187 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12893_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14030_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14024 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11559 ;
    wire REG_mem_5_12;
    wire REG_mem_26_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12878_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12881_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13094_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12354 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13100_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12372 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12293 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12298 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13220 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14189 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11670_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13223 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11576_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13097 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11577_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14054 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13208 ;
    wire REG_mem_26_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_12 ;
    wire REG_mem_55_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12292 ;
    wire FIFO_D10_c_10;
    wire \usb3_if_inst.usb3_data_in_latched_10 ;
    wire \usb3_if_inst.usb3_data_in_latched_11 ;
    wire \usb3_if_inst.usb3_data_in_latched_12 ;
    wire \usb3_if_inst.usb3_data_in_latched_13 ;
    wire \INVusb3_if_inst.state_FSM_i5C_net ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12461 ;
    wire REG_mem_55_9;
    wire REG_mem_26_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13028_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12463 ;
    wire REG_mem_16_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12833_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12070 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12788_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12791 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12460 ;
    wire REG_mem_17_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11530 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12190 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_15 ;
    wire REG_mem_23_3;
    wire REG_mem_18_3;
    wire REG_mem_17_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12247 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13484 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11647_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11648 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13487 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_10 ;
    wire REG_mem_16_3;
    wire REG_mem_17_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13814 ;
    wire REG_mem_11_14;
    wire REG_mem_5_14;
    wire REG_mem_6_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13022 ;
    wire REG_mem_49_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13244_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13247 ;
    wire REG_mem_51_3;
    wire REG_mem_51_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_3 ;
    wire REG_mem_63_0;
    wire REG_mem_6_3;
    wire REG_mem_43_3;
    wire REG_mem_41_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13454_cascade_ ;
    wire REG_mem_42_3;
    wire REG_mem_44_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12800_cascade_ ;
    wire REG_mem_45_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12803 ;
    wire REG_mem_58_15;
    wire REG_mem_12_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11625 ;
    wire REG_mem_43_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13457 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11990 ;
    wire REG_mem_10_3;
    wire REG_mem_11_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_11 ;
    wire REG_mem_10_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_12 ;
    wire REG_mem_42_7;
    wire REG_mem_42_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12494_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14252_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12481 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12476 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13292_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12475 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13295_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14255 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11643 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12487 ;
    wire REG_mem_42_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12488 ;
    wire REG_mem_43_12;
    wire REG_mem_31_12;
    wire REG_mem_44_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12493 ;
    wire REG_mem_45_12;
    wire REG_mem_9_10;
    wire REG_mem_43_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_12 ;
    wire REG_mem_41_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13397_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11630 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13142_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13145 ;
    wire REG_mem_42_10;
    wire REG_mem_43_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13394 ;
    wire REG_mem_45_10;
    wire REG_mem_44_10;
    wire REG_mem_46_10;
    wire REG_mem_10_13;
    wire pll_clk_unbuf;
    wire GB_BUFFER_pll_clk_unbuf_THRU_CO;
    wire FIFO_D9_c_9;
    wire \usb3_if_inst.usb3_data_in_latched_9 ;
    wire REG_mem_63_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12044 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12860_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_0 ;
    wire REG_mem_42_15;
    wire REG_mem_43_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13400_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13403_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12068_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12017 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12016 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12935 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12983 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13031 ;
    wire REG_mem_37_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13235_cascade_ ;
    wire REG_mem_47_0;
    wire REG_mem_4_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12343 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12923_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12059 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12896_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12899 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12812 ;
    wire REG_mem_13_15;
    wire REG_mem_44_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12830 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13916_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12168_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13922_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12165 ;
    wire REG_mem_31_7;
    wire REG_mem_26_7;
    wire REG_mem_14_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_7 ;
    wire REG_mem_40_14;
    wire REG_mem_8_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_0 ;
    wire REG_mem_45_14;
    wire REG_mem_50_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_12 ;
    wire REG_mem_16_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_7 ;
    wire REG_mem_15_10;
    wire REG_mem_13_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14162_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14165 ;
    wire REG_mem_12_10;
    wire REG_mem_14_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_13 ;
    wire REG_mem_4_10;
    wire REG_mem_4_14;
    wire REG_mem_48_3;
    wire REG_mem_40_3;
    wire REG_mem_51_14;
    wire REG_mem_17_10;
    wire REG_mem_63_7;
    wire REG_mem_5_3;
    wire REG_mem_50_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13700 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13652 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12237_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12228 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_3 ;
    wire REG_mem_58_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_7 ;
    wire REG_mem_8_7;
    wire REG_mem_4_3;
    wire REG_mem_15_7;
    wire REG_mem_9_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13088 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11598 ;
    wire REG_mem_11_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13334_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13337 ;
    wire REG_mem_45_3;
    wire REG_mem_46_3;
    wire REG_mem_23_10;
    wire REG_mem_10_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14354 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13757 ;
    wire REG_mem_23_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_3 ;
    wire REG_mem_47_12;
    wire REG_mem_63_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13820_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12198_cascade_ ;
    wire REG_mem_40_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13826 ;
    wire REG_mem_41_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12195 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_12 ;
    wire REG_mem_45_7;
    wire REG_mem_44_7;
    wire REG_mem_46_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12517 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12518 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12506 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13310_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13313 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13958 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12505 ;
    wire REG_mem_48_12;
    wire REG_mem_49_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12902 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12420 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12405_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12387 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12375_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12794 ;
    wire rd_addr_nxt_c_6_N_465_5_cascade_;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12153 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12138 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13034 ;
    wire bfn_7_19_0_;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10637 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10638 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10639 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10640 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10641 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10642 ;
    wire REG_mem_36_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11722 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11723_cascade_ ;
    wire REG_mem_48_0;
    wire REG_mem_50_15;
    wire REG_mem_44_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11495 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11492 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13172_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12863 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13505 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12067 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_0 ;
    wire REG_mem_39_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12932 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13151 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13148 ;
    wire REG_mem_8_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13586_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13589 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13502 ;
    wire REG_mem_23_0;
    wire REG_mem_17_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12920 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12445 ;
    wire REG_mem_40_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12941_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12815 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12095_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12094 ;
    wire REG_mem_45_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_15 ;
    wire REG_mem_12_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_0 ;
    wire REG_mem_7_14;
    wire REG_mem_40_9;
    wire REG_mem_48_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_0 ;
    wire REG_mem_41_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_12 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_13 ;
    wire n53_cascade_;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n63_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_0 ;
    wire REG_mem_50_14;
    wire REG_mem_44_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12340 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_12 ;
    wire REG_mem_46_9;
    wire REG_mem_8_3;
    wire REG_mem_40_11;
    wire REG_mem_47_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_3 ;
    wire REG_mem_44_3;
    wire REG_mem_36_12;
    wire REG_mem_37_12;
    wire REG_mem_17_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13406_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12312 ;
    wire REG_mem_16_12;
    wire REG_mem_38_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12482 ;
    wire REG_mem_4_12;
    wire REG_mem_37_11;
    wire REG_mem_36_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13427 ;
    wire REG_mem_40_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13802_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12204_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12968 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12225 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13712 ;
    wire REG_mem_44_13;
    wire REG_mem_46_13;
    wire REG_mem_55_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13508_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12276 ;
    wire REG_mem_40_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12123 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14174 ;
    wire REG_mem_8_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12075_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13076 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14126 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12102 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_12 ;
    wire REG_mem_13_13;
    wire REG_mem_12_13;
    wire REG_mem_14_13;
    wire REG_mem_7_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12884_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12887_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12953 ;
    wire REG_mem_23_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14066 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12950 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14366_cascade_ ;
    wire REG_mem_18_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14378_cascade_ ;
    wire REG_mem_16_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12471 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13436 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13439 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11986 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13670_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12013 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12020 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13676 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13679_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12083 ;
    wire REG_mem_40_15;
    wire REG_mem_7_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12344 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13706 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14156 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11998 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11999 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13673 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12080_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14114 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11732 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11731 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13565 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_14 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12184 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_0 ;
    wire REG_mem_49_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_9 ;
    wire REG_mem_23_9;
    wire REG_mem_55_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12938 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13112_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13115 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_0 ;
    wire REG_mem_23_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_0 ;
    wire REG_mem_55_0;
    wire REG_mem_41_0;
    wire REG_mem_42_0;
    wire REG_mem_9_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_15 ;
    wire REG_mem_38_14;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12356 ;
    wire REG_mem_16_0;
    wire REG_mem_39_14;
    wire REG_mem_43_0;
    wire REG_mem_43_14;
    wire REG_mem_8_14;
    wire dc32_fifo_data_in_14;
    wire REG_mem_42_14;
    wire REG_mem_7_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_nxt_c_0_cascade_ ;
    wire wr_addr_nxt_c_2_cascade_;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7612 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_0 ;
    wire REG_mem_39_12;
    wire REG_mem_41_15;
    wire n10_cascade_;
    wire REG_mem_55_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_11 ;
    wire REG_mem_41_11;
    wire REG_mem_17_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14102_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12108 ;
    wire REG_mem_16_13;
    wire REG_mem_18_13;
    wire REG_mem_19_13;
    wire REG_mem_4_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11481_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11420 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12527 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.full_max_w_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12 ;
    wire n7596_cascade_;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11831 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_13 ;
    wire REG_mem_42_13;
    wire REG_mem_40_12;
    wire REG_mem_17_11;
    wire REG_mem_47_3;
    wire REG_mem_19_12;
    wire REG_mem_41_12;
    wire REG_mem_11_13;
    wire REG_mem_9_13;
    wire REG_mem_51_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11400 ;
    wire REG_mem_23_11;
    wire rp_sync1_r_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_1 ;
    wire REG_mem_9_11;
    wire REG_mem_8_11;
    wire REG_mem_11_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14402 ;
    wire REG_mem_10_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12042 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_13 ;
    wire REG_mem_31_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13940_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13943 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14240 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_11 ;
    wire rd_grey_sync_r_1;
    wire rd_addr_nxt_c_6_N_465_3;
    wire rd_addr_nxt_c_6_N_465_5;
    wire rd_addr_nxt_c_6_N_465_1_cascade_;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13904_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12174 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_13 ;
    wire rd_grey_sync_r_0;
    wire rp_sync1_r_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_0 ;
    wire REG_mem_19_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12341 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11987 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11984 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11983 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11971 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13682_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14132 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12007 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11972 ;
    wire REG_mem_51_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_5 ;
    wire REG_mem_19_0;
    wire REG_mem_11_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13232 ;
    wire REG_mem_18_0;
    wire REG_mem_10_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12383 ;
    wire REG_mem_31_0;
    wire REG_mem_18_15;
    wire REG_mem_16_9;
    wire REG_mem_26_0;
    wire REG_mem_49_9;
    wire REG_mem_19_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12908 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12361 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12362_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12911 ;
    wire REG_mem_9_9;
    wire REG_mem_43_9;
    wire REG_mem_51_15;
    wire REG_mem_7_10;
    wire REG_mem_36_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11995 ;
    wire REG_mem_9_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_7 ;
    wire REG_mem_11_15;
    wire n26_cascade_;
    wire REG_mem_39_3;
    wire REG_mem_17_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n16_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n16 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n20_adj_1160_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12_adj_1156_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n20_adj_1160 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n36 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12_adj_1156 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.full_o ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n9_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n9 ;
    wire \INVusb3_if_inst.state_timeout_counter_i0_i2C_net ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n25 ;
    wire REG_mem_47_7;
    wire REG_mem_55_11;
    wire REG_mem_47_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11447 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10784_cascade_ ;
    wire DEBUG_3_c;
    wire afull_flag_impl_af_flag_p_w_N_603_3;
    wire afull_flag_impl_af_flag_p_w_N_603_3_cascade_;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n6_adj_1172 ;
    wire FT_OE_c;
    wire \usb3_if_inst.n551 ;
    wire \INVusb3_if_inst.FT_RD_internal_75C_net ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_sig_diff0_w_0 ;
    wire bfn_10_14_0_;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_sig_diff0_w_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10625 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_sig_diff0_w_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10626 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_sig_diff0_w_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10627 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n3_adj_1166 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11436 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10628 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11463 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10629 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11475 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10630 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_3_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11384 ;
    wire rd_grey_sync_r_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11402 ;
    wire rp_sync1_r_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_2 ;
    wire rd_grey_sync_r_3;
    wire REG_mem_9_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13430_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13433 ;
    wire REG_mem_8_12;
    wire REG_mem_10_12;
    wire REG_mem_41_13;
    wire REG_mem_7_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12299 ;
    wire rp_sync1_r_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_3 ;
    wire REG_mem_11_12;
    wire REG_mem_19_11;
    wire REG_mem_4_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12051 ;
    wire REG_mem_38_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13424 ;
    wire REG_mem_7_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14222 ;
    wire REG_mem_39_11;
    wire rd_addr_r_6;
    wire REG_mem_51_13;
    wire REG_mem_49_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13592_cascade_ ;
    wire REG_mem_48_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12255 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12453 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13154 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_13 ;
    wire REG_mem_18_12;
    wire REG_mem_26_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14144 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_13 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13874 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13877 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13043_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12058 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12926_cascade_ ;
    wire REG_mem_4_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12929 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13040 ;
    wire REG_mem_5_15;
    wire REG_mem_42_5;
    wire REG_mem_6_15;
    wire REG_mem_50_0;
    wire DEBUG_1_c_0_c;
    wire \usb3_if_inst.usb3_data_in_latched_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_7 ;
    wire REG_mem_12_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13835_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12038 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12019 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13832 ;
    wire REG_mem_13_0;
    wire REG_mem_14_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12014 ;
    wire REG_mem_47_15;
    wire REG_mem_45_15;
    wire REG_mem_15_0;
    wire REG_mem_49_2;
    wire REG_mem_10_15;
    wire REG_mem_49_15;
    wire REG_mem_48_15;
    wire REG_mem_45_11;
    wire REG_mem_50_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13976 ;
    wire REG_mem_7_15;
    wire REG_mem_51_2;
    wire REG_mem_38_9;
    wire REG_mem_41_9;
    wire REG_mem_37_15;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13202_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13205 ;
    wire REG_mem_12_9;
    wire REG_mem_5_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n15 ;
    wire REG_mem_63_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_w_6 ;
    wire wr_addr_nxt_c_4_cascade_;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n35 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n26_adj_1146 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14306 ;
    wire REG_mem_14_3;
    wire REG_mem_13_3;
    wire REG_mem_15_13;
    wire REG_mem_43_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n17 ;
    wire REG_mem_47_11;
    wire REG_mem_38_3;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13754 ;
    wire REG_mem_14_7;
    wire REG_mem_46_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_11 ;
    wire REG_mem_58_3;
    wire REG_mem_31_13;
    wire REG_mem_46_11;
    wire REG_mem_13_12;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13412_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13415 ;
    wire REG_mem_12_12;
    wire REG_mem_14_12;
    wire REG_mem_15_12;
    wire REG_mem_50_11;
    wire REG_mem_49_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14204_cascade_ ;
    wire REG_mem_48_11;
    wire REG_mem_50_13;
    wire REG_mem_47_13;
    wire REG_mem_51_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_11 ;
    wire REG_mem_5_11;
    wire REG_mem_37_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13838_cascade_ ;
    wire REG_mem_36_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12189 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_4 ;
    wire REG_mem_38_13;
    wire REG_mem_39_13;
    wire REG_mem_50_12;
    wire dc32_fifo_data_in_12;
    wire REG_mem_6_12;
    wire REG_mem_5_13;
    wire rd_grey_sync_r_4;
    wire rp_sync1_r_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_5 ;
    wire rd_grey_sync_r_5;
    wire rp_sync1_r_5;
    wire REG_mem_6_13;
    wire rp_sync1_r_6;
    wire REG_mem_13_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14396_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12456 ;
    wire REG_mem_12_11;
    wire REG_mem_14_11;
    wire REG_mem_15_11;
    wire dc32_fifo_data_in_11;
    wire REG_mem_6_11;
    wire dc32_fifo_data_in_13;
    wire REG_mem_45_13;
    wire bfn_11_18_0_;
    wire \spi0.n10694 ;
    wire \spi0.n10695 ;
    wire \spi0.n10696 ;
    wire \spi0.n10697 ;
    wire \spi0.n10698 ;
    wire \spi0.n10699 ;
    wire \spi0.n10700 ;
    wire \spi0.n10701 ;
    wire bfn_11_19_0_;
    wire \spi0.n10702 ;
    wire REG_mem_58_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13748_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_11 ;
    wire REG_mem_63_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13616_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_11 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13619_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13751 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14147 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14324_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14207 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14123_cascade_ ;
    wire REG_mem_7_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13886_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13889 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14120 ;
    wire REG_mem_5_2;
    wire REG_mem_4_2;
    wire REG_mem_48_1;
    wire REG_mem_49_1;
    wire REG_mem_47_1;
    wire REG_mem_46_1;
    wire REG_mem_41_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13742 ;
    wire REG_mem_6_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_5 ;
    wire REG_mem_45_1;
    wire REG_mem_46_15;
    wire REG_mem_40_5;
    wire REG_mem_55_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_5 ;
    wire REG_mem_4_1;
    wire REG_mem_5_1;
    wire REG_mem_36_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_0 ;
    wire REG_mem_48_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13685 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12098 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14078 ;
    wire REG_mem_10_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_9 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12382 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_9 ;
    wire REG_mem_49_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12304 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12305 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12295 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13214_cascade_ ;
    wire REG_mem_50_5;
    wire REG_mem_51_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12296 ;
    wire REG_mem_48_5;
    wire REG_mem_39_7;
    wire REG_mem_37_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13862_cascade_ ;
    wire REG_mem_36_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11762 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13562 ;
    wire REG_mem_7_0;
    wire REG_mem_14_9;
    wire REG_mem_9_7;
    wire REG_mem_13_9;
    wire REG_mem_18_9;
    wire REG_mem_15_15;
    wire dc32_fifo_data_in_10;
    wire REG_mem_47_10;
    wire REG_mem_15_3;
    wire n7596;
    wire wr_addr_nxt_c_2;
    wire wr_addr_nxt_c_4;
    wire wr_addr_r_0;
    wire wr_addr_p1_w_0;
    wire bfn_12_12_0_;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10631 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10632 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10633 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10634 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10635 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10636 ;
    wire wr_addr_p1_w_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13301 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14231 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12486 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12498 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13157 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14318_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12480 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14117 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13691 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13709 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14081 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14303 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13175 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13229 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13631 ;
    wire wr_grey_sync_r_1;
    wire REG_out_raw_10;
    wire wr_grey_sync_r_4;
    wire wp_sync1_r_4;
    wire wr_grey_sync_r_3;
    wire wp_sync1_r_3;
    wire wr_grey_sync_r_5;
    wire wp_sync1_r_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_4_cascade_ ;
    wire wp_sync1_r_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n4027 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_3_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n8_adj_1152 ;
    wire bfn_12_16_0_;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10619 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n6_adj_1150 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10620 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10621 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10622 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_sig_diff0_w_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10623 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n2_adj_1149 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_sig_diff0_w_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10624 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n8_adj_1157_cascade_ ;
    wire REG_mem_39_10;
    wire REG_mem_38_10;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11585 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n4025_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12_adj_1158 ;
    wire wr_grey_sync_r_0;
    wire wp_sync1_r_0;
    wire \spi0.counter_5 ;
    wire \spi0.counter_9 ;
    wire \spi0.counter_8 ;
    wire \spi0.counter_6 ;
    wire \spi0.counter_7 ;
    wire \spi0.counter_3 ;
    wire \spi0.counter_1 ;
    wire \spi0.counter_2 ;
    wire \spi0.counter_0 ;
    wire \spi0.n9 ;
    wire \spi0.n3909_cascade_ ;
    wire \spi0.n14 ;
    wire \spi0.n19_cascade_ ;
    wire \spi0.n88 ;
    wire \spi0.n8 ;
    wire \spi0.n12566 ;
    wire \spi0.n12567_cascade_ ;
    wire \spi0.SCLK_N_977 ;
    wire \spi0.n11351 ;
    wire \spi0.n2_cascade_ ;
    wire \spi0.n4409 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13844_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11750 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13847 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11713 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11714 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13970 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11698 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13358_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13361 ;
    wire REG_mem_43_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11705 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13745 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11489_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13217 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14258 ;
    wire REG_mem_38_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12131_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12130 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12088 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12818_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12821 ;
    wire REG_mem_7_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11507_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11506 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14276 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12509_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12508 ;
    wire REG_mem_44_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_1 ;
    wire REG_mem_40_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11704 ;
    wire REG_mem_8_1;
    wire REG_mem_9_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14288 ;
    wire REG_mem_8_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13859 ;
    wire REG_mem_44_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13577 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13574 ;
    wire REG_mem_6_0;
    wire REG_mem_6_5;
    wire REG_mem_47_5;
    wire REG_mem_38_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_2 ;
    wire REG_mem_5_5;
    wire REG_mem_5_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11761 ;
    wire REG_mem_9_0;
    wire REG_mem_19_15;
    wire REG_mem_46_5;
    wire REG_mem_11_0;
    wire REG_mem_10_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13856 ;
    wire REG_mem_43_5;
    wire REG_mem_17_7;
    wire REG_mem_11_1;
    wire REG_mem_16_7;
    wire REG_mem_7_7;
    wire REG_mem_6_7;
    wire REG_mem_4_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14072_cascade_ ;
    wire REG_mem_5_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13478 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12144 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13316 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12222 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12330_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12180 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13466 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12288 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13580 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12120 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12282 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12258_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13286 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13880_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12177 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_7 ;
    wire REG_mem_15_4;
    wire \usb3_if_inst.n2912_cascade_ ;
    wire \usb3_if_inst.n7_cascade_ ;
    wire \usb3_if_inst.n137 ;
    wire \usb3_if_inst.n3684 ;
    wire \usb3_if_inst.n138_cascade_ ;
    wire \usb3_if_inst.n2739_cascade_ ;
    wire \INVusb3_if_inst.state_timeout_counter_i0_i1C_net ;
    wire wr_grey_sync_r_6;
    wire wp_sync1_r_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6 ;
    wire wr_grey_sync_r_2;
    wire wp_sync1_r_2;
    wire REG_out_raw_7;
    wire REG_out_raw_14;
    wire REG_out_raw_13;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11445 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11408 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11483_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10760 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_fifo_en_w ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n8 ;
    wire rd_sig_diff0_w_0;
    wire rd_sig_diff0_w_1;
    wire n5_cascade_;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.genblk16_rd_prev_r ;
    wire REG_out_raw_11;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11430 ;
    wire REG_out_raw_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_0 ;
    wire rd_addr_nxt_c_6_N_465_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7_adj_1151 ;
    wire \spi0.tx_shift_reg_1 ;
    wire \spi0.tx_shift_reg_2 ;
    wire \spi0.tx_shift_reg_3 ;
    wire \spi0.tx_shift_reg_4 ;
    wire \spi0.tx_shift_reg_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n2 ;
    wire \spi0.n11317 ;
    wire \spi0.counter_4 ;
    wire \spi0.n24_cascade_ ;
    wire \spi0.n16 ;
    wire \spi0.n4105_cascade_ ;
    wire \spi0.n14442_cascade_ ;
    wire \spi0.n10119 ;
    wire \spi0.n11345 ;
    wire \spi0.n12594_cascade_ ;
    wire \spi0.n3295_cascade_ ;
    wire \spi0.n11346 ;
    wire \spi0.n11311 ;
    wire \spi0.n11311_cascade_ ;
    wire \spi0.n11344 ;
    wire \spi0.n4105 ;
    wire \spi0.n12607_cascade_ ;
    wire \spi0.n4120 ;
    wire \spi0.n12702 ;
    wire \spi0.n10106 ;
    wire \spi0.n12598_cascade_ ;
    wire \spi0.n14442 ;
    wire \spi0.CS_N_974 ;
    wire \spi0.n10082 ;
    wire \spi0.n10076_cascade_ ;
    wire \spi0.n10081 ;
    wire \spi0.n11398 ;
    wire \spi0.n11350 ;
    wire \spi0.n11398_cascade_ ;
    wire \spi0.n81 ;
    wire \spi0.n81_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11699 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12089 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_0 ;
    wire REG_mem_14_1;
    wire REG_mem_18_1;
    wire REG_mem_19_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11555 ;
    wire REG_mem_36_1;
    wire REG_mem_37_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11701 ;
    wire REG_mem_58_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13340_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13343 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_15 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11656 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11654 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11653 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13346_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11672 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11660 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11659 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13994_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11744_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13349 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13379 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11678 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13355_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13376 ;
    wire REG_mem_45_5;
    wire REG_mem_37_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13550_cascade_ ;
    wire REG_mem_36_6;
    wire REG_mem_38_6;
    wire REG_mem_39_6;
    wire REG_mem_37_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11671 ;
    wire REG_mem_12_1;
    wire REG_mem_13_1;
    wire REG_mem_42_1;
    wire REG_mem_38_1;
    wire REG_mem_39_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11702 ;
    wire REG_mem_15_1;
    wire REG_mem_39_0;
    wire REG_mem_37_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13016_cascade_ ;
    wire REG_mem_36_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13019 ;
    wire REG_mem_38_0;
    wire REG_mem_14_4;
    wire REG_mem_4_0;
    wire REG_mem_46_0;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_1 ;
    wire REG_mem_41_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14192_cascade_ ;
    wire REG_mem_14_8;
    wire REG_mem_15_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11996 ;
    wire REG_mem_38_15;
    wire REG_mem_39_15;
    wire n29;
    wire REG_mem_13_8;
    wire REG_mem_4_5;
    wire REG_mem_12_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14090_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12111 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_7 ;
    wire REG_mem_23_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13964_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12150 ;
    wire REG_mem_31_15;
    wire REG_mem_18_4;
    wire REG_mem_19_4;
    wire REG_mem_16_4;
    wire REG_mem_17_4;
    wire \usb3_if_inst.n3686_cascade_ ;
    wire \usb3_if_inst.state_timeout_counter_1 ;
    wire \usb3_if_inst.state_timeout_counter_0 ;
    wire \usb3_if_inst.n4_cascade_ ;
    wire \usb3_if_inst.n4403_cascade_ ;
    wire \usb3_if_inst.n6904 ;
    wire \usb3_if_inst.n135 ;
    wire \usb3_if_inst.n3686 ;
    wire \usb3_if_inst.state_timeout_counter_3 ;
    wire \INVusb3_if_inst.state_timeout_counter_i0_i3C_net ;
    wire \usb3_if_inst.n12582_cascade_ ;
    wire \usb3_if_inst.n4061 ;
    wire \usb3_if_inst.empty_o_N_599 ;
    wire \usb3_if_inst.num_lines_clocked_out_0 ;
    wire bfn_14_13_0_;
    wire \usb3_if_inst.n10660 ;
    wire \usb3_if_inst.num_lines_clocked_out_2 ;
    wire \usb3_if_inst.n10661 ;
    wire \usb3_if_inst.n10662 ;
    wire \usb3_if_inst.n10663 ;
    wire \usb3_if_inst.n10664 ;
    wire \usb3_if_inst.n10665 ;
    wire \usb3_if_inst.num_lines_clocked_out_7 ;
    wire \usb3_if_inst.n10666 ;
    wire \usb3_if_inst.n10667 ;
    wire \INVusb3_if_inst.num_lines_clocked_out_i0C_net ;
    wire bfn_14_14_0_;
    wire \usb3_if_inst.num_lines_clocked_out_9 ;
    wire \usb3_if_inst.n10668 ;
    wire \usb3_if_inst.n10669 ;
    wire \INVusb3_if_inst.num_lines_clocked_out_i8C_net ;
    wire \spi0.tx_shift_reg_9 ;
    wire \spi0.tx_shift_reg_10 ;
    wire \spi0.tx_shift_reg_11 ;
    wire \spi0.tx_shift_reg_12 ;
    wire \spi0.tx_shift_reg_13 ;
    wire \spi0.tx_shift_reg_8 ;
    wire \spi0.tx_shift_reg_6 ;
    wire \spi0.tx_shift_reg_7 ;
    wire tx_addr_byte_5;
    wire tx_addr_byte_1;
    wire pc_data_rx_5;
    wire tx_addr_byte_6;
    wire n10847_cascade_;
    wire pc_data_rx_0;
    wire tx_addr_byte_0;
    wire tx_addr_byte_3;
    wire tx_data_byte_5;
    wire tx_data_byte_3;
    wire n11412_cascade_;
    wire tx_data_byte_6;
    wire n11471_cascade_;
    wire tx_data_byte_1;
    wire \spi0.n12605 ;
    wire \spi0.n10090 ;
    wire multi_byte_spi_trans_flag_r;
    wire \spi0.n3 ;
    wire \spi0.state_0 ;
    wire \spi0.n12576_cascade_ ;
    wire \spi0.n37 ;
    wire \spi0.n2768 ;
    wire \spi0.n6 ;
    wire \spi0.n2768_cascade_ ;
    wire \spi0.n4260 ;
    wire \spi0.n14414 ;
    wire \spi0.state_2 ;
    wire \spi0.n19 ;
    wire \spi0.n21 ;
    wire \spi0.n10_cascade_ ;
    wire \spi0.state_1 ;
    wire \spi0.n1979_cascade_ ;
    wire \spi0.n12586 ;
    wire \spi0.state_3 ;
    wire \spi0.n19_adj_1139 ;
    wire \spi0.multi_byte_counter_0 ;
    wire bfn_14_20_0_;
    wire \spi0.n10653 ;
    wire \spi0.multi_byte_counter_2 ;
    wire \spi0.n10654 ;
    wire \spi0.n10655 ;
    wire \spi0.multi_byte_counter_4 ;
    wire \spi0.n10656 ;
    wire \spi0.n10657 ;
    wire \spi0.multi_byte_counter_6 ;
    wire \spi0.n10658 ;
    wire \spi0.n1979 ;
    wire \spi0.n10659 ;
    wire \spi0.n4281 ;
    wire \spi0.n4455 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13364 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11719 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13367 ;
    wire REG_mem_50_1;
    wire REG_mem_51_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11720 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13853 ;
    wire REG_mem_18_5;
    wire REG_mem_23_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12872_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12875_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12511_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12500 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13250_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12499 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13514 ;
    wire REG_mem_16_5;
    wire REG_mem_17_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13517 ;
    wire REG_mem_16_1;
    wire REG_mem_17_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11677 ;
    wire REG_mem_11_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13850 ;
    wire REG_mem_17_2;
    wire REG_mem_16_2;
    wire REG_mem_9_5;
    wire REG_mem_8_5;
    wire REG_mem_10_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12026_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11980 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14282_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12512 ;
    wire REG_mem_26_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11981 ;
    wire dc32_fifo_data_in_9;
    wire REG_mem_6_9;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12025 ;
    wire REG_mem_63_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13604_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_2 ;
    wire REG_mem_31_5;
    wire REG_mem_47_2;
    wire REG_mem_44_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14084_cascade_ ;
    wire REG_mem_46_2;
    wire REG_mem_19_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13982 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14168 ;
    wire REG_mem_41_2;
    wire REG_mem_40_2;
    wire REG_mem_43_2;
    wire REG_mem_63_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12986_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12989 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_5 ;
    wire REG_mem_45_2;
    wire REG_mem_47_4;
    wire REG_mem_46_4;
    wire REG_mem_45_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12992_cascade_ ;
    wire REG_mem_44_4;
    wire REG_mem_42_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13118_cascade_ ;
    wire REG_mem_40_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12995 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13121_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13622_cascade_ ;
    wire REG_mem_36_4;
    wire REG_mem_37_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13181 ;
    wire REG_mem_11_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11639 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13934_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11552 ;
    wire REG_mem_10_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13796 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11663 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11662 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11551 ;
    wire REG_mem_8_4;
    wire REG_mem_9_4;
    wire \usb3_if_inst.n2755_cascade_ ;
    wire \usb3_if_inst.n5_cascade_ ;
    wire \usb3_if_inst.n552 ;
    wire \usb3_if_inst.n554 ;
    wire \usb3_if_inst.n2798 ;
    wire \usb3_if_inst.n3973 ;
    wire \usb3_if_inst.n3973_cascade_ ;
    wire \INVusb3_if_inst.state_FSM_i2C_net ;
    wire \usb3_if_inst.n10751 ;
    wire \bluejay_data_inst.n6_cascade_ ;
    wire \usb3_if_inst.n10869 ;
    wire DEBUG_5_c;
    wire \usb3_if_inst.n555 ;
    wire \usb3_if_inst.n10746 ;
    wire DEBUG_2_c_c;
    wire \usb3_if_inst.n7360 ;
    wire \usb3_if_inst.state_timeout_counter_2 ;
    wire \usb3_if_inst.n4 ;
    wire \usb3_if_inst.n7360_cascade_ ;
    wire \usb3_if_inst.n7505 ;
    wire DATA15_c;
    wire \bluejay_data_inst.valid_N_707 ;
    wire \usb3_if_inst.n7 ;
    wire \usb3_if_inst.n4178 ;
    wire fifo_data_out_0;
    wire DATA16_c;
    wire \bluejay_data_inst.n4522 ;
    wire fifo_data_out_11;
    wire DATA11_c;
    wire fifo_data_out_10;
    wire DATA10_c;
    wire DATA9_c;
    wire \INVbluejay_data_inst.bluejay_data_out_i16C_net ;
    wire tx_data_byte_0;
    wire n4070;
    wire tx_shift_reg_0;
    wire n1928;
    wire \spi0.tx_shift_reg_14 ;
    wire \spi0.n1930 ;
    wire REG_out_raw_12;
    wire pc_data_rx_7;
    wire REG_out_raw_9;
    wire fifo_data_out_9;
    wire REG_out_raw_3;
    wire REG_out_raw_15;
    wire fifo_data_out_15;
    wire pc_data_rx_6;
    wire tx_data_byte_2;
    wire tx_addr_byte_2;
    wire n3997;
    wire pc_data_rx_2;
    wire pc_data_rx_1;
    wire pc_data_rx_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14261 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13253 ;
    wire REG_out_raw_5;
    wire n4_adj_1205;
    wire n4_adj_1206;
    wire n7455;
    wire \pc_rx.n149 ;
    wire \pc_rx.n149_cascade_ ;
    wire debug_led3;
    wire uart_rx_complete_prev;
    wire n4443;
    wire even_byte_flag;
    wire spi_start_transfer_r;
    wire tx_data_byte_7;
    wire tx_addr_byte_7;
    wire bfn_15_19_0_;
    wire \pc_rx.n10703 ;
    wire \pc_rx.n10704 ;
    wire \pc_rx.n10705 ;
    wire \pc_rx.n10706 ;
    wire \pc_rx.n10707 ;
    wire \pc_rx.n10708 ;
    wire \pc_rx.n10709 ;
    wire \pc_rx.n10710 ;
    wire bfn_15_20_0_;
    wire \pc_rx.n10711 ;
    wire \pc_rx.n6481 ;
    wire FIFO_D7_c_7;
    wire REG_mem_12_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14021 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11695 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11696_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_1 ;
    wire REG_mem_63_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11740 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11741 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11726 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13892_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11765 ;
    wire REG_mem_58_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_1 ;
    wire REG_mem_15_5;
    wire REG_mem_14_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14018 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13988 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11747 ;
    wire REG_mem_6_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11657 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13064_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13280 ;
    wire REG_mem_23_2;
    wire REG_mem_31_1;
    wire REG_mem_26_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11684 ;
    wire REG_mem_19_5;
    wire REG_mem_55_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13910_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13283 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13067 ;
    wire REG_mem_26_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13868_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_0 ;
    wire REG_mem_39_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13178 ;
    wire n27;
    wire REG_mem_38_4;
    wire REG_mem_39_5;
    wire n53;
    wire REG_mem_12_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11638 ;
    wire REG_mem_12_2;
    wire REG_mem_50_7;
    wire REG_mem_49_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13760_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12210 ;
    wire REG_mem_48_7;
    wire REG_mem_11_8;
    wire REG_mem_10_8;
    wire REG_mem_51_7;
    wire REG_mem_15_8;
    wire REG_mem_13_5;
    wire REG_mem_49_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13532_cascade_ ;
    wire REG_mem_48_8;
    wire REG_mem_51_8;
    wire REG_mem_55_7;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13718 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_7 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13736_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_4 ;
    wire bfn_16_11_0_;
    wire \bluejay_data_inst.state_timeout_counter_1 ;
    wire \bluejay_data_inst.n10581 ;
    wire \bluejay_data_inst.state_timeout_counter_2 ;
    wire \bluejay_data_inst.n86 ;
    wire \bluejay_data_inst.n10582 ;
    wire \bluejay_data_inst.n10583 ;
    wire \bluejay_data_inst.n10583_THRU_CRY_0_THRU_CO ;
    wire \bluejay_data_inst.n10583_THRU_CRY_1_THRU_CO ;
    wire \bluejay_data_inst.n10583_THRU_CRY_2_THRU_CO ;
    wire \bluejay_data_inst.n10583_THRU_CRY_3_THRU_CO ;
    wire \bluejay_data_inst.n10583_THRU_CRY_4_THRU_CO ;
    wire bfn_16_12_0_;
    wire \bluejay_data_inst.n10584 ;
    wire \bluejay_data_inst.n10584_THRU_CRY_0_THRU_CO ;
    wire \bluejay_data_inst.n10584_THRU_CRY_1_THRU_CO ;
    wire \bluejay_data_inst.n10584_THRU_CRY_2_THRU_CO ;
    wire \bluejay_data_inst.n10584_THRU_CRY_3_THRU_CO ;
    wire \bluejay_data_inst.n10584_THRU_CRY_4_THRU_CO ;
    wire \bluejay_data_inst.n10584_THRU_CRY_5_THRU_CO ;
    wire \bluejay_data_inst.n10584_THRU_CRY_6_THRU_CO ;
    wire bfn_16_13_0_;
    wire \bluejay_data_inst.n11177 ;
    wire \bluejay_data_inst.n10585 ;
    wire \bluejay_data_inst.n10585_THRU_CRY_0_THRU_CO ;
    wire \bluejay_data_inst.n10585_THRU_CRY_1_THRU_CO ;
    wire \bluejay_data_inst.n10585_THRU_CRY_2_THRU_CO ;
    wire \bluejay_data_inst.n10585_THRU_CRY_3_THRU_CO ;
    wire \bluejay_data_inst.n10585_THRU_CRY_4_THRU_CO ;
    wire \bluejay_data_inst.n10585_THRU_CRY_5_THRU_CO ;
    wire \bluejay_data_inst.n10585_THRU_CRY_6_THRU_CO ;
    wire \bluejay_data_inst.state_timeout_counter_5 ;
    wire bfn_16_14_0_;
    wire \bluejay_data_inst.n10586 ;
    wire \bluejay_data_inst.n10586_THRU_CRY_0_THRU_CO ;
    wire \bluejay_data_inst.n10586_THRU_CRY_1_THRU_CO ;
    wire \bluejay_data_inst.n10586_THRU_CRY_2_THRU_CO ;
    wire \bluejay_data_inst.n10586_THRU_CRY_3_THRU_CO ;
    wire \bluejay_data_inst.n10586_THRU_CRY_4_THRU_CO ;
    wire GNDG0;
    wire \bluejay_data_inst.n10586_THRU_CRY_5_THRU_CO ;
    wire \bluejay_data_inst.n10586_THRU_CRY_6_THRU_CO ;
    wire \bluejay_data_inst.state_timeout_counter_6 ;
    wire bfn_16_15_0_;
    wire \bluejay_data_inst.n10587 ;
    wire \bluejay_data_inst.state_timeout_counter_7 ;
    wire \pc_rx.r_Rx_Data_R ;
    wire n4002;
    wire n4002_cascade_;
    wire n4;
    wire pc_data_rx_3;
    wire REG_out_raw_1;
    wire \pc_rx.r_Bit_Index_2 ;
    wire \pc_rx.r_Bit_Index_0 ;
    wire \pc_rx.r_Bit_Index_1 ;
    wire \pc_rx.n4470 ;
    wire \pc_rx.n55_adj_1144_cascade_ ;
    wire \pc_rx.n145 ;
    wire \pc_rx.n145_cascade_ ;
    wire \pc_rx.n6490 ;
    wire \pc_rx.n4081 ;
    wire \pc_rx.n4140 ;
    wire \pc_rx.n151 ;
    wire \pc_rx.r_SM_Main_1 ;
    wire \pc_rx.n6515 ;
    wire \pc_rx.r_SM_Main_2 ;
    wire \pc_rx.r_Clock_Count_9 ;
    wire \pc_rx.r_Clock_Count_6 ;
    wire \pc_rx.r_Clock_Count_5 ;
    wire \pc_rx.n4_adj_1145_cascade_ ;
    wire \pc_rx.r_SM_Main_2_N_732_2 ;
    wire \pc_rx.r_Clock_Count_8 ;
    wire \pc_rx.r_Clock_Count_7 ;
    wire \pc_rx.n6 ;
    wire \pc_rx.r_Clock_Count_4 ;
    wire \pc_rx.r_Clock_Count_1 ;
    wire \pc_rx.r_Clock_Count_0 ;
    wire \pc_rx.r_Clock_Count_3 ;
    wire \pc_rx.n140 ;
    wire \pc_rx.n8_cascade_ ;
    wire \pc_rx.r_Clock_Count_2 ;
    wire \pc_rx.n13_cascade_ ;
    wire \pc_rx.n6500 ;
    wire n10562_cascade_;
    wire reset_clk_counter_1;
    wire reset_clk_counter_3;
    wire reset_clk_counter_2;
    wire reset_all_w_N_61;
    wire reset_all_w_N_61_cascade_;
    wire reset_clk_counter_0;
    wire \pc_rx.r_SM_Main_0 ;
    wire r_Rx_Data;
    wire \pc_rx.n13 ;
    wire \pc_rx.n125 ;
    wire FIFO_D4_c_4;
    wire FIFO_D5_c_5;
    wire FIFO_D6_c_6;
    wire FIFO_D3_c_3;
    wire \usb3_if_inst.usb3_data_in_latched_3 ;
    wire dc32_fifo_data_in_3;
    wire \usb3_if_inst.usb3_data_in_latched_4 ;
    wire \usb3_if_inst.usb3_data_in_latched_5 ;
    wire \usb3_if_inst.usb3_data_in_latched_6 ;
    wire \usb3_if_inst.usb3_data_in_latched_7 ;
    wire \INVusb3_if_inst.dc32_fifo_data_in_i2C_net ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12030 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12114 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12078 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12944 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13607 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13979 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14408_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13913 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14411_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12947 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11498_cascade_ ;
    wire REG_out_raw_2;
    wire REG_mem_36_2;
    wire REG_mem_37_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12057 ;
    wire REG_mem_58_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14198_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_4 ;
    wire REG_mem_42_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14360 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12848_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12851_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14363 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12377_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12376 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12346 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13010_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13013 ;
    wire REG_mem_38_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14210 ;
    wire REG_mem_41_4;
    wire n26;
    wire REG_mem_39_2;
    wire REG_mem_18_2;
    wire REG_mem_19_2;
    wire REG_mem_26_2;
    wire REG_mem_31_2;
    wire REG_mem_48_4;
    wire n16;
    wire REG_mem_49_4;
    wire dc32_fifo_data_in_5;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_5 ;
    wire dc32_fifo_data_in_15;
    wire REG_mem_26_15;
    wire REG_mem_7_4;
    wire REG_mem_6_4;
    wire REG_mem_13_2;
    wire REG_mem_39_8;
    wire REG_mem_38_8;
    wire n28;
    wire REG_mem_13_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_7 ;
    wire dc32_fifo_data_in_7;
    wire REG_mem_18_7;
    wire REG_mem_63_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14138 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11755 ;
    wire n50;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11756 ;
    wire REG_mem_23_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13418_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13421 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_4 ;
    wire \usb3_if_inst.n534 ;
    wire \usb3_if_inst.n550 ;
    wire \usb3_if_inst.n553 ;
    wire \INVusb3_if_inst.state_FSM_i3C_net ;
    wire \bluejay_data_inst.n8_cascade_ ;
    wire \bluejay_data_inst.n12_adj_1179 ;
    wire \bluejay_data_inst.state_timeout_counter_0 ;
    wire \bluejay_data_inst.state_timeout_counter_4 ;
    wire \bluejay_data_inst.n12 ;
    wire n7_cascade_;
    wire state_timeout_counter_3;
    wire n7;
    wire \bluejay_data_inst.n10745 ;
    wire DEBUG_9_c;
    wire dc32_fifo_almost_empty;
    wire \bluejay_data_inst.n714 ;
    wire \bluejay_data_inst.n717 ;
    wire \bluejay_data_inst.n108_cascade_ ;
    wire \bluejay_data_inst.n4062_cascade_ ;
    wire \bluejay_data_inst.n108 ;
    wire \bluejay_data_inst.n4519 ;
    wire \tx_fifo.lscc_fifo_inst.n13952 ;
    wire \usb3_if_inst.num_lines_clocked_out_3 ;
    wire \usb3_if_inst.num_lines_clocked_out_6 ;
    wire \usb3_if_inst.num_lines_clocked_out_10 ;
    wire \usb3_if_inst.n18 ;
    wire \usb3_if_inst.num_lines_clocked_out_8 ;
    wire \usb3_if_inst.num_lines_clocked_out_4 ;
    wire \usb3_if_inst.n20_cascade_ ;
    wire \usb3_if_inst.n21 ;
    wire \usb3_if_inst.num_lines_clocked_out_5 ;
    wire \usb3_if_inst.num_lines_clocked_out_1 ;
    wire \usb3_if_inst.n16 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_6 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_6 ;
    wire rx_shift_reg_5;
    wire rx_shift_reg_4;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_7 ;
    wire rx_shift_reg_7;
    wire rx_shift_reg_6;
    wire rx_buf_byte_6;
    wire rx_shift_reg_0;
    wire rx_shift_reg_1;
    wire rx_shift_reg_2;
    wire n4093;
    wire n3204;
    wire rx_shift_reg_3;
    wire fifo_data_out_8;
    wire DATA8_c;
    wire fifo_data_out_7;
    wire DATA7_c;
    wire fifo_data_out_4;
    wire DATA20_c;
    wire fifo_data_out_3;
    wire DATA19_c;
    wire fifo_data_out_2;
    wire DATA18_c;
    wire fifo_data_out_1;
    wire DATA17_c;
    wire fifo_data_out_5;
    wire DATA5_c;
    wire fifo_data_out_6;
    wire DATA6_c;
    wire \INVbluejay_data_inst.bluejay_data_out_i9C_net ;
    wire wr_addr_p1_w_2_cascade_;
    wire FIFO_D8_c_8;
    wire FIFO_D2_c_2;
    wire \usb3_if_inst.usb3_data_in_latched_2 ;
    wire FIFO_D1_c_1;
    wire \usb3_if_inst.usb3_data_in_latched_1 ;
    wire \usb3_if_inst.usb3_data_in_latched_8 ;
    wire \INVusb3_if_inst.dc32_fifo_data_in_i9C_net ;
    wire REG_mem_17_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13658_cascade_ ;
    wire n49;
    wire REG_mem_16_6;
    wire REG_mem_18_6;
    wire REG_mem_19_6;
    wire REG_mem_10_6;
    wire REG_mem_11_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_2 ;
    wire n24_adj_1185;
    wire n25;
    wire n59;
    wire n18;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11681_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13352 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11857 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13238_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11807 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12347 ;
    wire n55;
    wire REG_mem_10_2;
    wire n54;
    wire REG_mem_11_2;
    wire REG_mem_8_2;
    wire REG_mem_9_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11806 ;
    wire REG_mem_50_4;
    wire REG_mem_51_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14348 ;
    wire n48;
    wire REG_mem_17_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14108_cascade_ ;
    wire REG_mem_16_8;
    wire n47;
    wire REG_mem_18_8;
    wire n57;
    wire n56;
    wire REG_mem_37_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13808 ;
    wire REG_mem_36_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12521 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12515 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13784_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12514 ;
    wire n60;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_4 ;
    wire n2;
    wire REG_mem_63_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13382_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_8 ;
    wire n22;
    wire REG_mem_43_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_8 ;
    wire REG_mem_5_4;
    wire REG_mem_4_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12520 ;
    wire n23;
    wire bfn_18_11_0_;
    wire \bluejay_data_inst.n10643 ;
    wire \bluejay_data_inst.n10644 ;
    wire \bluejay_data_inst.n10645 ;
    wire \bluejay_data_inst.n10646 ;
    wire \bluejay_data_inst.n10647 ;
    wire \bluejay_data_inst.n10648 ;
    wire \bluejay_data_inst.n10649 ;
    wire \bluejay_data_inst.n10650 ;
    wire bfn_18_12_0_;
    wire \bluejay_data_inst.n10651 ;
    wire \bluejay_data_inst.n10652 ;
    wire \bluejay_data_inst.v_counter_10 ;
    wire \bluejay_data_inst.v_counter_9 ;
    wire \bluejay_data_inst.v_counter_7 ;
    wire \bluejay_data_inst.v_counter_1 ;
    wire \bluejay_data_inst.n11418_cascade_ ;
    wire \bluejay_data_inst.n11330 ;
    wire \bluejay_data_inst.v_counter_2 ;
    wire \bluejay_data_inst.v_counter_4 ;
    wire \bluejay_data_inst.v_counter_8 ;
    wire \bluejay_data_inst.v_counter_0 ;
    wire \bluejay_data_inst.n10_adj_1180_cascade_ ;
    wire \bluejay_data_inst.n14 ;
    wire \bluejay_data_inst.n10 ;
    wire \bluejay_data_inst.v_counter_5 ;
    wire \bluejay_data_inst.v_counter_3 ;
    wire \bluejay_data_inst.n10_cascade_ ;
    wire \bluejay_data_inst.v_counter_6 ;
    wire \bluejay_data_inst.n10781 ;
    wire \bluejay_data_inst.n4162 ;
    wire buffer_switch_done_latched;
    wire \bluejay_data_inst.n21 ;
    wire fifo_data_out_13;
    wire DATA13_c;
    wire fifo_data_out_12;
    wire DATA12_c;
    wire \bluejay_data_inst.n7424 ;
    wire \bluejay_data_inst.n4062 ;
    wire \bluejay_data_inst.bluejay_data_out_31__N_701 ;
    wire \bluejay_data_inst.n4442 ;
    wire \bluejay_data_inst.bluejay_data_out_31__N_702 ;
    wire get_next_word;
    wire bluejay_data_out_31__N_704;
    wire fifo_data_out_14;
    wire bluejay_data_out_31__N_703;
    wire DATA14_c;
    wire \INVbluejay_data_inst.bluejay_data_out_i14C_net ;
    wire \tx_fifo.lscc_fifo_inst.n13544_cascade_ ;
    wire \tx_fifo.lscc_fifo_inst.n13694_cascade_ ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_5 ;
    wire \tx_fifo.lscc_fifo_inst.n13766_cascade_ ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_2 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_2 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_4 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4 ;
    wire rx_buf_byte_7;
    wire tx_data_byte_4;
    wire uart_rx_complete_rising_edge;
    wire tx_addr_byte_4;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_5 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5 ;
    wire rx_buf_byte_5;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_4 ;
    wire \tx_fifo.lscc_fifo_inst.n3_adj_1136_cascade_ ;
    wire \tx_fifo.lscc_fifo_inst.n4_cascade_ ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0 ;
    wire \tx_fifo.lscc_fifo_inst.n3_adj_1136 ;
    wire rx_buf_byte_0;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_0 ;
    wire n11424_cascade_;
    wire n15_cascade_;
    wire full_nxt_r;
    wire rx_buf_byte_4;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4 ;
    wire spi_rx_byte_ready;
    wire is_tx_fifo_full_flag;
    wire rd_addr_p1_w_1;
    wire rd_addr_p1_w_2;
    wire rd_addr_p1_w_2_cascade_;
    wire RESET_c;
    wire \tx_fifo.lscc_fifo_inst.wr_addr_p1_w_1_cascade_ ;
    wire n1;
    wire n10727;
    wire wr_addr_r_2;
    wire rd_addr_r_2;
    wire \tx_fifo.lscc_fifo_inst.n3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13598_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13634_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13637_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13601 ;
    wire REG_mem_31_6;
    wire REG_mem_26_6;
    wire REG_mem_31_4;
    wire n39;
    wire REG_mem_26_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13778 ;
    wire REG_mem_8_6;
    wire REG_mem_9_6;
    wire n52;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12008 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11680 ;
    wire REG_mem_63_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14294_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n63 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n61_adj_1154 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_6 ;
    wire REG_mem_23_1;
    wire dc32_fifo_data_in_0;
    wire REG_mem_58_0;
    wire REG_mem_5_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_6 ;
    wire REG_mem_58_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_2 ;
    wire REG_mem_15_2;
    wire REG_mem_14_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11858 ;
    wire n14;
    wire n46;
    wire REG_mem_19_8;
    wire REG_mem_47_6;
    wire n20;
    wire n21;
    wire REG_mem_46_6;
    wire n61;
    wire REG_mem_4_6;
    wire n34;
    wire REG_mem_31_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_8 ;
    wire REG_mem_23_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14060_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_8 ;
    wire n15_adj_1184;
    wire REG_mem_50_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13871 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13739 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12182_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13799 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13787 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13937 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12066 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12093 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12006 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13610_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12240 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12246_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12183 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13442_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12162 ;
    wire REG_out_raw_4;
    wire \timing_controller_inst.n11375_cascade_ ;
    wire \timing_controller_inst.n4200 ;
    wire n11376;
    wire n11376_cascade_;
    wire \timing_controller_inst.invert_N_309 ;
    wire \usb3_if_inst.reset_per_frame_latched ;
    wire reset_per_frame;
    wire buffer_switch_done;
    wire reset_all;
    wire mem_LUT_data_raw_r_4;
    wire fifo_temp_output_4;
    wire mem_LUT_data_raw_r_5;
    wire fifo_temp_output_5;
    wire mem_LUT_data_raw_r_6;
    wire fifo_temp_output_6;
    wire mem_LUT_data_raw_r_7;
    wire fifo_temp_output_7;
    wire rx_buf_byte_2;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2 ;
    wire \spi0.multi_byte_counter_7 ;
    wire \spi0.multi_byte_counter_5 ;
    wire \spi0.multi_byte_counter_3 ;
    wire \spi0.multi_byte_counter_1 ;
    wire \spi0.n14_adj_1140 ;
    wire \timing_controller_inst.n62 ;
    wire \timing_controller_inst.n49 ;
    wire rx_buf_byte_3;
    wire \tx_fifo.lscc_fifo_inst.n4 ;
    wire rx_buf_byte_1;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_3 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3 ;
    wire wr_addr_r_1;
    wire n32_cascade_;
    wire fifo_write_cmd;
    wire \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r ;
    wire n2207;
    wire empty_o_N_1116;
    wire fifo_read_cmd;
    wire wr_addr_r_0_adj_1181;
    wire n11410;
    wire n4_adj_1186_cascade_;
    wire n24;
    wire is_fifo_empty_flag;
    wire REG_mem_12_6;
    wire REG_mem_13_6;
    wire REG_mem_15_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13772 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_8 ;
    wire n51;
    wire REG_mem_14_6;
    wire REG_mem_43_6;
    wire REG_mem_42_6;
    wire REG_mem_41_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13520_cascade_ ;
    wire REG_mem_40_6;
    wire REG_mem_51_6;
    wire REG_mem_50_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12782_cascade_ ;
    wire REG_mem_49_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12785 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14390_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12459 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11634 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13004 ;
    wire REG_mem_55_6;
    wire n42;
    wire REG_mem_23_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13646_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_6 ;
    wire REG_mem_58_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13730_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13733 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14372 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12474 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_2 ;
    wire dc32_fifo_data_in_2;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_2 ;
    wire n17;
    wire REG_mem_48_6;
    wire REG_mem_44_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13388 ;
    wire REG_mem_45_6;
    wire REG_mem_55_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14216_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12054 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n45 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_4 ;
    wire n10;
    wire REG_mem_55_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13460_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n47 ;
    wire dc32_fifo_data_in_4;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n49 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n65 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_6 ;
    wire REG_mem_5_8;
    wire REG_mem_4_8;
    wire \pc_tx.n12133_cascade_ ;
    wire \pc_tx.o_Tx_Serial_N_840_cascade_ ;
    wire UART_TX_c;
    wire r_Tx_Data_3;
    wire \pc_tx.n12134 ;
    wire r_Tx_Data_5;
    wire r_Tx_Data_4;
    wire \pc_tx.n12139_cascade_ ;
    wire \pc_tx.n13790 ;
    wire r_Tx_Data_7;
    wire r_Tx_Data_6;
    wire \pc_tx.n12140 ;
    wire \bluejay_data_inst.n710 ;
    wire n718;
    wire \bluejay_data_inst.n715 ;
    wire \bluejay_data_inst.n1137 ;
    wire n4_adj_1182;
    wire n3514;
    wire n4_adj_1182_cascade_;
    wire n12601;
    wire \timing_controller_inst.n53 ;
    wire \timing_controller_inst.n1740 ;
    wire \timing_controller_inst.n1742 ;
    wire \timing_controller_inst.n1739 ;
    wire \timing_controller_inst.n1736 ;
    wire \timing_controller_inst.n1754 ;
    wire \timing_controller_inst.n1735 ;
    wire \timing_controller_inst.n1734 ;
    wire fifo_temp_output_0;
    wire r_Tx_Data_0;
    wire fifo_temp_output_1;
    wire r_Tx_Data_1;
    wire mem_LUT_data_raw_r_2;
    wire fifo_temp_output_2;
    wire r_Tx_Data_2;
    wire reset_all_w;
    wire n4249;
    wire fifo_temp_output_3;
    wire \timing_controller_inst.n55 ;
    wire \timing_controller_inst.n56 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_1 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_1 ;
    wire \tx_fifo.lscc_fifo_inst.n13538_cascade_ ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1 ;
    wire mem_LUT_data_raw_r_1;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_7 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7 ;
    wire rd_addr_r_0;
    wire \tx_fifo.lscc_fifo_inst.n14234 ;
    wire \tx_fifo.lscc_fifo_inst.n13556 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_3 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3 ;
    wire mem_LUT_data_raw_r_3;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0 ;
    wire \tx_fifo.lscc_fifo_inst.n13496 ;
    wire \tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_0 ;
    wire rd_addr_r_1;
    wire mem_LUT_data_raw_r_0;
    wire rd_fifo_en_w;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13649 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13946 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13661 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13949 ;
    wire REG_out_raw_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13007 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14342 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12315 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11844 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11838 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13370_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13373 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13775 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13781 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12002_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12003 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13568_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11835 ;
    wire REG_mem_6_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11789 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11788 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11785 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13526 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11786_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13529 ;
    wire REG_mem_7_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_6 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_6 ;
    wire n7_adj_1183;
    wire REG_mem_58_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13448_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n59 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14042 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13928_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n42 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n40 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11718 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11709 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13136_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11691 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11874 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11862 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11853 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13082_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11841 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11913_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11898 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13058_cascade_ ;
    wire REG_out_raw_8;
    wire t_rd_fifo_en_w;
    wire n11339_cascade_;
    wire tx_uart_active_flag;
    wire n3710;
    wire r_SM_Main_2_N_811_0;
    wire \timing_controller_inst.n50 ;
    wire UPDATE_c_3;
    wire \timing_controller_inst.n5 ;
    wire n7495_cascade_;
    wire \timing_controller_inst.n1875 ;
    wire n7566;
    wire n63;
    wire n1876;
    wire n1721_cascade_;
    wire \timing_controller_inst.n11347_cascade_ ;
    wire \timing_controller_inst.n4586 ;
    wire state_2;
    wire n3929;
    wire \timing_controller_inst.n54 ;
    wire \timing_controller_inst.n1751_cascade_ ;
    wire \timing_controller_inst.n1732_cascade_ ;
    wire \timing_controller_inst.n1731 ;
    wire \timing_controller_inst.n1730_cascade_ ;
    wire \timing_controller_inst.n1745_cascade_ ;
    wire n1721;
    wire state_1;
    wire \timing_controller_inst.n1793 ;
    wire \timing_controller_inst.n1744_cascade_ ;
    wire \timing_controller_inst.n11368 ;
    wire \timing_controller_inst.n52 ;
    wire \timing_controller_inst.n38_cascade_ ;
    wire \timing_controller_inst.n58 ;
    wire n25_adj_1187;
    wire bfn_23_5_0_;
    wire n24_adj_1188;
    wire n10670;
    wire n23_adj_1189;
    wire n10671;
    wire n22_adj_1190;
    wire n10672;
    wire n21_adj_1191;
    wire n10673;
    wire n20_adj_1192;
    wire n10674;
    wire n19_adj_1193;
    wire n10675;
    wire n18_adj_1194;
    wire n10676;
    wire n10677;
    wire n17_adj_1195;
    wire bfn_23_6_0_;
    wire n16_adj_1196;
    wire n10678;
    wire n15_adj_1197;
    wire n10679;
    wire n14_adj_1198;
    wire n10680;
    wire n13;
    wire n10681;
    wire n12;
    wire n10682;
    wire n11;
    wire n10683;
    wire n10_adj_1199;
    wire n10684;
    wire n10685;
    wire n9;
    wire bfn_23_7_0_;
    wire n8;
    wire n10686;
    wire n7_adj_1200;
    wire n10687;
    wire n6;
    wire n10688;
    wire n5_adj_1201;
    wire n10689;
    wire n4_adj_1202;
    wire n10690;
    wire n3;
    wire n10691;
    wire n2_adj_1203;
    wire n10692;
    wire n10693;
    wire bfn_23_8_0_;
    wire DEBUG_0_c_24;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n44 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13070_cascade_ ;
    wire REG_mem_6_8;
    wire REG_mem_7_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12824 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14246 ;
    wire REG_mem_9_8;
    wire REG_mem_8_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11646_cascade_ ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11667 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_8 ;
    wire n4133;
    wire \pc_tx.n4468 ;
    wire \pc_tx.n4_cascade_ ;
    wire \pc_tx.n8 ;
    wire \pc_tx.n7 ;
    wire \pc_tx.n2813 ;
    wire r_SM_Main_2_N_808_1_cascade_;
    wire r_SM_Main_0;
    wire r_SM_Main_1;
    wire r_SM_Main_2_N_808_1;
    wire \pc_tx.r_SM_Main_2_N_805_0 ;
    wire \pc_tx.r_Bit_Index_1 ;
    wire \pc_tx.r_Bit_Index_2 ;
    wire r_Bit_Index_0;
    wire n11319;
    wire \timing_controller_inst.n7592 ;
    wire \timing_controller_inst.n7 ;
    wire state_3;
    wire state_0;
    wire \timing_controller_inst.n11377 ;
    wire r_SM_Main_2;
    wire GB_BUFFER_DEBUG_6_c_c_THRU_CO;
    wire GB_BUFFER_SLM_CLK_c_THRU_CO;
    wire \timing_controller_inst.state_timeout_counter_0 ;
    wire \timing_controller_inst.n12532 ;
    wire bfn_23_13_0_;
    wire \timing_controller_inst.state_timeout_counter_1 ;
    wire \timing_controller_inst.n12554 ;
    wire \timing_controller_inst.n10588 ;
    wire n7383;
    wire \timing_controller_inst.state_timeout_counter_2 ;
    wire \timing_controller_inst.n12553 ;
    wire \timing_controller_inst.n10589 ;
    wire \timing_controller_inst.state_timeout_counter_3 ;
    wire \timing_controller_inst.n12552 ;
    wire \timing_controller_inst.n10590 ;
    wire \timing_controller_inst.state_timeout_counter_4 ;
    wire \timing_controller_inst.n12604 ;
    wire \timing_controller_inst.n10591 ;
    wire \timing_controller_inst.n11347 ;
    wire \timing_controller_inst.state_timeout_counter_5 ;
    wire \timing_controller_inst.n12555 ;
    wire \timing_controller_inst.n10592 ;
    wire \timing_controller_inst.state_timeout_counter_6 ;
    wire \timing_controller_inst.n10593 ;
    wire \timing_controller_inst.state_timeout_counter_7 ;
    wire \timing_controller_inst.n10594 ;
    wire \timing_controller_inst.n10595 ;
    wire \timing_controller_inst.state_timeout_counter_8 ;
    wire bfn_23_14_0_;
    wire \timing_controller_inst.state_timeout_counter_9 ;
    wire \timing_controller_inst.n12551 ;
    wire \timing_controller_inst.n10596 ;
    wire \timing_controller_inst.state_timeout_counter_10 ;
    wire \timing_controller_inst.n12550 ;
    wire \timing_controller_inst.n10597 ;
    wire \timing_controller_inst.state_timeout_counter_11 ;
    wire \timing_controller_inst.n10598 ;
    wire \timing_controller_inst.state_timeout_counter_12 ;
    wire \timing_controller_inst.n12549 ;
    wire \timing_controller_inst.n10599 ;
    wire \timing_controller_inst.state_timeout_counter_13 ;
    wire \timing_controller_inst.n10600 ;
    wire \timing_controller_inst.state_timeout_counter_14 ;
    wire \timing_controller_inst.n12548 ;
    wire \timing_controller_inst.n10601 ;
    wire \timing_controller_inst.state_timeout_counter_15 ;
    wire \timing_controller_inst.n12547 ;
    wire \timing_controller_inst.n10602 ;
    wire \timing_controller_inst.n10603 ;
    wire \timing_controller_inst.state_timeout_counter_16 ;
    wire bfn_23_15_0_;
    wire \timing_controller_inst.state_timeout_counter_17 ;
    wire \timing_controller_inst.n10604 ;
    wire \timing_controller_inst.state_timeout_counter_18 ;
    wire \timing_controller_inst.n12545 ;
    wire \timing_controller_inst.n10605 ;
    wire \timing_controller_inst.state_timeout_counter_19 ;
    wire \timing_controller_inst.n12544 ;
    wire \timing_controller_inst.n10606 ;
    wire \timing_controller_inst.state_timeout_counter_20 ;
    wire \timing_controller_inst.n12542 ;
    wire \timing_controller_inst.n10607 ;
    wire \timing_controller_inst.state_timeout_counter_21 ;
    wire \timing_controller_inst.n10608 ;
    wire \timing_controller_inst.state_timeout_counter_22 ;
    wire \timing_controller_inst.n12541 ;
    wire \timing_controller_inst.n10609 ;
    wire \timing_controller_inst.state_timeout_counter_23 ;
    wire \timing_controller_inst.n12540 ;
    wire \timing_controller_inst.n10610 ;
    wire \timing_controller_inst.n10611 ;
    wire n1616;
    wire \timing_controller_inst.state_timeout_counter_24 ;
    wire \timing_controller_inst.n12539 ;
    wire bfn_23_16_0_;
    wire \timing_controller_inst.state_timeout_counter_25 ;
    wire \timing_controller_inst.n10612 ;
    wire \timing_controller_inst.state_timeout_counter_26 ;
    wire \timing_controller_inst.n10613 ;
    wire \timing_controller_inst.state_timeout_counter_27 ;
    wire \timing_controller_inst.n10614 ;
    wire \timing_controller_inst.state_timeout_counter_28 ;
    wire \timing_controller_inst.n10615 ;
    wire \timing_controller_inst.state_timeout_counter_29 ;
    wire \timing_controller_inst.n10616 ;
    wire \timing_controller_inst.state_timeout_counter_30 ;
    wire \timing_controller_inst.n10617 ;
    wire CONSTANT_ONE_NET;
    wire \timing_controller_inst.n10618 ;
    wire \timing_controller_inst.state_timeout_counter_31 ;
    wire \timing_controller_inst.n4301 ;
    wire \timing_controller_inst.n4589 ;
    wire REG_mem_43_8;
    wire REG_mem_42_8;
    wire REG_mem_40_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13724_cascade_ ;
    wire REG_mem_41_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11811_cascade_ ;
    wire REG_mem_47_8;
    wire REG_mem_44_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13640_cascade_ ;
    wire REG_mem_45_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11820 ;
    wire n58;
    wire REG_mem_7_1;
    wire dc32_fifo_data_in_8;
    wire n19;
    wire REG_mem_46_8;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11683 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11725 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n55 ;
    wire dc32_fifo_data_in_1;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_6 ;
    wire dc32_fifo_data_in_6;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_6 ;
    wire DEBUG_6_c_c;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11784 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13130 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11760 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11901 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14012 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_8 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11736 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13304 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13073 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12827 ;
    wire \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11880 ;
    wire \pc_tx.r_Clock_Count_0 ;
    wire bfn_24_11_0_;
    wire \pc_tx.r_Clock_Count_1 ;
    wire \pc_tx.n10712 ;
    wire \pc_tx.r_Clock_Count_2 ;
    wire \pc_tx.n10713 ;
    wire \pc_tx.r_Clock_Count_3 ;
    wire \pc_tx.n10714 ;
    wire \pc_tx.r_Clock_Count_4 ;
    wire \pc_tx.n10715 ;
    wire \pc_tx.r_Clock_Count_5 ;
    wire \pc_tx.n10716 ;
    wire \pc_tx.r_Clock_Count_6 ;
    wire \pc_tx.n10717 ;
    wire \pc_tx.r_Clock_Count_7 ;
    wire \pc_tx.n10718 ;
    wire \pc_tx.n10719 ;
    wire \pc_tx.r_Clock_Count_8 ;
    wire bfn_24_12_0_;
    wire \pc_tx.n10720 ;
    wire \pc_tx.r_Clock_Count_9 ;
    wire _gnd_net_;
    wire SLM_CLK_c;
    wire \pc_tx.n1 ;
    wire \pc_tx.n4577 ;

    defparam \clock_inst.pll_config .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \clock_inst.pll_config .TEST_MODE=1'b0;
    defparam \clock_inst.pll_config .SHIFTREG_DIV_MODE=2'b00;
    defparam \clock_inst.pll_config .PLLOUT_SELECT="GENCLK";
    defparam \clock_inst.pll_config .FILTER_RANGE=3'b001;
    defparam \clock_inst.pll_config .FEEDBACK_PATH="SIMPLE";
    defparam \clock_inst.pll_config .FDA_RELATIVE=4'b0000;
    defparam \clock_inst.pll_config .FDA_FEEDBACK=4'b0000;
    defparam \clock_inst.pll_config .ENABLE_ICEGATE=1'b0;
    defparam \clock_inst.pll_config .DIVR=4'b0001;
    defparam \clock_inst.pll_config .DIVQ=3'b100;
    defparam \clock_inst.pll_config .DIVF=7'b1010010;
    defparam \clock_inst.pll_config .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \clock_inst.pll_config  (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__32914),
            .RESETB(N__86663),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7}),
            .PLLOUTGLOBAL(pll_clk_unbuf));
    PRE_IO_GBUF DEBUG_6_c_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__98336),
            .GLOBALBUFFEROUTPUT(DEBUG_6_c_c));
    defparam DEBUG_6_c_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_6_c_pad_iopad.PULLUP=1'b0;
    IO_PAD DEBUG_6_c_pad_iopad (
            .OE(N__98338),
            .DIN(N__98337),
            .DOUT(N__98336),
            .PACKAGEPIN(FIFO_CLK));
    defparam DEBUG_6_c_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_6_c_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_6_c_pad_preio (
            .PADOEN(N__98338),
            .PADOUT(N__98337),
            .PADIN(N__98336),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA4_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA4_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA4_pad_iopad (
            .OE(N__98327),
            .DIN(N__98326),
            .DOUT(N__98325),
            .PACKAGEPIN(DATA4));
    defparam DATA4_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA4_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA4_pad_preio (
            .PADOEN(N__98327),
            .PADOUT(N__98326),
            .PADIN(N__98325),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__64968),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA17_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA17_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA17_pad_iopad (
            .OE(N__98318),
            .DIN(N__98317),
            .DOUT(N__98316),
            .PACKAGEPIN(DATA17));
    defparam DATA17_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA17_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA17_pad_preio (
            .PADOEN(N__98318),
            .PADOUT(N__98317),
            .PADIN(N__98316),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65413),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D10_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D10_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D10_pad_iopad (
            .OE(N__98309),
            .DIN(N__98308),
            .DOUT(N__98307),
            .PACKAGEPIN(FIFO_D10));
    defparam FIFO_D10_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D10_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D10_pad_preio (
            .PADOEN(N__98309),
            .PADOUT(N__98308),
            .PADIN(N__98307),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D10_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D13_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D13_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D13_pad_iopad (
            .OE(N__98300),
            .DIN(N__98299),
            .DOUT(N__98298),
            .PACKAGEPIN(FIFO_D13));
    defparam FIFO_D13_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D13_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D13_pad_preio (
            .PADOEN(N__98300),
            .PADOUT(N__98299),
            .PADIN(N__98298),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D13_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_3_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_3_pad_iopad.PULLUP=1'b0;
    IO_PAD DEBUG_3_pad_iopad (
            .OE(N__98291),
            .DIN(N__98290),
            .DOUT(N__98289),
            .PACKAGEPIN(DEBUG_3));
    defparam DEBUG_3_pad_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_3_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_3_pad_preio (
            .PADOEN(N__98291),
            .PADOUT(N__98290),
            .PADIN(N__98289),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__44017),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA20_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA20_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA20_pad_iopad (
            .OE(N__98282),
            .DIN(N__98281),
            .DOUT(N__98280),
            .PACKAGEPIN(DATA20));
    defparam DATA20_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA20_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA20_pad_preio (
            .PADOEN(N__98282),
            .PADOUT(N__98281),
            .PADIN(N__98280),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__64972),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D7_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D7_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D7_pad_iopad (
            .OE(N__98273),
            .DIN(N__98272),
            .DOUT(N__98271),
            .PACKAGEPIN(FIFO_D7));
    defparam FIFO_D7_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D7_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D7_pad_preio (
            .PADOEN(N__98273),
            .PADOUT(N__98272),
            .PADIN(N__98271),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D7_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam RST_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam RST_pad_iopad.PULLUP=1'b0;
    IO_PAD RST_pad_iopad (
            .OE(N__98264),
            .DIN(N__98263),
            .DOUT(N__98262),
            .PACKAGEPIN(RST));
    defparam RST_pad_preio.PIN_TYPE=6'b011001;
    defparam RST_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO RST_pad_preio (
            .PADOEN(N__98264),
            .PADOUT(N__98263),
            .PADIN(N__98262),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D12_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D12_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D12_pad_iopad (
            .OE(N__98255),
            .DIN(N__98254),
            .DOUT(N__98253),
            .PACKAGEPIN(FIFO_D12));
    defparam FIFO_D12_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D12_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D12_pad_preio (
            .PADOEN(N__98255),
            .PADOUT(N__98254),
            .PADIN(N__98253),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D12_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam UART_TX_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam UART_TX_pad_iopad.PULLUP=1'b0;
    IO_PAD UART_TX_pad_iopad (
            .OE(N__98246),
            .DIN(N__98245),
            .DOUT(N__98244),
            .PACKAGEPIN(UART_TX));
    defparam UART_TX_pad_preio.PIN_TYPE=6'b011001;
    defparam UART_TX_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO UART_TX_pad_preio (
            .PADOEN(N__98246),
            .PADOUT(N__98245),
            .PADIN(N__98244),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__77590),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_8_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_8_pad_iopad.PULLUP=1'b0;
    IO_PAD DEBUG_8_pad_iopad (
            .OE(N__98237),
            .DIN(N__98236),
            .DOUT(N__98235),
            .PACKAGEPIN(DEBUG_8));
    defparam DEBUG_8_pad_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_8_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_8_pad_preio (
            .PADOEN(N__98237),
            .PADOUT(N__98236),
            .PADIN(N__98235),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__43957),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA13_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA13_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA13_pad_iopad (
            .OE(N__98228),
            .DIN(N__98227),
            .DOUT(N__98226),
            .PACKAGEPIN(DATA13));
    defparam DATA13_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA13_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA13_pad_preio (
            .PADOEN(N__98228),
            .PADOUT(N__98227),
            .PADIN(N__98226),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__68481),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam UPDATE_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam UPDATE_pad_iopad.PULLUP=1'b0;
    IO_PAD UPDATE_pad_iopad (
            .OE(N__98219),
            .DIN(N__98218),
            .DOUT(N__98217),
            .PACKAGEPIN(UPDATE));
    defparam UPDATE_pad_preio.PIN_TYPE=6'b011001;
    defparam UPDATE_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO UPDATE_pad_preio (
            .PADOEN(N__98219),
            .PADOUT(N__98218),
            .PADIN(N__98217),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__81589),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ICE_CDONE_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ICE_CDONE_pad_iopad.PULLUP=1'b0;
    IO_PAD ICE_CDONE_pad_iopad (
            .OE(N__98210),
            .DIN(N__98209),
            .DOUT(N__98208),
            .PACKAGEPIN(ICE_CDONE));
    defparam ICE_CDONE_pad_preio.PIN_TYPE=6'b101001;
    defparam ICE_CDONE_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ICE_CDONE_pad_preio (
            .PADOEN(N__98210),
            .PADOUT(N__98209),
            .PADIN(N__98208),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D8_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D8_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D8_pad_iopad (
            .OE(N__98201),
            .DIN(N__98200),
            .DOUT(N__98199),
            .PACKAGEPIN(FIFO_D8));
    defparam FIFO_D8_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D8_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D8_pad_preio (
            .PADOEN(N__98201),
            .PADOUT(N__98200),
            .PADIN(N__98199),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D8_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_6_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_6_pad_iopad.PULLUP=1'b0;
    IO_PAD DEBUG_6_pad_iopad (
            .OE(N__98192),
            .DIN(N__98191),
            .DOUT(N__98190),
            .PACKAGEPIN(DEBUG_6));
    defparam DEBUG_6_pad_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_6_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_6_pad_preio (
            .PADOEN(N__98192),
            .PADOUT(N__98191),
            .PADIN(N__98190),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__83878),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_5_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_5_pad_iopad.PULLUP=1'b0;
    IO_PAD DEBUG_5_pad_iopad (
            .OE(N__98183),
            .DIN(N__98182),
            .DOUT(N__98181),
            .PACKAGEPIN(DEBUG_5));
    defparam DEBUG_5_pad_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_5_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_5_pad_preio (
            .PADOEN(N__98183),
            .PADOUT(N__98182),
            .PADIN(N__98181),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__57766),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_2_c_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_2_c_pad_iopad.PULLUP=1'b0;
    IO_PAD DEBUG_2_c_pad_iopad (
            .OE(N__98174),
            .DIN(N__98173),
            .DOUT(N__98172),
            .PACKAGEPIN(FR_RXF));
    defparam DEBUG_2_c_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_2_c_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_2_c_pad_preio (
            .PADOEN(N__98174),
            .PADOUT(N__98173),
            .PADIN(N__98172),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_2_c_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA5_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA5_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA5_pad_iopad (
            .OE(N__98165),
            .DIN(N__98164),
            .DOUT(N__98163),
            .PACKAGEPIN(DATA5));
    defparam DATA5_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA5_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA5_pad_preio (
            .PADOEN(N__98165),
            .PADOUT(N__98164),
            .PADIN(N__98163),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65362),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA15_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA15_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA15_pad_iopad (
            .OE(N__98156),
            .DIN(N__98155),
            .DOUT(N__98154),
            .PACKAGEPIN(DATA15));
    defparam DATA15_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA15_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA15_pad_preio (
            .PADOEN(N__98156),
            .PADOUT(N__98155),
            .PADIN(N__98154),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__57448),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA16_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA16_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA16_pad_iopad (
            .OE(N__98147),
            .DIN(N__98146),
            .DOUT(N__98145),
            .PACKAGEPIN(DATA16));
    defparam DATA16_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA16_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA16_pad_preio (
            .PADOEN(N__98147),
            .PADOUT(N__98146),
            .PADIN(N__98145),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__57303),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam CTS_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CTS_pad_iopad.PULLUP=1'b0;
    IO_PAD CTS_pad_iopad (
            .OE(N__98138),
            .DIN(N__98137),
            .DOUT(N__98136),
            .PACKAGEPIN(CTS));
    defparam CTS_pad_preio.PIN_TYPE=6'b011001;
    defparam CTS_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CTS_pad_preio (
            .PADOEN(N__98138),
            .PADOUT(N__98137),
            .PADIN(N__98136),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_1_c_0_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_1_c_0_pad_iopad.PULLUP=1'b0;
    IO_PAD DEBUG_1_c_0_pad_iopad (
            .OE(N__98129),
            .DIN(N__98128),
            .DOUT(N__98127),
            .PACKAGEPIN(FIFO_D0));
    defparam DEBUG_1_c_0_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_1_c_0_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_1_c_0_pad_preio (
            .PADOEN(N__98129),
            .PADOUT(N__98128),
            .PADIN(N__98127),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_1_c_0_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA19_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA19_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA19_pad_iopad (
            .OE(N__98120),
            .DIN(N__98119),
            .DOUT(N__98118),
            .PACKAGEPIN(DATA19));
    defparam DATA19_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA19_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA19_pad_preio (
            .PADOEN(N__98120),
            .PADOUT(N__98119),
            .PADIN(N__98118),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65515),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA14_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA14_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA14_pad_iopad (
            .OE(N__98111),
            .DIN(N__98110),
            .DOUT(N__98109),
            .PACKAGEPIN(DATA14));
    defparam DATA14_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA14_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA14_pad_preio (
            .PADOEN(N__98111),
            .PADOUT(N__98110),
            .PADIN(N__98109),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__68830),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D5_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D5_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D5_pad_iopad (
            .OE(N__98102),
            .DIN(N__98101),
            .DOUT(N__98100),
            .PACKAGEPIN(FIFO_D5));
    defparam FIFO_D5_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D5_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D5_pad_preio (
            .PADOEN(N__98102),
            .PADOUT(N__98101),
            .PADIN(N__98100),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D5_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ICE_SYSCLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ICE_SYSCLK_pad_iopad.PULLUP=1'b0;
    IO_PAD ICE_SYSCLK_pad_iopad (
            .OE(N__98093),
            .DIN(N__98092),
            .DOUT(N__98091),
            .PACKAGEPIN(ICE_SYSCLK));
    defparam ICE_SYSCLK_pad_preio.PIN_TYPE=6'b000001;
    defparam ICE_SYSCLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ICE_SYSCLK_pad_preio (
            .PADOEN(N__98093),
            .PADOUT(N__98092),
            .PADIN(N__98091),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ICE_SYSCLK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam SYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD SYNC_pad_iopad (
            .OE(N__98084),
            .DIN(N__98083),
            .DOUT(N__98082),
            .PACKAGEPIN(SYNC));
    defparam SYNC_pad_preio.PIN_TYPE=6'b010101;
    defparam SYNC_pad_preio.NEG_TRIGGER=1'b1;
    PRE_IO SYNC_pad_preio (
            .PADOEN(N__98084),
            .PADOUT(N__98083),
            .PADIN(N__98082),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__69106),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__97451));
    defparam DATA12_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA12_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA12_pad_iopad (
            .OE(N__98075),
            .DIN(N__98074),
            .DOUT(N__98073),
            .PACKAGEPIN(DATA12));
    defparam DATA12_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA12_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA12_pad_preio (
            .PADOEN(N__98075),
            .PADOUT(N__98074),
            .PADIN(N__98073),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__68406),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA11_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA11_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA11_pad_iopad (
            .OE(N__98066),
            .DIN(N__98065),
            .DOUT(N__98064),
            .PACKAGEPIN(DATA11));
    defparam DATA11_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA11_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA11_pad_preio (
            .PADOEN(N__98066),
            .PADOUT(N__98065),
            .PADIN(N__98064),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__58134),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ICE_CREST_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ICE_CREST_pad_iopad.PULLUP=1'b0;
    IO_PAD ICE_CREST_pad_iopad (
            .OE(N__98057),
            .DIN(N__98056),
            .DOUT(N__98055),
            .PACKAGEPIN(ICE_CREST));
    defparam ICE_CREST_pad_preio.PIN_TYPE=6'b101001;
    defparam ICE_CREST_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ICE_CREST_pad_preio (
            .PADOEN(N__98057),
            .PADOUT(N__98056),
            .PADIN(N__98055),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ICE_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ICE_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD ICE_CLK_pad_iopad (
            .OE(N__98048),
            .DIN(N__98047),
            .DOUT(N__98046),
            .PACKAGEPIN(ICE_CLK));
    defparam ICE_CLK_pad_preio.PIN_TYPE=6'b101001;
    defparam ICE_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ICE_CLK_pad_preio (
            .PADOEN(N__98048),
            .PADOUT(N__98047),
            .PADIN(N__98046),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VALID_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam VALID_pad_iopad.PULLUP=1'b0;
    IO_PAD VALID_pad_iopad (
            .OE(N__98039),
            .DIN(N__98038),
            .DOUT(N__98037),
            .PACKAGEPIN(VALID));
    defparam VALID_pad_preio.PIN_TYPE=6'b010101;
    defparam VALID_pad_preio.NEG_TRIGGER=1'b1;
    PRE_IO VALID_pad_preio (
            .PADOEN(N__98039),
            .PADOUT(N__98038),
            .PADIN(N__98037),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__57415),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__97448));
    defparam FT_SIWU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FT_SIWU_pad_iopad.PULLUP=1'b0;
    IO_PAD FT_SIWU_pad_iopad (
            .OE(N__98030),
            .DIN(N__98029),
            .DOUT(N__98028),
            .PACKAGEPIN(FT_SIWU));
    defparam FT_SIWU_pad_preio.PIN_TYPE=6'b011001;
    defparam FT_SIWU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FT_SIWU_pad_preio (
            .PADOEN(N__98030),
            .PADOUT(N__98029),
            .PADIN(N__98028),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__86664),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA21_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA21_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA21_pad_iopad (
            .OE(N__98021),
            .DIN(N__98020),
            .DOUT(N__98019),
            .PACKAGEPIN(DATA21));
    defparam DATA21_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA21_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA21_pad_preio (
            .PADOEN(N__98021),
            .PADOUT(N__98020),
            .PADIN(N__98019),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65358),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA22_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA22_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA22_pad_iopad (
            .OE(N__98012),
            .DIN(N__98011),
            .DOUT(N__98010),
            .PACKAGEPIN(DATA22));
    defparam DATA22_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA22_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA22_pad_preio (
            .PADOEN(N__98012),
            .PADOUT(N__98011),
            .PADIN(N__98010),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65317),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA26_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA26_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA26_pad_iopad (
            .OE(N__98003),
            .DIN(N__98002),
            .DOUT(N__98001),
            .PACKAGEPIN(DATA26));
    defparam DATA26_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA26_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA26_pad_preio (
            .PADOEN(N__98003),
            .PADOUT(N__98002),
            .PADIN(N__98001),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__58083),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam INVERT_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INVERT_pad_iopad.PULLUP=1'b0;
    IO_PAD INVERT_pad_iopad (
            .OE(N__97994),
            .DIN(N__97993),
            .DOUT(N__97992),
            .PACKAGEPIN(INVERT));
    defparam INVERT_pad_preio.PIN_TYPE=6'b010101;
    defparam INVERT_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INVERT_pad_preio (
            .PADOEN(N__97994),
            .PADOUT(N__97993),
            .PADIN(N__97992),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__73072),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__97450));
    defparam DATA28_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA28_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA28_pad_iopad (
            .OE(N__97985),
            .DIN(N__97984),
            .DOUT(N__97983),
            .PACKAGEPIN(DATA28));
    defparam DATA28_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA28_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA28_pad_preio (
            .PADOEN(N__97985),
            .PADOUT(N__97984),
            .PADIN(N__97983),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__68422),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SLM_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam SLM_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD SLM_CLK_pad_iopad (
            .OE(N__97976),
            .DIN(N__97975),
            .DOUT(N__97974),
            .PACKAGEPIN(SLM_CLK));
    defparam SLM_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam SLM_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO SLM_CLK_pad_preio (
            .PADOEN(N__97976),
            .PADOUT(N__97975),
            .PADIN(N__97974),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__83863),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam UART_RX_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam UART_RX_pad_iopad.PULLUP=1'b0;
    IO_PAD UART_RX_pad_iopad (
            .OE(N__97967),
            .DIN(N__97966),
            .DOUT(N__97965),
            .PACKAGEPIN(UART_RX));
    defparam UART_RX_pad_preio.PIN_TYPE=6'b000000;
    defparam UART_RX_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO UART_RX_pad_preio (
            .PADOEN(N__97967),
            .PADOUT(N__97966),
            .PADIN(N__97965),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(\pc_rx.r_Rx_Data_R ),
            .DOUT0(),
            .INPUTCLK(N__97452),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA9_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA9_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA9_pad_iopad (
            .OE(N__97958),
            .DIN(N__97957),
            .DOUT(N__97956),
            .PACKAGEPIN(DATA9));
    defparam DATA9_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA9_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA9_pad_preio (
            .PADOEN(N__97958),
            .PADOUT(N__97957),
            .PADIN(N__97956),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__58060),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA27_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA27_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA27_pad_iopad (
            .OE(N__97949),
            .DIN(N__97948),
            .DOUT(N__97947),
            .PACKAGEPIN(DATA27));
    defparam DATA27_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA27_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA27_pad_preio (
            .PADOEN(N__97949),
            .PADOUT(N__97948),
            .PADIN(N__97947),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__58135),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_0_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_0_pad_iopad.PULLUP=1'b0;
    IO_PAD DEBUG_0_pad_iopad (
            .OE(N__97940),
            .DIN(N__97939),
            .DOUT(N__97938),
            .PACKAGEPIN(DEBUG_0));
    defparam DEBUG_0_pad_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_0_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_0_pad_preio (
            .PADOEN(N__97940),
            .PADOUT(N__97939),
            .PADIN(N__97938),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__82609),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA2_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA2_pad_iopad (
            .OE(N__97931),
            .DIN(N__97930),
            .DOUT(N__97929),
            .PACKAGEPIN(DATA2));
    defparam DATA2_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA2_pad_preio (
            .PADOEN(N__97931),
            .PADOUT(N__97930),
            .PADIN(N__97929),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65457),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D4_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D4_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D4_pad_iopad (
            .OE(N__97922),
            .DIN(N__97921),
            .DOUT(N__97920),
            .PACKAGEPIN(FIFO_D4));
    defparam FIFO_D4_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D4_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D4_pad_preio (
            .PADOEN(N__97922),
            .PADOUT(N__97921),
            .PADIN(N__97920),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D4_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA18_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA18_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA18_pad_iopad (
            .OE(N__97913),
            .DIN(N__97912),
            .DOUT(N__97911),
            .PACKAGEPIN(DATA18));
    defparam DATA18_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA18_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA18_pad_preio (
            .PADOEN(N__97913),
            .PADOUT(N__97912),
            .PADIN(N__97911),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65464),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam RESET_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam RESET_pad_iopad.PULLUP=1'b0;
    IO_PAD RESET_pad_iopad (
            .OE(N__97904),
            .DIN(N__97903),
            .DOUT(N__97902),
            .PACKAGEPIN(RESET));
    defparam RESET_pad_preio.PIN_TYPE=6'b011001;
    defparam RESET_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO RESET_pad_preio (
            .PADOEN(N__97904),
            .PADOUT(N__97903),
            .PADIN(N__97902),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__69961),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D1_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D1_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D1_pad_iopad (
            .OE(N__97895),
            .DIN(N__97894),
            .DOUT(N__97893),
            .PACKAGEPIN(FIFO_D1));
    defparam FIFO_D1_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D1_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D1_pad_preio (
            .PADOEN(N__97895),
            .PADOUT(N__97894),
            .PADIN(N__97893),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D1_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SDAT_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam SDAT_pad_iopad.PULLUP=1'b0;
    IO_PAD SDAT_pad_iopad (
            .OE(N__97886),
            .DIN(N__97885),
            .DOUT(N__97884),
            .PACKAGEPIN(SDAT));
    defparam SDAT_pad_preio.PIN_TYPE=6'b010101;
    defparam SDAT_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO SDAT_pad_preio (
            .PADOEN(N__97886),
            .PADOUT(N__97885),
            .PADIN(N__97884),
            .CLOCKENABLE(N__58000),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__57856),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__97355));
    defparam DATA10_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA10_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA10_pad_iopad (
            .OE(N__97877),
            .DIN(N__97876),
            .DOUT(N__97875),
            .PACKAGEPIN(DATA10));
    defparam DATA10_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA10_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA10_pad_preio (
            .PADOEN(N__97877),
            .PADOUT(N__97876),
            .PADIN(N__97875),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__58084),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA6_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA6_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA6_pad_iopad (
            .OE(N__97868),
            .DIN(N__97867),
            .DOUT(N__97866),
            .PACKAGEPIN(DATA6));
    defparam DATA6_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA6_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA6_pad_preio (
            .PADOEN(N__97868),
            .PADOUT(N__97867),
            .PADIN(N__97866),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65313),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SEN_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam SEN_pad_iopad.PULLUP=1'b0;
    IO_PAD SEN_pad_iopad (
            .OE(N__97859),
            .DIN(N__97858),
            .DOUT(N__97857),
            .PACKAGEPIN(SEN));
    defparam SEN_pad_preio.PIN_TYPE=6'b010101;
    defparam SEN_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO SEN_pad_preio (
            .PADOEN(N__97859),
            .PADOUT(N__97858),
            .PADIN(N__97857),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__53047),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__97361));
    defparam DCD_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DCD_pad_iopad.PULLUP=1'b0;
    IO_PAD DCD_pad_iopad (
            .OE(N__97850),
            .DIN(N__97849),
            .DOUT(N__97848),
            .PACKAGEPIN(DCD));
    defparam DCD_pad_preio.PIN_TYPE=6'b011001;
    defparam DCD_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DCD_pad_preio (
            .PADOEN(N__97850),
            .PADOUT(N__97849),
            .PADIN(N__97848),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D14_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D14_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D14_pad_iopad (
            .OE(N__97841),
            .DIN(N__97840),
            .DOUT(N__97839),
            .PACKAGEPIN(FIFO_D14));
    defparam FIFO_D14_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D14_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D14_pad_preio (
            .PADOEN(N__97841),
            .PADOUT(N__97840),
            .PADIN(N__97839),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D14_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA30_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA30_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA30_pad_iopad (
            .OE(N__97832),
            .DIN(N__97831),
            .DOUT(N__97830),
            .PACKAGEPIN(DATA30));
    defparam DATA30_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA30_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA30_pad_preio (
            .PADOEN(N__97832),
            .PADOUT(N__97831),
            .PADIN(N__97830),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__68829),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_9_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_9_pad_iopad.PULLUP=1'b0;
    IO_PAD DEBUG_9_pad_iopad (
            .OE(N__97823),
            .DIN(N__97822),
            .DOUT(N__97821),
            .PACKAGEPIN(DEBUG_9));
    defparam DEBUG_9_pad_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_9_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_9_pad_preio (
            .PADOEN(N__97823),
            .PADOUT(N__97822),
            .PADIN(N__97821),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__64375),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA24_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA24_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA24_pad_iopad (
            .OE(N__97814),
            .DIN(N__97813),
            .DOUT(N__97812),
            .PACKAGEPIN(DATA24));
    defparam DATA24_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA24_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA24_pad_preio (
            .PADOEN(N__97814),
            .PADOUT(N__97813),
            .PADIN(N__97812),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65073),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DTR_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DTR_pad_iopad.PULLUP=1'b0;
    IO_PAD DTR_pad_iopad (
            .OE(N__97805),
            .DIN(N__97804),
            .DOUT(N__97803),
            .PACKAGEPIN(DTR));
    defparam DTR_pad_preio.PIN_TYPE=6'b011001;
    defparam DTR_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DTR_pad_preio (
            .PADOEN(N__97805),
            .PADOUT(N__97804),
            .PADIN(N__97803),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA29_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA29_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA29_pad_iopad (
            .OE(N__97796),
            .DIN(N__97795),
            .DOUT(N__97794),
            .PACKAGEPIN(DATA29));
    defparam DATA29_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA29_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA29_pad_preio (
            .PADOEN(N__97796),
            .PADOUT(N__97795),
            .PADIN(N__97794),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__68485),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DSR_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DSR_pad_iopad.PULLUP=1'b0;
    IO_PAD DSR_pad_iopad (
            .OE(N__97787),
            .DIN(N__97786),
            .DOUT(N__97785),
            .PACKAGEPIN(DSR));
    defparam DSR_pad_preio.PIN_TYPE=6'b011001;
    defparam DSR_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DSR_pad_preio (
            .PADOEN(N__97787),
            .PADOUT(N__97786),
            .PADIN(N__97785),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FT_WR_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FT_WR_pad_iopad.PULLUP=1'b0;
    IO_PAD FT_WR_pad_iopad (
            .OE(N__97778),
            .DIN(N__97777),
            .DOUT(N__97776),
            .PACKAGEPIN(FT_WR));
    defparam FT_WR_pad_preio.PIN_TYPE=6'b011001;
    defparam FT_WR_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FT_WR_pad_preio (
            .PADOEN(N__97778),
            .PADOUT(N__97777),
            .PADIN(N__97776),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__86668),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FT_RD_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FT_RD_pad_iopad.PULLUP=1'b0;
    IO_PAD FT_RD_pad_iopad (
            .OE(N__97769),
            .DIN(N__97768),
            .DOUT(N__97767),
            .PACKAGEPIN(FT_RD));
    defparam FT_RD_pad_preio.PIN_TYPE=6'b011001;
    defparam FT_RD_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FT_RD_pad_preio (
            .PADOEN(N__97769),
            .PADOUT(N__97768),
            .PADIN(N__97767),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__44013),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA31_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA31_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA31_pad_iopad (
            .OE(N__97760),
            .DIN(N__97759),
            .DOUT(N__97758),
            .PACKAGEPIN(DATA31));
    defparam DATA31_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA31_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA31_pad_preio (
            .PADOEN(N__97760),
            .PADOUT(N__97759),
            .PADIN(N__97758),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__57444),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA8_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA8_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA8_pad_iopad (
            .OE(N__97751),
            .DIN(N__97750),
            .DOUT(N__97749),
            .PACKAGEPIN(DATA8));
    defparam DATA8_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA8_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA8_pad_preio (
            .PADOEN(N__97751),
            .PADOUT(N__97750),
            .PADIN(N__97749),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65077),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D6_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D6_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D6_pad_iopad (
            .OE(N__97742),
            .DIN(N__97741),
            .DOUT(N__97740),
            .PACKAGEPIN(FIFO_D6));
    defparam FIFO_D6_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D6_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D6_pad_preio (
            .PADOEN(N__97742),
            .PADOUT(N__97741),
            .PADIN(N__97740),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D6_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D11_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D11_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D11_pad_iopad (
            .OE(N__97733),
            .DIN(N__97732),
            .DOUT(N__97731),
            .PACKAGEPIN(FIFO_D11));
    defparam FIFO_D11_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D11_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D11_pad_preio (
            .PADOEN(N__97733),
            .PADOUT(N__97732),
            .PADIN(N__97731),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D11_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D2_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D2_pad_iopad (
            .OE(N__97724),
            .DIN(N__97723),
            .DOUT(N__97722),
            .PACKAGEPIN(FIFO_D2));
    defparam FIFO_D2_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D2_pad_preio (
            .PADOEN(N__97724),
            .PADOUT(N__97723),
            .PADIN(N__97722),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D2_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D15_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D15_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D15_pad_iopad (
            .OE(N__97715),
            .DIN(N__97714),
            .DOUT(N__97713),
            .PACKAGEPIN(FIFO_D15));
    defparam FIFO_D15_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D15_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D15_pad_preio (
            .PADOEN(N__97715),
            .PADOUT(N__97714),
            .PADIN(N__97713),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D15_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_2_pad_iopad.PULLUP=1'b0;
    IO_PAD DEBUG_2_pad_iopad (
            .OE(N__97706),
            .DIN(N__97705),
            .DOUT(N__97704),
            .PACKAGEPIN(DEBUG_2));
    defparam DEBUG_2_pad_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_2_pad_preio (
            .PADOEN(N__97706),
            .PADOUT(N__97705),
            .PADIN(N__97704),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__57649),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA23_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA23_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA23_pad_iopad (
            .OE(N__97697),
            .DIN(N__97696),
            .DOUT(N__97695),
            .PACKAGEPIN(DATA23));
    defparam DATA23_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA23_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA23_pad_preio (
            .PADOEN(N__97697),
            .PADOUT(N__97696),
            .PADIN(N__97695),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65019),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA0_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA0_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA0_pad_iopad (
            .OE(N__97688),
            .DIN(N__97687),
            .DOUT(N__97686),
            .PACKAGEPIN(DATA0));
    defparam DATA0_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA0_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA0_pad_preio (
            .PADOEN(N__97688),
            .PADOUT(N__97687),
            .PADIN(N__97686),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__57304),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SCK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam SCK_pad_iopad.PULLUP=1'b0;
    IO_PAD SCK_pad_iopad (
            .OE(N__97679),
            .DIN(N__97678),
            .DOUT(N__97677),
            .PACKAGEPIN(SCK));
    defparam SCK_pad_preio.PIN_TYPE=6'b010101;
    defparam SCK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO SCK_pad_preio (
            .PADOEN(N__97679),
            .PADOUT(N__97678),
            .PADIN(N__97677),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__51160),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__97350));
    defparam DATA3_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA3_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA3_pad_iopad (
            .OE(N__97670),
            .DIN(N__97669),
            .DOUT(N__97668),
            .PACKAGEPIN(DATA3));
    defparam DATA3_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA3_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA3_pad_preio (
            .PADOEN(N__97670),
            .PADOUT(N__97669),
            .PADIN(N__97668),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65508),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA25_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA25_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA25_pad_iopad (
            .OE(N__97661),
            .DIN(N__97660),
            .DOUT(N__97659),
            .PACKAGEPIN(DATA25));
    defparam DATA25_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA25_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA25_pad_preio (
            .PADOEN(N__97661),
            .PADOUT(N__97660),
            .PADIN(N__97659),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__58056),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SOUT_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam SOUT_pad_iopad.PULLUP=1'b0;
    IO_PAD SOUT_pad_iopad (
            .OE(N__97652),
            .DIN(N__97651),
            .DOUT(N__97650),
            .PACKAGEPIN(SOUT));
    defparam SOUT_pad_preio.PIN_TYPE=6'b000000;
    defparam SOUT_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO SOUT_pad_preio (
            .PADOEN(N__97652),
            .PADOUT(N__97651),
            .PADIN(N__97650),
            .CLOCKENABLE(N__65230),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(rx_shift_reg_0),
            .DOUT0(),
            .INPUTCLK(N__97369),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA1_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA1_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA1_pad_iopad (
            .OE(N__97643),
            .DIN(N__97642),
            .DOUT(N__97641),
            .PACKAGEPIN(DATA1));
    defparam DATA1_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA1_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA1_pad_preio (
            .PADOEN(N__97643),
            .PADOUT(N__97642),
            .PADIN(N__97641),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65412),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FT_OE_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FT_OE_pad_iopad.PULLUP=1'b0;
    IO_PAD FT_OE_pad_iopad (
            .OE(N__97634),
            .DIN(N__97633),
            .DOUT(N__97632),
            .PACKAGEPIN(FT_OE));
    defparam FT_OE_pad_preio.PIN_TYPE=6'b011001;
    defparam FT_OE_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FT_OE_pad_preio (
            .PADOEN(N__97634),
            .PADOUT(N__97633),
            .PADIN(N__97632),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__43897),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D3_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D3_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D3_pad_iopad (
            .OE(N__97625),
            .DIN(N__97624),
            .DOUT(N__97623),
            .PACKAGEPIN(FIFO_D3));
    defparam FIFO_D3_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D3_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D3_pad_preio (
            .PADOEN(N__97625),
            .PADOUT(N__97624),
            .PADIN(N__97623),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D3_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam FIFO_D9_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam FIFO_D9_pad_iopad.PULLUP=1'b0;
    IO_PAD FIFO_D9_pad_iopad (
            .OE(N__97616),
            .DIN(N__97615),
            .DOUT(N__97614),
            .PACKAGEPIN(FIFO_D9));
    defparam FIFO_D9_pad_preio.PIN_TYPE=6'b000001;
    defparam FIFO_D9_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO FIFO_D9_pad_preio (
            .PADOEN(N__97616),
            .PADOUT(N__97615),
            .PADIN(N__97614),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(FIFO_D9_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DATA7_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DATA7_pad_iopad.PULLUP=1'b0;
    IO_PAD DATA7_pad_iopad (
            .OE(N__97607),
            .DIN(N__97606),
            .DOUT(N__97605),
            .PACKAGEPIN(DATA7));
    defparam DATA7_pad_preio.PIN_TYPE=6'b011001;
    defparam DATA7_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DATA7_pad_preio (
            .PADOEN(N__97607),
            .PADOUT(N__97606),
            .PADIN(N__97605),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__65026),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_1_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_1_pad_iopad.PULLUP=1'b0;
    IO_PAD DEBUG_1_pad_iopad (
            .OE(N__97598),
            .DIN(N__97597),
            .DOUT(N__97596),
            .PACKAGEPIN(DEBUG_1));
    defparam DEBUG_1_pad_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_1_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_1_pad_preio (
            .PADOEN(N__97598),
            .PADOUT(N__97597),
            .PADIN(N__97596),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__44916),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__24326 (
            .O(N__97579),
            .I(N__97575));
    InMux I__24325 (
            .O(N__97578),
            .I(N__97572));
    LocalMux I__24324 (
            .O(N__97575),
            .I(\pc_tx.r_Clock_Count_2 ));
    LocalMux I__24323 (
            .O(N__97572),
            .I(\pc_tx.r_Clock_Count_2 ));
    InMux I__24322 (
            .O(N__97567),
            .I(\pc_tx.n10713 ));
    InMux I__24321 (
            .O(N__97564),
            .I(N__97560));
    InMux I__24320 (
            .O(N__97563),
            .I(N__97557));
    LocalMux I__24319 (
            .O(N__97560),
            .I(\pc_tx.r_Clock_Count_3 ));
    LocalMux I__24318 (
            .O(N__97557),
            .I(\pc_tx.r_Clock_Count_3 ));
    InMux I__24317 (
            .O(N__97552),
            .I(\pc_tx.n10714 ));
    InMux I__24316 (
            .O(N__97549),
            .I(N__97545));
    InMux I__24315 (
            .O(N__97548),
            .I(N__97542));
    LocalMux I__24314 (
            .O(N__97545),
            .I(\pc_tx.r_Clock_Count_4 ));
    LocalMux I__24313 (
            .O(N__97542),
            .I(\pc_tx.r_Clock_Count_4 ));
    InMux I__24312 (
            .O(N__97537),
            .I(\pc_tx.n10715 ));
    CascadeMux I__24311 (
            .O(N__97534),
            .I(N__97531));
    InMux I__24310 (
            .O(N__97531),
            .I(N__97527));
    InMux I__24309 (
            .O(N__97530),
            .I(N__97524));
    LocalMux I__24308 (
            .O(N__97527),
            .I(\pc_tx.r_Clock_Count_5 ));
    LocalMux I__24307 (
            .O(N__97524),
            .I(\pc_tx.r_Clock_Count_5 ));
    InMux I__24306 (
            .O(N__97519),
            .I(\pc_tx.n10716 ));
    InMux I__24305 (
            .O(N__97516),
            .I(N__97512));
    InMux I__24304 (
            .O(N__97515),
            .I(N__97509));
    LocalMux I__24303 (
            .O(N__97512),
            .I(\pc_tx.r_Clock_Count_6 ));
    LocalMux I__24302 (
            .O(N__97509),
            .I(\pc_tx.r_Clock_Count_6 ));
    InMux I__24301 (
            .O(N__97504),
            .I(\pc_tx.n10717 ));
    InMux I__24300 (
            .O(N__97501),
            .I(N__97497));
    InMux I__24299 (
            .O(N__97500),
            .I(N__97494));
    LocalMux I__24298 (
            .O(N__97497),
            .I(\pc_tx.r_Clock_Count_7 ));
    LocalMux I__24297 (
            .O(N__97494),
            .I(\pc_tx.r_Clock_Count_7 ));
    InMux I__24296 (
            .O(N__97489),
            .I(\pc_tx.n10718 ));
    InMux I__24295 (
            .O(N__97486),
            .I(N__97482));
    InMux I__24294 (
            .O(N__97485),
            .I(N__97479));
    LocalMux I__24293 (
            .O(N__97482),
            .I(\pc_tx.r_Clock_Count_8 ));
    LocalMux I__24292 (
            .O(N__97479),
            .I(\pc_tx.r_Clock_Count_8 ));
    InMux I__24291 (
            .O(N__97474),
            .I(bfn_24_12_0_));
    InMux I__24290 (
            .O(N__97471),
            .I(\pc_tx.n10720 ));
    InMux I__24289 (
            .O(N__97468),
            .I(N__97464));
    InMux I__24288 (
            .O(N__97467),
            .I(N__97461));
    LocalMux I__24287 (
            .O(N__97464),
            .I(\pc_tx.r_Clock_Count_9 ));
    LocalMux I__24286 (
            .O(N__97461),
            .I(\pc_tx.r_Clock_Count_9 ));
    InMux I__24285 (
            .O(N__97456),
            .I(N__97453));
    LocalMux I__24284 (
            .O(N__97453),
            .I(N__97414));
    ClkMux I__24283 (
            .O(N__97452),
            .I(N__97123));
    ClkMux I__24282 (
            .O(N__97451),
            .I(N__97123));
    ClkMux I__24281 (
            .O(N__97450),
            .I(N__97123));
    ClkMux I__24280 (
            .O(N__97449),
            .I(N__97123));
    ClkMux I__24279 (
            .O(N__97448),
            .I(N__97123));
    ClkMux I__24278 (
            .O(N__97447),
            .I(N__97123));
    ClkMux I__24277 (
            .O(N__97446),
            .I(N__97123));
    ClkMux I__24276 (
            .O(N__97445),
            .I(N__97123));
    ClkMux I__24275 (
            .O(N__97444),
            .I(N__97123));
    ClkMux I__24274 (
            .O(N__97443),
            .I(N__97123));
    ClkMux I__24273 (
            .O(N__97442),
            .I(N__97123));
    ClkMux I__24272 (
            .O(N__97441),
            .I(N__97123));
    ClkMux I__24271 (
            .O(N__97440),
            .I(N__97123));
    ClkMux I__24270 (
            .O(N__97439),
            .I(N__97123));
    ClkMux I__24269 (
            .O(N__97438),
            .I(N__97123));
    ClkMux I__24268 (
            .O(N__97437),
            .I(N__97123));
    ClkMux I__24267 (
            .O(N__97436),
            .I(N__97123));
    ClkMux I__24266 (
            .O(N__97435),
            .I(N__97123));
    ClkMux I__24265 (
            .O(N__97434),
            .I(N__97123));
    ClkMux I__24264 (
            .O(N__97433),
            .I(N__97123));
    ClkMux I__24263 (
            .O(N__97432),
            .I(N__97123));
    ClkMux I__24262 (
            .O(N__97431),
            .I(N__97123));
    ClkMux I__24261 (
            .O(N__97430),
            .I(N__97123));
    ClkMux I__24260 (
            .O(N__97429),
            .I(N__97123));
    ClkMux I__24259 (
            .O(N__97428),
            .I(N__97123));
    ClkMux I__24258 (
            .O(N__97427),
            .I(N__97123));
    ClkMux I__24257 (
            .O(N__97426),
            .I(N__97123));
    ClkMux I__24256 (
            .O(N__97425),
            .I(N__97123));
    ClkMux I__24255 (
            .O(N__97424),
            .I(N__97123));
    ClkMux I__24254 (
            .O(N__97423),
            .I(N__97123));
    ClkMux I__24253 (
            .O(N__97422),
            .I(N__97123));
    ClkMux I__24252 (
            .O(N__97421),
            .I(N__97123));
    ClkMux I__24251 (
            .O(N__97420),
            .I(N__97123));
    ClkMux I__24250 (
            .O(N__97419),
            .I(N__97123));
    ClkMux I__24249 (
            .O(N__97418),
            .I(N__97123));
    ClkMux I__24248 (
            .O(N__97417),
            .I(N__97123));
    Glb2LocalMux I__24247 (
            .O(N__97414),
            .I(N__97123));
    ClkMux I__24246 (
            .O(N__97413),
            .I(N__97123));
    ClkMux I__24245 (
            .O(N__97412),
            .I(N__97123));
    ClkMux I__24244 (
            .O(N__97411),
            .I(N__97123));
    ClkMux I__24243 (
            .O(N__97410),
            .I(N__97123));
    ClkMux I__24242 (
            .O(N__97409),
            .I(N__97123));
    ClkMux I__24241 (
            .O(N__97408),
            .I(N__97123));
    ClkMux I__24240 (
            .O(N__97407),
            .I(N__97123));
    ClkMux I__24239 (
            .O(N__97406),
            .I(N__97123));
    ClkMux I__24238 (
            .O(N__97405),
            .I(N__97123));
    ClkMux I__24237 (
            .O(N__97404),
            .I(N__97123));
    ClkMux I__24236 (
            .O(N__97403),
            .I(N__97123));
    ClkMux I__24235 (
            .O(N__97402),
            .I(N__97123));
    ClkMux I__24234 (
            .O(N__97401),
            .I(N__97123));
    ClkMux I__24233 (
            .O(N__97400),
            .I(N__97123));
    ClkMux I__24232 (
            .O(N__97399),
            .I(N__97123));
    ClkMux I__24231 (
            .O(N__97398),
            .I(N__97123));
    ClkMux I__24230 (
            .O(N__97397),
            .I(N__97123));
    ClkMux I__24229 (
            .O(N__97396),
            .I(N__97123));
    ClkMux I__24228 (
            .O(N__97395),
            .I(N__97123));
    ClkMux I__24227 (
            .O(N__97394),
            .I(N__97123));
    ClkMux I__24226 (
            .O(N__97393),
            .I(N__97123));
    ClkMux I__24225 (
            .O(N__97392),
            .I(N__97123));
    ClkMux I__24224 (
            .O(N__97391),
            .I(N__97123));
    ClkMux I__24223 (
            .O(N__97390),
            .I(N__97123));
    ClkMux I__24222 (
            .O(N__97389),
            .I(N__97123));
    ClkMux I__24221 (
            .O(N__97388),
            .I(N__97123));
    ClkMux I__24220 (
            .O(N__97387),
            .I(N__97123));
    ClkMux I__24219 (
            .O(N__97386),
            .I(N__97123));
    ClkMux I__24218 (
            .O(N__97385),
            .I(N__97123));
    ClkMux I__24217 (
            .O(N__97384),
            .I(N__97123));
    ClkMux I__24216 (
            .O(N__97383),
            .I(N__97123));
    ClkMux I__24215 (
            .O(N__97382),
            .I(N__97123));
    ClkMux I__24214 (
            .O(N__97381),
            .I(N__97123));
    ClkMux I__24213 (
            .O(N__97380),
            .I(N__97123));
    ClkMux I__24212 (
            .O(N__97379),
            .I(N__97123));
    ClkMux I__24211 (
            .O(N__97378),
            .I(N__97123));
    ClkMux I__24210 (
            .O(N__97377),
            .I(N__97123));
    ClkMux I__24209 (
            .O(N__97376),
            .I(N__97123));
    ClkMux I__24208 (
            .O(N__97375),
            .I(N__97123));
    ClkMux I__24207 (
            .O(N__97374),
            .I(N__97123));
    ClkMux I__24206 (
            .O(N__97373),
            .I(N__97123));
    ClkMux I__24205 (
            .O(N__97372),
            .I(N__97123));
    ClkMux I__24204 (
            .O(N__97371),
            .I(N__97123));
    ClkMux I__24203 (
            .O(N__97370),
            .I(N__97123));
    ClkMux I__24202 (
            .O(N__97369),
            .I(N__97123));
    ClkMux I__24201 (
            .O(N__97368),
            .I(N__97123));
    ClkMux I__24200 (
            .O(N__97367),
            .I(N__97123));
    ClkMux I__24199 (
            .O(N__97366),
            .I(N__97123));
    ClkMux I__24198 (
            .O(N__97365),
            .I(N__97123));
    ClkMux I__24197 (
            .O(N__97364),
            .I(N__97123));
    ClkMux I__24196 (
            .O(N__97363),
            .I(N__97123));
    ClkMux I__24195 (
            .O(N__97362),
            .I(N__97123));
    ClkMux I__24194 (
            .O(N__97361),
            .I(N__97123));
    ClkMux I__24193 (
            .O(N__97360),
            .I(N__97123));
    ClkMux I__24192 (
            .O(N__97359),
            .I(N__97123));
    ClkMux I__24191 (
            .O(N__97358),
            .I(N__97123));
    ClkMux I__24190 (
            .O(N__97357),
            .I(N__97123));
    ClkMux I__24189 (
            .O(N__97356),
            .I(N__97123));
    ClkMux I__24188 (
            .O(N__97355),
            .I(N__97123));
    ClkMux I__24187 (
            .O(N__97354),
            .I(N__97123));
    ClkMux I__24186 (
            .O(N__97353),
            .I(N__97123));
    ClkMux I__24185 (
            .O(N__97352),
            .I(N__97123));
    ClkMux I__24184 (
            .O(N__97351),
            .I(N__97123));
    ClkMux I__24183 (
            .O(N__97350),
            .I(N__97123));
    ClkMux I__24182 (
            .O(N__97349),
            .I(N__97123));
    ClkMux I__24181 (
            .O(N__97348),
            .I(N__97123));
    ClkMux I__24180 (
            .O(N__97347),
            .I(N__97123));
    ClkMux I__24179 (
            .O(N__97346),
            .I(N__97123));
    ClkMux I__24178 (
            .O(N__97345),
            .I(N__97123));
    ClkMux I__24177 (
            .O(N__97344),
            .I(N__97123));
    ClkMux I__24176 (
            .O(N__97343),
            .I(N__97123));
    ClkMux I__24175 (
            .O(N__97342),
            .I(N__97123));
    GlobalMux I__24174 (
            .O(N__97123),
            .I(N__97120));
    gio2CtrlBuf I__24173 (
            .O(N__97120),
            .I(SLM_CLK_c));
    CEMux I__24172 (
            .O(N__97117),
            .I(N__97114));
    LocalMux I__24171 (
            .O(N__97114),
            .I(N__97111));
    Span4Mux_v I__24170 (
            .O(N__97111),
            .I(N__97107));
    CEMux I__24169 (
            .O(N__97110),
            .I(N__97104));
    Span4Mux_h I__24168 (
            .O(N__97107),
            .I(N__97099));
    LocalMux I__24167 (
            .O(N__97104),
            .I(N__97099));
    Span4Mux_v I__24166 (
            .O(N__97099),
            .I(N__97095));
    CEMux I__24165 (
            .O(N__97098),
            .I(N__97092));
    Span4Mux_v I__24164 (
            .O(N__97095),
            .I(N__97087));
    LocalMux I__24163 (
            .O(N__97092),
            .I(N__97087));
    Odrv4 I__24162 (
            .O(N__97087),
            .I(\pc_tx.n1 ));
    SRMux I__24161 (
            .O(N__97084),
            .I(N__97081));
    LocalMux I__24160 (
            .O(N__97081),
            .I(N__97078));
    Span4Mux_v I__24159 (
            .O(N__97078),
            .I(N__97074));
    SRMux I__24158 (
            .O(N__97077),
            .I(N__97071));
    Span4Mux_s3_h I__24157 (
            .O(N__97074),
            .I(N__97066));
    LocalMux I__24156 (
            .O(N__97071),
            .I(N__97066));
    Sp12to4 I__24155 (
            .O(N__97066),
            .I(N__97063));
    Odrv12 I__24154 (
            .O(N__97063),
            .I(\pc_tx.n4577 ));
    CascadeMux I__24153 (
            .O(N__97060),
            .I(N__97056));
    InMux I__24152 (
            .O(N__97059),
            .I(N__97050));
    InMux I__24151 (
            .O(N__97056),
            .I(N__97042));
    InMux I__24150 (
            .O(N__97055),
            .I(N__97031));
    InMux I__24149 (
            .O(N__97054),
            .I(N__97026));
    InMux I__24148 (
            .O(N__97053),
            .I(N__97026));
    LocalMux I__24147 (
            .O(N__97050),
            .I(N__97018));
    InMux I__24146 (
            .O(N__97049),
            .I(N__97013));
    InMux I__24145 (
            .O(N__97048),
            .I(N__97013));
    InMux I__24144 (
            .O(N__97047),
            .I(N__97010));
    InMux I__24143 (
            .O(N__97046),
            .I(N__97005));
    InMux I__24142 (
            .O(N__97045),
            .I(N__97005));
    LocalMux I__24141 (
            .O(N__97042),
            .I(N__97002));
    InMux I__24140 (
            .O(N__97041),
            .I(N__96991));
    InMux I__24139 (
            .O(N__97040),
            .I(N__96991));
    InMux I__24138 (
            .O(N__97039),
            .I(N__96991));
    InMux I__24137 (
            .O(N__97038),
            .I(N__96991));
    InMux I__24136 (
            .O(N__97037),
            .I(N__96991));
    InMux I__24135 (
            .O(N__97036),
            .I(N__96985));
    InMux I__24134 (
            .O(N__97035),
            .I(N__96982));
    InMux I__24133 (
            .O(N__97034),
            .I(N__96977));
    LocalMux I__24132 (
            .O(N__97031),
            .I(N__96974));
    LocalMux I__24131 (
            .O(N__97026),
            .I(N__96971));
    InMux I__24130 (
            .O(N__97025),
            .I(N__96964));
    InMux I__24129 (
            .O(N__97024),
            .I(N__96964));
    InMux I__24128 (
            .O(N__97023),
            .I(N__96964));
    InMux I__24127 (
            .O(N__97022),
            .I(N__96959));
    InMux I__24126 (
            .O(N__97021),
            .I(N__96959));
    Span4Mux_h I__24125 (
            .O(N__97018),
            .I(N__96954));
    LocalMux I__24124 (
            .O(N__97013),
            .I(N__96954));
    LocalMux I__24123 (
            .O(N__97010),
            .I(N__96949));
    LocalMux I__24122 (
            .O(N__97005),
            .I(N__96949));
    Span4Mux_h I__24121 (
            .O(N__97002),
            .I(N__96944));
    LocalMux I__24120 (
            .O(N__96991),
            .I(N__96944));
    InMux I__24119 (
            .O(N__96990),
            .I(N__96938));
    InMux I__24118 (
            .O(N__96989),
            .I(N__96935));
    InMux I__24117 (
            .O(N__96988),
            .I(N__96931));
    LocalMux I__24116 (
            .O(N__96985),
            .I(N__96928));
    LocalMux I__24115 (
            .O(N__96982),
            .I(N__96925));
    InMux I__24114 (
            .O(N__96981),
            .I(N__96920));
    InMux I__24113 (
            .O(N__96980),
            .I(N__96920));
    LocalMux I__24112 (
            .O(N__96977),
            .I(N__96917));
    Span4Mux_h I__24111 (
            .O(N__96974),
            .I(N__96910));
    Span4Mux_h I__24110 (
            .O(N__96971),
            .I(N__96910));
    LocalMux I__24109 (
            .O(N__96964),
            .I(N__96910));
    LocalMux I__24108 (
            .O(N__96959),
            .I(N__96905));
    Span4Mux_h I__24107 (
            .O(N__96954),
            .I(N__96905));
    Span4Mux_h I__24106 (
            .O(N__96949),
            .I(N__96900));
    Span4Mux_v I__24105 (
            .O(N__96944),
            .I(N__96900));
    InMux I__24104 (
            .O(N__96943),
            .I(N__96895));
    InMux I__24103 (
            .O(N__96942),
            .I(N__96895));
    InMux I__24102 (
            .O(N__96941),
            .I(N__96892));
    LocalMux I__24101 (
            .O(N__96938),
            .I(N__96889));
    LocalMux I__24100 (
            .O(N__96935),
            .I(N__96886));
    InMux I__24099 (
            .O(N__96934),
            .I(N__96883));
    LocalMux I__24098 (
            .O(N__96931),
            .I(N__96880));
    Span4Mux_v I__24097 (
            .O(N__96928),
            .I(N__96877));
    Sp12to4 I__24096 (
            .O(N__96925),
            .I(N__96874));
    LocalMux I__24095 (
            .O(N__96920),
            .I(N__96871));
    Span4Mux_h I__24094 (
            .O(N__96917),
            .I(N__96868));
    Span4Mux_h I__24093 (
            .O(N__96910),
            .I(N__96863));
    Span4Mux_v I__24092 (
            .O(N__96905),
            .I(N__96863));
    Span4Mux_h I__24091 (
            .O(N__96900),
            .I(N__96860));
    LocalMux I__24090 (
            .O(N__96895),
            .I(N__96857));
    LocalMux I__24089 (
            .O(N__96892),
            .I(N__96852));
    Span4Mux_h I__24088 (
            .O(N__96889),
            .I(N__96852));
    Span4Mux_v I__24087 (
            .O(N__96886),
            .I(N__96849));
    LocalMux I__24086 (
            .O(N__96883),
            .I(N__96842));
    Span4Mux_v I__24085 (
            .O(N__96880),
            .I(N__96842));
    Span4Mux_h I__24084 (
            .O(N__96877),
            .I(N__96842));
    Span12Mux_h I__24083 (
            .O(N__96874),
            .I(N__96837));
    Span12Mux_s11_v I__24082 (
            .O(N__96871),
            .I(N__96837));
    Span4Mux_v I__24081 (
            .O(N__96868),
            .I(N__96830));
    Span4Mux_h I__24080 (
            .O(N__96863),
            .I(N__96830));
    Span4Mux_v I__24079 (
            .O(N__96860),
            .I(N__96830));
    Odrv12 I__24078 (
            .O(N__96857),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n55 ));
    Odrv4 I__24077 (
            .O(N__96852),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n55 ));
    Odrv4 I__24076 (
            .O(N__96849),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n55 ));
    Odrv4 I__24075 (
            .O(N__96842),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n55 ));
    Odrv12 I__24074 (
            .O(N__96837),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n55 ));
    Odrv4 I__24073 (
            .O(N__96830),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n55 ));
    InMux I__24072 (
            .O(N__96817),
            .I(N__96808));
    InMux I__24071 (
            .O(N__96816),
            .I(N__96801));
    InMux I__24070 (
            .O(N__96815),
            .I(N__96801));
    InMux I__24069 (
            .O(N__96814),
            .I(N__96794));
    InMux I__24068 (
            .O(N__96813),
            .I(N__96794));
    InMux I__24067 (
            .O(N__96812),
            .I(N__96794));
    InMux I__24066 (
            .O(N__96811),
            .I(N__96791));
    LocalMux I__24065 (
            .O(N__96808),
            .I(N__96788));
    InMux I__24064 (
            .O(N__96807),
            .I(N__96785));
    InMux I__24063 (
            .O(N__96806),
            .I(N__96779));
    LocalMux I__24062 (
            .O(N__96801),
            .I(N__96764));
    LocalMux I__24061 (
            .O(N__96794),
            .I(N__96764));
    LocalMux I__24060 (
            .O(N__96791),
            .I(N__96757));
    Span4Mux_h I__24059 (
            .O(N__96788),
            .I(N__96757));
    LocalMux I__24058 (
            .O(N__96785),
            .I(N__96757));
    InMux I__24057 (
            .O(N__96784),
            .I(N__96754));
    InMux I__24056 (
            .O(N__96783),
            .I(N__96751));
    InMux I__24055 (
            .O(N__96782),
            .I(N__96747));
    LocalMux I__24054 (
            .O(N__96779),
            .I(N__96744));
    InMux I__24053 (
            .O(N__96778),
            .I(N__96741));
    InMux I__24052 (
            .O(N__96777),
            .I(N__96724));
    InMux I__24051 (
            .O(N__96776),
            .I(N__96721));
    InMux I__24050 (
            .O(N__96775),
            .I(N__96718));
    InMux I__24049 (
            .O(N__96774),
            .I(N__96713));
    InMux I__24048 (
            .O(N__96773),
            .I(N__96713));
    InMux I__24047 (
            .O(N__96772),
            .I(N__96706));
    InMux I__24046 (
            .O(N__96771),
            .I(N__96703));
    InMux I__24045 (
            .O(N__96770),
            .I(N__96700));
    InMux I__24044 (
            .O(N__96769),
            .I(N__96691));
    Span4Mux_v I__24043 (
            .O(N__96764),
            .I(N__96682));
    Span4Mux_v I__24042 (
            .O(N__96757),
            .I(N__96682));
    LocalMux I__24041 (
            .O(N__96754),
            .I(N__96682));
    LocalMux I__24040 (
            .O(N__96751),
            .I(N__96682));
    InMux I__24039 (
            .O(N__96750),
            .I(N__96679));
    LocalMux I__24038 (
            .O(N__96747),
            .I(N__96676));
    Span4Mux_v I__24037 (
            .O(N__96744),
            .I(N__96671));
    LocalMux I__24036 (
            .O(N__96741),
            .I(N__96671));
    InMux I__24035 (
            .O(N__96740),
            .I(N__96666));
    InMux I__24034 (
            .O(N__96739),
            .I(N__96666));
    InMux I__24033 (
            .O(N__96738),
            .I(N__96661));
    InMux I__24032 (
            .O(N__96737),
            .I(N__96654));
    InMux I__24031 (
            .O(N__96736),
            .I(N__96654));
    InMux I__24030 (
            .O(N__96735),
            .I(N__96654));
    InMux I__24029 (
            .O(N__96734),
            .I(N__96651));
    InMux I__24028 (
            .O(N__96733),
            .I(N__96646));
    InMux I__24027 (
            .O(N__96732),
            .I(N__96646));
    InMux I__24026 (
            .O(N__96731),
            .I(N__96643));
    InMux I__24025 (
            .O(N__96730),
            .I(N__96640));
    InMux I__24024 (
            .O(N__96729),
            .I(N__96632));
    InMux I__24023 (
            .O(N__96728),
            .I(N__96629));
    InMux I__24022 (
            .O(N__96727),
            .I(N__96626));
    LocalMux I__24021 (
            .O(N__96724),
            .I(N__96623));
    LocalMux I__24020 (
            .O(N__96721),
            .I(N__96616));
    LocalMux I__24019 (
            .O(N__96718),
            .I(N__96616));
    LocalMux I__24018 (
            .O(N__96713),
            .I(N__96616));
    InMux I__24017 (
            .O(N__96712),
            .I(N__96607));
    InMux I__24016 (
            .O(N__96711),
            .I(N__96607));
    InMux I__24015 (
            .O(N__96710),
            .I(N__96607));
    InMux I__24014 (
            .O(N__96709),
            .I(N__96607));
    LocalMux I__24013 (
            .O(N__96706),
            .I(N__96604));
    LocalMux I__24012 (
            .O(N__96703),
            .I(N__96599));
    LocalMux I__24011 (
            .O(N__96700),
            .I(N__96599));
    InMux I__24010 (
            .O(N__96699),
            .I(N__96588));
    InMux I__24009 (
            .O(N__96698),
            .I(N__96588));
    InMux I__24008 (
            .O(N__96697),
            .I(N__96588));
    InMux I__24007 (
            .O(N__96696),
            .I(N__96588));
    InMux I__24006 (
            .O(N__96695),
            .I(N__96588));
    InMux I__24005 (
            .O(N__96694),
            .I(N__96585));
    LocalMux I__24004 (
            .O(N__96691),
            .I(N__96577));
    Span4Mux_h I__24003 (
            .O(N__96682),
            .I(N__96568));
    LocalMux I__24002 (
            .O(N__96679),
            .I(N__96568));
    Span4Mux_h I__24001 (
            .O(N__96676),
            .I(N__96561));
    Span4Mux_v I__24000 (
            .O(N__96671),
            .I(N__96561));
    LocalMux I__23999 (
            .O(N__96666),
            .I(N__96561));
    InMux I__23998 (
            .O(N__96665),
            .I(N__96558));
    InMux I__23997 (
            .O(N__96664),
            .I(N__96555));
    LocalMux I__23996 (
            .O(N__96661),
            .I(N__96548));
    LocalMux I__23995 (
            .O(N__96654),
            .I(N__96548));
    LocalMux I__23994 (
            .O(N__96651),
            .I(N__96548));
    LocalMux I__23993 (
            .O(N__96646),
            .I(N__96541));
    LocalMux I__23992 (
            .O(N__96643),
            .I(N__96541));
    LocalMux I__23991 (
            .O(N__96640),
            .I(N__96541));
    InMux I__23990 (
            .O(N__96639),
            .I(N__96538));
    InMux I__23989 (
            .O(N__96638),
            .I(N__96529));
    InMux I__23988 (
            .O(N__96637),
            .I(N__96529));
    InMux I__23987 (
            .O(N__96636),
            .I(N__96529));
    InMux I__23986 (
            .O(N__96635),
            .I(N__96529));
    LocalMux I__23985 (
            .O(N__96632),
            .I(N__96525));
    LocalMux I__23984 (
            .O(N__96629),
            .I(N__96520));
    LocalMux I__23983 (
            .O(N__96626),
            .I(N__96520));
    Span4Mux_h I__23982 (
            .O(N__96623),
            .I(N__96513));
    Span4Mux_v I__23981 (
            .O(N__96616),
            .I(N__96513));
    LocalMux I__23980 (
            .O(N__96607),
            .I(N__96513));
    Span4Mux_h I__23979 (
            .O(N__96604),
            .I(N__96504));
    Span4Mux_v I__23978 (
            .O(N__96599),
            .I(N__96504));
    LocalMux I__23977 (
            .O(N__96588),
            .I(N__96504));
    LocalMux I__23976 (
            .O(N__96585),
            .I(N__96504));
    InMux I__23975 (
            .O(N__96584),
            .I(N__96493));
    InMux I__23974 (
            .O(N__96583),
            .I(N__96493));
    InMux I__23973 (
            .O(N__96582),
            .I(N__96493));
    InMux I__23972 (
            .O(N__96581),
            .I(N__96493));
    InMux I__23971 (
            .O(N__96580),
            .I(N__96493));
    Sp12to4 I__23970 (
            .O(N__96577),
            .I(N__96490));
    InMux I__23969 (
            .O(N__96576),
            .I(N__96485));
    InMux I__23968 (
            .O(N__96575),
            .I(N__96485));
    InMux I__23967 (
            .O(N__96574),
            .I(N__96480));
    InMux I__23966 (
            .O(N__96573),
            .I(N__96480));
    Span4Mux_h I__23965 (
            .O(N__96568),
            .I(N__96477));
    Span4Mux_h I__23964 (
            .O(N__96561),
            .I(N__96472));
    LocalMux I__23963 (
            .O(N__96558),
            .I(N__96472));
    LocalMux I__23962 (
            .O(N__96555),
            .I(N__96461));
    Span12Mux_v I__23961 (
            .O(N__96548),
            .I(N__96461));
    Span12Mux_v I__23960 (
            .O(N__96541),
            .I(N__96461));
    LocalMux I__23959 (
            .O(N__96538),
            .I(N__96461));
    LocalMux I__23958 (
            .O(N__96529),
            .I(N__96461));
    InMux I__23957 (
            .O(N__96528),
            .I(N__96458));
    Span4Mux_v I__23956 (
            .O(N__96525),
            .I(N__96447));
    Span4Mux_v I__23955 (
            .O(N__96520),
            .I(N__96447));
    Span4Mux_h I__23954 (
            .O(N__96513),
            .I(N__96447));
    Span4Mux_v I__23953 (
            .O(N__96504),
            .I(N__96447));
    LocalMux I__23952 (
            .O(N__96493),
            .I(N__96447));
    Odrv12 I__23951 (
            .O(N__96490),
            .I(dc32_fifo_data_in_1));
    LocalMux I__23950 (
            .O(N__96485),
            .I(dc32_fifo_data_in_1));
    LocalMux I__23949 (
            .O(N__96480),
            .I(dc32_fifo_data_in_1));
    Odrv4 I__23948 (
            .O(N__96477),
            .I(dc32_fifo_data_in_1));
    Odrv4 I__23947 (
            .O(N__96472),
            .I(dc32_fifo_data_in_1));
    Odrv12 I__23946 (
            .O(N__96461),
            .I(dc32_fifo_data_in_1));
    LocalMux I__23945 (
            .O(N__96458),
            .I(dc32_fifo_data_in_1));
    Odrv4 I__23944 (
            .O(N__96447),
            .I(dc32_fifo_data_in_1));
    CascadeMux I__23943 (
            .O(N__96430),
            .I(N__96426));
    InMux I__23942 (
            .O(N__96429),
            .I(N__96423));
    InMux I__23941 (
            .O(N__96426),
            .I(N__96420));
    LocalMux I__23940 (
            .O(N__96423),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_1 ));
    LocalMux I__23939 (
            .O(N__96420),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_1 ));
    InMux I__23938 (
            .O(N__96415),
            .I(N__96412));
    LocalMux I__23937 (
            .O(N__96412),
            .I(N__96409));
    Span4Mux_h I__23936 (
            .O(N__96409),
            .I(N__96405));
    CascadeMux I__23935 (
            .O(N__96408),
            .I(N__96402));
    Span4Mux_v I__23934 (
            .O(N__96405),
            .I(N__96399));
    InMux I__23933 (
            .O(N__96402),
            .I(N__96396));
    Odrv4 I__23932 (
            .O(N__96399),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_6 ));
    LocalMux I__23931 (
            .O(N__96396),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_6 ));
    InMux I__23930 (
            .O(N__96391),
            .I(N__96383));
    InMux I__23929 (
            .O(N__96390),
            .I(N__96371));
    InMux I__23928 (
            .O(N__96389),
            .I(N__96371));
    InMux I__23927 (
            .O(N__96388),
            .I(N__96371));
    InMux I__23926 (
            .O(N__96387),
            .I(N__96371));
    InMux I__23925 (
            .O(N__96386),
            .I(N__96371));
    LocalMux I__23924 (
            .O(N__96383),
            .I(N__96362));
    InMux I__23923 (
            .O(N__96382),
            .I(N__96359));
    LocalMux I__23922 (
            .O(N__96371),
            .I(N__96346));
    InMux I__23921 (
            .O(N__96370),
            .I(N__96337));
    InMux I__23920 (
            .O(N__96369),
            .I(N__96328));
    InMux I__23919 (
            .O(N__96368),
            .I(N__96328));
    InMux I__23918 (
            .O(N__96367),
            .I(N__96328));
    InMux I__23917 (
            .O(N__96366),
            .I(N__96328));
    InMux I__23916 (
            .O(N__96365),
            .I(N__96325));
    Span4Mux_v I__23915 (
            .O(N__96362),
            .I(N__96316));
    LocalMux I__23914 (
            .O(N__96359),
            .I(N__96316));
    InMux I__23913 (
            .O(N__96358),
            .I(N__96299));
    InMux I__23912 (
            .O(N__96357),
            .I(N__96299));
    InMux I__23911 (
            .O(N__96356),
            .I(N__96299));
    InMux I__23910 (
            .O(N__96355),
            .I(N__96299));
    InMux I__23909 (
            .O(N__96354),
            .I(N__96299));
    InMux I__23908 (
            .O(N__96353),
            .I(N__96299));
    InMux I__23907 (
            .O(N__96352),
            .I(N__96296));
    InMux I__23906 (
            .O(N__96351),
            .I(N__96289));
    InMux I__23905 (
            .O(N__96350),
            .I(N__96289));
    InMux I__23904 (
            .O(N__96349),
            .I(N__96289));
    Span4Mux_v I__23903 (
            .O(N__96346),
            .I(N__96286));
    InMux I__23902 (
            .O(N__96345),
            .I(N__96281));
    InMux I__23901 (
            .O(N__96344),
            .I(N__96281));
    InMux I__23900 (
            .O(N__96343),
            .I(N__96276));
    InMux I__23899 (
            .O(N__96342),
            .I(N__96276));
    CascadeMux I__23898 (
            .O(N__96341),
            .I(N__96273));
    CascadeMux I__23897 (
            .O(N__96340),
            .I(N__96270));
    LocalMux I__23896 (
            .O(N__96337),
            .I(N__96264));
    LocalMux I__23895 (
            .O(N__96328),
            .I(N__96264));
    LocalMux I__23894 (
            .O(N__96325),
            .I(N__96261));
    InMux I__23893 (
            .O(N__96324),
            .I(N__96257));
    InMux I__23892 (
            .O(N__96323),
            .I(N__96252));
    InMux I__23891 (
            .O(N__96322),
            .I(N__96252));
    CascadeMux I__23890 (
            .O(N__96321),
            .I(N__96248));
    Span4Mux_h I__23889 (
            .O(N__96316),
            .I(N__96240));
    InMux I__23888 (
            .O(N__96315),
            .I(N__96237));
    InMux I__23887 (
            .O(N__96314),
            .I(N__96232));
    InMux I__23886 (
            .O(N__96313),
            .I(N__96232));
    InMux I__23885 (
            .O(N__96312),
            .I(N__96222));
    LocalMux I__23884 (
            .O(N__96299),
            .I(N__96215));
    LocalMux I__23883 (
            .O(N__96296),
            .I(N__96215));
    LocalMux I__23882 (
            .O(N__96289),
            .I(N__96215));
    Span4Mux_h I__23881 (
            .O(N__96286),
            .I(N__96210));
    LocalMux I__23880 (
            .O(N__96281),
            .I(N__96210));
    LocalMux I__23879 (
            .O(N__96276),
            .I(N__96206));
    InMux I__23878 (
            .O(N__96273),
            .I(N__96199));
    InMux I__23877 (
            .O(N__96270),
            .I(N__96199));
    InMux I__23876 (
            .O(N__96269),
            .I(N__96199));
    Span4Mux_v I__23875 (
            .O(N__96264),
            .I(N__96194));
    Span4Mux_v I__23874 (
            .O(N__96261),
            .I(N__96194));
    InMux I__23873 (
            .O(N__96260),
            .I(N__96186));
    LocalMux I__23872 (
            .O(N__96257),
            .I(N__96183));
    LocalMux I__23871 (
            .O(N__96252),
            .I(N__96180));
    InMux I__23870 (
            .O(N__96251),
            .I(N__96177));
    InMux I__23869 (
            .O(N__96248),
            .I(N__96174));
    InMux I__23868 (
            .O(N__96247),
            .I(N__96163));
    InMux I__23867 (
            .O(N__96246),
            .I(N__96163));
    InMux I__23866 (
            .O(N__96245),
            .I(N__96163));
    InMux I__23865 (
            .O(N__96244),
            .I(N__96163));
    InMux I__23864 (
            .O(N__96243),
            .I(N__96163));
    Span4Mux_v I__23863 (
            .O(N__96240),
            .I(N__96158));
    LocalMux I__23862 (
            .O(N__96237),
            .I(N__96158));
    LocalMux I__23861 (
            .O(N__96232),
            .I(N__96149));
    InMux I__23860 (
            .O(N__96231),
            .I(N__96144));
    InMux I__23859 (
            .O(N__96230),
            .I(N__96144));
    InMux I__23858 (
            .O(N__96229),
            .I(N__96141));
    InMux I__23857 (
            .O(N__96228),
            .I(N__96132));
    InMux I__23856 (
            .O(N__96227),
            .I(N__96132));
    InMux I__23855 (
            .O(N__96226),
            .I(N__96132));
    InMux I__23854 (
            .O(N__96225),
            .I(N__96132));
    LocalMux I__23853 (
            .O(N__96222),
            .I(N__96125));
    Span4Mux_v I__23852 (
            .O(N__96215),
            .I(N__96125));
    Span4Mux_h I__23851 (
            .O(N__96210),
            .I(N__96125));
    InMux I__23850 (
            .O(N__96209),
            .I(N__96122));
    Span4Mux_h I__23849 (
            .O(N__96206),
            .I(N__96115));
    LocalMux I__23848 (
            .O(N__96199),
            .I(N__96115));
    Span4Mux_h I__23847 (
            .O(N__96194),
            .I(N__96115));
    InMux I__23846 (
            .O(N__96193),
            .I(N__96106));
    InMux I__23845 (
            .O(N__96192),
            .I(N__96106));
    InMux I__23844 (
            .O(N__96191),
            .I(N__96106));
    InMux I__23843 (
            .O(N__96190),
            .I(N__96106));
    InMux I__23842 (
            .O(N__96189),
            .I(N__96103));
    LocalMux I__23841 (
            .O(N__96186),
            .I(N__96100));
    Span4Mux_v I__23840 (
            .O(N__96183),
            .I(N__96089));
    Span4Mux_h I__23839 (
            .O(N__96180),
            .I(N__96089));
    LocalMux I__23838 (
            .O(N__96177),
            .I(N__96089));
    LocalMux I__23837 (
            .O(N__96174),
            .I(N__96089));
    LocalMux I__23836 (
            .O(N__96163),
            .I(N__96089));
    Span4Mux_v I__23835 (
            .O(N__96158),
            .I(N__96086));
    InMux I__23834 (
            .O(N__96157),
            .I(N__96083));
    InMux I__23833 (
            .O(N__96156),
            .I(N__96072));
    InMux I__23832 (
            .O(N__96155),
            .I(N__96072));
    InMux I__23831 (
            .O(N__96154),
            .I(N__96072));
    InMux I__23830 (
            .O(N__96153),
            .I(N__96072));
    InMux I__23829 (
            .O(N__96152),
            .I(N__96072));
    Span4Mux_v I__23828 (
            .O(N__96149),
            .I(N__96067));
    LocalMux I__23827 (
            .O(N__96144),
            .I(N__96067));
    LocalMux I__23826 (
            .O(N__96141),
            .I(N__96064));
    LocalMux I__23825 (
            .O(N__96132),
            .I(N__96053));
    Sp12to4 I__23824 (
            .O(N__96125),
            .I(N__96053));
    LocalMux I__23823 (
            .O(N__96122),
            .I(N__96053));
    Sp12to4 I__23822 (
            .O(N__96115),
            .I(N__96053));
    LocalMux I__23821 (
            .O(N__96106),
            .I(N__96053));
    LocalMux I__23820 (
            .O(N__96103),
            .I(N__96048));
    Span4Mux_v I__23819 (
            .O(N__96100),
            .I(N__96048));
    Span4Mux_v I__23818 (
            .O(N__96089),
            .I(N__96045));
    Span4Mux_v I__23817 (
            .O(N__96086),
            .I(N__96040));
    LocalMux I__23816 (
            .O(N__96083),
            .I(N__96040));
    LocalMux I__23815 (
            .O(N__96072),
            .I(N__96037));
    Span4Mux_h I__23814 (
            .O(N__96067),
            .I(N__96032));
    Span4Mux_h I__23813 (
            .O(N__96064),
            .I(N__96032));
    Span12Mux_v I__23812 (
            .O(N__96053),
            .I(N__96029));
    Span4Mux_v I__23811 (
            .O(N__96048),
            .I(N__96022));
    Span4Mux_h I__23810 (
            .O(N__96045),
            .I(N__96022));
    Span4Mux_h I__23809 (
            .O(N__96040),
            .I(N__96022));
    Odrv4 I__23808 (
            .O(N__96037),
            .I(dc32_fifo_data_in_6));
    Odrv4 I__23807 (
            .O(N__96032),
            .I(dc32_fifo_data_in_6));
    Odrv12 I__23806 (
            .O(N__96029),
            .I(dc32_fifo_data_in_6));
    Odrv4 I__23805 (
            .O(N__96022),
            .I(dc32_fifo_data_in_6));
    InMux I__23804 (
            .O(N__96013),
            .I(N__96000));
    InMux I__23803 (
            .O(N__96012),
            .I(N__95994));
    InMux I__23802 (
            .O(N__96011),
            .I(N__95991));
    InMux I__23801 (
            .O(N__96010),
            .I(N__95986));
    InMux I__23800 (
            .O(N__96009),
            .I(N__95973));
    InMux I__23799 (
            .O(N__96008),
            .I(N__95973));
    InMux I__23798 (
            .O(N__96007),
            .I(N__95970));
    InMux I__23797 (
            .O(N__96006),
            .I(N__95967));
    InMux I__23796 (
            .O(N__96005),
            .I(N__95962));
    InMux I__23795 (
            .O(N__96004),
            .I(N__95962));
    InMux I__23794 (
            .O(N__96003),
            .I(N__95959));
    LocalMux I__23793 (
            .O(N__96000),
            .I(N__95956));
    InMux I__23792 (
            .O(N__95999),
            .I(N__95950));
    InMux I__23791 (
            .O(N__95998),
            .I(N__95950));
    InMux I__23790 (
            .O(N__95997),
            .I(N__95947));
    LocalMux I__23789 (
            .O(N__95994),
            .I(N__95944));
    LocalMux I__23788 (
            .O(N__95991),
            .I(N__95941));
    CascadeMux I__23787 (
            .O(N__95990),
            .I(N__95938));
    InMux I__23786 (
            .O(N__95989),
            .I(N__95934));
    LocalMux I__23785 (
            .O(N__95986),
            .I(N__95931));
    InMux I__23784 (
            .O(N__95985),
            .I(N__95925));
    InMux I__23783 (
            .O(N__95984),
            .I(N__95925));
    InMux I__23782 (
            .O(N__95983),
            .I(N__95922));
    InMux I__23781 (
            .O(N__95982),
            .I(N__95915));
    InMux I__23780 (
            .O(N__95981),
            .I(N__95915));
    InMux I__23779 (
            .O(N__95980),
            .I(N__95915));
    InMux I__23778 (
            .O(N__95979),
            .I(N__95910));
    InMux I__23777 (
            .O(N__95978),
            .I(N__95910));
    LocalMux I__23776 (
            .O(N__95973),
            .I(N__95907));
    LocalMux I__23775 (
            .O(N__95970),
            .I(N__95902));
    LocalMux I__23774 (
            .O(N__95967),
            .I(N__95902));
    LocalMux I__23773 (
            .O(N__95962),
            .I(N__95899));
    LocalMux I__23772 (
            .O(N__95959),
            .I(N__95894));
    Span4Mux_h I__23771 (
            .O(N__95956),
            .I(N__95894));
    InMux I__23770 (
            .O(N__95955),
            .I(N__95887));
    LocalMux I__23769 (
            .O(N__95950),
            .I(N__95884));
    LocalMux I__23768 (
            .O(N__95947),
            .I(N__95881));
    Span4Mux_h I__23767 (
            .O(N__95944),
            .I(N__95876));
    Span4Mux_v I__23766 (
            .O(N__95941),
            .I(N__95876));
    InMux I__23765 (
            .O(N__95938),
            .I(N__95873));
    InMux I__23764 (
            .O(N__95937),
            .I(N__95870));
    LocalMux I__23763 (
            .O(N__95934),
            .I(N__95867));
    Span4Mux_v I__23762 (
            .O(N__95931),
            .I(N__95864));
    InMux I__23761 (
            .O(N__95930),
            .I(N__95861));
    LocalMux I__23760 (
            .O(N__95925),
            .I(N__95858));
    LocalMux I__23759 (
            .O(N__95922),
            .I(N__95851));
    LocalMux I__23758 (
            .O(N__95915),
            .I(N__95851));
    LocalMux I__23757 (
            .O(N__95910),
            .I(N__95851));
    Span4Mux_h I__23756 (
            .O(N__95907),
            .I(N__95844));
    Span4Mux_v I__23755 (
            .O(N__95902),
            .I(N__95844));
    Span4Mux_v I__23754 (
            .O(N__95899),
            .I(N__95844));
    Span4Mux_v I__23753 (
            .O(N__95894),
            .I(N__95841));
    InMux I__23752 (
            .O(N__95893),
            .I(N__95836));
    InMux I__23751 (
            .O(N__95892),
            .I(N__95836));
    InMux I__23750 (
            .O(N__95891),
            .I(N__95833));
    InMux I__23749 (
            .O(N__95890),
            .I(N__95830));
    LocalMux I__23748 (
            .O(N__95887),
            .I(N__95827));
    Span4Mux_h I__23747 (
            .O(N__95884),
            .I(N__95824));
    Span4Mux_h I__23746 (
            .O(N__95881),
            .I(N__95819));
    Span4Mux_h I__23745 (
            .O(N__95876),
            .I(N__95819));
    LocalMux I__23744 (
            .O(N__95873),
            .I(N__95810));
    LocalMux I__23743 (
            .O(N__95870),
            .I(N__95810));
    Span4Mux_v I__23742 (
            .O(N__95867),
            .I(N__95810));
    Span4Mux_h I__23741 (
            .O(N__95864),
            .I(N__95810));
    LocalMux I__23740 (
            .O(N__95861),
            .I(N__95803));
    Sp12to4 I__23739 (
            .O(N__95858),
            .I(N__95803));
    Span12Mux_s8_h I__23738 (
            .O(N__95851),
            .I(N__95803));
    Span4Mux_h I__23737 (
            .O(N__95844),
            .I(N__95798));
    Span4Mux_v I__23736 (
            .O(N__95841),
            .I(N__95798));
    LocalMux I__23735 (
            .O(N__95836),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53 ));
    LocalMux I__23734 (
            .O(N__95833),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53 ));
    LocalMux I__23733 (
            .O(N__95830),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53 ));
    Odrv12 I__23732 (
            .O(N__95827),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53 ));
    Odrv4 I__23731 (
            .O(N__95824),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53 ));
    Odrv4 I__23730 (
            .O(N__95819),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53 ));
    Odrv4 I__23729 (
            .O(N__95810),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53 ));
    Odrv12 I__23728 (
            .O(N__95803),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53 ));
    Odrv4 I__23727 (
            .O(N__95798),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53 ));
    CascadeMux I__23726 (
            .O(N__95779),
            .I(N__95776));
    InMux I__23725 (
            .O(N__95776),
            .I(N__95763));
    InMux I__23724 (
            .O(N__95775),
            .I(N__95763));
    InMux I__23723 (
            .O(N__95774),
            .I(N__95763));
    InMux I__23722 (
            .O(N__95773),
            .I(N__95756));
    InMux I__23721 (
            .O(N__95772),
            .I(N__95753));
    CascadeMux I__23720 (
            .O(N__95771),
            .I(N__95737));
    CascadeMux I__23719 (
            .O(N__95770),
            .I(N__95732));
    LocalMux I__23718 (
            .O(N__95763),
            .I(N__95714));
    InMux I__23717 (
            .O(N__95762),
            .I(N__95709));
    InMux I__23716 (
            .O(N__95761),
            .I(N__95709));
    CascadeMux I__23715 (
            .O(N__95760),
            .I(N__95695));
    CascadeMux I__23714 (
            .O(N__95759),
            .I(N__95692));
    LocalMux I__23713 (
            .O(N__95756),
            .I(N__95677));
    LocalMux I__23712 (
            .O(N__95753),
            .I(N__95677));
    InMux I__23711 (
            .O(N__95752),
            .I(N__95672));
    InMux I__23710 (
            .O(N__95751),
            .I(N__95672));
    InMux I__23709 (
            .O(N__95750),
            .I(N__95669));
    InMux I__23708 (
            .O(N__95749),
            .I(N__95658));
    InMux I__23707 (
            .O(N__95748),
            .I(N__95658));
    InMux I__23706 (
            .O(N__95747),
            .I(N__95658));
    InMux I__23705 (
            .O(N__95746),
            .I(N__95658));
    InMux I__23704 (
            .O(N__95745),
            .I(N__95658));
    InMux I__23703 (
            .O(N__95744),
            .I(N__95651));
    InMux I__23702 (
            .O(N__95743),
            .I(N__95651));
    InMux I__23701 (
            .O(N__95742),
            .I(N__95651));
    InMux I__23700 (
            .O(N__95741),
            .I(N__95645));
    InMux I__23699 (
            .O(N__95740),
            .I(N__95645));
    InMux I__23698 (
            .O(N__95737),
            .I(N__95635));
    InMux I__23697 (
            .O(N__95736),
            .I(N__95635));
    InMux I__23696 (
            .O(N__95735),
            .I(N__95635));
    InMux I__23695 (
            .O(N__95732),
            .I(N__95613));
    InMux I__23694 (
            .O(N__95731),
            .I(N__95608));
    InMux I__23693 (
            .O(N__95730),
            .I(N__95608));
    InMux I__23692 (
            .O(N__95729),
            .I(N__95595));
    InMux I__23691 (
            .O(N__95728),
            .I(N__95595));
    InMux I__23690 (
            .O(N__95727),
            .I(N__95595));
    InMux I__23689 (
            .O(N__95726),
            .I(N__95595));
    InMux I__23688 (
            .O(N__95725),
            .I(N__95595));
    InMux I__23687 (
            .O(N__95724),
            .I(N__95595));
    CascadeMux I__23686 (
            .O(N__95723),
            .I(N__95591));
    CascadeMux I__23685 (
            .O(N__95722),
            .I(N__95588));
    CascadeMux I__23684 (
            .O(N__95721),
            .I(N__95585));
    InMux I__23683 (
            .O(N__95720),
            .I(N__95579));
    InMux I__23682 (
            .O(N__95719),
            .I(N__95572));
    InMux I__23681 (
            .O(N__95718),
            .I(N__95572));
    InMux I__23680 (
            .O(N__95717),
            .I(N__95572));
    Span4Mux_v I__23679 (
            .O(N__95714),
            .I(N__95567));
    LocalMux I__23678 (
            .O(N__95709),
            .I(N__95567));
    InMux I__23677 (
            .O(N__95708),
            .I(N__95562));
    InMux I__23676 (
            .O(N__95707),
            .I(N__95562));
    CascadeMux I__23675 (
            .O(N__95706),
            .I(N__95559));
    CascadeMux I__23674 (
            .O(N__95705),
            .I(N__95556));
    CascadeMux I__23673 (
            .O(N__95704),
            .I(N__95550));
    CascadeMux I__23672 (
            .O(N__95703),
            .I(N__95542));
    InMux I__23671 (
            .O(N__95702),
            .I(N__95517));
    InMux I__23670 (
            .O(N__95701),
            .I(N__95517));
    InMux I__23669 (
            .O(N__95700),
            .I(N__95517));
    InMux I__23668 (
            .O(N__95699),
            .I(N__95517));
    InMux I__23667 (
            .O(N__95698),
            .I(N__95517));
    InMux I__23666 (
            .O(N__95695),
            .I(N__95504));
    InMux I__23665 (
            .O(N__95692),
            .I(N__95504));
    InMux I__23664 (
            .O(N__95691),
            .I(N__95504));
    InMux I__23663 (
            .O(N__95690),
            .I(N__95504));
    InMux I__23662 (
            .O(N__95689),
            .I(N__95504));
    InMux I__23661 (
            .O(N__95688),
            .I(N__95504));
    CascadeMux I__23660 (
            .O(N__95687),
            .I(N__95498));
    InMux I__23659 (
            .O(N__95686),
            .I(N__95481));
    InMux I__23658 (
            .O(N__95685),
            .I(N__95481));
    InMux I__23657 (
            .O(N__95684),
            .I(N__95481));
    InMux I__23656 (
            .O(N__95683),
            .I(N__95481));
    InMux I__23655 (
            .O(N__95682),
            .I(N__95481));
    Span4Mux_v I__23654 (
            .O(N__95677),
            .I(N__95478));
    LocalMux I__23653 (
            .O(N__95672),
            .I(N__95475));
    LocalMux I__23652 (
            .O(N__95669),
            .I(N__95470));
    LocalMux I__23651 (
            .O(N__95658),
            .I(N__95470));
    LocalMux I__23650 (
            .O(N__95651),
            .I(N__95467));
    CascadeMux I__23649 (
            .O(N__95650),
            .I(N__95453));
    LocalMux I__23648 (
            .O(N__95645),
            .I(N__95439));
    InMux I__23647 (
            .O(N__95644),
            .I(N__95436));
    InMux I__23646 (
            .O(N__95643),
            .I(N__95431));
    InMux I__23645 (
            .O(N__95642),
            .I(N__95431));
    LocalMux I__23644 (
            .O(N__95635),
            .I(N__95428));
    CascadeMux I__23643 (
            .O(N__95634),
            .I(N__95404));
    InMux I__23642 (
            .O(N__95633),
            .I(N__95364));
    InMux I__23641 (
            .O(N__95632),
            .I(N__95359));
    InMux I__23640 (
            .O(N__95631),
            .I(N__95359));
    InMux I__23639 (
            .O(N__95630),
            .I(N__95356));
    InMux I__23638 (
            .O(N__95629),
            .I(N__95349));
    InMux I__23637 (
            .O(N__95628),
            .I(N__95349));
    InMux I__23636 (
            .O(N__95627),
            .I(N__95349));
    CascadeMux I__23635 (
            .O(N__95626),
            .I(N__95339));
    CascadeMux I__23634 (
            .O(N__95625),
            .I(N__95330));
    CascadeMux I__23633 (
            .O(N__95624),
            .I(N__95327));
    InMux I__23632 (
            .O(N__95623),
            .I(N__95305));
    InMux I__23631 (
            .O(N__95622),
            .I(N__95305));
    InMux I__23630 (
            .O(N__95621),
            .I(N__95305));
    InMux I__23629 (
            .O(N__95620),
            .I(N__95305));
    InMux I__23628 (
            .O(N__95619),
            .I(N__95300));
    InMux I__23627 (
            .O(N__95618),
            .I(N__95300));
    CascadeMux I__23626 (
            .O(N__95617),
            .I(N__95295));
    CascadeMux I__23625 (
            .O(N__95616),
            .I(N__95291));
    LocalMux I__23624 (
            .O(N__95613),
            .I(N__95276));
    LocalMux I__23623 (
            .O(N__95608),
            .I(N__95276));
    LocalMux I__23622 (
            .O(N__95595),
            .I(N__95276));
    InMux I__23621 (
            .O(N__95594),
            .I(N__95273));
    InMux I__23620 (
            .O(N__95591),
            .I(N__95262));
    InMux I__23619 (
            .O(N__95588),
            .I(N__95262));
    InMux I__23618 (
            .O(N__95585),
            .I(N__95262));
    InMux I__23617 (
            .O(N__95584),
            .I(N__95262));
    InMux I__23616 (
            .O(N__95583),
            .I(N__95262));
    InMux I__23615 (
            .O(N__95582),
            .I(N__95259));
    LocalMux I__23614 (
            .O(N__95579),
            .I(N__95254));
    LocalMux I__23613 (
            .O(N__95572),
            .I(N__95254));
    Span4Mux_h I__23612 (
            .O(N__95567),
            .I(N__95249));
    LocalMux I__23611 (
            .O(N__95562),
            .I(N__95249));
    InMux I__23610 (
            .O(N__95559),
            .I(N__95238));
    InMux I__23609 (
            .O(N__95556),
            .I(N__95238));
    InMux I__23608 (
            .O(N__95555),
            .I(N__95238));
    InMux I__23607 (
            .O(N__95554),
            .I(N__95238));
    InMux I__23606 (
            .O(N__95553),
            .I(N__95238));
    InMux I__23605 (
            .O(N__95550),
            .I(N__95225));
    InMux I__23604 (
            .O(N__95549),
            .I(N__95225));
    InMux I__23603 (
            .O(N__95548),
            .I(N__95225));
    InMux I__23602 (
            .O(N__95547),
            .I(N__95225));
    InMux I__23601 (
            .O(N__95546),
            .I(N__95225));
    InMux I__23600 (
            .O(N__95545),
            .I(N__95225));
    InMux I__23599 (
            .O(N__95542),
            .I(N__95211));
    InMux I__23598 (
            .O(N__95541),
            .I(N__95211));
    InMux I__23597 (
            .O(N__95540),
            .I(N__95211));
    InMux I__23596 (
            .O(N__95539),
            .I(N__95206));
    InMux I__23595 (
            .O(N__95538),
            .I(N__95206));
    InMux I__23594 (
            .O(N__95537),
            .I(N__95197));
    InMux I__23593 (
            .O(N__95536),
            .I(N__95197));
    InMux I__23592 (
            .O(N__95535),
            .I(N__95197));
    InMux I__23591 (
            .O(N__95534),
            .I(N__95197));
    InMux I__23590 (
            .O(N__95533),
            .I(N__95186));
    InMux I__23589 (
            .O(N__95532),
            .I(N__95186));
    InMux I__23588 (
            .O(N__95531),
            .I(N__95186));
    InMux I__23587 (
            .O(N__95530),
            .I(N__95186));
    InMux I__23586 (
            .O(N__95529),
            .I(N__95186));
    InMux I__23585 (
            .O(N__95528),
            .I(N__95183));
    LocalMux I__23584 (
            .O(N__95517),
            .I(N__95178));
    LocalMux I__23583 (
            .O(N__95504),
            .I(N__95178));
    InMux I__23582 (
            .O(N__95503),
            .I(N__95166));
    InMux I__23581 (
            .O(N__95502),
            .I(N__95166));
    InMux I__23580 (
            .O(N__95501),
            .I(N__95166));
    InMux I__23579 (
            .O(N__95498),
            .I(N__95157));
    InMux I__23578 (
            .O(N__95497),
            .I(N__95157));
    InMux I__23577 (
            .O(N__95496),
            .I(N__95157));
    InMux I__23576 (
            .O(N__95495),
            .I(N__95157));
    InMux I__23575 (
            .O(N__95494),
            .I(N__95139));
    InMux I__23574 (
            .O(N__95493),
            .I(N__95139));
    InMux I__23573 (
            .O(N__95492),
            .I(N__95139));
    LocalMux I__23572 (
            .O(N__95481),
            .I(N__95132));
    Span4Mux_h I__23571 (
            .O(N__95478),
            .I(N__95132));
    Span4Mux_v I__23570 (
            .O(N__95475),
            .I(N__95132));
    Span4Mux_v I__23569 (
            .O(N__95470),
            .I(N__95127));
    Span4Mux_v I__23568 (
            .O(N__95467),
            .I(N__95127));
    InMux I__23567 (
            .O(N__95466),
            .I(N__95122));
    InMux I__23566 (
            .O(N__95465),
            .I(N__95122));
    InMux I__23565 (
            .O(N__95464),
            .I(N__95119));
    InMux I__23564 (
            .O(N__95463),
            .I(N__95106));
    InMux I__23563 (
            .O(N__95462),
            .I(N__95106));
    InMux I__23562 (
            .O(N__95461),
            .I(N__95106));
    InMux I__23561 (
            .O(N__95460),
            .I(N__95106));
    InMux I__23560 (
            .O(N__95459),
            .I(N__95106));
    InMux I__23559 (
            .O(N__95458),
            .I(N__95106));
    CascadeMux I__23558 (
            .O(N__95457),
            .I(N__95084));
    CascadeMux I__23557 (
            .O(N__95456),
            .I(N__95081));
    InMux I__23556 (
            .O(N__95453),
            .I(N__95070));
    InMux I__23555 (
            .O(N__95452),
            .I(N__95070));
    InMux I__23554 (
            .O(N__95451),
            .I(N__95067));
    InMux I__23553 (
            .O(N__95450),
            .I(N__95058));
    InMux I__23552 (
            .O(N__95449),
            .I(N__95058));
    InMux I__23551 (
            .O(N__95448),
            .I(N__95058));
    InMux I__23550 (
            .O(N__95447),
            .I(N__95058));
    InMux I__23549 (
            .O(N__95446),
            .I(N__95055));
    InMux I__23548 (
            .O(N__95445),
            .I(N__95039));
    InMux I__23547 (
            .O(N__95444),
            .I(N__95039));
    InMux I__23546 (
            .O(N__95443),
            .I(N__95039));
    InMux I__23545 (
            .O(N__95442),
            .I(N__95039));
    Span4Mux_v I__23544 (
            .O(N__95439),
            .I(N__95030));
    LocalMux I__23543 (
            .O(N__95436),
            .I(N__95030));
    LocalMux I__23542 (
            .O(N__95431),
            .I(N__95030));
    Span4Mux_v I__23541 (
            .O(N__95428),
            .I(N__95030));
    InMux I__23540 (
            .O(N__95427),
            .I(N__95019));
    InMux I__23539 (
            .O(N__95426),
            .I(N__95019));
    InMux I__23538 (
            .O(N__95425),
            .I(N__95019));
    InMux I__23537 (
            .O(N__95424),
            .I(N__95019));
    InMux I__23536 (
            .O(N__95423),
            .I(N__95019));
    InMux I__23535 (
            .O(N__95422),
            .I(N__95010));
    InMux I__23534 (
            .O(N__95421),
            .I(N__95010));
    InMux I__23533 (
            .O(N__95420),
            .I(N__95010));
    InMux I__23532 (
            .O(N__95419),
            .I(N__95010));
    InMux I__23531 (
            .O(N__95418),
            .I(N__95002));
    InMux I__23530 (
            .O(N__95417),
            .I(N__94993));
    InMux I__23529 (
            .O(N__95416),
            .I(N__94993));
    InMux I__23528 (
            .O(N__95415),
            .I(N__94993));
    InMux I__23527 (
            .O(N__95414),
            .I(N__94993));
    CascadeMux I__23526 (
            .O(N__95413),
            .I(N__94990));
    CascadeMux I__23525 (
            .O(N__95412),
            .I(N__94987));
    CascadeMux I__23524 (
            .O(N__95411),
            .I(N__94984));
    CascadeMux I__23523 (
            .O(N__95410),
            .I(N__94981));
    InMux I__23522 (
            .O(N__95409),
            .I(N__94975));
    InMux I__23521 (
            .O(N__95408),
            .I(N__94967));
    InMux I__23520 (
            .O(N__95407),
            .I(N__94964));
    InMux I__23519 (
            .O(N__95404),
            .I(N__94957));
    InMux I__23518 (
            .O(N__95403),
            .I(N__94957));
    InMux I__23517 (
            .O(N__95402),
            .I(N__94957));
    InMux I__23516 (
            .O(N__95401),
            .I(N__94944));
    InMux I__23515 (
            .O(N__95400),
            .I(N__94944));
    InMux I__23514 (
            .O(N__95399),
            .I(N__94944));
    InMux I__23513 (
            .O(N__95398),
            .I(N__94944));
    InMux I__23512 (
            .O(N__95397),
            .I(N__94944));
    InMux I__23511 (
            .O(N__95396),
            .I(N__94944));
    InMux I__23510 (
            .O(N__95395),
            .I(N__94931));
    InMux I__23509 (
            .O(N__95394),
            .I(N__94931));
    InMux I__23508 (
            .O(N__95393),
            .I(N__94931));
    InMux I__23507 (
            .O(N__95392),
            .I(N__94931));
    InMux I__23506 (
            .O(N__95391),
            .I(N__94931));
    InMux I__23505 (
            .O(N__95390),
            .I(N__94931));
    InMux I__23504 (
            .O(N__95389),
            .I(N__94920));
    InMux I__23503 (
            .O(N__95388),
            .I(N__94920));
    InMux I__23502 (
            .O(N__95387),
            .I(N__94920));
    InMux I__23501 (
            .O(N__95386),
            .I(N__94920));
    InMux I__23500 (
            .O(N__95385),
            .I(N__94920));
    InMux I__23499 (
            .O(N__95384),
            .I(N__94915));
    InMux I__23498 (
            .O(N__95383),
            .I(N__94915));
    InMux I__23497 (
            .O(N__95382),
            .I(N__94904));
    InMux I__23496 (
            .O(N__95381),
            .I(N__94904));
    InMux I__23495 (
            .O(N__95380),
            .I(N__94904));
    InMux I__23494 (
            .O(N__95379),
            .I(N__94904));
    InMux I__23493 (
            .O(N__95378),
            .I(N__94904));
    InMux I__23492 (
            .O(N__95377),
            .I(N__94899));
    InMux I__23491 (
            .O(N__95376),
            .I(N__94899));
    InMux I__23490 (
            .O(N__95375),
            .I(N__94894));
    InMux I__23489 (
            .O(N__95374),
            .I(N__94894));
    InMux I__23488 (
            .O(N__95373),
            .I(N__94889));
    InMux I__23487 (
            .O(N__95372),
            .I(N__94889));
    InMux I__23486 (
            .O(N__95371),
            .I(N__94878));
    InMux I__23485 (
            .O(N__95370),
            .I(N__94878));
    InMux I__23484 (
            .O(N__95369),
            .I(N__94878));
    InMux I__23483 (
            .O(N__95368),
            .I(N__94878));
    InMux I__23482 (
            .O(N__95367),
            .I(N__94878));
    LocalMux I__23481 (
            .O(N__95364),
            .I(N__94871));
    LocalMux I__23480 (
            .O(N__95359),
            .I(N__94868));
    LocalMux I__23479 (
            .O(N__95356),
            .I(N__94863));
    LocalMux I__23478 (
            .O(N__95349),
            .I(N__94863));
    InMux I__23477 (
            .O(N__95348),
            .I(N__94858));
    InMux I__23476 (
            .O(N__95347),
            .I(N__94858));
    InMux I__23475 (
            .O(N__95346),
            .I(N__94849));
    InMux I__23474 (
            .O(N__95345),
            .I(N__94849));
    InMux I__23473 (
            .O(N__95344),
            .I(N__94849));
    InMux I__23472 (
            .O(N__95343),
            .I(N__94849));
    InMux I__23471 (
            .O(N__95342),
            .I(N__94846));
    InMux I__23470 (
            .O(N__95339),
            .I(N__94835));
    InMux I__23469 (
            .O(N__95338),
            .I(N__94835));
    InMux I__23468 (
            .O(N__95337),
            .I(N__94835));
    InMux I__23467 (
            .O(N__95336),
            .I(N__94835));
    InMux I__23466 (
            .O(N__95335),
            .I(N__94835));
    InMux I__23465 (
            .O(N__95334),
            .I(N__94832));
    InMux I__23464 (
            .O(N__95333),
            .I(N__94819));
    InMux I__23463 (
            .O(N__95330),
            .I(N__94810));
    InMux I__23462 (
            .O(N__95327),
            .I(N__94810));
    InMux I__23461 (
            .O(N__95326),
            .I(N__94810));
    InMux I__23460 (
            .O(N__95325),
            .I(N__94810));
    InMux I__23459 (
            .O(N__95324),
            .I(N__94805));
    InMux I__23458 (
            .O(N__95323),
            .I(N__94805));
    InMux I__23457 (
            .O(N__95322),
            .I(N__94794));
    InMux I__23456 (
            .O(N__95321),
            .I(N__94794));
    InMux I__23455 (
            .O(N__95320),
            .I(N__94794));
    InMux I__23454 (
            .O(N__95319),
            .I(N__94794));
    InMux I__23453 (
            .O(N__95318),
            .I(N__94794));
    InMux I__23452 (
            .O(N__95317),
            .I(N__94785));
    InMux I__23451 (
            .O(N__95316),
            .I(N__94785));
    InMux I__23450 (
            .O(N__95315),
            .I(N__94785));
    InMux I__23449 (
            .O(N__95314),
            .I(N__94785));
    LocalMux I__23448 (
            .O(N__95305),
            .I(N__94780));
    LocalMux I__23447 (
            .O(N__95300),
            .I(N__94780));
    CascadeMux I__23446 (
            .O(N__95299),
            .I(N__94777));
    CascadeMux I__23445 (
            .O(N__95298),
            .I(N__94773));
    InMux I__23444 (
            .O(N__95295),
            .I(N__94760));
    InMux I__23443 (
            .O(N__95294),
            .I(N__94757));
    InMux I__23442 (
            .O(N__95291),
            .I(N__94752));
    InMux I__23441 (
            .O(N__95290),
            .I(N__94752));
    InMux I__23440 (
            .O(N__95289),
            .I(N__94743));
    InMux I__23439 (
            .O(N__95288),
            .I(N__94743));
    InMux I__23438 (
            .O(N__95287),
            .I(N__94743));
    InMux I__23437 (
            .O(N__95286),
            .I(N__94743));
    InMux I__23436 (
            .O(N__95285),
            .I(N__94736));
    InMux I__23435 (
            .O(N__95284),
            .I(N__94736));
    InMux I__23434 (
            .O(N__95283),
            .I(N__94736));
    Span4Mux_v I__23433 (
            .O(N__95276),
            .I(N__94723));
    LocalMux I__23432 (
            .O(N__95273),
            .I(N__94723));
    LocalMux I__23431 (
            .O(N__95262),
            .I(N__94723));
    LocalMux I__23430 (
            .O(N__95259),
            .I(N__94723));
    Span4Mux_h I__23429 (
            .O(N__95254),
            .I(N__94723));
    Span4Mux_h I__23428 (
            .O(N__95249),
            .I(N__94723));
    LocalMux I__23427 (
            .O(N__95238),
            .I(N__94720));
    LocalMux I__23426 (
            .O(N__95225),
            .I(N__94717));
    InMux I__23425 (
            .O(N__95224),
            .I(N__94712));
    InMux I__23424 (
            .O(N__95223),
            .I(N__94712));
    InMux I__23423 (
            .O(N__95222),
            .I(N__94701));
    InMux I__23422 (
            .O(N__95221),
            .I(N__94701));
    InMux I__23421 (
            .O(N__95220),
            .I(N__94701));
    InMux I__23420 (
            .O(N__95219),
            .I(N__94701));
    InMux I__23419 (
            .O(N__95218),
            .I(N__94701));
    LocalMux I__23418 (
            .O(N__95211),
            .I(N__94692));
    LocalMux I__23417 (
            .O(N__95206),
            .I(N__94692));
    LocalMux I__23416 (
            .O(N__95197),
            .I(N__94692));
    LocalMux I__23415 (
            .O(N__95186),
            .I(N__94692));
    LocalMux I__23414 (
            .O(N__95183),
            .I(N__94687));
    Span4Mux_v I__23413 (
            .O(N__95178),
            .I(N__94687));
    CascadeMux I__23412 (
            .O(N__95177),
            .I(N__94682));
    CascadeMux I__23411 (
            .O(N__95176),
            .I(N__94678));
    CascadeMux I__23410 (
            .O(N__95175),
            .I(N__94675));
    CascadeMux I__23409 (
            .O(N__95174),
            .I(N__94672));
    InMux I__23408 (
            .O(N__95173),
            .I(N__94657));
    LocalMux I__23407 (
            .O(N__95166),
            .I(N__94654));
    LocalMux I__23406 (
            .O(N__95157),
            .I(N__94651));
    InMux I__23405 (
            .O(N__95156),
            .I(N__94648));
    InMux I__23404 (
            .O(N__95155),
            .I(N__94645));
    InMux I__23403 (
            .O(N__95154),
            .I(N__94636));
    InMux I__23402 (
            .O(N__95153),
            .I(N__94636));
    InMux I__23401 (
            .O(N__95152),
            .I(N__94636));
    InMux I__23400 (
            .O(N__95151),
            .I(N__94636));
    InMux I__23399 (
            .O(N__95150),
            .I(N__94633));
    InMux I__23398 (
            .O(N__95149),
            .I(N__94624));
    InMux I__23397 (
            .O(N__95148),
            .I(N__94624));
    InMux I__23396 (
            .O(N__95147),
            .I(N__94624));
    InMux I__23395 (
            .O(N__95146),
            .I(N__94624));
    LocalMux I__23394 (
            .O(N__95139),
            .I(N__94613));
    Span4Mux_h I__23393 (
            .O(N__95132),
            .I(N__94613));
    Span4Mux_h I__23392 (
            .O(N__95127),
            .I(N__94613));
    LocalMux I__23391 (
            .O(N__95122),
            .I(N__94613));
    LocalMux I__23390 (
            .O(N__95119),
            .I(N__94613));
    LocalMux I__23389 (
            .O(N__95106),
            .I(N__94610));
    InMux I__23388 (
            .O(N__95105),
            .I(N__94605));
    InMux I__23387 (
            .O(N__95104),
            .I(N__94605));
    InMux I__23386 (
            .O(N__95103),
            .I(N__94585));
    InMux I__23385 (
            .O(N__95102),
            .I(N__94585));
    InMux I__23384 (
            .O(N__95101),
            .I(N__94574));
    InMux I__23383 (
            .O(N__95100),
            .I(N__94565));
    InMux I__23382 (
            .O(N__95099),
            .I(N__94565));
    InMux I__23381 (
            .O(N__95098),
            .I(N__94565));
    InMux I__23380 (
            .O(N__95097),
            .I(N__94565));
    InMux I__23379 (
            .O(N__95096),
            .I(N__94556));
    InMux I__23378 (
            .O(N__95095),
            .I(N__94556));
    InMux I__23377 (
            .O(N__95094),
            .I(N__94556));
    InMux I__23376 (
            .O(N__95093),
            .I(N__94556));
    InMux I__23375 (
            .O(N__95092),
            .I(N__94553));
    InMux I__23374 (
            .O(N__95091),
            .I(N__94542));
    InMux I__23373 (
            .O(N__95090),
            .I(N__94542));
    InMux I__23372 (
            .O(N__95089),
            .I(N__94542));
    InMux I__23371 (
            .O(N__95088),
            .I(N__94542));
    InMux I__23370 (
            .O(N__95087),
            .I(N__94542));
    InMux I__23369 (
            .O(N__95084),
            .I(N__94531));
    InMux I__23368 (
            .O(N__95081),
            .I(N__94531));
    InMux I__23367 (
            .O(N__95080),
            .I(N__94531));
    InMux I__23366 (
            .O(N__95079),
            .I(N__94531));
    InMux I__23365 (
            .O(N__95078),
            .I(N__94531));
    InMux I__23364 (
            .O(N__95077),
            .I(N__94524));
    InMux I__23363 (
            .O(N__95076),
            .I(N__94524));
    InMux I__23362 (
            .O(N__95075),
            .I(N__94524));
    LocalMux I__23361 (
            .O(N__95070),
            .I(N__94521));
    LocalMux I__23360 (
            .O(N__95067),
            .I(N__94516));
    LocalMux I__23359 (
            .O(N__95058),
            .I(N__94516));
    LocalMux I__23358 (
            .O(N__95055),
            .I(N__94513));
    InMux I__23357 (
            .O(N__95054),
            .I(N__94510));
    InMux I__23356 (
            .O(N__95053),
            .I(N__94505));
    InMux I__23355 (
            .O(N__95052),
            .I(N__94505));
    InMux I__23354 (
            .O(N__95051),
            .I(N__94496));
    InMux I__23353 (
            .O(N__95050),
            .I(N__94496));
    InMux I__23352 (
            .O(N__95049),
            .I(N__94496));
    InMux I__23351 (
            .O(N__95048),
            .I(N__94496));
    LocalMux I__23350 (
            .O(N__95039),
            .I(N__94493));
    Span4Mux_v I__23349 (
            .O(N__95030),
            .I(N__94486));
    LocalMux I__23348 (
            .O(N__95019),
            .I(N__94486));
    LocalMux I__23347 (
            .O(N__95010),
            .I(N__94486));
    CascadeMux I__23346 (
            .O(N__95009),
            .I(N__94477));
    CascadeMux I__23345 (
            .O(N__95008),
            .I(N__94474));
    InMux I__23344 (
            .O(N__95007),
            .I(N__94464));
    InMux I__23343 (
            .O(N__95006),
            .I(N__94464));
    InMux I__23342 (
            .O(N__95005),
            .I(N__94464));
    LocalMux I__23341 (
            .O(N__95002),
            .I(N__94459));
    LocalMux I__23340 (
            .O(N__94993),
            .I(N__94459));
    InMux I__23339 (
            .O(N__94990),
            .I(N__94441));
    InMux I__23338 (
            .O(N__94987),
            .I(N__94441));
    InMux I__23337 (
            .O(N__94984),
            .I(N__94441));
    InMux I__23336 (
            .O(N__94981),
            .I(N__94441));
    InMux I__23335 (
            .O(N__94980),
            .I(N__94441));
    InMux I__23334 (
            .O(N__94979),
            .I(N__94441));
    InMux I__23333 (
            .O(N__94978),
            .I(N__94441));
    LocalMux I__23332 (
            .O(N__94975),
            .I(N__94438));
    InMux I__23331 (
            .O(N__94974),
            .I(N__94433));
    InMux I__23330 (
            .O(N__94973),
            .I(N__94433));
    InMux I__23329 (
            .O(N__94972),
            .I(N__94426));
    InMux I__23328 (
            .O(N__94971),
            .I(N__94426));
    InMux I__23327 (
            .O(N__94970),
            .I(N__94426));
    LocalMux I__23326 (
            .O(N__94967),
            .I(N__94411));
    LocalMux I__23325 (
            .O(N__94964),
            .I(N__94411));
    LocalMux I__23324 (
            .O(N__94957),
            .I(N__94411));
    LocalMux I__23323 (
            .O(N__94944),
            .I(N__94411));
    LocalMux I__23322 (
            .O(N__94931),
            .I(N__94411));
    LocalMux I__23321 (
            .O(N__94920),
            .I(N__94411));
    LocalMux I__23320 (
            .O(N__94915),
            .I(N__94411));
    LocalMux I__23319 (
            .O(N__94904),
            .I(N__94406));
    LocalMux I__23318 (
            .O(N__94899),
            .I(N__94406));
    LocalMux I__23317 (
            .O(N__94894),
            .I(N__94399));
    LocalMux I__23316 (
            .O(N__94889),
            .I(N__94399));
    LocalMux I__23315 (
            .O(N__94878),
            .I(N__94399));
    InMux I__23314 (
            .O(N__94877),
            .I(N__94396));
    InMux I__23313 (
            .O(N__94876),
            .I(N__94393));
    InMux I__23312 (
            .O(N__94875),
            .I(N__94390));
    InMux I__23311 (
            .O(N__94874),
            .I(N__94387));
    Span4Mux_v I__23310 (
            .O(N__94871),
            .I(N__94376));
    Span4Mux_h I__23309 (
            .O(N__94868),
            .I(N__94376));
    Span4Mux_v I__23308 (
            .O(N__94863),
            .I(N__94376));
    LocalMux I__23307 (
            .O(N__94858),
            .I(N__94376));
    LocalMux I__23306 (
            .O(N__94849),
            .I(N__94376));
    LocalMux I__23305 (
            .O(N__94846),
            .I(N__94369));
    LocalMux I__23304 (
            .O(N__94835),
            .I(N__94369));
    LocalMux I__23303 (
            .O(N__94832),
            .I(N__94369));
    InMux I__23302 (
            .O(N__94831),
            .I(N__94364));
    InMux I__23301 (
            .O(N__94830),
            .I(N__94364));
    InMux I__23300 (
            .O(N__94829),
            .I(N__94359));
    InMux I__23299 (
            .O(N__94828),
            .I(N__94359));
    InMux I__23298 (
            .O(N__94827),
            .I(N__94354));
    InMux I__23297 (
            .O(N__94826),
            .I(N__94354));
    InMux I__23296 (
            .O(N__94825),
            .I(N__94351));
    InMux I__23295 (
            .O(N__94824),
            .I(N__94344));
    InMux I__23294 (
            .O(N__94823),
            .I(N__94344));
    InMux I__23293 (
            .O(N__94822),
            .I(N__94344));
    LocalMux I__23292 (
            .O(N__94819),
            .I(N__94337));
    LocalMux I__23291 (
            .O(N__94810),
            .I(N__94337));
    LocalMux I__23290 (
            .O(N__94805),
            .I(N__94337));
    LocalMux I__23289 (
            .O(N__94794),
            .I(N__94330));
    LocalMux I__23288 (
            .O(N__94785),
            .I(N__94330));
    Span4Mux_v I__23287 (
            .O(N__94780),
            .I(N__94330));
    InMux I__23286 (
            .O(N__94777),
            .I(N__94325));
    InMux I__23285 (
            .O(N__94776),
            .I(N__94318));
    InMux I__23284 (
            .O(N__94773),
            .I(N__94318));
    InMux I__23283 (
            .O(N__94772),
            .I(N__94318));
    InMux I__23282 (
            .O(N__94771),
            .I(N__94315));
    InMux I__23281 (
            .O(N__94770),
            .I(N__94308));
    InMux I__23280 (
            .O(N__94769),
            .I(N__94308));
    InMux I__23279 (
            .O(N__94768),
            .I(N__94308));
    InMux I__23278 (
            .O(N__94767),
            .I(N__94297));
    InMux I__23277 (
            .O(N__94766),
            .I(N__94297));
    InMux I__23276 (
            .O(N__94765),
            .I(N__94297));
    InMux I__23275 (
            .O(N__94764),
            .I(N__94297));
    InMux I__23274 (
            .O(N__94763),
            .I(N__94297));
    LocalMux I__23273 (
            .O(N__94760),
            .I(N__94279));
    LocalMux I__23272 (
            .O(N__94757),
            .I(N__94279));
    LocalMux I__23271 (
            .O(N__94752),
            .I(N__94279));
    LocalMux I__23270 (
            .O(N__94743),
            .I(N__94279));
    LocalMux I__23269 (
            .O(N__94736),
            .I(N__94279));
    Span4Mux_h I__23268 (
            .O(N__94723),
            .I(N__94279));
    Span4Mux_v I__23267 (
            .O(N__94720),
            .I(N__94279));
    Span4Mux_v I__23266 (
            .O(N__94717),
            .I(N__94279));
    LocalMux I__23265 (
            .O(N__94712),
            .I(N__94270));
    LocalMux I__23264 (
            .O(N__94701),
            .I(N__94270));
    Span4Mux_v I__23263 (
            .O(N__94692),
            .I(N__94270));
    Span4Mux_h I__23262 (
            .O(N__94687),
            .I(N__94270));
    InMux I__23261 (
            .O(N__94686),
            .I(N__94259));
    InMux I__23260 (
            .O(N__94685),
            .I(N__94259));
    InMux I__23259 (
            .O(N__94682),
            .I(N__94259));
    InMux I__23258 (
            .O(N__94681),
            .I(N__94259));
    InMux I__23257 (
            .O(N__94678),
            .I(N__94259));
    InMux I__23256 (
            .O(N__94675),
            .I(N__94252));
    InMux I__23255 (
            .O(N__94672),
            .I(N__94252));
    InMux I__23254 (
            .O(N__94671),
            .I(N__94252));
    InMux I__23253 (
            .O(N__94670),
            .I(N__94245));
    InMux I__23252 (
            .O(N__94669),
            .I(N__94245));
    InMux I__23251 (
            .O(N__94668),
            .I(N__94245));
    InMux I__23250 (
            .O(N__94667),
            .I(N__94224));
    InMux I__23249 (
            .O(N__94666),
            .I(N__94224));
    InMux I__23248 (
            .O(N__94665),
            .I(N__94224));
    InMux I__23247 (
            .O(N__94664),
            .I(N__94224));
    InMux I__23246 (
            .O(N__94663),
            .I(N__94212));
    InMux I__23245 (
            .O(N__94662),
            .I(N__94212));
    InMux I__23244 (
            .O(N__94661),
            .I(N__94212));
    InMux I__23243 (
            .O(N__94660),
            .I(N__94212));
    LocalMux I__23242 (
            .O(N__94657),
            .I(N__94203));
    Span4Mux_v I__23241 (
            .O(N__94654),
            .I(N__94203));
    Span4Mux_h I__23240 (
            .O(N__94651),
            .I(N__94203));
    LocalMux I__23239 (
            .O(N__94648),
            .I(N__94203));
    LocalMux I__23238 (
            .O(N__94645),
            .I(N__94192));
    LocalMux I__23237 (
            .O(N__94636),
            .I(N__94192));
    LocalMux I__23236 (
            .O(N__94633),
            .I(N__94192));
    LocalMux I__23235 (
            .O(N__94624),
            .I(N__94192));
    Span4Mux_h I__23234 (
            .O(N__94613),
            .I(N__94192));
    Span4Mux_v I__23233 (
            .O(N__94610),
            .I(N__94187));
    LocalMux I__23232 (
            .O(N__94605),
            .I(N__94187));
    InMux I__23231 (
            .O(N__94604),
            .I(N__94182));
    InMux I__23230 (
            .O(N__94603),
            .I(N__94182));
    CascadeMux I__23229 (
            .O(N__94602),
            .I(N__94173));
    InMux I__23228 (
            .O(N__94601),
            .I(N__94163));
    InMux I__23227 (
            .O(N__94600),
            .I(N__94163));
    CascadeMux I__23226 (
            .O(N__94599),
            .I(N__94157));
    CascadeMux I__23225 (
            .O(N__94598),
            .I(N__94154));
    CascadeMux I__23224 (
            .O(N__94597),
            .I(N__94151));
    CascadeMux I__23223 (
            .O(N__94596),
            .I(N__94146));
    CascadeMux I__23222 (
            .O(N__94595),
            .I(N__94143));
    InMux I__23221 (
            .O(N__94594),
            .I(N__94132));
    InMux I__23220 (
            .O(N__94593),
            .I(N__94132));
    InMux I__23219 (
            .O(N__94592),
            .I(N__94132));
    InMux I__23218 (
            .O(N__94591),
            .I(N__94129));
    CascadeMux I__23217 (
            .O(N__94590),
            .I(N__94126));
    LocalMux I__23216 (
            .O(N__94585),
            .I(N__94123));
    InMux I__23215 (
            .O(N__94584),
            .I(N__94109));
    InMux I__23214 (
            .O(N__94583),
            .I(N__94109));
    InMux I__23213 (
            .O(N__94582),
            .I(N__94109));
    InMux I__23212 (
            .O(N__94581),
            .I(N__94109));
    InMux I__23211 (
            .O(N__94580),
            .I(N__94109));
    InMux I__23210 (
            .O(N__94579),
            .I(N__94104));
    InMux I__23209 (
            .O(N__94578),
            .I(N__94104));
    InMux I__23208 (
            .O(N__94577),
            .I(N__94097));
    LocalMux I__23207 (
            .O(N__94574),
            .I(N__94090));
    LocalMux I__23206 (
            .O(N__94565),
            .I(N__94090));
    LocalMux I__23205 (
            .O(N__94556),
            .I(N__94090));
    LocalMux I__23204 (
            .O(N__94553),
            .I(N__94085));
    LocalMux I__23203 (
            .O(N__94542),
            .I(N__94085));
    LocalMux I__23202 (
            .O(N__94531),
            .I(N__94074));
    LocalMux I__23201 (
            .O(N__94524),
            .I(N__94074));
    Span4Mux_v I__23200 (
            .O(N__94521),
            .I(N__94074));
    Span4Mux_v I__23199 (
            .O(N__94516),
            .I(N__94074));
    Span4Mux_v I__23198 (
            .O(N__94513),
            .I(N__94074));
    LocalMux I__23197 (
            .O(N__94510),
            .I(N__94069));
    LocalMux I__23196 (
            .O(N__94505),
            .I(N__94069));
    LocalMux I__23195 (
            .O(N__94496),
            .I(N__94062));
    Span4Mux_v I__23194 (
            .O(N__94493),
            .I(N__94062));
    Span4Mux_v I__23193 (
            .O(N__94486),
            .I(N__94062));
    InMux I__23192 (
            .O(N__94485),
            .I(N__94055));
    InMux I__23191 (
            .O(N__94484),
            .I(N__94055));
    InMux I__23190 (
            .O(N__94483),
            .I(N__94055));
    CascadeMux I__23189 (
            .O(N__94482),
            .I(N__94052));
    CascadeMux I__23188 (
            .O(N__94481),
            .I(N__94045));
    CascadeMux I__23187 (
            .O(N__94480),
            .I(N__94042));
    InMux I__23186 (
            .O(N__94477),
            .I(N__94037));
    InMux I__23185 (
            .O(N__94474),
            .I(N__94037));
    InMux I__23184 (
            .O(N__94473),
            .I(N__94034));
    InMux I__23183 (
            .O(N__94472),
            .I(N__94029));
    InMux I__23182 (
            .O(N__94471),
            .I(N__94029));
    LocalMux I__23181 (
            .O(N__94464),
            .I(N__94024));
    Span4Mux_v I__23180 (
            .O(N__94459),
            .I(N__94024));
    InMux I__23179 (
            .O(N__94458),
            .I(N__94021));
    InMux I__23178 (
            .O(N__94457),
            .I(N__94016));
    InMux I__23177 (
            .O(N__94456),
            .I(N__94016));
    LocalMux I__23176 (
            .O(N__94441),
            .I(N__94013));
    Span4Mux_v I__23175 (
            .O(N__94438),
            .I(N__94010));
    LocalMux I__23174 (
            .O(N__94433),
            .I(N__93999));
    LocalMux I__23173 (
            .O(N__94426),
            .I(N__93999));
    Span4Mux_v I__23172 (
            .O(N__94411),
            .I(N__93999));
    Span4Mux_v I__23171 (
            .O(N__94406),
            .I(N__93999));
    Span4Mux_v I__23170 (
            .O(N__94399),
            .I(N__93999));
    LocalMux I__23169 (
            .O(N__94396),
            .I(N__93990));
    LocalMux I__23168 (
            .O(N__94393),
            .I(N__93990));
    LocalMux I__23167 (
            .O(N__94390),
            .I(N__93990));
    LocalMux I__23166 (
            .O(N__94387),
            .I(N__93990));
    Span4Mux_v I__23165 (
            .O(N__94376),
            .I(N__93983));
    Span4Mux_v I__23164 (
            .O(N__94369),
            .I(N__93983));
    LocalMux I__23163 (
            .O(N__94364),
            .I(N__93983));
    LocalMux I__23162 (
            .O(N__94359),
            .I(N__93972));
    LocalMux I__23161 (
            .O(N__94354),
            .I(N__93972));
    LocalMux I__23160 (
            .O(N__94351),
            .I(N__93972));
    LocalMux I__23159 (
            .O(N__94344),
            .I(N__93972));
    Span4Mux_v I__23158 (
            .O(N__94337),
            .I(N__93972));
    Span4Mux_v I__23157 (
            .O(N__94330),
            .I(N__93969));
    InMux I__23156 (
            .O(N__94329),
            .I(N__93961));
    InMux I__23155 (
            .O(N__94328),
            .I(N__93958));
    LocalMux I__23154 (
            .O(N__94325),
            .I(N__93947));
    LocalMux I__23153 (
            .O(N__94318),
            .I(N__93947));
    LocalMux I__23152 (
            .O(N__94315),
            .I(N__93947));
    LocalMux I__23151 (
            .O(N__94308),
            .I(N__93947));
    LocalMux I__23150 (
            .O(N__94297),
            .I(N__93947));
    InMux I__23149 (
            .O(N__94296),
            .I(N__93944));
    Span4Mux_v I__23148 (
            .O(N__94279),
            .I(N__93933));
    Span4Mux_h I__23147 (
            .O(N__94270),
            .I(N__93933));
    LocalMux I__23146 (
            .O(N__94259),
            .I(N__93933));
    LocalMux I__23145 (
            .O(N__94252),
            .I(N__93933));
    LocalMux I__23144 (
            .O(N__94245),
            .I(N__93933));
    InMux I__23143 (
            .O(N__94244),
            .I(N__93920));
    InMux I__23142 (
            .O(N__94243),
            .I(N__93909));
    InMux I__23141 (
            .O(N__94242),
            .I(N__93909));
    InMux I__23140 (
            .O(N__94241),
            .I(N__93909));
    InMux I__23139 (
            .O(N__94240),
            .I(N__93909));
    InMux I__23138 (
            .O(N__94239),
            .I(N__93909));
    InMux I__23137 (
            .O(N__94238),
            .I(N__93906));
    InMux I__23136 (
            .O(N__94237),
            .I(N__93899));
    InMux I__23135 (
            .O(N__94236),
            .I(N__93899));
    InMux I__23134 (
            .O(N__94235),
            .I(N__93899));
    InMux I__23133 (
            .O(N__94234),
            .I(N__93894));
    InMux I__23132 (
            .O(N__94233),
            .I(N__93894));
    LocalMux I__23131 (
            .O(N__94224),
            .I(N__93891));
    InMux I__23130 (
            .O(N__94223),
            .I(N__93886));
    InMux I__23129 (
            .O(N__94222),
            .I(N__93886));
    InMux I__23128 (
            .O(N__94221),
            .I(N__93883));
    LocalMux I__23127 (
            .O(N__94212),
            .I(N__93872));
    Span4Mux_h I__23126 (
            .O(N__94203),
            .I(N__93872));
    Span4Mux_v I__23125 (
            .O(N__94192),
            .I(N__93872));
    Span4Mux_h I__23124 (
            .O(N__94187),
            .I(N__93872));
    LocalMux I__23123 (
            .O(N__94182),
            .I(N__93872));
    InMux I__23122 (
            .O(N__94181),
            .I(N__93865));
    InMux I__23121 (
            .O(N__94180),
            .I(N__93865));
    InMux I__23120 (
            .O(N__94179),
            .I(N__93865));
    InMux I__23119 (
            .O(N__94178),
            .I(N__93858));
    InMux I__23118 (
            .O(N__94177),
            .I(N__93858));
    InMux I__23117 (
            .O(N__94176),
            .I(N__93858));
    InMux I__23116 (
            .O(N__94173),
            .I(N__93845));
    InMux I__23115 (
            .O(N__94172),
            .I(N__93845));
    InMux I__23114 (
            .O(N__94171),
            .I(N__93845));
    InMux I__23113 (
            .O(N__94170),
            .I(N__93845));
    InMux I__23112 (
            .O(N__94169),
            .I(N__93845));
    InMux I__23111 (
            .O(N__94168),
            .I(N__93845));
    LocalMux I__23110 (
            .O(N__94163),
            .I(N__93842));
    InMux I__23109 (
            .O(N__94162),
            .I(N__93829));
    InMux I__23108 (
            .O(N__94161),
            .I(N__93829));
    InMux I__23107 (
            .O(N__94160),
            .I(N__93829));
    InMux I__23106 (
            .O(N__94157),
            .I(N__93829));
    InMux I__23105 (
            .O(N__94154),
            .I(N__93829));
    InMux I__23104 (
            .O(N__94151),
            .I(N__93829));
    InMux I__23103 (
            .O(N__94150),
            .I(N__93816));
    InMux I__23102 (
            .O(N__94149),
            .I(N__93816));
    InMux I__23101 (
            .O(N__94146),
            .I(N__93816));
    InMux I__23100 (
            .O(N__94143),
            .I(N__93816));
    InMux I__23099 (
            .O(N__94142),
            .I(N__93816));
    InMux I__23098 (
            .O(N__94141),
            .I(N__93816));
    CascadeMux I__23097 (
            .O(N__94140),
            .I(N__93812));
    InMux I__23096 (
            .O(N__94139),
            .I(N__93801));
    LocalMux I__23095 (
            .O(N__94132),
            .I(N__93798));
    LocalMux I__23094 (
            .O(N__94129),
            .I(N__93795));
    InMux I__23093 (
            .O(N__94126),
            .I(N__93792));
    Span4Mux_v I__23092 (
            .O(N__94123),
            .I(N__93789));
    InMux I__23091 (
            .O(N__94122),
            .I(N__93782));
    InMux I__23090 (
            .O(N__94121),
            .I(N__93782));
    InMux I__23089 (
            .O(N__94120),
            .I(N__93782));
    LocalMux I__23088 (
            .O(N__94109),
            .I(N__93777));
    LocalMux I__23087 (
            .O(N__94104),
            .I(N__93777));
    CascadeMux I__23086 (
            .O(N__94103),
            .I(N__93774));
    CascadeMux I__23085 (
            .O(N__94102),
            .I(N__93765));
    InMux I__23084 (
            .O(N__94101),
            .I(N__93760));
    InMux I__23083 (
            .O(N__94100),
            .I(N__93760));
    LocalMux I__23082 (
            .O(N__94097),
            .I(N__93753));
    Span4Mux_v I__23081 (
            .O(N__94090),
            .I(N__93753));
    Span4Mux_v I__23080 (
            .O(N__94085),
            .I(N__93753));
    Span4Mux_v I__23079 (
            .O(N__94074),
            .I(N__93744));
    Span4Mux_v I__23078 (
            .O(N__94069),
            .I(N__93744));
    Span4Mux_h I__23077 (
            .O(N__94062),
            .I(N__93744));
    LocalMux I__23076 (
            .O(N__94055),
            .I(N__93744));
    InMux I__23075 (
            .O(N__94052),
            .I(N__93729));
    InMux I__23074 (
            .O(N__94051),
            .I(N__93729));
    InMux I__23073 (
            .O(N__94050),
            .I(N__93729));
    InMux I__23072 (
            .O(N__94049),
            .I(N__93729));
    InMux I__23071 (
            .O(N__94048),
            .I(N__93729));
    InMux I__23070 (
            .O(N__94045),
            .I(N__93729));
    InMux I__23069 (
            .O(N__94042),
            .I(N__93729));
    LocalMux I__23068 (
            .O(N__94037),
            .I(N__93722));
    LocalMux I__23067 (
            .O(N__94034),
            .I(N__93722));
    LocalMux I__23066 (
            .O(N__94029),
            .I(N__93722));
    Span4Mux_v I__23065 (
            .O(N__94024),
            .I(N__93717));
    LocalMux I__23064 (
            .O(N__94021),
            .I(N__93717));
    LocalMux I__23063 (
            .O(N__94016),
            .I(N__93704));
    Span4Mux_v I__23062 (
            .O(N__94013),
            .I(N__93704));
    Span4Mux_h I__23061 (
            .O(N__94010),
            .I(N__93704));
    Span4Mux_h I__23060 (
            .O(N__93999),
            .I(N__93704));
    Span4Mux_v I__23059 (
            .O(N__93990),
            .I(N__93704));
    Span4Mux_v I__23058 (
            .O(N__93983),
            .I(N__93704));
    Span4Mux_v I__23057 (
            .O(N__93972),
            .I(N__93699));
    Span4Mux_h I__23056 (
            .O(N__93969),
            .I(N__93699));
    InMux I__23055 (
            .O(N__93968),
            .I(N__93696));
    InMux I__23054 (
            .O(N__93967),
            .I(N__93687));
    InMux I__23053 (
            .O(N__93966),
            .I(N__93687));
    InMux I__23052 (
            .O(N__93965),
            .I(N__93687));
    InMux I__23051 (
            .O(N__93964),
            .I(N__93687));
    LocalMux I__23050 (
            .O(N__93961),
            .I(N__93676));
    LocalMux I__23049 (
            .O(N__93958),
            .I(N__93676));
    Span4Mux_v I__23048 (
            .O(N__93947),
            .I(N__93676));
    LocalMux I__23047 (
            .O(N__93944),
            .I(N__93676));
    Span4Mux_v I__23046 (
            .O(N__93933),
            .I(N__93676));
    InMux I__23045 (
            .O(N__93932),
            .I(N__93665));
    InMux I__23044 (
            .O(N__93931),
            .I(N__93665));
    InMux I__23043 (
            .O(N__93930),
            .I(N__93665));
    InMux I__23042 (
            .O(N__93929),
            .I(N__93665));
    InMux I__23041 (
            .O(N__93928),
            .I(N__93665));
    InMux I__23040 (
            .O(N__93927),
            .I(N__93654));
    InMux I__23039 (
            .O(N__93926),
            .I(N__93654));
    InMux I__23038 (
            .O(N__93925),
            .I(N__93654));
    InMux I__23037 (
            .O(N__93924),
            .I(N__93654));
    InMux I__23036 (
            .O(N__93923),
            .I(N__93654));
    LocalMux I__23035 (
            .O(N__93920),
            .I(N__93643));
    LocalMux I__23034 (
            .O(N__93909),
            .I(N__93643));
    LocalMux I__23033 (
            .O(N__93906),
            .I(N__93643));
    LocalMux I__23032 (
            .O(N__93899),
            .I(N__93643));
    LocalMux I__23031 (
            .O(N__93894),
            .I(N__93643));
    Sp12to4 I__23030 (
            .O(N__93891),
            .I(N__93638));
    LocalMux I__23029 (
            .O(N__93886),
            .I(N__93638));
    LocalMux I__23028 (
            .O(N__93883),
            .I(N__93635));
    Sp12to4 I__23027 (
            .O(N__93872),
            .I(N__93632));
    LocalMux I__23026 (
            .O(N__93865),
            .I(N__93619));
    LocalMux I__23025 (
            .O(N__93858),
            .I(N__93619));
    LocalMux I__23024 (
            .O(N__93845),
            .I(N__93619));
    Sp12to4 I__23023 (
            .O(N__93842),
            .I(N__93619));
    LocalMux I__23022 (
            .O(N__93829),
            .I(N__93619));
    LocalMux I__23021 (
            .O(N__93816),
            .I(N__93619));
    InMux I__23020 (
            .O(N__93815),
            .I(N__93615));
    InMux I__23019 (
            .O(N__93812),
            .I(N__93608));
    InMux I__23018 (
            .O(N__93811),
            .I(N__93608));
    InMux I__23017 (
            .O(N__93810),
            .I(N__93608));
    InMux I__23016 (
            .O(N__93809),
            .I(N__93599));
    InMux I__23015 (
            .O(N__93808),
            .I(N__93599));
    InMux I__23014 (
            .O(N__93807),
            .I(N__93599));
    InMux I__23013 (
            .O(N__93806),
            .I(N__93599));
    InMux I__23012 (
            .O(N__93805),
            .I(N__93594));
    InMux I__23011 (
            .O(N__93804),
            .I(N__93594));
    LocalMux I__23010 (
            .O(N__93801),
            .I(N__93591));
    Span4Mux_h I__23009 (
            .O(N__93798),
            .I(N__93588));
    Span4Mux_v I__23008 (
            .O(N__93795),
            .I(N__93585));
    LocalMux I__23007 (
            .O(N__93792),
            .I(N__93580));
    Span4Mux_h I__23006 (
            .O(N__93789),
            .I(N__93580));
    LocalMux I__23005 (
            .O(N__93782),
            .I(N__93575));
    Span4Mux_v I__23004 (
            .O(N__93777),
            .I(N__93575));
    InMux I__23003 (
            .O(N__93774),
            .I(N__93564));
    InMux I__23002 (
            .O(N__93773),
            .I(N__93564));
    InMux I__23001 (
            .O(N__93772),
            .I(N__93564));
    InMux I__23000 (
            .O(N__93771),
            .I(N__93564));
    InMux I__22999 (
            .O(N__93770),
            .I(N__93564));
    InMux I__22998 (
            .O(N__93769),
            .I(N__93559));
    InMux I__22997 (
            .O(N__93768),
            .I(N__93559));
    InMux I__22996 (
            .O(N__93765),
            .I(N__93556));
    LocalMux I__22995 (
            .O(N__93760),
            .I(N__93547));
    Span4Mux_h I__22994 (
            .O(N__93753),
            .I(N__93547));
    Span4Mux_h I__22993 (
            .O(N__93744),
            .I(N__93547));
    LocalMux I__22992 (
            .O(N__93729),
            .I(N__93547));
    Span4Mux_v I__22991 (
            .O(N__93722),
            .I(N__93532));
    Span4Mux_v I__22990 (
            .O(N__93717),
            .I(N__93532));
    Span4Mux_h I__22989 (
            .O(N__93704),
            .I(N__93532));
    Span4Mux_h I__22988 (
            .O(N__93699),
            .I(N__93532));
    LocalMux I__22987 (
            .O(N__93696),
            .I(N__93532));
    LocalMux I__22986 (
            .O(N__93687),
            .I(N__93532));
    Span4Mux_v I__22985 (
            .O(N__93676),
            .I(N__93532));
    LocalMux I__22984 (
            .O(N__93665),
            .I(N__93517));
    LocalMux I__22983 (
            .O(N__93654),
            .I(N__93517));
    Span12Mux_v I__22982 (
            .O(N__93643),
            .I(N__93517));
    Span12Mux_v I__22981 (
            .O(N__93638),
            .I(N__93517));
    Span12Mux_s11_h I__22980 (
            .O(N__93635),
            .I(N__93517));
    Span12Mux_v I__22979 (
            .O(N__93632),
            .I(N__93517));
    Span12Mux_v I__22978 (
            .O(N__93619),
            .I(N__93517));
    InMux I__22977 (
            .O(N__93618),
            .I(N__93514));
    LocalMux I__22976 (
            .O(N__93615),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    LocalMux I__22975 (
            .O(N__93608),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    LocalMux I__22974 (
            .O(N__93599),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    LocalMux I__22973 (
            .O(N__93594),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    Odrv12 I__22972 (
            .O(N__93591),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    Odrv4 I__22971 (
            .O(N__93588),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    Odrv4 I__22970 (
            .O(N__93585),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    Odrv4 I__22969 (
            .O(N__93580),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    Odrv4 I__22968 (
            .O(N__93575),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    LocalMux I__22967 (
            .O(N__93564),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    LocalMux I__22966 (
            .O(N__93559),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    LocalMux I__22965 (
            .O(N__93556),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    Odrv4 I__22964 (
            .O(N__93547),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    Odrv4 I__22963 (
            .O(N__93532),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    Odrv12 I__22962 (
            .O(N__93517),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    LocalMux I__22961 (
            .O(N__93514),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ));
    InMux I__22960 (
            .O(N__93481),
            .I(N__93478));
    LocalMux I__22959 (
            .O(N__93478),
            .I(N__93474));
    CascadeMux I__22958 (
            .O(N__93477),
            .I(N__93471));
    Span4Mux_h I__22957 (
            .O(N__93474),
            .I(N__93468));
    InMux I__22956 (
            .O(N__93471),
            .I(N__93465));
    Odrv4 I__22955 (
            .O(N__93468),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_6 ));
    LocalMux I__22954 (
            .O(N__93465),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_6 ));
    InMux I__22953 (
            .O(N__93460),
            .I(N__93457));
    LocalMux I__22952 (
            .O(N__93457),
            .I(N__93443));
    ClkMux I__22951 (
            .O(N__93456),
            .I(N__92746));
    ClkMux I__22950 (
            .O(N__93455),
            .I(N__92746));
    ClkMux I__22949 (
            .O(N__93454),
            .I(N__92746));
    ClkMux I__22948 (
            .O(N__93453),
            .I(N__92746));
    ClkMux I__22947 (
            .O(N__93452),
            .I(N__92746));
    ClkMux I__22946 (
            .O(N__93451),
            .I(N__92746));
    ClkMux I__22945 (
            .O(N__93450),
            .I(N__92746));
    ClkMux I__22944 (
            .O(N__93449),
            .I(N__92746));
    ClkMux I__22943 (
            .O(N__93448),
            .I(N__92746));
    ClkMux I__22942 (
            .O(N__93447),
            .I(N__92746));
    ClkMux I__22941 (
            .O(N__93446),
            .I(N__92746));
    Glb2LocalMux I__22940 (
            .O(N__93443),
            .I(N__92746));
    ClkMux I__22939 (
            .O(N__93442),
            .I(N__92746));
    ClkMux I__22938 (
            .O(N__93441),
            .I(N__92746));
    ClkMux I__22937 (
            .O(N__93440),
            .I(N__92746));
    ClkMux I__22936 (
            .O(N__93439),
            .I(N__92746));
    ClkMux I__22935 (
            .O(N__93438),
            .I(N__92746));
    ClkMux I__22934 (
            .O(N__93437),
            .I(N__92746));
    ClkMux I__22933 (
            .O(N__93436),
            .I(N__92746));
    ClkMux I__22932 (
            .O(N__93435),
            .I(N__92746));
    ClkMux I__22931 (
            .O(N__93434),
            .I(N__92746));
    ClkMux I__22930 (
            .O(N__93433),
            .I(N__92746));
    ClkMux I__22929 (
            .O(N__93432),
            .I(N__92746));
    ClkMux I__22928 (
            .O(N__93431),
            .I(N__92746));
    ClkMux I__22927 (
            .O(N__93430),
            .I(N__92746));
    ClkMux I__22926 (
            .O(N__93429),
            .I(N__92746));
    ClkMux I__22925 (
            .O(N__93428),
            .I(N__92746));
    ClkMux I__22924 (
            .O(N__93427),
            .I(N__92746));
    ClkMux I__22923 (
            .O(N__93426),
            .I(N__92746));
    ClkMux I__22922 (
            .O(N__93425),
            .I(N__92746));
    ClkMux I__22921 (
            .O(N__93424),
            .I(N__92746));
    ClkMux I__22920 (
            .O(N__93423),
            .I(N__92746));
    ClkMux I__22919 (
            .O(N__93422),
            .I(N__92746));
    ClkMux I__22918 (
            .O(N__93421),
            .I(N__92746));
    ClkMux I__22917 (
            .O(N__93420),
            .I(N__92746));
    ClkMux I__22916 (
            .O(N__93419),
            .I(N__92746));
    ClkMux I__22915 (
            .O(N__93418),
            .I(N__92746));
    ClkMux I__22914 (
            .O(N__93417),
            .I(N__92746));
    ClkMux I__22913 (
            .O(N__93416),
            .I(N__92746));
    ClkMux I__22912 (
            .O(N__93415),
            .I(N__92746));
    ClkMux I__22911 (
            .O(N__93414),
            .I(N__92746));
    ClkMux I__22910 (
            .O(N__93413),
            .I(N__92746));
    ClkMux I__22909 (
            .O(N__93412),
            .I(N__92746));
    ClkMux I__22908 (
            .O(N__93411),
            .I(N__92746));
    ClkMux I__22907 (
            .O(N__93410),
            .I(N__92746));
    ClkMux I__22906 (
            .O(N__93409),
            .I(N__92746));
    ClkMux I__22905 (
            .O(N__93408),
            .I(N__92746));
    ClkMux I__22904 (
            .O(N__93407),
            .I(N__92746));
    ClkMux I__22903 (
            .O(N__93406),
            .I(N__92746));
    ClkMux I__22902 (
            .O(N__93405),
            .I(N__92746));
    ClkMux I__22901 (
            .O(N__93404),
            .I(N__92746));
    ClkMux I__22900 (
            .O(N__93403),
            .I(N__92746));
    ClkMux I__22899 (
            .O(N__93402),
            .I(N__92746));
    ClkMux I__22898 (
            .O(N__93401),
            .I(N__92746));
    ClkMux I__22897 (
            .O(N__93400),
            .I(N__92746));
    ClkMux I__22896 (
            .O(N__93399),
            .I(N__92746));
    ClkMux I__22895 (
            .O(N__93398),
            .I(N__92746));
    ClkMux I__22894 (
            .O(N__93397),
            .I(N__92746));
    ClkMux I__22893 (
            .O(N__93396),
            .I(N__92746));
    ClkMux I__22892 (
            .O(N__93395),
            .I(N__92746));
    ClkMux I__22891 (
            .O(N__93394),
            .I(N__92746));
    ClkMux I__22890 (
            .O(N__93393),
            .I(N__92746));
    ClkMux I__22889 (
            .O(N__93392),
            .I(N__92746));
    ClkMux I__22888 (
            .O(N__93391),
            .I(N__92746));
    ClkMux I__22887 (
            .O(N__93390),
            .I(N__92746));
    ClkMux I__22886 (
            .O(N__93389),
            .I(N__92746));
    ClkMux I__22885 (
            .O(N__93388),
            .I(N__92746));
    ClkMux I__22884 (
            .O(N__93387),
            .I(N__92746));
    ClkMux I__22883 (
            .O(N__93386),
            .I(N__92746));
    ClkMux I__22882 (
            .O(N__93385),
            .I(N__92746));
    ClkMux I__22881 (
            .O(N__93384),
            .I(N__92746));
    ClkMux I__22880 (
            .O(N__93383),
            .I(N__92746));
    ClkMux I__22879 (
            .O(N__93382),
            .I(N__92746));
    ClkMux I__22878 (
            .O(N__93381),
            .I(N__92746));
    ClkMux I__22877 (
            .O(N__93380),
            .I(N__92746));
    ClkMux I__22876 (
            .O(N__93379),
            .I(N__92746));
    ClkMux I__22875 (
            .O(N__93378),
            .I(N__92746));
    ClkMux I__22874 (
            .O(N__93377),
            .I(N__92746));
    ClkMux I__22873 (
            .O(N__93376),
            .I(N__92746));
    ClkMux I__22872 (
            .O(N__93375),
            .I(N__92746));
    ClkMux I__22871 (
            .O(N__93374),
            .I(N__92746));
    ClkMux I__22870 (
            .O(N__93373),
            .I(N__92746));
    ClkMux I__22869 (
            .O(N__93372),
            .I(N__92746));
    ClkMux I__22868 (
            .O(N__93371),
            .I(N__92746));
    ClkMux I__22867 (
            .O(N__93370),
            .I(N__92746));
    ClkMux I__22866 (
            .O(N__93369),
            .I(N__92746));
    ClkMux I__22865 (
            .O(N__93368),
            .I(N__92746));
    ClkMux I__22864 (
            .O(N__93367),
            .I(N__92746));
    ClkMux I__22863 (
            .O(N__93366),
            .I(N__92746));
    ClkMux I__22862 (
            .O(N__93365),
            .I(N__92746));
    ClkMux I__22861 (
            .O(N__93364),
            .I(N__92746));
    ClkMux I__22860 (
            .O(N__93363),
            .I(N__92746));
    ClkMux I__22859 (
            .O(N__93362),
            .I(N__92746));
    ClkMux I__22858 (
            .O(N__93361),
            .I(N__92746));
    ClkMux I__22857 (
            .O(N__93360),
            .I(N__92746));
    ClkMux I__22856 (
            .O(N__93359),
            .I(N__92746));
    ClkMux I__22855 (
            .O(N__93358),
            .I(N__92746));
    ClkMux I__22854 (
            .O(N__93357),
            .I(N__92746));
    ClkMux I__22853 (
            .O(N__93356),
            .I(N__92746));
    ClkMux I__22852 (
            .O(N__93355),
            .I(N__92746));
    ClkMux I__22851 (
            .O(N__93354),
            .I(N__92746));
    ClkMux I__22850 (
            .O(N__93353),
            .I(N__92746));
    ClkMux I__22849 (
            .O(N__93352),
            .I(N__92746));
    ClkMux I__22848 (
            .O(N__93351),
            .I(N__92746));
    ClkMux I__22847 (
            .O(N__93350),
            .I(N__92746));
    ClkMux I__22846 (
            .O(N__93349),
            .I(N__92746));
    ClkMux I__22845 (
            .O(N__93348),
            .I(N__92746));
    ClkMux I__22844 (
            .O(N__93347),
            .I(N__92746));
    ClkMux I__22843 (
            .O(N__93346),
            .I(N__92746));
    ClkMux I__22842 (
            .O(N__93345),
            .I(N__92746));
    ClkMux I__22841 (
            .O(N__93344),
            .I(N__92746));
    ClkMux I__22840 (
            .O(N__93343),
            .I(N__92746));
    ClkMux I__22839 (
            .O(N__93342),
            .I(N__92746));
    ClkMux I__22838 (
            .O(N__93341),
            .I(N__92746));
    ClkMux I__22837 (
            .O(N__93340),
            .I(N__92746));
    ClkMux I__22836 (
            .O(N__93339),
            .I(N__92746));
    ClkMux I__22835 (
            .O(N__93338),
            .I(N__92746));
    ClkMux I__22834 (
            .O(N__93337),
            .I(N__92746));
    ClkMux I__22833 (
            .O(N__93336),
            .I(N__92746));
    ClkMux I__22832 (
            .O(N__93335),
            .I(N__92746));
    ClkMux I__22831 (
            .O(N__93334),
            .I(N__92746));
    ClkMux I__22830 (
            .O(N__93333),
            .I(N__92746));
    ClkMux I__22829 (
            .O(N__93332),
            .I(N__92746));
    ClkMux I__22828 (
            .O(N__93331),
            .I(N__92746));
    ClkMux I__22827 (
            .O(N__93330),
            .I(N__92746));
    ClkMux I__22826 (
            .O(N__93329),
            .I(N__92746));
    ClkMux I__22825 (
            .O(N__93328),
            .I(N__92746));
    ClkMux I__22824 (
            .O(N__93327),
            .I(N__92746));
    ClkMux I__22823 (
            .O(N__93326),
            .I(N__92746));
    ClkMux I__22822 (
            .O(N__93325),
            .I(N__92746));
    ClkMux I__22821 (
            .O(N__93324),
            .I(N__92746));
    ClkMux I__22820 (
            .O(N__93323),
            .I(N__92746));
    ClkMux I__22819 (
            .O(N__93322),
            .I(N__92746));
    ClkMux I__22818 (
            .O(N__93321),
            .I(N__92746));
    ClkMux I__22817 (
            .O(N__93320),
            .I(N__92746));
    ClkMux I__22816 (
            .O(N__93319),
            .I(N__92746));
    ClkMux I__22815 (
            .O(N__93318),
            .I(N__92746));
    ClkMux I__22814 (
            .O(N__93317),
            .I(N__92746));
    ClkMux I__22813 (
            .O(N__93316),
            .I(N__92746));
    ClkMux I__22812 (
            .O(N__93315),
            .I(N__92746));
    ClkMux I__22811 (
            .O(N__93314),
            .I(N__92746));
    ClkMux I__22810 (
            .O(N__93313),
            .I(N__92746));
    ClkMux I__22809 (
            .O(N__93312),
            .I(N__92746));
    ClkMux I__22808 (
            .O(N__93311),
            .I(N__92746));
    ClkMux I__22807 (
            .O(N__93310),
            .I(N__92746));
    ClkMux I__22806 (
            .O(N__93309),
            .I(N__92746));
    ClkMux I__22805 (
            .O(N__93308),
            .I(N__92746));
    ClkMux I__22804 (
            .O(N__93307),
            .I(N__92746));
    ClkMux I__22803 (
            .O(N__93306),
            .I(N__92746));
    ClkMux I__22802 (
            .O(N__93305),
            .I(N__92746));
    ClkMux I__22801 (
            .O(N__93304),
            .I(N__92746));
    ClkMux I__22800 (
            .O(N__93303),
            .I(N__92746));
    ClkMux I__22799 (
            .O(N__93302),
            .I(N__92746));
    ClkMux I__22798 (
            .O(N__93301),
            .I(N__92746));
    ClkMux I__22797 (
            .O(N__93300),
            .I(N__92746));
    ClkMux I__22796 (
            .O(N__93299),
            .I(N__92746));
    ClkMux I__22795 (
            .O(N__93298),
            .I(N__92746));
    ClkMux I__22794 (
            .O(N__93297),
            .I(N__92746));
    ClkMux I__22793 (
            .O(N__93296),
            .I(N__92746));
    ClkMux I__22792 (
            .O(N__93295),
            .I(N__92746));
    ClkMux I__22791 (
            .O(N__93294),
            .I(N__92746));
    ClkMux I__22790 (
            .O(N__93293),
            .I(N__92746));
    ClkMux I__22789 (
            .O(N__93292),
            .I(N__92746));
    ClkMux I__22788 (
            .O(N__93291),
            .I(N__92746));
    ClkMux I__22787 (
            .O(N__93290),
            .I(N__92746));
    ClkMux I__22786 (
            .O(N__93289),
            .I(N__92746));
    ClkMux I__22785 (
            .O(N__93288),
            .I(N__92746));
    ClkMux I__22784 (
            .O(N__93287),
            .I(N__92746));
    ClkMux I__22783 (
            .O(N__93286),
            .I(N__92746));
    ClkMux I__22782 (
            .O(N__93285),
            .I(N__92746));
    ClkMux I__22781 (
            .O(N__93284),
            .I(N__92746));
    ClkMux I__22780 (
            .O(N__93283),
            .I(N__92746));
    ClkMux I__22779 (
            .O(N__93282),
            .I(N__92746));
    ClkMux I__22778 (
            .O(N__93281),
            .I(N__92746));
    ClkMux I__22777 (
            .O(N__93280),
            .I(N__92746));
    ClkMux I__22776 (
            .O(N__93279),
            .I(N__92746));
    ClkMux I__22775 (
            .O(N__93278),
            .I(N__92746));
    ClkMux I__22774 (
            .O(N__93277),
            .I(N__92746));
    ClkMux I__22773 (
            .O(N__93276),
            .I(N__92746));
    ClkMux I__22772 (
            .O(N__93275),
            .I(N__92746));
    ClkMux I__22771 (
            .O(N__93274),
            .I(N__92746));
    ClkMux I__22770 (
            .O(N__93273),
            .I(N__92746));
    ClkMux I__22769 (
            .O(N__93272),
            .I(N__92746));
    ClkMux I__22768 (
            .O(N__93271),
            .I(N__92746));
    ClkMux I__22767 (
            .O(N__93270),
            .I(N__92746));
    ClkMux I__22766 (
            .O(N__93269),
            .I(N__92746));
    ClkMux I__22765 (
            .O(N__93268),
            .I(N__92746));
    ClkMux I__22764 (
            .O(N__93267),
            .I(N__92746));
    ClkMux I__22763 (
            .O(N__93266),
            .I(N__92746));
    ClkMux I__22762 (
            .O(N__93265),
            .I(N__92746));
    ClkMux I__22761 (
            .O(N__93264),
            .I(N__92746));
    ClkMux I__22760 (
            .O(N__93263),
            .I(N__92746));
    ClkMux I__22759 (
            .O(N__93262),
            .I(N__92746));
    ClkMux I__22758 (
            .O(N__93261),
            .I(N__92746));
    ClkMux I__22757 (
            .O(N__93260),
            .I(N__92746));
    ClkMux I__22756 (
            .O(N__93259),
            .I(N__92746));
    ClkMux I__22755 (
            .O(N__93258),
            .I(N__92746));
    ClkMux I__22754 (
            .O(N__93257),
            .I(N__92746));
    ClkMux I__22753 (
            .O(N__93256),
            .I(N__92746));
    ClkMux I__22752 (
            .O(N__93255),
            .I(N__92746));
    ClkMux I__22751 (
            .O(N__93254),
            .I(N__92746));
    ClkMux I__22750 (
            .O(N__93253),
            .I(N__92746));
    ClkMux I__22749 (
            .O(N__93252),
            .I(N__92746));
    ClkMux I__22748 (
            .O(N__93251),
            .I(N__92746));
    ClkMux I__22747 (
            .O(N__93250),
            .I(N__92746));
    ClkMux I__22746 (
            .O(N__93249),
            .I(N__92746));
    ClkMux I__22745 (
            .O(N__93248),
            .I(N__92746));
    ClkMux I__22744 (
            .O(N__93247),
            .I(N__92746));
    ClkMux I__22743 (
            .O(N__93246),
            .I(N__92746));
    ClkMux I__22742 (
            .O(N__93245),
            .I(N__92746));
    ClkMux I__22741 (
            .O(N__93244),
            .I(N__92746));
    ClkMux I__22740 (
            .O(N__93243),
            .I(N__92746));
    ClkMux I__22739 (
            .O(N__93242),
            .I(N__92746));
    ClkMux I__22738 (
            .O(N__93241),
            .I(N__92746));
    ClkMux I__22737 (
            .O(N__93240),
            .I(N__92746));
    ClkMux I__22736 (
            .O(N__93239),
            .I(N__92746));
    ClkMux I__22735 (
            .O(N__93238),
            .I(N__92746));
    ClkMux I__22734 (
            .O(N__93237),
            .I(N__92746));
    ClkMux I__22733 (
            .O(N__93236),
            .I(N__92746));
    ClkMux I__22732 (
            .O(N__93235),
            .I(N__92746));
    ClkMux I__22731 (
            .O(N__93234),
            .I(N__92746));
    ClkMux I__22730 (
            .O(N__93233),
            .I(N__92746));
    ClkMux I__22729 (
            .O(N__93232),
            .I(N__92746));
    ClkMux I__22728 (
            .O(N__93231),
            .I(N__92746));
    ClkMux I__22727 (
            .O(N__93230),
            .I(N__92746));
    ClkMux I__22726 (
            .O(N__93229),
            .I(N__92746));
    ClkMux I__22725 (
            .O(N__93228),
            .I(N__92746));
    ClkMux I__22724 (
            .O(N__93227),
            .I(N__92746));
    ClkMux I__22723 (
            .O(N__93226),
            .I(N__92746));
    ClkMux I__22722 (
            .O(N__93225),
            .I(N__92746));
    ClkMux I__22721 (
            .O(N__93224),
            .I(N__92746));
    ClkMux I__22720 (
            .O(N__93223),
            .I(N__92746));
    ClkMux I__22719 (
            .O(N__93222),
            .I(N__92746));
    ClkMux I__22718 (
            .O(N__93221),
            .I(N__92746));
    ClkMux I__22717 (
            .O(N__93220),
            .I(N__92746));
    ClkMux I__22716 (
            .O(N__93219),
            .I(N__92746));
    GlobalMux I__22715 (
            .O(N__92746),
            .I(N__92743));
    gio2CtrlBuf I__22714 (
            .O(N__92743),
            .I(DEBUG_6_c_c));
    InMux I__22713 (
            .O(N__92740),
            .I(N__92737));
    LocalMux I__22712 (
            .O(N__92737),
            .I(N__92734));
    Span4Mux_h I__22711 (
            .O(N__92734),
            .I(N__92731));
    Odrv4 I__22710 (
            .O(N__92731),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11784 ));
    CascadeMux I__22709 (
            .O(N__92728),
            .I(N__92725));
    InMux I__22708 (
            .O(N__92725),
            .I(N__92722));
    LocalMux I__22707 (
            .O(N__92722),
            .I(N__92719));
    Odrv4 I__22706 (
            .O(N__92719),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13130 ));
    InMux I__22705 (
            .O(N__92716),
            .I(N__92713));
    LocalMux I__22704 (
            .O(N__92713),
            .I(N__92710));
    Odrv12 I__22703 (
            .O(N__92710),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11760 ));
    InMux I__22702 (
            .O(N__92707),
            .I(N__92704));
    LocalMux I__22701 (
            .O(N__92704),
            .I(N__92701));
    Span4Mux_v I__22700 (
            .O(N__92701),
            .I(N__92698));
    Odrv4 I__22699 (
            .O(N__92698),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11901 ));
    InMux I__22698 (
            .O(N__92695),
            .I(N__92691));
    CascadeMux I__22697 (
            .O(N__92694),
            .I(N__92688));
    LocalMux I__22696 (
            .O(N__92691),
            .I(N__92685));
    InMux I__22695 (
            .O(N__92688),
            .I(N__92682));
    Odrv12 I__22694 (
            .O(N__92685),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_8 ));
    LocalMux I__22693 (
            .O(N__92682),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_8 ));
    InMux I__22692 (
            .O(N__92677),
            .I(N__92669));
    InMux I__22691 (
            .O(N__92676),
            .I(N__92637));
    InMux I__22690 (
            .O(N__92675),
            .I(N__92637));
    InMux I__22689 (
            .O(N__92674),
            .I(N__92637));
    InMux I__22688 (
            .O(N__92673),
            .I(N__92637));
    CascadeMux I__22687 (
            .O(N__92672),
            .I(N__92630));
    LocalMux I__22686 (
            .O(N__92669),
            .I(N__92613));
    CascadeMux I__22685 (
            .O(N__92668),
            .I(N__92606));
    InMux I__22684 (
            .O(N__92667),
            .I(N__92600));
    InMux I__22683 (
            .O(N__92666),
            .I(N__92600));
    CascadeMux I__22682 (
            .O(N__92665),
            .I(N__92590));
    CascadeMux I__22681 (
            .O(N__92664),
            .I(N__92577));
    InMux I__22680 (
            .O(N__92663),
            .I(N__92568));
    InMux I__22679 (
            .O(N__92662),
            .I(N__92568));
    InMux I__22678 (
            .O(N__92661),
            .I(N__92568));
    InMux I__22677 (
            .O(N__92660),
            .I(N__92568));
    CascadeMux I__22676 (
            .O(N__92659),
            .I(N__92557));
    InMux I__22675 (
            .O(N__92658),
            .I(N__92546));
    InMux I__22674 (
            .O(N__92657),
            .I(N__92546));
    InMux I__22673 (
            .O(N__92656),
            .I(N__92546));
    InMux I__22672 (
            .O(N__92655),
            .I(N__92546));
    CascadeMux I__22671 (
            .O(N__92654),
            .I(N__92542));
    InMux I__22670 (
            .O(N__92653),
            .I(N__92531));
    InMux I__22669 (
            .O(N__92652),
            .I(N__92531));
    InMux I__22668 (
            .O(N__92651),
            .I(N__92531));
    InMux I__22667 (
            .O(N__92650),
            .I(N__92531));
    InMux I__22666 (
            .O(N__92649),
            .I(N__92522));
    InMux I__22665 (
            .O(N__92648),
            .I(N__92522));
    InMux I__22664 (
            .O(N__92647),
            .I(N__92522));
    InMux I__22663 (
            .O(N__92646),
            .I(N__92522));
    LocalMux I__22662 (
            .O(N__92637),
            .I(N__92514));
    InMux I__22661 (
            .O(N__92636),
            .I(N__92511));
    InMux I__22660 (
            .O(N__92635),
            .I(N__92504));
    InMux I__22659 (
            .O(N__92634),
            .I(N__92504));
    InMux I__22658 (
            .O(N__92633),
            .I(N__92504));
    InMux I__22657 (
            .O(N__92630),
            .I(N__92499));
    InMux I__22656 (
            .O(N__92629),
            .I(N__92499));
    CascadeMux I__22655 (
            .O(N__92628),
            .I(N__92496));
    InMux I__22654 (
            .O(N__92627),
            .I(N__92482));
    InMux I__22653 (
            .O(N__92626),
            .I(N__92482));
    InMux I__22652 (
            .O(N__92625),
            .I(N__92482));
    InMux I__22651 (
            .O(N__92624),
            .I(N__92482));
    InMux I__22650 (
            .O(N__92623),
            .I(N__92477));
    InMux I__22649 (
            .O(N__92622),
            .I(N__92477));
    InMux I__22648 (
            .O(N__92621),
            .I(N__92470));
    InMux I__22647 (
            .O(N__92620),
            .I(N__92470));
    InMux I__22646 (
            .O(N__92619),
            .I(N__92470));
    InMux I__22645 (
            .O(N__92618),
            .I(N__92465));
    InMux I__22644 (
            .O(N__92617),
            .I(N__92465));
    InMux I__22643 (
            .O(N__92616),
            .I(N__92462));
    Span4Mux_v I__22642 (
            .O(N__92613),
            .I(N__92459));
    InMux I__22641 (
            .O(N__92612),
            .I(N__92450));
    InMux I__22640 (
            .O(N__92611),
            .I(N__92450));
    InMux I__22639 (
            .O(N__92610),
            .I(N__92450));
    InMux I__22638 (
            .O(N__92609),
            .I(N__92450));
    InMux I__22637 (
            .O(N__92606),
            .I(N__92436));
    InMux I__22636 (
            .O(N__92605),
            .I(N__92436));
    LocalMux I__22635 (
            .O(N__92600),
            .I(N__92433));
    InMux I__22634 (
            .O(N__92599),
            .I(N__92427));
    CascadeMux I__22633 (
            .O(N__92598),
            .I(N__92421));
    CascadeMux I__22632 (
            .O(N__92597),
            .I(N__92416));
    CascadeMux I__22631 (
            .O(N__92596),
            .I(N__92410));
    InMux I__22630 (
            .O(N__92595),
            .I(N__92402));
    InMux I__22629 (
            .O(N__92594),
            .I(N__92402));
    InMux I__22628 (
            .O(N__92593),
            .I(N__92393));
    InMux I__22627 (
            .O(N__92590),
            .I(N__92393));
    InMux I__22626 (
            .O(N__92589),
            .I(N__92390));
    CascadeMux I__22625 (
            .O(N__92588),
            .I(N__92381));
    InMux I__22624 (
            .O(N__92587),
            .I(N__92377));
    CascadeMux I__22623 (
            .O(N__92586),
            .I(N__92374));
    InMux I__22622 (
            .O(N__92585),
            .I(N__92367));
    InMux I__22621 (
            .O(N__92584),
            .I(N__92367));
    InMux I__22620 (
            .O(N__92583),
            .I(N__92364));
    InMux I__22619 (
            .O(N__92582),
            .I(N__92361));
    InMux I__22618 (
            .O(N__92581),
            .I(N__92358));
    InMux I__22617 (
            .O(N__92580),
            .I(N__92353));
    InMux I__22616 (
            .O(N__92577),
            .I(N__92353));
    LocalMux I__22615 (
            .O(N__92568),
            .I(N__92347));
    InMux I__22614 (
            .O(N__92567),
            .I(N__92344));
    InMux I__22613 (
            .O(N__92566),
            .I(N__92341));
    InMux I__22612 (
            .O(N__92565),
            .I(N__92334));
    InMux I__22611 (
            .O(N__92564),
            .I(N__92334));
    InMux I__22610 (
            .O(N__92563),
            .I(N__92334));
    InMux I__22609 (
            .O(N__92562),
            .I(N__92329));
    InMux I__22608 (
            .O(N__92561),
            .I(N__92329));
    InMux I__22607 (
            .O(N__92560),
            .I(N__92322));
    InMux I__22606 (
            .O(N__92557),
            .I(N__92322));
    InMux I__22605 (
            .O(N__92556),
            .I(N__92322));
    InMux I__22604 (
            .O(N__92555),
            .I(N__92313));
    LocalMux I__22603 (
            .O(N__92546),
            .I(N__92310));
    InMux I__22602 (
            .O(N__92545),
            .I(N__92307));
    InMux I__22601 (
            .O(N__92542),
            .I(N__92304));
    InMux I__22600 (
            .O(N__92541),
            .I(N__92299));
    InMux I__22599 (
            .O(N__92540),
            .I(N__92299));
    LocalMux I__22598 (
            .O(N__92531),
            .I(N__92294));
    LocalMux I__22597 (
            .O(N__92522),
            .I(N__92294));
    InMux I__22596 (
            .O(N__92521),
            .I(N__92289));
    InMux I__22595 (
            .O(N__92520),
            .I(N__92289));
    InMux I__22594 (
            .O(N__92519),
            .I(N__92276));
    InMux I__22593 (
            .O(N__92518),
            .I(N__92276));
    InMux I__22592 (
            .O(N__92517),
            .I(N__92273));
    Span4Mux_h I__22591 (
            .O(N__92514),
            .I(N__92263));
    LocalMux I__22590 (
            .O(N__92511),
            .I(N__92263));
    LocalMux I__22589 (
            .O(N__92504),
            .I(N__92260));
    LocalMux I__22588 (
            .O(N__92499),
            .I(N__92257));
    InMux I__22587 (
            .O(N__92496),
            .I(N__92252));
    InMux I__22586 (
            .O(N__92495),
            .I(N__92252));
    InMux I__22585 (
            .O(N__92494),
            .I(N__92249));
    InMux I__22584 (
            .O(N__92493),
            .I(N__92246));
    InMux I__22583 (
            .O(N__92492),
            .I(N__92243));
    InMux I__22582 (
            .O(N__92491),
            .I(N__92240));
    LocalMux I__22581 (
            .O(N__92482),
            .I(N__92237));
    LocalMux I__22580 (
            .O(N__92477),
            .I(N__92228));
    LocalMux I__22579 (
            .O(N__92470),
            .I(N__92228));
    LocalMux I__22578 (
            .O(N__92465),
            .I(N__92228));
    LocalMux I__22577 (
            .O(N__92462),
            .I(N__92228));
    Span4Mux_h I__22576 (
            .O(N__92459),
            .I(N__92223));
    LocalMux I__22575 (
            .O(N__92450),
            .I(N__92223));
    InMux I__22574 (
            .O(N__92449),
            .I(N__92220));
    InMux I__22573 (
            .O(N__92448),
            .I(N__92217));
    InMux I__22572 (
            .O(N__92447),
            .I(N__92206));
    InMux I__22571 (
            .O(N__92446),
            .I(N__92197));
    InMux I__22570 (
            .O(N__92445),
            .I(N__92197));
    InMux I__22569 (
            .O(N__92444),
            .I(N__92197));
    InMux I__22568 (
            .O(N__92443),
            .I(N__92197));
    InMux I__22567 (
            .O(N__92442),
            .I(N__92192));
    InMux I__22566 (
            .O(N__92441),
            .I(N__92192));
    LocalMux I__22565 (
            .O(N__92436),
            .I(N__92188));
    Span4Mux_h I__22564 (
            .O(N__92433),
            .I(N__92185));
    InMux I__22563 (
            .O(N__92432),
            .I(N__92180));
    InMux I__22562 (
            .O(N__92431),
            .I(N__92180));
    CascadeMux I__22561 (
            .O(N__92430),
            .I(N__92177));
    LocalMux I__22560 (
            .O(N__92427),
            .I(N__92166));
    InMux I__22559 (
            .O(N__92426),
            .I(N__92159));
    InMux I__22558 (
            .O(N__92425),
            .I(N__92159));
    InMux I__22557 (
            .O(N__92424),
            .I(N__92159));
    InMux I__22556 (
            .O(N__92421),
            .I(N__92152));
    InMux I__22555 (
            .O(N__92420),
            .I(N__92152));
    InMux I__22554 (
            .O(N__92419),
            .I(N__92152));
    InMux I__22553 (
            .O(N__92416),
            .I(N__92143));
    InMux I__22552 (
            .O(N__92415),
            .I(N__92143));
    InMux I__22551 (
            .O(N__92414),
            .I(N__92143));
    InMux I__22550 (
            .O(N__92413),
            .I(N__92143));
    InMux I__22549 (
            .O(N__92410),
            .I(N__92136));
    CascadeMux I__22548 (
            .O(N__92409),
            .I(N__92132));
    InMux I__22547 (
            .O(N__92408),
            .I(N__92124));
    InMux I__22546 (
            .O(N__92407),
            .I(N__92124));
    LocalMux I__22545 (
            .O(N__92402),
            .I(N__92121));
    InMux I__22544 (
            .O(N__92401),
            .I(N__92116));
    InMux I__22543 (
            .O(N__92400),
            .I(N__92116));
    CascadeMux I__22542 (
            .O(N__92399),
            .I(N__92101));
    CascadeMux I__22541 (
            .O(N__92398),
            .I(N__92098));
    LocalMux I__22540 (
            .O(N__92393),
            .I(N__92092));
    LocalMux I__22539 (
            .O(N__92390),
            .I(N__92092));
    InMux I__22538 (
            .O(N__92389),
            .I(N__92083));
    InMux I__22537 (
            .O(N__92388),
            .I(N__92083));
    InMux I__22536 (
            .O(N__92387),
            .I(N__92083));
    InMux I__22535 (
            .O(N__92386),
            .I(N__92083));
    InMux I__22534 (
            .O(N__92385),
            .I(N__92078));
    InMux I__22533 (
            .O(N__92384),
            .I(N__92078));
    InMux I__22532 (
            .O(N__92381),
            .I(N__92073));
    InMux I__22531 (
            .O(N__92380),
            .I(N__92073));
    LocalMux I__22530 (
            .O(N__92377),
            .I(N__92070));
    InMux I__22529 (
            .O(N__92374),
            .I(N__92063));
    InMux I__22528 (
            .O(N__92373),
            .I(N__92063));
    InMux I__22527 (
            .O(N__92372),
            .I(N__92063));
    LocalMux I__22526 (
            .O(N__92367),
            .I(N__92057));
    LocalMux I__22525 (
            .O(N__92364),
            .I(N__92057));
    LocalMux I__22524 (
            .O(N__92361),
            .I(N__92052));
    LocalMux I__22523 (
            .O(N__92358),
            .I(N__92052));
    LocalMux I__22522 (
            .O(N__92353),
            .I(N__92049));
    InMux I__22521 (
            .O(N__92352),
            .I(N__92042));
    InMux I__22520 (
            .O(N__92351),
            .I(N__92042));
    InMux I__22519 (
            .O(N__92350),
            .I(N__92042));
    Span4Mux_h I__22518 (
            .O(N__92347),
            .I(N__92032));
    LocalMux I__22517 (
            .O(N__92344),
            .I(N__92032));
    LocalMux I__22516 (
            .O(N__92341),
            .I(N__92032));
    LocalMux I__22515 (
            .O(N__92334),
            .I(N__92022));
    LocalMux I__22514 (
            .O(N__92329),
            .I(N__92022));
    LocalMux I__22513 (
            .O(N__92322),
            .I(N__92019));
    InMux I__22512 (
            .O(N__92321),
            .I(N__92016));
    InMux I__22511 (
            .O(N__92320),
            .I(N__92011));
    InMux I__22510 (
            .O(N__92319),
            .I(N__92011));
    InMux I__22509 (
            .O(N__92318),
            .I(N__91996));
    InMux I__22508 (
            .O(N__92317),
            .I(N__91996));
    InMux I__22507 (
            .O(N__92316),
            .I(N__91996));
    LocalMux I__22506 (
            .O(N__92313),
            .I(N__91982));
    Span4Mux_v I__22505 (
            .O(N__92310),
            .I(N__91977));
    LocalMux I__22504 (
            .O(N__92307),
            .I(N__91977));
    LocalMux I__22503 (
            .O(N__92304),
            .I(N__91972));
    LocalMux I__22502 (
            .O(N__92299),
            .I(N__91972));
    Span4Mux_v I__22501 (
            .O(N__92294),
            .I(N__91967));
    LocalMux I__22500 (
            .O(N__92289),
            .I(N__91967));
    InMux I__22499 (
            .O(N__92288),
            .I(N__91956));
    InMux I__22498 (
            .O(N__92287),
            .I(N__91956));
    InMux I__22497 (
            .O(N__92286),
            .I(N__91956));
    InMux I__22496 (
            .O(N__92285),
            .I(N__91956));
    InMux I__22495 (
            .O(N__92284),
            .I(N__91956));
    InMux I__22494 (
            .O(N__92283),
            .I(N__91949));
    InMux I__22493 (
            .O(N__92282),
            .I(N__91949));
    InMux I__22492 (
            .O(N__92281),
            .I(N__91949));
    LocalMux I__22491 (
            .O(N__92276),
            .I(N__91942));
    LocalMux I__22490 (
            .O(N__92273),
            .I(N__91942));
    InMux I__22489 (
            .O(N__92272),
            .I(N__91939));
    InMux I__22488 (
            .O(N__92271),
            .I(N__91936));
    InMux I__22487 (
            .O(N__92270),
            .I(N__91931));
    InMux I__22486 (
            .O(N__92269),
            .I(N__91931));
    InMux I__22485 (
            .O(N__92268),
            .I(N__91928));
    Span4Mux_h I__22484 (
            .O(N__92263),
            .I(N__91917));
    Span4Mux_v I__22483 (
            .O(N__92260),
            .I(N__91917));
    Span4Mux_h I__22482 (
            .O(N__92257),
            .I(N__91917));
    LocalMux I__22481 (
            .O(N__92252),
            .I(N__91917));
    LocalMux I__22480 (
            .O(N__92249),
            .I(N__91912));
    LocalMux I__22479 (
            .O(N__92246),
            .I(N__91912));
    LocalMux I__22478 (
            .O(N__92243),
            .I(N__91907));
    LocalMux I__22477 (
            .O(N__92240),
            .I(N__91907));
    Span4Mux_v I__22476 (
            .O(N__92237),
            .I(N__91896));
    Span4Mux_v I__22475 (
            .O(N__92228),
            .I(N__91896));
    Span4Mux_h I__22474 (
            .O(N__92223),
            .I(N__91896));
    LocalMux I__22473 (
            .O(N__92220),
            .I(N__91896));
    LocalMux I__22472 (
            .O(N__92217),
            .I(N__91896));
    InMux I__22471 (
            .O(N__92216),
            .I(N__91887));
    InMux I__22470 (
            .O(N__92215),
            .I(N__91887));
    InMux I__22469 (
            .O(N__92214),
            .I(N__91887));
    InMux I__22468 (
            .O(N__92213),
            .I(N__91887));
    CascadeMux I__22467 (
            .O(N__92212),
            .I(N__91880));
    InMux I__22466 (
            .O(N__92211),
            .I(N__91873));
    InMux I__22465 (
            .O(N__92210),
            .I(N__91873));
    CascadeMux I__22464 (
            .O(N__92209),
            .I(N__91865));
    LocalMux I__22463 (
            .O(N__92206),
            .I(N__91854));
    LocalMux I__22462 (
            .O(N__92197),
            .I(N__91854));
    LocalMux I__22461 (
            .O(N__92192),
            .I(N__91854));
    InMux I__22460 (
            .O(N__92191),
            .I(N__91851));
    Span4Mux_h I__22459 (
            .O(N__92188),
            .I(N__91844));
    Span4Mux_v I__22458 (
            .O(N__92185),
            .I(N__91844));
    LocalMux I__22457 (
            .O(N__92180),
            .I(N__91844));
    InMux I__22456 (
            .O(N__92177),
            .I(N__91837));
    InMux I__22455 (
            .O(N__92176),
            .I(N__91837));
    InMux I__22454 (
            .O(N__92175),
            .I(N__91837));
    InMux I__22453 (
            .O(N__92174),
            .I(N__91828));
    InMux I__22452 (
            .O(N__92173),
            .I(N__91828));
    InMux I__22451 (
            .O(N__92172),
            .I(N__91821));
    InMux I__22450 (
            .O(N__92171),
            .I(N__91821));
    InMux I__22449 (
            .O(N__92170),
            .I(N__91821));
    CascadeMux I__22448 (
            .O(N__92169),
            .I(N__91817));
    Span4Mux_h I__22447 (
            .O(N__92166),
            .I(N__91803));
    LocalMux I__22446 (
            .O(N__92159),
            .I(N__91803));
    LocalMux I__22445 (
            .O(N__92152),
            .I(N__91798));
    LocalMux I__22444 (
            .O(N__92143),
            .I(N__91798));
    InMux I__22443 (
            .O(N__92142),
            .I(N__91787));
    InMux I__22442 (
            .O(N__92141),
            .I(N__91787));
    InMux I__22441 (
            .O(N__92140),
            .I(N__91787));
    InMux I__22440 (
            .O(N__92139),
            .I(N__91787));
    LocalMux I__22439 (
            .O(N__92136),
            .I(N__91781));
    InMux I__22438 (
            .O(N__92135),
            .I(N__91776));
    InMux I__22437 (
            .O(N__92132),
            .I(N__91776));
    CascadeMux I__22436 (
            .O(N__92131),
            .I(N__91772));
    CascadeMux I__22435 (
            .O(N__92130),
            .I(N__91769));
    InMux I__22434 (
            .O(N__92129),
            .I(N__91760));
    LocalMux I__22433 (
            .O(N__92124),
            .I(N__91753));
    Span4Mux_v I__22432 (
            .O(N__92121),
            .I(N__91753));
    LocalMux I__22431 (
            .O(N__92116),
            .I(N__91753));
    InMux I__22430 (
            .O(N__92115),
            .I(N__91748));
    InMux I__22429 (
            .O(N__92114),
            .I(N__91748));
    CascadeMux I__22428 (
            .O(N__92113),
            .I(N__91740));
    InMux I__22427 (
            .O(N__92112),
            .I(N__91723));
    InMux I__22426 (
            .O(N__92111),
            .I(N__91723));
    InMux I__22425 (
            .O(N__92110),
            .I(N__91723));
    InMux I__22424 (
            .O(N__92109),
            .I(N__91720));
    InMux I__22423 (
            .O(N__92108),
            .I(N__91717));
    InMux I__22422 (
            .O(N__92107),
            .I(N__91712));
    InMux I__22421 (
            .O(N__92106),
            .I(N__91712));
    InMux I__22420 (
            .O(N__92105),
            .I(N__91707));
    InMux I__22419 (
            .O(N__92104),
            .I(N__91707));
    InMux I__22418 (
            .O(N__92101),
            .I(N__91700));
    InMux I__22417 (
            .O(N__92098),
            .I(N__91700));
    InMux I__22416 (
            .O(N__92097),
            .I(N__91700));
    Span4Mux_v I__22415 (
            .O(N__92092),
            .I(N__91694));
    LocalMux I__22414 (
            .O(N__92083),
            .I(N__91694));
    LocalMux I__22413 (
            .O(N__92078),
            .I(N__91689));
    LocalMux I__22412 (
            .O(N__92073),
            .I(N__91689));
    Span4Mux_h I__22411 (
            .O(N__92070),
            .I(N__91684));
    LocalMux I__22410 (
            .O(N__92063),
            .I(N__91684));
    InMux I__22409 (
            .O(N__92062),
            .I(N__91681));
    Span4Mux_h I__22408 (
            .O(N__92057),
            .I(N__91670));
    Span4Mux_h I__22407 (
            .O(N__92052),
            .I(N__91670));
    Span4Mux_v I__22406 (
            .O(N__92049),
            .I(N__91670));
    LocalMux I__22405 (
            .O(N__92042),
            .I(N__91670));
    InMux I__22404 (
            .O(N__92041),
            .I(N__91663));
    InMux I__22403 (
            .O(N__92040),
            .I(N__91663));
    InMux I__22402 (
            .O(N__92039),
            .I(N__91663));
    Span4Mux_h I__22401 (
            .O(N__92032),
            .I(N__91658));
    InMux I__22400 (
            .O(N__92031),
            .I(N__91655));
    InMux I__22399 (
            .O(N__92030),
            .I(N__91650));
    InMux I__22398 (
            .O(N__92029),
            .I(N__91650));
    InMux I__22397 (
            .O(N__92028),
            .I(N__91647));
    InMux I__22396 (
            .O(N__92027),
            .I(N__91644));
    Span4Mux_v I__22395 (
            .O(N__92022),
            .I(N__91633));
    Span4Mux_v I__22394 (
            .O(N__92019),
            .I(N__91633));
    LocalMux I__22393 (
            .O(N__92016),
            .I(N__91633));
    LocalMux I__22392 (
            .O(N__92011),
            .I(N__91633));
    InMux I__22391 (
            .O(N__92010),
            .I(N__91630));
    InMux I__22390 (
            .O(N__92009),
            .I(N__91625));
    InMux I__22389 (
            .O(N__92008),
            .I(N__91625));
    InMux I__22388 (
            .O(N__92007),
            .I(N__91614));
    InMux I__22387 (
            .O(N__92006),
            .I(N__91614));
    InMux I__22386 (
            .O(N__92005),
            .I(N__91614));
    InMux I__22385 (
            .O(N__92004),
            .I(N__91614));
    InMux I__22384 (
            .O(N__92003),
            .I(N__91614));
    LocalMux I__22383 (
            .O(N__91996),
            .I(N__91611));
    InMux I__22382 (
            .O(N__91995),
            .I(N__91606));
    InMux I__22381 (
            .O(N__91994),
            .I(N__91606));
    InMux I__22380 (
            .O(N__91993),
            .I(N__91603));
    InMux I__22379 (
            .O(N__91992),
            .I(N__91597));
    InMux I__22378 (
            .O(N__91991),
            .I(N__91594));
    CascadeMux I__22377 (
            .O(N__91990),
            .I(N__91591));
    CascadeMux I__22376 (
            .O(N__91989),
            .I(N__91584));
    InMux I__22375 (
            .O(N__91988),
            .I(N__91575));
    InMux I__22374 (
            .O(N__91987),
            .I(N__91575));
    InMux I__22373 (
            .O(N__91986),
            .I(N__91575));
    InMux I__22372 (
            .O(N__91985),
            .I(N__91575));
    Span4Mux_v I__22371 (
            .O(N__91982),
            .I(N__91564));
    Span4Mux_v I__22370 (
            .O(N__91977),
            .I(N__91553));
    Span4Mux_h I__22369 (
            .O(N__91972),
            .I(N__91553));
    Span4Mux_v I__22368 (
            .O(N__91967),
            .I(N__91553));
    LocalMux I__22367 (
            .O(N__91956),
            .I(N__91553));
    LocalMux I__22366 (
            .O(N__91949),
            .I(N__91553));
    InMux I__22365 (
            .O(N__91948),
            .I(N__91548));
    InMux I__22364 (
            .O(N__91947),
            .I(N__91548));
    Span4Mux_v I__22363 (
            .O(N__91942),
            .I(N__91537));
    LocalMux I__22362 (
            .O(N__91939),
            .I(N__91537));
    LocalMux I__22361 (
            .O(N__91936),
            .I(N__91537));
    LocalMux I__22360 (
            .O(N__91931),
            .I(N__91537));
    LocalMux I__22359 (
            .O(N__91928),
            .I(N__91537));
    InMux I__22358 (
            .O(N__91927),
            .I(N__91532));
    InMux I__22357 (
            .O(N__91926),
            .I(N__91532));
    Span4Mux_h I__22356 (
            .O(N__91917),
            .I(N__91521));
    Span4Mux_v I__22355 (
            .O(N__91912),
            .I(N__91521));
    Span4Mux_v I__22354 (
            .O(N__91907),
            .I(N__91521));
    Span4Mux_v I__22353 (
            .O(N__91896),
            .I(N__91521));
    LocalMux I__22352 (
            .O(N__91887),
            .I(N__91521));
    InMux I__22351 (
            .O(N__91886),
            .I(N__91518));
    InMux I__22350 (
            .O(N__91885),
            .I(N__91511));
    InMux I__22349 (
            .O(N__91884),
            .I(N__91511));
    InMux I__22348 (
            .O(N__91883),
            .I(N__91511));
    InMux I__22347 (
            .O(N__91880),
            .I(N__91506));
    InMux I__22346 (
            .O(N__91879),
            .I(N__91506));
    CascadeMux I__22345 (
            .O(N__91878),
            .I(N__91503));
    LocalMux I__22344 (
            .O(N__91873),
            .I(N__91499));
    InMux I__22343 (
            .O(N__91872),
            .I(N__91492));
    InMux I__22342 (
            .O(N__91871),
            .I(N__91492));
    InMux I__22341 (
            .O(N__91870),
            .I(N__91492));
    InMux I__22340 (
            .O(N__91869),
            .I(N__91483));
    InMux I__22339 (
            .O(N__91868),
            .I(N__91483));
    InMux I__22338 (
            .O(N__91865),
            .I(N__91483));
    InMux I__22337 (
            .O(N__91864),
            .I(N__91483));
    CascadeMux I__22336 (
            .O(N__91863),
            .I(N__91480));
    InMux I__22335 (
            .O(N__91862),
            .I(N__91474));
    InMux I__22334 (
            .O(N__91861),
            .I(N__91471));
    Span4Mux_h I__22333 (
            .O(N__91854),
            .I(N__91462));
    LocalMux I__22332 (
            .O(N__91851),
            .I(N__91462));
    Span4Mux_h I__22331 (
            .O(N__91844),
            .I(N__91462));
    LocalMux I__22330 (
            .O(N__91837),
            .I(N__91462));
    InMux I__22329 (
            .O(N__91836),
            .I(N__91453));
    InMux I__22328 (
            .O(N__91835),
            .I(N__91453));
    InMux I__22327 (
            .O(N__91834),
            .I(N__91453));
    InMux I__22326 (
            .O(N__91833),
            .I(N__91453));
    LocalMux I__22325 (
            .O(N__91828),
            .I(N__91450));
    LocalMux I__22324 (
            .O(N__91821),
            .I(N__91447));
    InMux I__22323 (
            .O(N__91820),
            .I(N__91440));
    InMux I__22322 (
            .O(N__91817),
            .I(N__91440));
    InMux I__22321 (
            .O(N__91816),
            .I(N__91440));
    InMux I__22320 (
            .O(N__91815),
            .I(N__91435));
    InMux I__22319 (
            .O(N__91814),
            .I(N__91435));
    CascadeMux I__22318 (
            .O(N__91813),
            .I(N__91432));
    InMux I__22317 (
            .O(N__91812),
            .I(N__91427));
    InMux I__22316 (
            .O(N__91811),
            .I(N__91427));
    InMux I__22315 (
            .O(N__91810),
            .I(N__91422));
    InMux I__22314 (
            .O(N__91809),
            .I(N__91422));
    InMux I__22313 (
            .O(N__91808),
            .I(N__91419));
    Span4Mux_h I__22312 (
            .O(N__91803),
            .I(N__91411));
    Span4Mux_v I__22311 (
            .O(N__91798),
            .I(N__91411));
    InMux I__22310 (
            .O(N__91797),
            .I(N__91406));
    InMux I__22309 (
            .O(N__91796),
            .I(N__91406));
    LocalMux I__22308 (
            .O(N__91787),
            .I(N__91400));
    InMux I__22307 (
            .O(N__91786),
            .I(N__91397));
    InMux I__22306 (
            .O(N__91785),
            .I(N__91394));
    InMux I__22305 (
            .O(N__91784),
            .I(N__91391));
    Span4Mux_v I__22304 (
            .O(N__91781),
            .I(N__91386));
    LocalMux I__22303 (
            .O(N__91776),
            .I(N__91386));
    InMux I__22302 (
            .O(N__91775),
            .I(N__91381));
    InMux I__22301 (
            .O(N__91772),
            .I(N__91381));
    InMux I__22300 (
            .O(N__91769),
            .I(N__91378));
    InMux I__22299 (
            .O(N__91768),
            .I(N__91369));
    InMux I__22298 (
            .O(N__91767),
            .I(N__91369));
    InMux I__22297 (
            .O(N__91766),
            .I(N__91369));
    InMux I__22296 (
            .O(N__91765),
            .I(N__91369));
    InMux I__22295 (
            .O(N__91764),
            .I(N__91357));
    InMux I__22294 (
            .O(N__91763),
            .I(N__91357));
    LocalMux I__22293 (
            .O(N__91760),
            .I(N__91340));
    Span4Mux_h I__22292 (
            .O(N__91753),
            .I(N__91340));
    LocalMux I__22291 (
            .O(N__91748),
            .I(N__91340));
    InMux I__22290 (
            .O(N__91747),
            .I(N__91331));
    InMux I__22289 (
            .O(N__91746),
            .I(N__91331));
    InMux I__22288 (
            .O(N__91745),
            .I(N__91331));
    InMux I__22287 (
            .O(N__91744),
            .I(N__91331));
    InMux I__22286 (
            .O(N__91743),
            .I(N__91322));
    InMux I__22285 (
            .O(N__91740),
            .I(N__91319));
    InMux I__22284 (
            .O(N__91739),
            .I(N__91316));
    InMux I__22283 (
            .O(N__91738),
            .I(N__91309));
    InMux I__22282 (
            .O(N__91737),
            .I(N__91309));
    InMux I__22281 (
            .O(N__91736),
            .I(N__91309));
    InMux I__22280 (
            .O(N__91735),
            .I(N__91302));
    InMux I__22279 (
            .O(N__91734),
            .I(N__91302));
    InMux I__22278 (
            .O(N__91733),
            .I(N__91302));
    InMux I__22277 (
            .O(N__91732),
            .I(N__91299));
    InMux I__22276 (
            .O(N__91731),
            .I(N__91296));
    CascadeMux I__22275 (
            .O(N__91730),
            .I(N__91285));
    LocalMux I__22274 (
            .O(N__91723),
            .I(N__91275));
    LocalMux I__22273 (
            .O(N__91720),
            .I(N__91275));
    LocalMux I__22272 (
            .O(N__91717),
            .I(N__91275));
    LocalMux I__22271 (
            .O(N__91712),
            .I(N__91268));
    LocalMux I__22270 (
            .O(N__91707),
            .I(N__91268));
    LocalMux I__22269 (
            .O(N__91700),
            .I(N__91268));
    InMux I__22268 (
            .O(N__91699),
            .I(N__91265));
    Span4Mux_h I__22267 (
            .O(N__91694),
            .I(N__91256));
    Span4Mux_v I__22266 (
            .O(N__91689),
            .I(N__91256));
    Span4Mux_v I__22265 (
            .O(N__91684),
            .I(N__91256));
    LocalMux I__22264 (
            .O(N__91681),
            .I(N__91256));
    InMux I__22263 (
            .O(N__91680),
            .I(N__91251));
    InMux I__22262 (
            .O(N__91679),
            .I(N__91251));
    Span4Mux_v I__22261 (
            .O(N__91670),
            .I(N__91246));
    LocalMux I__22260 (
            .O(N__91663),
            .I(N__91246));
    InMux I__22259 (
            .O(N__91662),
            .I(N__91243));
    CascadeMux I__22258 (
            .O(N__91661),
            .I(N__91231));
    Span4Mux_h I__22257 (
            .O(N__91658),
            .I(N__91214));
    LocalMux I__22256 (
            .O(N__91655),
            .I(N__91214));
    LocalMux I__22255 (
            .O(N__91650),
            .I(N__91214));
    LocalMux I__22254 (
            .O(N__91647),
            .I(N__91209));
    LocalMux I__22253 (
            .O(N__91644),
            .I(N__91209));
    InMux I__22252 (
            .O(N__91643),
            .I(N__91204));
    InMux I__22251 (
            .O(N__91642),
            .I(N__91204));
    Span4Mux_h I__22250 (
            .O(N__91633),
            .I(N__91195));
    LocalMux I__22249 (
            .O(N__91630),
            .I(N__91195));
    LocalMux I__22248 (
            .O(N__91625),
            .I(N__91195));
    LocalMux I__22247 (
            .O(N__91614),
            .I(N__91195));
    Span4Mux_v I__22246 (
            .O(N__91611),
            .I(N__91188));
    LocalMux I__22245 (
            .O(N__91606),
            .I(N__91188));
    LocalMux I__22244 (
            .O(N__91603),
            .I(N__91188));
    InMux I__22243 (
            .O(N__91602),
            .I(N__91185));
    InMux I__22242 (
            .O(N__91601),
            .I(N__91180));
    InMux I__22241 (
            .O(N__91600),
            .I(N__91180));
    LocalMux I__22240 (
            .O(N__91597),
            .I(N__91175));
    LocalMux I__22239 (
            .O(N__91594),
            .I(N__91175));
    InMux I__22238 (
            .O(N__91591),
            .I(N__91164));
    InMux I__22237 (
            .O(N__91590),
            .I(N__91164));
    InMux I__22236 (
            .O(N__91589),
            .I(N__91164));
    InMux I__22235 (
            .O(N__91588),
            .I(N__91164));
    InMux I__22234 (
            .O(N__91587),
            .I(N__91164));
    InMux I__22233 (
            .O(N__91584),
            .I(N__91161));
    LocalMux I__22232 (
            .O(N__91575),
            .I(N__91158));
    InMux I__22231 (
            .O(N__91574),
            .I(N__91155));
    InMux I__22230 (
            .O(N__91573),
            .I(N__91146));
    InMux I__22229 (
            .O(N__91572),
            .I(N__91146));
    InMux I__22228 (
            .O(N__91571),
            .I(N__91146));
    InMux I__22227 (
            .O(N__91570),
            .I(N__91146));
    InMux I__22226 (
            .O(N__91569),
            .I(N__91139));
    InMux I__22225 (
            .O(N__91568),
            .I(N__91139));
    InMux I__22224 (
            .O(N__91567),
            .I(N__91139));
    Span4Mux_h I__22223 (
            .O(N__91564),
            .I(N__91132));
    Span4Mux_h I__22222 (
            .O(N__91553),
            .I(N__91132));
    LocalMux I__22221 (
            .O(N__91548),
            .I(N__91132));
    Span4Mux_v I__22220 (
            .O(N__91537),
            .I(N__91127));
    LocalMux I__22219 (
            .O(N__91532),
            .I(N__91127));
    Span4Mux_h I__22218 (
            .O(N__91521),
            .I(N__91118));
    LocalMux I__22217 (
            .O(N__91518),
            .I(N__91118));
    LocalMux I__22216 (
            .O(N__91511),
            .I(N__91118));
    LocalMux I__22215 (
            .O(N__91506),
            .I(N__91118));
    InMux I__22214 (
            .O(N__91503),
            .I(N__91115));
    InMux I__22213 (
            .O(N__91502),
            .I(N__91112));
    Span4Mux_v I__22212 (
            .O(N__91499),
            .I(N__91103));
    LocalMux I__22211 (
            .O(N__91492),
            .I(N__91103));
    LocalMux I__22210 (
            .O(N__91483),
            .I(N__91103));
    InMux I__22209 (
            .O(N__91480),
            .I(N__91096));
    InMux I__22208 (
            .O(N__91479),
            .I(N__91096));
    InMux I__22207 (
            .O(N__91478),
            .I(N__91096));
    InMux I__22206 (
            .O(N__91477),
            .I(N__91093));
    LocalMux I__22205 (
            .O(N__91474),
            .I(N__91084));
    LocalMux I__22204 (
            .O(N__91471),
            .I(N__91084));
    Span4Mux_h I__22203 (
            .O(N__91462),
            .I(N__91084));
    LocalMux I__22202 (
            .O(N__91453),
            .I(N__91084));
    Span4Mux_v I__22201 (
            .O(N__91450),
            .I(N__91075));
    Span4Mux_h I__22200 (
            .O(N__91447),
            .I(N__91075));
    LocalMux I__22199 (
            .O(N__91440),
            .I(N__91075));
    LocalMux I__22198 (
            .O(N__91435),
            .I(N__91075));
    InMux I__22197 (
            .O(N__91432),
            .I(N__91072));
    LocalMux I__22196 (
            .O(N__91427),
            .I(N__91069));
    LocalMux I__22195 (
            .O(N__91422),
            .I(N__91064));
    LocalMux I__22194 (
            .O(N__91419),
            .I(N__91064));
    InMux I__22193 (
            .O(N__91418),
            .I(N__91057));
    InMux I__22192 (
            .O(N__91417),
            .I(N__91057));
    InMux I__22191 (
            .O(N__91416),
            .I(N__91057));
    Span4Mux_h I__22190 (
            .O(N__91411),
            .I(N__91052));
    LocalMux I__22189 (
            .O(N__91406),
            .I(N__91052));
    InMux I__22188 (
            .O(N__91405),
            .I(N__91047));
    InMux I__22187 (
            .O(N__91404),
            .I(N__91047));
    CascadeMux I__22186 (
            .O(N__91403),
            .I(N__91044));
    Span4Mux_v I__22185 (
            .O(N__91400),
            .I(N__91039));
    LocalMux I__22184 (
            .O(N__91397),
            .I(N__91039));
    LocalMux I__22183 (
            .O(N__91394),
            .I(N__91034));
    LocalMux I__22182 (
            .O(N__91391),
            .I(N__91034));
    Span4Mux_v I__22181 (
            .O(N__91386),
            .I(N__91027));
    LocalMux I__22180 (
            .O(N__91381),
            .I(N__91027));
    LocalMux I__22179 (
            .O(N__91378),
            .I(N__91027));
    LocalMux I__22178 (
            .O(N__91369),
            .I(N__91024));
    InMux I__22177 (
            .O(N__91368),
            .I(N__91019));
    InMux I__22176 (
            .O(N__91367),
            .I(N__91019));
    InMux I__22175 (
            .O(N__91366),
            .I(N__91012));
    InMux I__22174 (
            .O(N__91365),
            .I(N__91012));
    InMux I__22173 (
            .O(N__91364),
            .I(N__91012));
    InMux I__22172 (
            .O(N__91363),
            .I(N__91007));
    InMux I__22171 (
            .O(N__91362),
            .I(N__91007));
    LocalMux I__22170 (
            .O(N__91357),
            .I(N__91004));
    InMux I__22169 (
            .O(N__91356),
            .I(N__91001));
    InMux I__22168 (
            .O(N__91355),
            .I(N__90998));
    InMux I__22167 (
            .O(N__91354),
            .I(N__90991));
    InMux I__22166 (
            .O(N__91353),
            .I(N__90991));
    InMux I__22165 (
            .O(N__91352),
            .I(N__90991));
    InMux I__22164 (
            .O(N__91351),
            .I(N__90982));
    InMux I__22163 (
            .O(N__91350),
            .I(N__90982));
    InMux I__22162 (
            .O(N__91349),
            .I(N__90982));
    InMux I__22161 (
            .O(N__91348),
            .I(N__90982));
    InMux I__22160 (
            .O(N__91347),
            .I(N__90979));
    Span4Mux_v I__22159 (
            .O(N__91340),
            .I(N__90968));
    LocalMux I__22158 (
            .O(N__91331),
            .I(N__90968));
    InMux I__22157 (
            .O(N__91330),
            .I(N__90963));
    InMux I__22156 (
            .O(N__91329),
            .I(N__90963));
    InMux I__22155 (
            .O(N__91328),
            .I(N__90960));
    InMux I__22154 (
            .O(N__91327),
            .I(N__90953));
    InMux I__22153 (
            .O(N__91326),
            .I(N__90953));
    InMux I__22152 (
            .O(N__91325),
            .I(N__90953));
    LocalMux I__22151 (
            .O(N__91322),
            .I(N__90946));
    LocalMux I__22150 (
            .O(N__91319),
            .I(N__90946));
    LocalMux I__22149 (
            .O(N__91316),
            .I(N__90946));
    LocalMux I__22148 (
            .O(N__91309),
            .I(N__90937));
    LocalMux I__22147 (
            .O(N__91302),
            .I(N__90937));
    LocalMux I__22146 (
            .O(N__91299),
            .I(N__90937));
    LocalMux I__22145 (
            .O(N__91296),
            .I(N__90937));
    InMux I__22144 (
            .O(N__91295),
            .I(N__90930));
    InMux I__22143 (
            .O(N__91294),
            .I(N__90930));
    InMux I__22142 (
            .O(N__91293),
            .I(N__90930));
    InMux I__22141 (
            .O(N__91292),
            .I(N__90919));
    InMux I__22140 (
            .O(N__91291),
            .I(N__90919));
    InMux I__22139 (
            .O(N__91290),
            .I(N__90919));
    InMux I__22138 (
            .O(N__91289),
            .I(N__90919));
    InMux I__22137 (
            .O(N__91288),
            .I(N__90919));
    InMux I__22136 (
            .O(N__91285),
            .I(N__90910));
    InMux I__22135 (
            .O(N__91284),
            .I(N__90910));
    InMux I__22134 (
            .O(N__91283),
            .I(N__90910));
    InMux I__22133 (
            .O(N__91282),
            .I(N__90910));
    Span4Mux_h I__22132 (
            .O(N__91275),
            .I(N__90895));
    Span4Mux_v I__22131 (
            .O(N__91268),
            .I(N__90895));
    LocalMux I__22130 (
            .O(N__91265),
            .I(N__90895));
    Span4Mux_h I__22129 (
            .O(N__91256),
            .I(N__90895));
    LocalMux I__22128 (
            .O(N__91251),
            .I(N__90895));
    Span4Mux_v I__22127 (
            .O(N__91246),
            .I(N__90895));
    LocalMux I__22126 (
            .O(N__91243),
            .I(N__90895));
    InMux I__22125 (
            .O(N__91242),
            .I(N__90892));
    InMux I__22124 (
            .O(N__91241),
            .I(N__90885));
    InMux I__22123 (
            .O(N__91240),
            .I(N__90885));
    InMux I__22122 (
            .O(N__91239),
            .I(N__90885));
    InMux I__22121 (
            .O(N__91238),
            .I(N__90882));
    CascadeMux I__22120 (
            .O(N__91237),
            .I(N__90879));
    InMux I__22119 (
            .O(N__91236),
            .I(N__90873));
    InMux I__22118 (
            .O(N__91235),
            .I(N__90873));
    InMux I__22117 (
            .O(N__91234),
            .I(N__90860));
    InMux I__22116 (
            .O(N__91231),
            .I(N__90860));
    InMux I__22115 (
            .O(N__91230),
            .I(N__90860));
    InMux I__22114 (
            .O(N__91229),
            .I(N__90860));
    InMux I__22113 (
            .O(N__91228),
            .I(N__90850));
    InMux I__22112 (
            .O(N__91227),
            .I(N__90841));
    InMux I__22111 (
            .O(N__91226),
            .I(N__90841));
    InMux I__22110 (
            .O(N__91225),
            .I(N__90841));
    InMux I__22109 (
            .O(N__91224),
            .I(N__90841));
    InMux I__22108 (
            .O(N__91223),
            .I(N__90836));
    InMux I__22107 (
            .O(N__91222),
            .I(N__90836));
    InMux I__22106 (
            .O(N__91221),
            .I(N__90833));
    Span4Mux_v I__22105 (
            .O(N__91214),
            .I(N__90830));
    Span4Mux_v I__22104 (
            .O(N__91209),
            .I(N__90825));
    LocalMux I__22103 (
            .O(N__91204),
            .I(N__90825));
    Span4Mux_v I__22102 (
            .O(N__91195),
            .I(N__90816));
    Span4Mux_h I__22101 (
            .O(N__91188),
            .I(N__90816));
    LocalMux I__22100 (
            .O(N__91185),
            .I(N__90816));
    LocalMux I__22099 (
            .O(N__91180),
            .I(N__90816));
    Span4Mux_h I__22098 (
            .O(N__91175),
            .I(N__90811));
    LocalMux I__22097 (
            .O(N__91164),
            .I(N__90811));
    LocalMux I__22096 (
            .O(N__91161),
            .I(N__90800));
    Span4Mux_v I__22095 (
            .O(N__91158),
            .I(N__90800));
    LocalMux I__22094 (
            .O(N__91155),
            .I(N__90800));
    LocalMux I__22093 (
            .O(N__91146),
            .I(N__90800));
    LocalMux I__22092 (
            .O(N__91139),
            .I(N__90800));
    Span4Mux_h I__22091 (
            .O(N__91132),
            .I(N__90791));
    Span4Mux_h I__22090 (
            .O(N__91127),
            .I(N__90791));
    Span4Mux_v I__22089 (
            .O(N__91118),
            .I(N__90791));
    LocalMux I__22088 (
            .O(N__91115),
            .I(N__90791));
    LocalMux I__22087 (
            .O(N__91112),
            .I(N__90788));
    InMux I__22086 (
            .O(N__91111),
            .I(N__90783));
    InMux I__22085 (
            .O(N__91110),
            .I(N__90783));
    Span4Mux_h I__22084 (
            .O(N__91103),
            .I(N__90776));
    LocalMux I__22083 (
            .O(N__91096),
            .I(N__90776));
    LocalMux I__22082 (
            .O(N__91093),
            .I(N__90776));
    Span4Mux_v I__22081 (
            .O(N__91084),
            .I(N__90759));
    Span4Mux_h I__22080 (
            .O(N__91075),
            .I(N__90759));
    LocalMux I__22079 (
            .O(N__91072),
            .I(N__90759));
    Span4Mux_v I__22078 (
            .O(N__91069),
            .I(N__90759));
    Span4Mux_v I__22077 (
            .O(N__91064),
            .I(N__90759));
    LocalMux I__22076 (
            .O(N__91057),
            .I(N__90759));
    Span4Mux_h I__22075 (
            .O(N__91052),
            .I(N__90759));
    LocalMux I__22074 (
            .O(N__91047),
            .I(N__90759));
    InMux I__22073 (
            .O(N__91044),
            .I(N__90756));
    Span4Mux_h I__22072 (
            .O(N__91039),
            .I(N__90741));
    Span4Mux_v I__22071 (
            .O(N__91034),
            .I(N__90741));
    Span4Mux_v I__22070 (
            .O(N__91027),
            .I(N__90741));
    Span4Mux_v I__22069 (
            .O(N__91024),
            .I(N__90741));
    LocalMux I__22068 (
            .O(N__91019),
            .I(N__90741));
    LocalMux I__22067 (
            .O(N__91012),
            .I(N__90741));
    LocalMux I__22066 (
            .O(N__91007),
            .I(N__90741));
    Span4Mux_h I__22065 (
            .O(N__91004),
            .I(N__90728));
    LocalMux I__22064 (
            .O(N__91001),
            .I(N__90728));
    LocalMux I__22063 (
            .O(N__90998),
            .I(N__90728));
    LocalMux I__22062 (
            .O(N__90991),
            .I(N__90728));
    LocalMux I__22061 (
            .O(N__90982),
            .I(N__90728));
    LocalMux I__22060 (
            .O(N__90979),
            .I(N__90728));
    InMux I__22059 (
            .O(N__90978),
            .I(N__90723));
    InMux I__22058 (
            .O(N__90977),
            .I(N__90723));
    InMux I__22057 (
            .O(N__90976),
            .I(N__90718));
    InMux I__22056 (
            .O(N__90975),
            .I(N__90718));
    InMux I__22055 (
            .O(N__90974),
            .I(N__90713));
    InMux I__22054 (
            .O(N__90973),
            .I(N__90713));
    Span4Mux_h I__22053 (
            .O(N__90968),
            .I(N__90696));
    LocalMux I__22052 (
            .O(N__90963),
            .I(N__90696));
    LocalMux I__22051 (
            .O(N__90960),
            .I(N__90696));
    LocalMux I__22050 (
            .O(N__90953),
            .I(N__90696));
    Span4Mux_v I__22049 (
            .O(N__90946),
            .I(N__90685));
    Span4Mux_h I__22048 (
            .O(N__90937),
            .I(N__90685));
    LocalMux I__22047 (
            .O(N__90930),
            .I(N__90685));
    LocalMux I__22046 (
            .O(N__90919),
            .I(N__90685));
    LocalMux I__22045 (
            .O(N__90910),
            .I(N__90685));
    Span4Mux_h I__22044 (
            .O(N__90895),
            .I(N__90676));
    LocalMux I__22043 (
            .O(N__90892),
            .I(N__90676));
    LocalMux I__22042 (
            .O(N__90885),
            .I(N__90676));
    LocalMux I__22041 (
            .O(N__90882),
            .I(N__90676));
    InMux I__22040 (
            .O(N__90879),
            .I(N__90671));
    InMux I__22039 (
            .O(N__90878),
            .I(N__90671));
    LocalMux I__22038 (
            .O(N__90873),
            .I(N__90668));
    InMux I__22037 (
            .O(N__90872),
            .I(N__90663));
    InMux I__22036 (
            .O(N__90871),
            .I(N__90663));
    InMux I__22035 (
            .O(N__90870),
            .I(N__90658));
    InMux I__22034 (
            .O(N__90869),
            .I(N__90658));
    LocalMux I__22033 (
            .O(N__90860),
            .I(N__90655));
    InMux I__22032 (
            .O(N__90859),
            .I(N__90652));
    InMux I__22031 (
            .O(N__90858),
            .I(N__90649));
    InMux I__22030 (
            .O(N__90857),
            .I(N__90646));
    InMux I__22029 (
            .O(N__90856),
            .I(N__90641));
    InMux I__22028 (
            .O(N__90855),
            .I(N__90641));
    InMux I__22027 (
            .O(N__90854),
            .I(N__90636));
    InMux I__22026 (
            .O(N__90853),
            .I(N__90636));
    LocalMux I__22025 (
            .O(N__90850),
            .I(N__90627));
    LocalMux I__22024 (
            .O(N__90841),
            .I(N__90627));
    LocalMux I__22023 (
            .O(N__90836),
            .I(N__90627));
    LocalMux I__22022 (
            .O(N__90833),
            .I(N__90624));
    Span4Mux_v I__22021 (
            .O(N__90830),
            .I(N__90619));
    Span4Mux_v I__22020 (
            .O(N__90825),
            .I(N__90619));
    Span4Mux_h I__22019 (
            .O(N__90816),
            .I(N__90616));
    Span4Mux_h I__22018 (
            .O(N__90811),
            .I(N__90611));
    Span4Mux_v I__22017 (
            .O(N__90800),
            .I(N__90611));
    Span4Mux_h I__22016 (
            .O(N__90791),
            .I(N__90608));
    Span4Mux_h I__22015 (
            .O(N__90788),
            .I(N__90603));
    LocalMux I__22014 (
            .O(N__90783),
            .I(N__90603));
    Span4Mux_h I__22013 (
            .O(N__90776),
            .I(N__90600));
    Span4Mux_h I__22012 (
            .O(N__90759),
            .I(N__90595));
    LocalMux I__22011 (
            .O(N__90756),
            .I(N__90595));
    Span4Mux_h I__22010 (
            .O(N__90741),
            .I(N__90588));
    Span4Mux_v I__22009 (
            .O(N__90728),
            .I(N__90588));
    LocalMux I__22008 (
            .O(N__90723),
            .I(N__90588));
    LocalMux I__22007 (
            .O(N__90718),
            .I(N__90583));
    LocalMux I__22006 (
            .O(N__90713),
            .I(N__90583));
    InMux I__22005 (
            .O(N__90712),
            .I(N__90576));
    InMux I__22004 (
            .O(N__90711),
            .I(N__90576));
    InMux I__22003 (
            .O(N__90710),
            .I(N__90576));
    InMux I__22002 (
            .O(N__90709),
            .I(N__90567));
    InMux I__22001 (
            .O(N__90708),
            .I(N__90567));
    InMux I__22000 (
            .O(N__90707),
            .I(N__90567));
    InMux I__21999 (
            .O(N__90706),
            .I(N__90567));
    InMux I__21998 (
            .O(N__90705),
            .I(N__90564));
    Span4Mux_h I__21997 (
            .O(N__90696),
            .I(N__90561));
    Span4Mux_h I__21996 (
            .O(N__90685),
            .I(N__90554));
    Span4Mux_v I__21995 (
            .O(N__90676),
            .I(N__90554));
    LocalMux I__21994 (
            .O(N__90671),
            .I(N__90554));
    Sp12to4 I__21993 (
            .O(N__90668),
            .I(N__90547));
    LocalMux I__21992 (
            .O(N__90663),
            .I(N__90547));
    LocalMux I__21991 (
            .O(N__90658),
            .I(N__90547));
    Span12Mux_h I__21990 (
            .O(N__90655),
            .I(N__90534));
    LocalMux I__21989 (
            .O(N__90652),
            .I(N__90534));
    LocalMux I__21988 (
            .O(N__90649),
            .I(N__90534));
    LocalMux I__21987 (
            .O(N__90646),
            .I(N__90534));
    LocalMux I__21986 (
            .O(N__90641),
            .I(N__90534));
    LocalMux I__21985 (
            .O(N__90636),
            .I(N__90534));
    InMux I__21984 (
            .O(N__90635),
            .I(N__90529));
    InMux I__21983 (
            .O(N__90634),
            .I(N__90529));
    Span12Mux_h I__21982 (
            .O(N__90627),
            .I(N__90522));
    Span12Mux_v I__21981 (
            .O(N__90624),
            .I(N__90522));
    Span4Mux_v I__21980 (
            .O(N__90619),
            .I(N__90517));
    Span4Mux_h I__21979 (
            .O(N__90616),
            .I(N__90517));
    Span4Mux_h I__21978 (
            .O(N__90611),
            .I(N__90510));
    Span4Mux_v I__21977 (
            .O(N__90608),
            .I(N__90510));
    Span4Mux_v I__21976 (
            .O(N__90603),
            .I(N__90510));
    Span4Mux_h I__21975 (
            .O(N__90600),
            .I(N__90503));
    Span4Mux_v I__21974 (
            .O(N__90595),
            .I(N__90503));
    Span4Mux_h I__21973 (
            .O(N__90588),
            .I(N__90503));
    Span12Mux_v I__21972 (
            .O(N__90583),
            .I(N__90494));
    LocalMux I__21971 (
            .O(N__90576),
            .I(N__90494));
    LocalMux I__21970 (
            .O(N__90567),
            .I(N__90494));
    LocalMux I__21969 (
            .O(N__90564),
            .I(N__90494));
    Span4Mux_h I__21968 (
            .O(N__90561),
            .I(N__90489));
    Span4Mux_v I__21967 (
            .O(N__90554),
            .I(N__90489));
    Span12Mux_s11_v I__21966 (
            .O(N__90547),
            .I(N__90482));
    Span12Mux_v I__21965 (
            .O(N__90534),
            .I(N__90482));
    LocalMux I__21964 (
            .O(N__90529),
            .I(N__90482));
    InMux I__21963 (
            .O(N__90528),
            .I(N__90477));
    InMux I__21962 (
            .O(N__90527),
            .I(N__90477));
    Odrv12 I__21961 (
            .O(N__90522),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1 ));
    Odrv4 I__21960 (
            .O(N__90517),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1 ));
    Odrv4 I__21959 (
            .O(N__90510),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1 ));
    Odrv4 I__21958 (
            .O(N__90503),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1 ));
    Odrv12 I__21957 (
            .O(N__90494),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1 ));
    Odrv4 I__21956 (
            .O(N__90489),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1 ));
    Odrv12 I__21955 (
            .O(N__90482),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1 ));
    LocalMux I__21954 (
            .O(N__90477),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1 ));
    CascadeMux I__21953 (
            .O(N__90460),
            .I(N__90457));
    InMux I__21952 (
            .O(N__90457),
            .I(N__90454));
    LocalMux I__21951 (
            .O(N__90454),
            .I(N__90451));
    Span4Mux_h I__21950 (
            .O(N__90451),
            .I(N__90448));
    Span4Mux_h I__21949 (
            .O(N__90448),
            .I(N__90445));
    Odrv4 I__21948 (
            .O(N__90445),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14012 ));
    InMux I__21947 (
            .O(N__90442),
            .I(N__90439));
    LocalMux I__21946 (
            .O(N__90439),
            .I(N__90436));
    Span4Mux_v I__21945 (
            .O(N__90436),
            .I(N__90432));
    CascadeMux I__21944 (
            .O(N__90435),
            .I(N__90429));
    Sp12to4 I__21943 (
            .O(N__90432),
            .I(N__90426));
    InMux I__21942 (
            .O(N__90429),
            .I(N__90423));
    Odrv12 I__21941 (
            .O(N__90426),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_8 ));
    LocalMux I__21940 (
            .O(N__90423),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_8 ));
    InMux I__21939 (
            .O(N__90418),
            .I(N__90415));
    LocalMux I__21938 (
            .O(N__90415),
            .I(N__90412));
    Span4Mux_v I__21937 (
            .O(N__90412),
            .I(N__90409));
    Odrv4 I__21936 (
            .O(N__90409),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11736 ));
    InMux I__21935 (
            .O(N__90406),
            .I(N__90403));
    LocalMux I__21934 (
            .O(N__90403),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13304 ));
    CascadeMux I__21933 (
            .O(N__90400),
            .I(N__90395));
    CascadeMux I__21932 (
            .O(N__90399),
            .I(N__90392));
    InMux I__21931 (
            .O(N__90398),
            .I(N__90382));
    InMux I__21930 (
            .O(N__90395),
            .I(N__90379));
    InMux I__21929 (
            .O(N__90392),
            .I(N__90370));
    InMux I__21928 (
            .O(N__90391),
            .I(N__90370));
    InMux I__21927 (
            .O(N__90390),
            .I(N__90370));
    InMux I__21926 (
            .O(N__90389),
            .I(N__90370));
    InMux I__21925 (
            .O(N__90388),
            .I(N__90366));
    InMux I__21924 (
            .O(N__90387),
            .I(N__90363));
    InMux I__21923 (
            .O(N__90386),
            .I(N__90359));
    CascadeMux I__21922 (
            .O(N__90385),
            .I(N__90356));
    LocalMux I__21921 (
            .O(N__90382),
            .I(N__90344));
    LocalMux I__21920 (
            .O(N__90379),
            .I(N__90336));
    LocalMux I__21919 (
            .O(N__90370),
            .I(N__90333));
    InMux I__21918 (
            .O(N__90369),
            .I(N__90330));
    LocalMux I__21917 (
            .O(N__90366),
            .I(N__90325));
    LocalMux I__21916 (
            .O(N__90363),
            .I(N__90325));
    InMux I__21915 (
            .O(N__90362),
            .I(N__90322));
    LocalMux I__21914 (
            .O(N__90359),
            .I(N__90319));
    InMux I__21913 (
            .O(N__90356),
            .I(N__90312));
    InMux I__21912 (
            .O(N__90355),
            .I(N__90312));
    InMux I__21911 (
            .O(N__90354),
            .I(N__90312));
    InMux I__21910 (
            .O(N__90353),
            .I(N__90309));
    InMux I__21909 (
            .O(N__90352),
            .I(N__90306));
    InMux I__21908 (
            .O(N__90351),
            .I(N__90303));
    CascadeMux I__21907 (
            .O(N__90350),
            .I(N__90297));
    InMux I__21906 (
            .O(N__90349),
            .I(N__90294));
    InMux I__21905 (
            .O(N__90348),
            .I(N__90291));
    InMux I__21904 (
            .O(N__90347),
            .I(N__90287));
    Span4Mux_h I__21903 (
            .O(N__90344),
            .I(N__90284));
    InMux I__21902 (
            .O(N__90343),
            .I(N__90279));
    InMux I__21901 (
            .O(N__90342),
            .I(N__90279));
    InMux I__21900 (
            .O(N__90341),
            .I(N__90276));
    InMux I__21899 (
            .O(N__90340),
            .I(N__90273));
    InMux I__21898 (
            .O(N__90339),
            .I(N__90270));
    Span4Mux_h I__21897 (
            .O(N__90336),
            .I(N__90267));
    Span4Mux_v I__21896 (
            .O(N__90333),
            .I(N__90262));
    LocalMux I__21895 (
            .O(N__90330),
            .I(N__90262));
    Span4Mux_v I__21894 (
            .O(N__90325),
            .I(N__90257));
    LocalMux I__21893 (
            .O(N__90322),
            .I(N__90257));
    Span4Mux_h I__21892 (
            .O(N__90319),
            .I(N__90254));
    LocalMux I__21891 (
            .O(N__90312),
            .I(N__90245));
    LocalMux I__21890 (
            .O(N__90309),
            .I(N__90245));
    LocalMux I__21889 (
            .O(N__90306),
            .I(N__90242));
    LocalMux I__21888 (
            .O(N__90303),
            .I(N__90239));
    InMux I__21887 (
            .O(N__90302),
            .I(N__90236));
    InMux I__21886 (
            .O(N__90301),
            .I(N__90233));
    InMux I__21885 (
            .O(N__90300),
            .I(N__90226));
    InMux I__21884 (
            .O(N__90297),
            .I(N__90223));
    LocalMux I__21883 (
            .O(N__90294),
            .I(N__90216));
    LocalMux I__21882 (
            .O(N__90291),
            .I(N__90216));
    CascadeMux I__21881 (
            .O(N__90290),
            .I(N__90213));
    LocalMux I__21880 (
            .O(N__90287),
            .I(N__90207));
    Span4Mux_h I__21879 (
            .O(N__90284),
            .I(N__90202));
    LocalMux I__21878 (
            .O(N__90279),
            .I(N__90202));
    LocalMux I__21877 (
            .O(N__90276),
            .I(N__90199));
    LocalMux I__21876 (
            .O(N__90273),
            .I(N__90196));
    LocalMux I__21875 (
            .O(N__90270),
            .I(N__90193));
    Span4Mux_h I__21874 (
            .O(N__90267),
            .I(N__90186));
    Span4Mux_h I__21873 (
            .O(N__90262),
            .I(N__90186));
    Span4Mux_v I__21872 (
            .O(N__90257),
            .I(N__90186));
    Span4Mux_v I__21871 (
            .O(N__90254),
            .I(N__90183));
    InMux I__21870 (
            .O(N__90253),
            .I(N__90174));
    InMux I__21869 (
            .O(N__90252),
            .I(N__90174));
    InMux I__21868 (
            .O(N__90251),
            .I(N__90174));
    InMux I__21867 (
            .O(N__90250),
            .I(N__90174));
    Span4Mux_h I__21866 (
            .O(N__90245),
            .I(N__90171));
    Span4Mux_v I__21865 (
            .O(N__90242),
            .I(N__90164));
    Span4Mux_h I__21864 (
            .O(N__90239),
            .I(N__90164));
    LocalMux I__21863 (
            .O(N__90236),
            .I(N__90164));
    LocalMux I__21862 (
            .O(N__90233),
            .I(N__90161));
    InMux I__21861 (
            .O(N__90232),
            .I(N__90158));
    InMux I__21860 (
            .O(N__90231),
            .I(N__90155));
    InMux I__21859 (
            .O(N__90230),
            .I(N__90152));
    CascadeMux I__21858 (
            .O(N__90229),
            .I(N__90149));
    LocalMux I__21857 (
            .O(N__90226),
            .I(N__90144));
    LocalMux I__21856 (
            .O(N__90223),
            .I(N__90144));
    InMux I__21855 (
            .O(N__90222),
            .I(N__90138));
    InMux I__21854 (
            .O(N__90221),
            .I(N__90135));
    Span4Mux_h I__21853 (
            .O(N__90216),
            .I(N__90131));
    InMux I__21852 (
            .O(N__90213),
            .I(N__90122));
    InMux I__21851 (
            .O(N__90212),
            .I(N__90122));
    InMux I__21850 (
            .O(N__90211),
            .I(N__90122));
    InMux I__21849 (
            .O(N__90210),
            .I(N__90122));
    Span4Mux_v I__21848 (
            .O(N__90207),
            .I(N__90119));
    Span4Mux_h I__21847 (
            .O(N__90202),
            .I(N__90116));
    Span4Mux_v I__21846 (
            .O(N__90199),
            .I(N__90109));
    Span4Mux_h I__21845 (
            .O(N__90196),
            .I(N__90109));
    Span4Mux_v I__21844 (
            .O(N__90193),
            .I(N__90109));
    Span4Mux_v I__21843 (
            .O(N__90186),
            .I(N__90102));
    Span4Mux_v I__21842 (
            .O(N__90183),
            .I(N__90102));
    LocalMux I__21841 (
            .O(N__90174),
            .I(N__90102));
    Span4Mux_v I__21840 (
            .O(N__90171),
            .I(N__90096));
    Span4Mux_h I__21839 (
            .O(N__90164),
            .I(N__90096));
    Span4Mux_v I__21838 (
            .O(N__90161),
            .I(N__90093));
    LocalMux I__21837 (
            .O(N__90158),
            .I(N__90090));
    LocalMux I__21836 (
            .O(N__90155),
            .I(N__90085));
    LocalMux I__21835 (
            .O(N__90152),
            .I(N__90085));
    InMux I__21834 (
            .O(N__90149),
            .I(N__90077));
    Span4Mux_v I__21833 (
            .O(N__90144),
            .I(N__90074));
    InMux I__21832 (
            .O(N__90143),
            .I(N__90067));
    InMux I__21831 (
            .O(N__90142),
            .I(N__90067));
    InMux I__21830 (
            .O(N__90141),
            .I(N__90067));
    LocalMux I__21829 (
            .O(N__90138),
            .I(N__90062));
    LocalMux I__21828 (
            .O(N__90135),
            .I(N__90059));
    InMux I__21827 (
            .O(N__90134),
            .I(N__90056));
    Span4Mux_v I__21826 (
            .O(N__90131),
            .I(N__90048));
    LocalMux I__21825 (
            .O(N__90122),
            .I(N__90048));
    Span4Mux_v I__21824 (
            .O(N__90119),
            .I(N__90039));
    Span4Mux_h I__21823 (
            .O(N__90116),
            .I(N__90039));
    Span4Mux_h I__21822 (
            .O(N__90109),
            .I(N__90039));
    Span4Mux_h I__21821 (
            .O(N__90102),
            .I(N__90039));
    InMux I__21820 (
            .O(N__90101),
            .I(N__90036));
    Span4Mux_h I__21819 (
            .O(N__90096),
            .I(N__90029));
    Span4Mux_v I__21818 (
            .O(N__90093),
            .I(N__90029));
    Span4Mux_v I__21817 (
            .O(N__90090),
            .I(N__90026));
    Span4Mux_v I__21816 (
            .O(N__90085),
            .I(N__90023));
    InMux I__21815 (
            .O(N__90084),
            .I(N__90019));
    InMux I__21814 (
            .O(N__90083),
            .I(N__90009));
    InMux I__21813 (
            .O(N__90082),
            .I(N__90009));
    InMux I__21812 (
            .O(N__90081),
            .I(N__90009));
    InMux I__21811 (
            .O(N__90080),
            .I(N__90009));
    LocalMux I__21810 (
            .O(N__90077),
            .I(N__90006));
    Span4Mux_v I__21809 (
            .O(N__90074),
            .I(N__90001));
    LocalMux I__21808 (
            .O(N__90067),
            .I(N__90001));
    InMux I__21807 (
            .O(N__90066),
            .I(N__89996));
    InMux I__21806 (
            .O(N__90065),
            .I(N__89996));
    Span4Mux_v I__21805 (
            .O(N__90062),
            .I(N__89993));
    Span4Mux_h I__21804 (
            .O(N__90059),
            .I(N__89988));
    LocalMux I__21803 (
            .O(N__90056),
            .I(N__89988));
    InMux I__21802 (
            .O(N__90055),
            .I(N__89985));
    InMux I__21801 (
            .O(N__90054),
            .I(N__89982));
    InMux I__21800 (
            .O(N__90053),
            .I(N__89979));
    Span4Mux_v I__21799 (
            .O(N__90048),
            .I(N__89975));
    Span4Mux_h I__21798 (
            .O(N__90039),
            .I(N__89970));
    LocalMux I__21797 (
            .O(N__90036),
            .I(N__89970));
    InMux I__21796 (
            .O(N__90035),
            .I(N__89965));
    InMux I__21795 (
            .O(N__90034),
            .I(N__89965));
    Span4Mux_h I__21794 (
            .O(N__90029),
            .I(N__89957));
    Span4Mux_v I__21793 (
            .O(N__90026),
            .I(N__89957));
    Span4Mux_v I__21792 (
            .O(N__90023),
            .I(N__89957));
    InMux I__21791 (
            .O(N__90022),
            .I(N__89954));
    LocalMux I__21790 (
            .O(N__90019),
            .I(N__89950));
    InMux I__21789 (
            .O(N__90018),
            .I(N__89947));
    LocalMux I__21788 (
            .O(N__90009),
            .I(N__89939));
    Span4Mux_v I__21787 (
            .O(N__90006),
            .I(N__89932));
    Span4Mux_v I__21786 (
            .O(N__90001),
            .I(N__89932));
    LocalMux I__21785 (
            .O(N__89996),
            .I(N__89932));
    Span4Mux_v I__21784 (
            .O(N__89993),
            .I(N__89921));
    Span4Mux_h I__21783 (
            .O(N__89988),
            .I(N__89921));
    LocalMux I__21782 (
            .O(N__89985),
            .I(N__89921));
    LocalMux I__21781 (
            .O(N__89982),
            .I(N__89921));
    LocalMux I__21780 (
            .O(N__89979),
            .I(N__89921));
    InMux I__21779 (
            .O(N__89978),
            .I(N__89918));
    Span4Mux_v I__21778 (
            .O(N__89975),
            .I(N__89915));
    Span4Mux_v I__21777 (
            .O(N__89970),
            .I(N__89910));
    LocalMux I__21776 (
            .O(N__89965),
            .I(N__89910));
    InMux I__21775 (
            .O(N__89964),
            .I(N__89907));
    Span4Mux_h I__21774 (
            .O(N__89957),
            .I(N__89900));
    LocalMux I__21773 (
            .O(N__89954),
            .I(N__89900));
    InMux I__21772 (
            .O(N__89953),
            .I(N__89897));
    Span4Mux_h I__21771 (
            .O(N__89950),
            .I(N__89892));
    LocalMux I__21770 (
            .O(N__89947),
            .I(N__89892));
    InMux I__21769 (
            .O(N__89946),
            .I(N__89883));
    InMux I__21768 (
            .O(N__89945),
            .I(N__89883));
    InMux I__21767 (
            .O(N__89944),
            .I(N__89883));
    InMux I__21766 (
            .O(N__89943),
            .I(N__89883));
    InMux I__21765 (
            .O(N__89942),
            .I(N__89877));
    Span12Mux_v I__21764 (
            .O(N__89939),
            .I(N__89873));
    Span4Mux_h I__21763 (
            .O(N__89932),
            .I(N__89868));
    Span4Mux_v I__21762 (
            .O(N__89921),
            .I(N__89868));
    LocalMux I__21761 (
            .O(N__89918),
            .I(N__89865));
    Span4Mux_v I__21760 (
            .O(N__89915),
            .I(N__89862));
    Sp12to4 I__21759 (
            .O(N__89910),
            .I(N__89857));
    LocalMux I__21758 (
            .O(N__89907),
            .I(N__89857));
    InMux I__21757 (
            .O(N__89906),
            .I(N__89854));
    InMux I__21756 (
            .O(N__89905),
            .I(N__89851));
    Span4Mux_v I__21755 (
            .O(N__89900),
            .I(N__89845));
    LocalMux I__21754 (
            .O(N__89897),
            .I(N__89845));
    Span4Mux_v I__21753 (
            .O(N__89892),
            .I(N__89840));
    LocalMux I__21752 (
            .O(N__89883),
            .I(N__89840));
    InMux I__21751 (
            .O(N__89882),
            .I(N__89833));
    InMux I__21750 (
            .O(N__89881),
            .I(N__89833));
    InMux I__21749 (
            .O(N__89880),
            .I(N__89833));
    LocalMux I__21748 (
            .O(N__89877),
            .I(N__89830));
    InMux I__21747 (
            .O(N__89876),
            .I(N__89827));
    Span12Mux_h I__21746 (
            .O(N__89873),
            .I(N__89822));
    Span4Mux_v I__21745 (
            .O(N__89868),
            .I(N__89817));
    Span4Mux_v I__21744 (
            .O(N__89865),
            .I(N__89817));
    Sp12to4 I__21743 (
            .O(N__89862),
            .I(N__89808));
    Span12Mux_v I__21742 (
            .O(N__89857),
            .I(N__89808));
    LocalMux I__21741 (
            .O(N__89854),
            .I(N__89808));
    LocalMux I__21740 (
            .O(N__89851),
            .I(N__89808));
    InMux I__21739 (
            .O(N__89850),
            .I(N__89805));
    Span4Mux_v I__21738 (
            .O(N__89845),
            .I(N__89794));
    Span4Mux_h I__21737 (
            .O(N__89840),
            .I(N__89794));
    LocalMux I__21736 (
            .O(N__89833),
            .I(N__89794));
    Span4Mux_h I__21735 (
            .O(N__89830),
            .I(N__89794));
    LocalMux I__21734 (
            .O(N__89827),
            .I(N__89794));
    InMux I__21733 (
            .O(N__89826),
            .I(N__89789));
    InMux I__21732 (
            .O(N__89825),
            .I(N__89789));
    Odrv12 I__21731 (
            .O(N__89822),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3 ));
    Odrv4 I__21730 (
            .O(N__89817),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3 ));
    Odrv12 I__21729 (
            .O(N__89808),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3 ));
    LocalMux I__21728 (
            .O(N__89805),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3 ));
    Odrv4 I__21727 (
            .O(N__89794),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3 ));
    LocalMux I__21726 (
            .O(N__89789),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3 ));
    CascadeMux I__21725 (
            .O(N__89776),
            .I(N__89773));
    InMux I__21724 (
            .O(N__89773),
            .I(N__89770));
    LocalMux I__21723 (
            .O(N__89770),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13073 ));
    InMux I__21722 (
            .O(N__89767),
            .I(N__89764));
    LocalMux I__21721 (
            .O(N__89764),
            .I(N__89761));
    Odrv12 I__21720 (
            .O(N__89761),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12827 ));
    InMux I__21719 (
            .O(N__89758),
            .I(N__89755));
    LocalMux I__21718 (
            .O(N__89755),
            .I(N__89752));
    Odrv4 I__21717 (
            .O(N__89752),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11880 ));
    InMux I__21716 (
            .O(N__89749),
            .I(N__89745));
    InMux I__21715 (
            .O(N__89748),
            .I(N__89742));
    LocalMux I__21714 (
            .O(N__89745),
            .I(\pc_tx.r_Clock_Count_0 ));
    LocalMux I__21713 (
            .O(N__89742),
            .I(\pc_tx.r_Clock_Count_0 ));
    InMux I__21712 (
            .O(N__89737),
            .I(bfn_24_11_0_));
    InMux I__21711 (
            .O(N__89734),
            .I(N__89730));
    InMux I__21710 (
            .O(N__89733),
            .I(N__89727));
    LocalMux I__21709 (
            .O(N__89730),
            .I(\pc_tx.r_Clock_Count_1 ));
    LocalMux I__21708 (
            .O(N__89727),
            .I(\pc_tx.r_Clock_Count_1 ));
    InMux I__21707 (
            .O(N__89722),
            .I(\pc_tx.n10712 ));
    InMux I__21706 (
            .O(N__89719),
            .I(N__89716));
    LocalMux I__21705 (
            .O(N__89716),
            .I(N__89712));
    InMux I__21704 (
            .O(N__89715),
            .I(N__89709));
    Odrv12 I__21703 (
            .O(N__89712),
            .I(REG_mem_44_8));
    LocalMux I__21702 (
            .O(N__89709),
            .I(REG_mem_44_8));
    CascadeMux I__21701 (
            .O(N__89704),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13640_cascade_ ));
    InMux I__21700 (
            .O(N__89701),
            .I(N__89698));
    LocalMux I__21699 (
            .O(N__89698),
            .I(N__89695));
    Span4Mux_v I__21698 (
            .O(N__89695),
            .I(N__89691));
    CascadeMux I__21697 (
            .O(N__89694),
            .I(N__89688));
    Span4Mux_h I__21696 (
            .O(N__89691),
            .I(N__89685));
    InMux I__21695 (
            .O(N__89688),
            .I(N__89682));
    Odrv4 I__21694 (
            .O(N__89685),
            .I(REG_mem_45_8));
    LocalMux I__21693 (
            .O(N__89682),
            .I(REG_mem_45_8));
    InMux I__21692 (
            .O(N__89677),
            .I(N__89674));
    LocalMux I__21691 (
            .O(N__89674),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11820 ));
    InMux I__21690 (
            .O(N__89671),
            .I(N__89667));
    InMux I__21689 (
            .O(N__89670),
            .I(N__89664));
    LocalMux I__21688 (
            .O(N__89667),
            .I(N__89658));
    LocalMux I__21687 (
            .O(N__89664),
            .I(N__89655));
    InMux I__21686 (
            .O(N__89663),
            .I(N__89652));
    InMux I__21685 (
            .O(N__89662),
            .I(N__89646));
    InMux I__21684 (
            .O(N__89661),
            .I(N__89643));
    Span4Mux_v I__21683 (
            .O(N__89658),
            .I(N__89639));
    Span4Mux_v I__21682 (
            .O(N__89655),
            .I(N__89636));
    LocalMux I__21681 (
            .O(N__89652),
            .I(N__89633));
    InMux I__21680 (
            .O(N__89651),
            .I(N__89630));
    InMux I__21679 (
            .O(N__89650),
            .I(N__89627));
    InMux I__21678 (
            .O(N__89649),
            .I(N__89621));
    LocalMux I__21677 (
            .O(N__89646),
            .I(N__89616));
    LocalMux I__21676 (
            .O(N__89643),
            .I(N__89616));
    InMux I__21675 (
            .O(N__89642),
            .I(N__89613));
    Span4Mux_v I__21674 (
            .O(N__89639),
            .I(N__89604));
    Span4Mux_h I__21673 (
            .O(N__89636),
            .I(N__89604));
    Span4Mux_h I__21672 (
            .O(N__89633),
            .I(N__89601));
    LocalMux I__21671 (
            .O(N__89630),
            .I(N__89596));
    LocalMux I__21670 (
            .O(N__89627),
            .I(N__89596));
    InMux I__21669 (
            .O(N__89626),
            .I(N__89589));
    InMux I__21668 (
            .O(N__89625),
            .I(N__89589));
    InMux I__21667 (
            .O(N__89624),
            .I(N__89589));
    LocalMux I__21666 (
            .O(N__89621),
            .I(N__89586));
    Span12Mux_h I__21665 (
            .O(N__89616),
            .I(N__89581));
    LocalMux I__21664 (
            .O(N__89613),
            .I(N__89581));
    InMux I__21663 (
            .O(N__89612),
            .I(N__89578));
    InMux I__21662 (
            .O(N__89611),
            .I(N__89573));
    InMux I__21661 (
            .O(N__89610),
            .I(N__89573));
    InMux I__21660 (
            .O(N__89609),
            .I(N__89570));
    Odrv4 I__21659 (
            .O(N__89604),
            .I(n58));
    Odrv4 I__21658 (
            .O(N__89601),
            .I(n58));
    Odrv12 I__21657 (
            .O(N__89596),
            .I(n58));
    LocalMux I__21656 (
            .O(N__89589),
            .I(n58));
    Odrv4 I__21655 (
            .O(N__89586),
            .I(n58));
    Odrv12 I__21654 (
            .O(N__89581),
            .I(n58));
    LocalMux I__21653 (
            .O(N__89578),
            .I(n58));
    LocalMux I__21652 (
            .O(N__89573),
            .I(n58));
    LocalMux I__21651 (
            .O(N__89570),
            .I(n58));
    InMux I__21650 (
            .O(N__89551),
            .I(N__89548));
    LocalMux I__21649 (
            .O(N__89548),
            .I(N__89545));
    Span4Mux_v I__21648 (
            .O(N__89545),
            .I(N__89542));
    Span4Mux_h I__21647 (
            .O(N__89542),
            .I(N__89538));
    InMux I__21646 (
            .O(N__89541),
            .I(N__89535));
    Odrv4 I__21645 (
            .O(N__89538),
            .I(REG_mem_7_1));
    LocalMux I__21644 (
            .O(N__89535),
            .I(REG_mem_7_1));
    CascadeMux I__21643 (
            .O(N__89530),
            .I(N__89523));
    CascadeMux I__21642 (
            .O(N__89529),
            .I(N__89511));
    CascadeMux I__21641 (
            .O(N__89528),
            .I(N__89508));
    InMux I__21640 (
            .O(N__89527),
            .I(N__89505));
    InMux I__21639 (
            .O(N__89526),
            .I(N__89501));
    InMux I__21638 (
            .O(N__89523),
            .I(N__89494));
    InMux I__21637 (
            .O(N__89522),
            .I(N__89494));
    InMux I__21636 (
            .O(N__89521),
            .I(N__89494));
    CascadeMux I__21635 (
            .O(N__89520),
            .I(N__89484));
    InMux I__21634 (
            .O(N__89519),
            .I(N__89479));
    CascadeMux I__21633 (
            .O(N__89518),
            .I(N__89476));
    CascadeMux I__21632 (
            .O(N__89517),
            .I(N__89469));
    CascadeMux I__21631 (
            .O(N__89516),
            .I(N__89465));
    InMux I__21630 (
            .O(N__89515),
            .I(N__89448));
    CascadeMux I__21629 (
            .O(N__89514),
            .I(N__89445));
    InMux I__21628 (
            .O(N__89511),
            .I(N__89440));
    InMux I__21627 (
            .O(N__89508),
            .I(N__89440));
    LocalMux I__21626 (
            .O(N__89505),
            .I(N__89431));
    InMux I__21625 (
            .O(N__89504),
            .I(N__89428));
    LocalMux I__21624 (
            .O(N__89501),
            .I(N__89423));
    LocalMux I__21623 (
            .O(N__89494),
            .I(N__89423));
    InMux I__21622 (
            .O(N__89493),
            .I(N__89412));
    InMux I__21621 (
            .O(N__89492),
            .I(N__89412));
    InMux I__21620 (
            .O(N__89491),
            .I(N__89412));
    InMux I__21619 (
            .O(N__89490),
            .I(N__89412));
    InMux I__21618 (
            .O(N__89489),
            .I(N__89412));
    InMux I__21617 (
            .O(N__89488),
            .I(N__89401));
    InMux I__21616 (
            .O(N__89487),
            .I(N__89401));
    InMux I__21615 (
            .O(N__89484),
            .I(N__89401));
    InMux I__21614 (
            .O(N__89483),
            .I(N__89401));
    InMux I__21613 (
            .O(N__89482),
            .I(N__89401));
    LocalMux I__21612 (
            .O(N__89479),
            .I(N__89395));
    InMux I__21611 (
            .O(N__89476),
            .I(N__89390));
    InMux I__21610 (
            .O(N__89475),
            .I(N__89390));
    InMux I__21609 (
            .O(N__89474),
            .I(N__89385));
    InMux I__21608 (
            .O(N__89473),
            .I(N__89382));
    InMux I__21607 (
            .O(N__89472),
            .I(N__89379));
    InMux I__21606 (
            .O(N__89469),
            .I(N__89374));
    InMux I__21605 (
            .O(N__89468),
            .I(N__89374));
    InMux I__21604 (
            .O(N__89465),
            .I(N__89367));
    InMux I__21603 (
            .O(N__89464),
            .I(N__89367));
    InMux I__21602 (
            .O(N__89463),
            .I(N__89367));
    InMux I__21601 (
            .O(N__89462),
            .I(N__89362));
    InMux I__21600 (
            .O(N__89461),
            .I(N__89362));
    InMux I__21599 (
            .O(N__89460),
            .I(N__89357));
    InMux I__21598 (
            .O(N__89459),
            .I(N__89357));
    InMux I__21597 (
            .O(N__89458),
            .I(N__89354));
    InMux I__21596 (
            .O(N__89457),
            .I(N__89351));
    InMux I__21595 (
            .O(N__89456),
            .I(N__89346));
    InMux I__21594 (
            .O(N__89455),
            .I(N__89346));
    InMux I__21593 (
            .O(N__89454),
            .I(N__89343));
    InMux I__21592 (
            .O(N__89453),
            .I(N__89336));
    InMux I__21591 (
            .O(N__89452),
            .I(N__89336));
    InMux I__21590 (
            .O(N__89451),
            .I(N__89336));
    LocalMux I__21589 (
            .O(N__89448),
            .I(N__89333));
    InMux I__21588 (
            .O(N__89445),
            .I(N__89330));
    LocalMux I__21587 (
            .O(N__89440),
            .I(N__89327));
    InMux I__21586 (
            .O(N__89439),
            .I(N__89322));
    InMux I__21585 (
            .O(N__89438),
            .I(N__89317));
    InMux I__21584 (
            .O(N__89437),
            .I(N__89317));
    InMux I__21583 (
            .O(N__89436),
            .I(N__89310));
    InMux I__21582 (
            .O(N__89435),
            .I(N__89310));
    InMux I__21581 (
            .O(N__89434),
            .I(N__89310));
    Span4Mux_h I__21580 (
            .O(N__89431),
            .I(N__89307));
    LocalMux I__21579 (
            .O(N__89428),
            .I(N__89304));
    Span4Mux_v I__21578 (
            .O(N__89423),
            .I(N__89296));
    LocalMux I__21577 (
            .O(N__89412),
            .I(N__89293));
    LocalMux I__21576 (
            .O(N__89401),
            .I(N__89290));
    InMux I__21575 (
            .O(N__89400),
            .I(N__89283));
    InMux I__21574 (
            .O(N__89399),
            .I(N__89283));
    InMux I__21573 (
            .O(N__89398),
            .I(N__89283));
    Span4Mux_v I__21572 (
            .O(N__89395),
            .I(N__89278));
    LocalMux I__21571 (
            .O(N__89390),
            .I(N__89278));
    InMux I__21570 (
            .O(N__89389),
            .I(N__89272));
    InMux I__21569 (
            .O(N__89388),
            .I(N__89269));
    LocalMux I__21568 (
            .O(N__89385),
            .I(N__89254));
    LocalMux I__21567 (
            .O(N__89382),
            .I(N__89254));
    LocalMux I__21566 (
            .O(N__89379),
            .I(N__89254));
    LocalMux I__21565 (
            .O(N__89374),
            .I(N__89254));
    LocalMux I__21564 (
            .O(N__89367),
            .I(N__89254));
    LocalMux I__21563 (
            .O(N__89362),
            .I(N__89254));
    LocalMux I__21562 (
            .O(N__89357),
            .I(N__89254));
    LocalMux I__21561 (
            .O(N__89354),
            .I(N__89241));
    LocalMux I__21560 (
            .O(N__89351),
            .I(N__89241));
    LocalMux I__21559 (
            .O(N__89346),
            .I(N__89241));
    LocalMux I__21558 (
            .O(N__89343),
            .I(N__89241));
    LocalMux I__21557 (
            .O(N__89336),
            .I(N__89241));
    Span4Mux_h I__21556 (
            .O(N__89333),
            .I(N__89241));
    LocalMux I__21555 (
            .O(N__89330),
            .I(N__89238));
    Span4Mux_v I__21554 (
            .O(N__89327),
            .I(N__89235));
    InMux I__21553 (
            .O(N__89326),
            .I(N__89230));
    InMux I__21552 (
            .O(N__89325),
            .I(N__89230));
    LocalMux I__21551 (
            .O(N__89322),
            .I(N__89227));
    LocalMux I__21550 (
            .O(N__89317),
            .I(N__89222));
    LocalMux I__21549 (
            .O(N__89310),
            .I(N__89222));
    Span4Mux_h I__21548 (
            .O(N__89307),
            .I(N__89217));
    Span4Mux_h I__21547 (
            .O(N__89304),
            .I(N__89217));
    InMux I__21546 (
            .O(N__89303),
            .I(N__89206));
    InMux I__21545 (
            .O(N__89302),
            .I(N__89206));
    InMux I__21544 (
            .O(N__89301),
            .I(N__89206));
    InMux I__21543 (
            .O(N__89300),
            .I(N__89206));
    InMux I__21542 (
            .O(N__89299),
            .I(N__89206));
    Span4Mux_h I__21541 (
            .O(N__89296),
            .I(N__89199));
    Span4Mux_v I__21540 (
            .O(N__89293),
            .I(N__89199));
    Span4Mux_h I__21539 (
            .O(N__89290),
            .I(N__89199));
    LocalMux I__21538 (
            .O(N__89283),
            .I(N__89194));
    Span4Mux_h I__21537 (
            .O(N__89278),
            .I(N__89194));
    InMux I__21536 (
            .O(N__89277),
            .I(N__89191));
    InMux I__21535 (
            .O(N__89276),
            .I(N__89186));
    InMux I__21534 (
            .O(N__89275),
            .I(N__89186));
    LocalMux I__21533 (
            .O(N__89272),
            .I(N__89179));
    LocalMux I__21532 (
            .O(N__89269),
            .I(N__89179));
    Span4Mux_v I__21531 (
            .O(N__89254),
            .I(N__89179));
    Span4Mux_v I__21530 (
            .O(N__89241),
            .I(N__89176));
    Span4Mux_v I__21529 (
            .O(N__89238),
            .I(N__89171));
    Span4Mux_h I__21528 (
            .O(N__89235),
            .I(N__89171));
    LocalMux I__21527 (
            .O(N__89230),
            .I(N__89162));
    Span4Mux_h I__21526 (
            .O(N__89227),
            .I(N__89162));
    Span4Mux_v I__21525 (
            .O(N__89222),
            .I(N__89162));
    Span4Mux_h I__21524 (
            .O(N__89217),
            .I(N__89162));
    LocalMux I__21523 (
            .O(N__89206),
            .I(N__89155));
    Span4Mux_h I__21522 (
            .O(N__89199),
            .I(N__89155));
    Span4Mux_h I__21521 (
            .O(N__89194),
            .I(N__89155));
    LocalMux I__21520 (
            .O(N__89191),
            .I(N__89150));
    LocalMux I__21519 (
            .O(N__89186),
            .I(N__89150));
    Span4Mux_v I__21518 (
            .O(N__89179),
            .I(N__89143));
    Span4Mux_v I__21517 (
            .O(N__89176),
            .I(N__89143));
    Span4Mux_v I__21516 (
            .O(N__89171),
            .I(N__89143));
    Span4Mux_v I__21515 (
            .O(N__89162),
            .I(N__89140));
    Span4Mux_v I__21514 (
            .O(N__89155),
            .I(N__89137));
    Odrv12 I__21513 (
            .O(N__89150),
            .I(dc32_fifo_data_in_8));
    Odrv4 I__21512 (
            .O(N__89143),
            .I(dc32_fifo_data_in_8));
    Odrv4 I__21511 (
            .O(N__89140),
            .I(dc32_fifo_data_in_8));
    Odrv4 I__21510 (
            .O(N__89137),
            .I(dc32_fifo_data_in_8));
    InMux I__21509 (
            .O(N__89128),
            .I(N__89125));
    LocalMux I__21508 (
            .O(N__89125),
            .I(N__89119));
    InMux I__21507 (
            .O(N__89124),
            .I(N__89116));
    InMux I__21506 (
            .O(N__89123),
            .I(N__89111));
    InMux I__21505 (
            .O(N__89122),
            .I(N__89108));
    Span4Mux_h I__21504 (
            .O(N__89119),
            .I(N__89105));
    LocalMux I__21503 (
            .O(N__89116),
            .I(N__89099));
    InMux I__21502 (
            .O(N__89115),
            .I(N__89096));
    InMux I__21501 (
            .O(N__89114),
            .I(N__89093));
    LocalMux I__21500 (
            .O(N__89111),
            .I(N__89090));
    LocalMux I__21499 (
            .O(N__89108),
            .I(N__89087));
    Span4Mux_h I__21498 (
            .O(N__89105),
            .I(N__89084));
    InMux I__21497 (
            .O(N__89104),
            .I(N__89081));
    InMux I__21496 (
            .O(N__89103),
            .I(N__89078));
    InMux I__21495 (
            .O(N__89102),
            .I(N__89075));
    Span4Mux_v I__21494 (
            .O(N__89099),
            .I(N__89069));
    LocalMux I__21493 (
            .O(N__89096),
            .I(N__89066));
    LocalMux I__21492 (
            .O(N__89093),
            .I(N__89063));
    Span4Mux_h I__21491 (
            .O(N__89090),
            .I(N__89058));
    Span4Mux_h I__21490 (
            .O(N__89087),
            .I(N__89058));
    Span4Mux_h I__21489 (
            .O(N__89084),
            .I(N__89049));
    LocalMux I__21488 (
            .O(N__89081),
            .I(N__89049));
    LocalMux I__21487 (
            .O(N__89078),
            .I(N__89049));
    LocalMux I__21486 (
            .O(N__89075),
            .I(N__89049));
    InMux I__21485 (
            .O(N__89074),
            .I(N__89046));
    InMux I__21484 (
            .O(N__89073),
            .I(N__89043));
    InMux I__21483 (
            .O(N__89072),
            .I(N__89040));
    Span4Mux_h I__21482 (
            .O(N__89069),
            .I(N__89035));
    Span4Mux_v I__21481 (
            .O(N__89066),
            .I(N__89032));
    Span4Mux_h I__21480 (
            .O(N__89063),
            .I(N__89029));
    Span4Mux_v I__21479 (
            .O(N__89058),
            .I(N__89024));
    Span4Mux_h I__21478 (
            .O(N__89049),
            .I(N__89024));
    LocalMux I__21477 (
            .O(N__89046),
            .I(N__89017));
    LocalMux I__21476 (
            .O(N__89043),
            .I(N__89017));
    LocalMux I__21475 (
            .O(N__89040),
            .I(N__89017));
    InMux I__21474 (
            .O(N__89039),
            .I(N__89012));
    InMux I__21473 (
            .O(N__89038),
            .I(N__89012));
    Span4Mux_h I__21472 (
            .O(N__89035),
            .I(N__89005));
    Span4Mux_h I__21471 (
            .O(N__89032),
            .I(N__89005));
    Span4Mux_h I__21470 (
            .O(N__89029),
            .I(N__89002));
    Span4Mux_v I__21469 (
            .O(N__89024),
            .I(N__88995));
    Span4Mux_v I__21468 (
            .O(N__89017),
            .I(N__88995));
    LocalMux I__21467 (
            .O(N__89012),
            .I(N__88995));
    InMux I__21466 (
            .O(N__89011),
            .I(N__88990));
    InMux I__21465 (
            .O(N__89010),
            .I(N__88990));
    Odrv4 I__21464 (
            .O(N__89005),
            .I(n19));
    Odrv4 I__21463 (
            .O(N__89002),
            .I(n19));
    Odrv4 I__21462 (
            .O(N__88995),
            .I(n19));
    LocalMux I__21461 (
            .O(N__88990),
            .I(n19));
    CascadeMux I__21460 (
            .O(N__88981),
            .I(N__88978));
    InMux I__21459 (
            .O(N__88978),
            .I(N__88972));
    InMux I__21458 (
            .O(N__88977),
            .I(N__88972));
    LocalMux I__21457 (
            .O(N__88972),
            .I(REG_mem_46_8));
    CascadeMux I__21456 (
            .O(N__88969),
            .I(N__88966));
    InMux I__21455 (
            .O(N__88966),
            .I(N__88963));
    LocalMux I__21454 (
            .O(N__88963),
            .I(N__88960));
    Span4Mux_v I__21453 (
            .O(N__88960),
            .I(N__88957));
    Span4Mux_h I__21452 (
            .O(N__88957),
            .I(N__88954));
    Span4Mux_h I__21451 (
            .O(N__88954),
            .I(N__88951));
    Odrv4 I__21450 (
            .O(N__88951),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11683 ));
    CascadeMux I__21449 (
            .O(N__88948),
            .I(N__88944));
    InMux I__21448 (
            .O(N__88947),
            .I(N__88939));
    InMux I__21447 (
            .O(N__88944),
            .I(N__88939));
    LocalMux I__21446 (
            .O(N__88939),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_1 ));
    CascadeMux I__21445 (
            .O(N__88936),
            .I(N__88932));
    InMux I__21444 (
            .O(N__88935),
            .I(N__88927));
    InMux I__21443 (
            .O(N__88932),
            .I(N__88927));
    LocalMux I__21442 (
            .O(N__88927),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_1 ));
    CascadeMux I__21441 (
            .O(N__88924),
            .I(N__88920));
    InMux I__21440 (
            .O(N__88923),
            .I(N__88915));
    InMux I__21439 (
            .O(N__88920),
            .I(N__88915));
    LocalMux I__21438 (
            .O(N__88915),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_1 ));
    CascadeMux I__21437 (
            .O(N__88912),
            .I(N__88908));
    CascadeMux I__21436 (
            .O(N__88911),
            .I(N__88902));
    InMux I__21435 (
            .O(N__88908),
            .I(N__88891));
    InMux I__21434 (
            .O(N__88907),
            .I(N__88891));
    InMux I__21433 (
            .O(N__88906),
            .I(N__88891));
    CascadeMux I__21432 (
            .O(N__88905),
            .I(N__88888));
    InMux I__21431 (
            .O(N__88902),
            .I(N__88872));
    InMux I__21430 (
            .O(N__88901),
            .I(N__88872));
    InMux I__21429 (
            .O(N__88900),
            .I(N__88869));
    InMux I__21428 (
            .O(N__88899),
            .I(N__88864));
    InMux I__21427 (
            .O(N__88898),
            .I(N__88864));
    LocalMux I__21426 (
            .O(N__88891),
            .I(N__88861));
    InMux I__21425 (
            .O(N__88888),
            .I(N__88858));
    CascadeMux I__21424 (
            .O(N__88887),
            .I(N__88846));
    CascadeMux I__21423 (
            .O(N__88886),
            .I(N__88838));
    InMux I__21422 (
            .O(N__88885),
            .I(N__88829));
    InMux I__21421 (
            .O(N__88884),
            .I(N__88829));
    InMux I__21420 (
            .O(N__88883),
            .I(N__88822));
    InMux I__21419 (
            .O(N__88882),
            .I(N__88822));
    InMux I__21418 (
            .O(N__88881),
            .I(N__88822));
    CascadeMux I__21417 (
            .O(N__88880),
            .I(N__88815));
    CascadeMux I__21416 (
            .O(N__88879),
            .I(N__88805));
    InMux I__21415 (
            .O(N__88878),
            .I(N__88799));
    InMux I__21414 (
            .O(N__88877),
            .I(N__88796));
    LocalMux I__21413 (
            .O(N__88872),
            .I(N__88793));
    LocalMux I__21412 (
            .O(N__88869),
            .I(N__88788));
    LocalMux I__21411 (
            .O(N__88864),
            .I(N__88788));
    Span4Mux_v I__21410 (
            .O(N__88861),
            .I(N__88783));
    LocalMux I__21409 (
            .O(N__88858),
            .I(N__88783));
    InMux I__21408 (
            .O(N__88857),
            .I(N__88780));
    InMux I__21407 (
            .O(N__88856),
            .I(N__88761));
    InMux I__21406 (
            .O(N__88855),
            .I(N__88761));
    InMux I__21405 (
            .O(N__88854),
            .I(N__88761));
    InMux I__21404 (
            .O(N__88853),
            .I(N__88761));
    CascadeMux I__21403 (
            .O(N__88852),
            .I(N__88750));
    InMux I__21402 (
            .O(N__88851),
            .I(N__88745));
    CascadeMux I__21401 (
            .O(N__88850),
            .I(N__88739));
    InMux I__21400 (
            .O(N__88849),
            .I(N__88734));
    InMux I__21399 (
            .O(N__88846),
            .I(N__88729));
    InMux I__21398 (
            .O(N__88845),
            .I(N__88729));
    InMux I__21397 (
            .O(N__88844),
            .I(N__88721));
    InMux I__21396 (
            .O(N__88843),
            .I(N__88721));
    InMux I__21395 (
            .O(N__88842),
            .I(N__88716));
    InMux I__21394 (
            .O(N__88841),
            .I(N__88716));
    InMux I__21393 (
            .O(N__88838),
            .I(N__88711));
    InMux I__21392 (
            .O(N__88837),
            .I(N__88711));
    InMux I__21391 (
            .O(N__88836),
            .I(N__88708));
    InMux I__21390 (
            .O(N__88835),
            .I(N__88705));
    CascadeMux I__21389 (
            .O(N__88834),
            .I(N__88702));
    LocalMux I__21388 (
            .O(N__88829),
            .I(N__88693));
    LocalMux I__21387 (
            .O(N__88822),
            .I(N__88693));
    InMux I__21386 (
            .O(N__88821),
            .I(N__88688));
    InMux I__21385 (
            .O(N__88820),
            .I(N__88688));
    InMux I__21384 (
            .O(N__88819),
            .I(N__88681));
    InMux I__21383 (
            .O(N__88818),
            .I(N__88681));
    InMux I__21382 (
            .O(N__88815),
            .I(N__88681));
    InMux I__21381 (
            .O(N__88814),
            .I(N__88676));
    InMux I__21380 (
            .O(N__88813),
            .I(N__88676));
    CascadeMux I__21379 (
            .O(N__88812),
            .I(N__88671));
    InMux I__21378 (
            .O(N__88811),
            .I(N__88666));
    InMux I__21377 (
            .O(N__88810),
            .I(N__88661));
    InMux I__21376 (
            .O(N__88809),
            .I(N__88661));
    InMux I__21375 (
            .O(N__88808),
            .I(N__88656));
    InMux I__21374 (
            .O(N__88805),
            .I(N__88656));
    InMux I__21373 (
            .O(N__88804),
            .I(N__88653));
    CascadeMux I__21372 (
            .O(N__88803),
            .I(N__88650));
    CascadeMux I__21371 (
            .O(N__88802),
            .I(N__88647));
    LocalMux I__21370 (
            .O(N__88799),
            .I(N__88644));
    LocalMux I__21369 (
            .O(N__88796),
            .I(N__88641));
    Span4Mux_h I__21368 (
            .O(N__88793),
            .I(N__88632));
    Span4Mux_v I__21367 (
            .O(N__88788),
            .I(N__88632));
    Span4Mux_v I__21366 (
            .O(N__88783),
            .I(N__88632));
    LocalMux I__21365 (
            .O(N__88780),
            .I(N__88632));
    InMux I__21364 (
            .O(N__88779),
            .I(N__88625));
    InMux I__21363 (
            .O(N__88778),
            .I(N__88625));
    InMux I__21362 (
            .O(N__88777),
            .I(N__88625));
    InMux I__21361 (
            .O(N__88776),
            .I(N__88620));
    InMux I__21360 (
            .O(N__88775),
            .I(N__88620));
    CascadeMux I__21359 (
            .O(N__88774),
            .I(N__88614));
    CascadeMux I__21358 (
            .O(N__88773),
            .I(N__88599));
    CascadeMux I__21357 (
            .O(N__88772),
            .I(N__88592));
    InMux I__21356 (
            .O(N__88771),
            .I(N__88576));
    InMux I__21355 (
            .O(N__88770),
            .I(N__88576));
    LocalMux I__21354 (
            .O(N__88761),
            .I(N__88572));
    InMux I__21353 (
            .O(N__88760),
            .I(N__88569));
    InMux I__21352 (
            .O(N__88759),
            .I(N__88560));
    InMux I__21351 (
            .O(N__88758),
            .I(N__88560));
    InMux I__21350 (
            .O(N__88757),
            .I(N__88560));
    InMux I__21349 (
            .O(N__88756),
            .I(N__88560));
    InMux I__21348 (
            .O(N__88755),
            .I(N__88555));
    InMux I__21347 (
            .O(N__88754),
            .I(N__88555));
    InMux I__21346 (
            .O(N__88753),
            .I(N__88550));
    InMux I__21345 (
            .O(N__88750),
            .I(N__88550));
    CascadeMux I__21344 (
            .O(N__88749),
            .I(N__88547));
    CascadeMux I__21343 (
            .O(N__88748),
            .I(N__88542));
    LocalMux I__21342 (
            .O(N__88745),
            .I(N__88531));
    InMux I__21341 (
            .O(N__88744),
            .I(N__88526));
    InMux I__21340 (
            .O(N__88743),
            .I(N__88526));
    InMux I__21339 (
            .O(N__88742),
            .I(N__88523));
    InMux I__21338 (
            .O(N__88739),
            .I(N__88518));
    InMux I__21337 (
            .O(N__88738),
            .I(N__88518));
    CascadeMux I__21336 (
            .O(N__88737),
            .I(N__88515));
    LocalMux I__21335 (
            .O(N__88734),
            .I(N__88504));
    LocalMux I__21334 (
            .O(N__88729),
            .I(N__88504));
    InMux I__21333 (
            .O(N__88728),
            .I(N__88497));
    InMux I__21332 (
            .O(N__88727),
            .I(N__88497));
    InMux I__21331 (
            .O(N__88726),
            .I(N__88497));
    LocalMux I__21330 (
            .O(N__88721),
            .I(N__88486));
    LocalMux I__21329 (
            .O(N__88716),
            .I(N__88486));
    LocalMux I__21328 (
            .O(N__88711),
            .I(N__88486));
    LocalMux I__21327 (
            .O(N__88708),
            .I(N__88486));
    LocalMux I__21326 (
            .O(N__88705),
            .I(N__88486));
    InMux I__21325 (
            .O(N__88702),
            .I(N__88483));
    InMux I__21324 (
            .O(N__88701),
            .I(N__88476));
    InMux I__21323 (
            .O(N__88700),
            .I(N__88476));
    InMux I__21322 (
            .O(N__88699),
            .I(N__88476));
    InMux I__21321 (
            .O(N__88698),
            .I(N__88470));
    Span4Mux_v I__21320 (
            .O(N__88693),
            .I(N__88465));
    LocalMux I__21319 (
            .O(N__88688),
            .I(N__88465));
    LocalMux I__21318 (
            .O(N__88681),
            .I(N__88460));
    LocalMux I__21317 (
            .O(N__88676),
            .I(N__88460));
    InMux I__21316 (
            .O(N__88675),
            .I(N__88455));
    InMux I__21315 (
            .O(N__88674),
            .I(N__88455));
    InMux I__21314 (
            .O(N__88671),
            .I(N__88452));
    InMux I__21313 (
            .O(N__88670),
            .I(N__88449));
    CascadeMux I__21312 (
            .O(N__88669),
            .I(N__88439));
    LocalMux I__21311 (
            .O(N__88666),
            .I(N__88436));
    LocalMux I__21310 (
            .O(N__88661),
            .I(N__88433));
    LocalMux I__21309 (
            .O(N__88656),
            .I(N__88428));
    LocalMux I__21308 (
            .O(N__88653),
            .I(N__88428));
    InMux I__21307 (
            .O(N__88650),
            .I(N__88423));
    InMux I__21306 (
            .O(N__88647),
            .I(N__88423));
    Span4Mux_h I__21305 (
            .O(N__88644),
            .I(N__88412));
    Span4Mux_v I__21304 (
            .O(N__88641),
            .I(N__88412));
    Span4Mux_h I__21303 (
            .O(N__88632),
            .I(N__88412));
    LocalMux I__21302 (
            .O(N__88625),
            .I(N__88412));
    LocalMux I__21301 (
            .O(N__88620),
            .I(N__88412));
    InMux I__21300 (
            .O(N__88619),
            .I(N__88409));
    CascadeMux I__21299 (
            .O(N__88618),
            .I(N__88405));
    InMux I__21298 (
            .O(N__88617),
            .I(N__88402));
    InMux I__21297 (
            .O(N__88614),
            .I(N__88395));
    InMux I__21296 (
            .O(N__88613),
            .I(N__88395));
    InMux I__21295 (
            .O(N__88612),
            .I(N__88395));
    InMux I__21294 (
            .O(N__88611),
            .I(N__88392));
    InMux I__21293 (
            .O(N__88610),
            .I(N__88385));
    InMux I__21292 (
            .O(N__88609),
            .I(N__88385));
    InMux I__21291 (
            .O(N__88608),
            .I(N__88385));
    InMux I__21290 (
            .O(N__88607),
            .I(N__88378));
    InMux I__21289 (
            .O(N__88606),
            .I(N__88378));
    InMux I__21288 (
            .O(N__88605),
            .I(N__88378));
    InMux I__21287 (
            .O(N__88604),
            .I(N__88375));
    InMux I__21286 (
            .O(N__88603),
            .I(N__88366));
    InMux I__21285 (
            .O(N__88602),
            .I(N__88366));
    InMux I__21284 (
            .O(N__88599),
            .I(N__88363));
    InMux I__21283 (
            .O(N__88598),
            .I(N__88360));
    InMux I__21282 (
            .O(N__88597),
            .I(N__88355));
    InMux I__21281 (
            .O(N__88596),
            .I(N__88355));
    InMux I__21280 (
            .O(N__88595),
            .I(N__88351));
    InMux I__21279 (
            .O(N__88592),
            .I(N__88348));
    InMux I__21278 (
            .O(N__88591),
            .I(N__88343));
    InMux I__21277 (
            .O(N__88590),
            .I(N__88343));
    InMux I__21276 (
            .O(N__88589),
            .I(N__88338));
    CascadeMux I__21275 (
            .O(N__88588),
            .I(N__88327));
    InMux I__21274 (
            .O(N__88587),
            .I(N__88322));
    InMux I__21273 (
            .O(N__88586),
            .I(N__88311));
    InMux I__21272 (
            .O(N__88585),
            .I(N__88311));
    InMux I__21271 (
            .O(N__88584),
            .I(N__88311));
    InMux I__21270 (
            .O(N__88583),
            .I(N__88304));
    InMux I__21269 (
            .O(N__88582),
            .I(N__88304));
    InMux I__21268 (
            .O(N__88581),
            .I(N__88304));
    LocalMux I__21267 (
            .O(N__88576),
            .I(N__88297));
    InMux I__21266 (
            .O(N__88575),
            .I(N__88294));
    Span4Mux_v I__21265 (
            .O(N__88572),
            .I(N__88287));
    LocalMux I__21264 (
            .O(N__88569),
            .I(N__88287));
    LocalMux I__21263 (
            .O(N__88560),
            .I(N__88287));
    LocalMux I__21262 (
            .O(N__88555),
            .I(N__88282));
    LocalMux I__21261 (
            .O(N__88550),
            .I(N__88282));
    InMux I__21260 (
            .O(N__88547),
            .I(N__88279));
    InMux I__21259 (
            .O(N__88546),
            .I(N__88276));
    InMux I__21258 (
            .O(N__88545),
            .I(N__88273));
    InMux I__21257 (
            .O(N__88542),
            .I(N__88268));
    InMux I__21256 (
            .O(N__88541),
            .I(N__88268));
    InMux I__21255 (
            .O(N__88540),
            .I(N__88265));
    CascadeMux I__21254 (
            .O(N__88539),
            .I(N__88258));
    CascadeMux I__21253 (
            .O(N__88538),
            .I(N__88255));
    InMux I__21252 (
            .O(N__88537),
            .I(N__88248));
    InMux I__21251 (
            .O(N__88536),
            .I(N__88248));
    CascadeMux I__21250 (
            .O(N__88535),
            .I(N__88235));
    CascadeMux I__21249 (
            .O(N__88534),
            .I(N__88229));
    Span4Mux_v I__21248 (
            .O(N__88531),
            .I(N__88219));
    LocalMux I__21247 (
            .O(N__88526),
            .I(N__88219));
    LocalMux I__21246 (
            .O(N__88523),
            .I(N__88219));
    LocalMux I__21245 (
            .O(N__88518),
            .I(N__88219));
    InMux I__21244 (
            .O(N__88515),
            .I(N__88216));
    InMux I__21243 (
            .O(N__88514),
            .I(N__88213));
    InMux I__21242 (
            .O(N__88513),
            .I(N__88208));
    InMux I__21241 (
            .O(N__88512),
            .I(N__88208));
    InMux I__21240 (
            .O(N__88511),
            .I(N__88205));
    InMux I__21239 (
            .O(N__88510),
            .I(N__88200));
    InMux I__21238 (
            .O(N__88509),
            .I(N__88200));
    Span4Mux_v I__21237 (
            .O(N__88504),
            .I(N__88195));
    LocalMux I__21236 (
            .O(N__88497),
            .I(N__88195));
    Span4Mux_v I__21235 (
            .O(N__88486),
            .I(N__88188));
    LocalMux I__21234 (
            .O(N__88483),
            .I(N__88188));
    LocalMux I__21233 (
            .O(N__88476),
            .I(N__88188));
    InMux I__21232 (
            .O(N__88475),
            .I(N__88185));
    InMux I__21231 (
            .O(N__88474),
            .I(N__88180));
    InMux I__21230 (
            .O(N__88473),
            .I(N__88180));
    LocalMux I__21229 (
            .O(N__88470),
            .I(N__88177));
    Span4Mux_h I__21228 (
            .O(N__88465),
            .I(N__88166));
    Span4Mux_v I__21227 (
            .O(N__88460),
            .I(N__88166));
    LocalMux I__21226 (
            .O(N__88455),
            .I(N__88166));
    LocalMux I__21225 (
            .O(N__88452),
            .I(N__88166));
    LocalMux I__21224 (
            .O(N__88449),
            .I(N__88166));
    InMux I__21223 (
            .O(N__88448),
            .I(N__88163));
    InMux I__21222 (
            .O(N__88447),
            .I(N__88160));
    InMux I__21221 (
            .O(N__88446),
            .I(N__88157));
    InMux I__21220 (
            .O(N__88445),
            .I(N__88152));
    InMux I__21219 (
            .O(N__88444),
            .I(N__88152));
    InMux I__21218 (
            .O(N__88443),
            .I(N__88149));
    InMux I__21217 (
            .O(N__88442),
            .I(N__88143));
    InMux I__21216 (
            .O(N__88439),
            .I(N__88143));
    Span4Mux_h I__21215 (
            .O(N__88436),
            .I(N__88134));
    Span4Mux_h I__21214 (
            .O(N__88433),
            .I(N__88134));
    Span4Mux_v I__21213 (
            .O(N__88428),
            .I(N__88134));
    LocalMux I__21212 (
            .O(N__88423),
            .I(N__88134));
    Span4Mux_h I__21211 (
            .O(N__88412),
            .I(N__88129));
    LocalMux I__21210 (
            .O(N__88409),
            .I(N__88129));
    CascadeMux I__21209 (
            .O(N__88408),
            .I(N__88126));
    InMux I__21208 (
            .O(N__88405),
            .I(N__88122));
    LocalMux I__21207 (
            .O(N__88402),
            .I(N__88109));
    LocalMux I__21206 (
            .O(N__88395),
            .I(N__88109));
    LocalMux I__21205 (
            .O(N__88392),
            .I(N__88109));
    LocalMux I__21204 (
            .O(N__88385),
            .I(N__88109));
    LocalMux I__21203 (
            .O(N__88378),
            .I(N__88109));
    LocalMux I__21202 (
            .O(N__88375),
            .I(N__88109));
    InMux I__21201 (
            .O(N__88374),
            .I(N__88104));
    InMux I__21200 (
            .O(N__88373),
            .I(N__88104));
    CascadeMux I__21199 (
            .O(N__88372),
            .I(N__88101));
    CascadeMux I__21198 (
            .O(N__88371),
            .I(N__88098));
    LocalMux I__21197 (
            .O(N__88366),
            .I(N__88086));
    LocalMux I__21196 (
            .O(N__88363),
            .I(N__88086));
    LocalMux I__21195 (
            .O(N__88360),
            .I(N__88086));
    LocalMux I__21194 (
            .O(N__88355),
            .I(N__88086));
    InMux I__21193 (
            .O(N__88354),
            .I(N__88083));
    LocalMux I__21192 (
            .O(N__88351),
            .I(N__88076));
    LocalMux I__21191 (
            .O(N__88348),
            .I(N__88076));
    LocalMux I__21190 (
            .O(N__88343),
            .I(N__88076));
    InMux I__21189 (
            .O(N__88342),
            .I(N__88071));
    InMux I__21188 (
            .O(N__88341),
            .I(N__88071));
    LocalMux I__21187 (
            .O(N__88338),
            .I(N__88066));
    InMux I__21186 (
            .O(N__88337),
            .I(N__88063));
    InMux I__21185 (
            .O(N__88336),
            .I(N__88060));
    InMux I__21184 (
            .O(N__88335),
            .I(N__88055));
    InMux I__21183 (
            .O(N__88334),
            .I(N__88055));
    CascadeMux I__21182 (
            .O(N__88333),
            .I(N__88047));
    CascadeMux I__21181 (
            .O(N__88332),
            .I(N__88037));
    InMux I__21180 (
            .O(N__88331),
            .I(N__88033));
    InMux I__21179 (
            .O(N__88330),
            .I(N__88024));
    InMux I__21178 (
            .O(N__88327),
            .I(N__88024));
    InMux I__21177 (
            .O(N__88326),
            .I(N__88019));
    InMux I__21176 (
            .O(N__88325),
            .I(N__88019));
    LocalMux I__21175 (
            .O(N__88322),
            .I(N__88016));
    InMux I__21174 (
            .O(N__88321),
            .I(N__88009));
    InMux I__21173 (
            .O(N__88320),
            .I(N__88009));
    InMux I__21172 (
            .O(N__88319),
            .I(N__88009));
    InMux I__21171 (
            .O(N__88318),
            .I(N__87993));
    LocalMux I__21170 (
            .O(N__88311),
            .I(N__87988));
    LocalMux I__21169 (
            .O(N__88304),
            .I(N__87988));
    InMux I__21168 (
            .O(N__88303),
            .I(N__87985));
    InMux I__21167 (
            .O(N__88302),
            .I(N__87978));
    InMux I__21166 (
            .O(N__88301),
            .I(N__87978));
    InMux I__21165 (
            .O(N__88300),
            .I(N__87978));
    Span4Mux_v I__21164 (
            .O(N__88297),
            .I(N__87974));
    LocalMux I__21163 (
            .O(N__88294),
            .I(N__87971));
    Span4Mux_v I__21162 (
            .O(N__88287),
            .I(N__87968));
    Span4Mux_v I__21161 (
            .O(N__88282),
            .I(N__87961));
    LocalMux I__21160 (
            .O(N__88279),
            .I(N__87961));
    LocalMux I__21159 (
            .O(N__88276),
            .I(N__87961));
    LocalMux I__21158 (
            .O(N__88273),
            .I(N__87954));
    LocalMux I__21157 (
            .O(N__88268),
            .I(N__87954));
    LocalMux I__21156 (
            .O(N__88265),
            .I(N__87954));
    InMux I__21155 (
            .O(N__88264),
            .I(N__87951));
    InMux I__21154 (
            .O(N__88263),
            .I(N__87944));
    InMux I__21153 (
            .O(N__88262),
            .I(N__87944));
    InMux I__21152 (
            .O(N__88261),
            .I(N__87944));
    InMux I__21151 (
            .O(N__88258),
            .I(N__87941));
    InMux I__21150 (
            .O(N__88255),
            .I(N__87936));
    InMux I__21149 (
            .O(N__88254),
            .I(N__87936));
    InMux I__21148 (
            .O(N__88253),
            .I(N__87933));
    LocalMux I__21147 (
            .O(N__88248),
            .I(N__87930));
    InMux I__21146 (
            .O(N__88247),
            .I(N__87925));
    InMux I__21145 (
            .O(N__88246),
            .I(N__87925));
    InMux I__21144 (
            .O(N__88245),
            .I(N__87920));
    InMux I__21143 (
            .O(N__88244),
            .I(N__87920));
    InMux I__21142 (
            .O(N__88243),
            .I(N__87915));
    InMux I__21141 (
            .O(N__88242),
            .I(N__87915));
    InMux I__21140 (
            .O(N__88241),
            .I(N__87911));
    InMux I__21139 (
            .O(N__88240),
            .I(N__87904));
    InMux I__21138 (
            .O(N__88239),
            .I(N__87904));
    InMux I__21137 (
            .O(N__88238),
            .I(N__87904));
    InMux I__21136 (
            .O(N__88235),
            .I(N__87897));
    InMux I__21135 (
            .O(N__88234),
            .I(N__87897));
    InMux I__21134 (
            .O(N__88233),
            .I(N__87892));
    InMux I__21133 (
            .O(N__88232),
            .I(N__87892));
    InMux I__21132 (
            .O(N__88229),
            .I(N__87887));
    InMux I__21131 (
            .O(N__88228),
            .I(N__87887));
    Span4Mux_v I__21130 (
            .O(N__88219),
            .I(N__87883));
    LocalMux I__21129 (
            .O(N__88216),
            .I(N__87880));
    LocalMux I__21128 (
            .O(N__88213),
            .I(N__87871));
    LocalMux I__21127 (
            .O(N__88208),
            .I(N__87871));
    LocalMux I__21126 (
            .O(N__88205),
            .I(N__87871));
    LocalMux I__21125 (
            .O(N__88200),
            .I(N__87871));
    Span4Mux_v I__21124 (
            .O(N__88195),
            .I(N__87862));
    Span4Mux_h I__21123 (
            .O(N__88188),
            .I(N__87862));
    LocalMux I__21122 (
            .O(N__88185),
            .I(N__87862));
    LocalMux I__21121 (
            .O(N__88180),
            .I(N__87862));
    Span4Mux_v I__21120 (
            .O(N__88177),
            .I(N__87847));
    Span4Mux_h I__21119 (
            .O(N__88166),
            .I(N__87847));
    LocalMux I__21118 (
            .O(N__88163),
            .I(N__87847));
    LocalMux I__21117 (
            .O(N__88160),
            .I(N__87847));
    LocalMux I__21116 (
            .O(N__88157),
            .I(N__87847));
    LocalMux I__21115 (
            .O(N__88152),
            .I(N__87847));
    LocalMux I__21114 (
            .O(N__88149),
            .I(N__87847));
    InMux I__21113 (
            .O(N__88148),
            .I(N__87844));
    LocalMux I__21112 (
            .O(N__88143),
            .I(N__87841));
    Span4Mux_h I__21111 (
            .O(N__88134),
            .I(N__87836));
    Span4Mux_h I__21110 (
            .O(N__88129),
            .I(N__87836));
    InMux I__21109 (
            .O(N__88126),
            .I(N__87833));
    InMux I__21108 (
            .O(N__88125),
            .I(N__87830));
    LocalMux I__21107 (
            .O(N__88122),
            .I(N__87823));
    Span4Mux_v I__21106 (
            .O(N__88109),
            .I(N__87823));
    LocalMux I__21105 (
            .O(N__88104),
            .I(N__87823));
    InMux I__21104 (
            .O(N__88101),
            .I(N__87820));
    InMux I__21103 (
            .O(N__88098),
            .I(N__87815));
    InMux I__21102 (
            .O(N__88097),
            .I(N__87815));
    InMux I__21101 (
            .O(N__88096),
            .I(N__87810));
    InMux I__21100 (
            .O(N__88095),
            .I(N__87810));
    Span4Mux_v I__21099 (
            .O(N__88086),
            .I(N__87805));
    LocalMux I__21098 (
            .O(N__88083),
            .I(N__87805));
    Span4Mux_v I__21097 (
            .O(N__88076),
            .I(N__87800));
    LocalMux I__21096 (
            .O(N__88071),
            .I(N__87800));
    InMux I__21095 (
            .O(N__88070),
            .I(N__87797));
    CascadeMux I__21094 (
            .O(N__88069),
            .I(N__87794));
    Span4Mux_v I__21093 (
            .O(N__88066),
            .I(N__87784));
    LocalMux I__21092 (
            .O(N__88063),
            .I(N__87784));
    LocalMux I__21091 (
            .O(N__88060),
            .I(N__87784));
    LocalMux I__21090 (
            .O(N__88055),
            .I(N__87781));
    InMux I__21089 (
            .O(N__88054),
            .I(N__87776));
    InMux I__21088 (
            .O(N__88053),
            .I(N__87776));
    InMux I__21087 (
            .O(N__88052),
            .I(N__87771));
    InMux I__21086 (
            .O(N__88051),
            .I(N__87771));
    InMux I__21085 (
            .O(N__88050),
            .I(N__87768));
    InMux I__21084 (
            .O(N__88047),
            .I(N__87763));
    InMux I__21083 (
            .O(N__88046),
            .I(N__87763));
    InMux I__21082 (
            .O(N__88045),
            .I(N__87760));
    InMux I__21081 (
            .O(N__88044),
            .I(N__87757));
    InMux I__21080 (
            .O(N__88043),
            .I(N__87742));
    InMux I__21079 (
            .O(N__88042),
            .I(N__87742));
    InMux I__21078 (
            .O(N__88041),
            .I(N__87742));
    InMux I__21077 (
            .O(N__88040),
            .I(N__87742));
    InMux I__21076 (
            .O(N__88037),
            .I(N__87737));
    InMux I__21075 (
            .O(N__88036),
            .I(N__87737));
    LocalMux I__21074 (
            .O(N__88033),
            .I(N__87730));
    InMux I__21073 (
            .O(N__88032),
            .I(N__87727));
    InMux I__21072 (
            .O(N__88031),
            .I(N__87723));
    InMux I__21071 (
            .O(N__88030),
            .I(N__87718));
    InMux I__21070 (
            .O(N__88029),
            .I(N__87718));
    LocalMux I__21069 (
            .O(N__88024),
            .I(N__87709));
    LocalMux I__21068 (
            .O(N__88019),
            .I(N__87702));
    Span4Mux_v I__21067 (
            .O(N__88016),
            .I(N__87702));
    LocalMux I__21066 (
            .O(N__88009),
            .I(N__87702));
    InMux I__21065 (
            .O(N__88008),
            .I(N__87699));
    InMux I__21064 (
            .O(N__88007),
            .I(N__87694));
    InMux I__21063 (
            .O(N__88006),
            .I(N__87694));
    InMux I__21062 (
            .O(N__88005),
            .I(N__87689));
    InMux I__21061 (
            .O(N__88004),
            .I(N__87689));
    InMux I__21060 (
            .O(N__88003),
            .I(N__87684));
    InMux I__21059 (
            .O(N__88002),
            .I(N__87684));
    InMux I__21058 (
            .O(N__88001),
            .I(N__87679));
    InMux I__21057 (
            .O(N__88000),
            .I(N__87679));
    InMux I__21056 (
            .O(N__87999),
            .I(N__87667));
    InMux I__21055 (
            .O(N__87998),
            .I(N__87667));
    InMux I__21054 (
            .O(N__87997),
            .I(N__87667));
    InMux I__21053 (
            .O(N__87996),
            .I(N__87667));
    LocalMux I__21052 (
            .O(N__87993),
            .I(N__87658));
    Span4Mux_v I__21051 (
            .O(N__87988),
            .I(N__87651));
    LocalMux I__21050 (
            .O(N__87985),
            .I(N__87651));
    LocalMux I__21049 (
            .O(N__87978),
            .I(N__87651));
    InMux I__21048 (
            .O(N__87977),
            .I(N__87643));
    Span4Mux_h I__21047 (
            .O(N__87974),
            .I(N__87634));
    Span4Mux_v I__21046 (
            .O(N__87971),
            .I(N__87634));
    Span4Mux_v I__21045 (
            .O(N__87968),
            .I(N__87634));
    Span4Mux_v I__21044 (
            .O(N__87961),
            .I(N__87634));
    Span4Mux_v I__21043 (
            .O(N__87954),
            .I(N__87627));
    LocalMux I__21042 (
            .O(N__87951),
            .I(N__87627));
    LocalMux I__21041 (
            .O(N__87944),
            .I(N__87627));
    LocalMux I__21040 (
            .O(N__87941),
            .I(N__87620));
    LocalMux I__21039 (
            .O(N__87936),
            .I(N__87620));
    LocalMux I__21038 (
            .O(N__87933),
            .I(N__87620));
    Span4Mux_v I__21037 (
            .O(N__87930),
            .I(N__87615));
    LocalMux I__21036 (
            .O(N__87925),
            .I(N__87615));
    LocalMux I__21035 (
            .O(N__87920),
            .I(N__87610));
    LocalMux I__21034 (
            .O(N__87915),
            .I(N__87610));
    InMux I__21033 (
            .O(N__87914),
            .I(N__87607));
    LocalMux I__21032 (
            .O(N__87911),
            .I(N__87604));
    LocalMux I__21031 (
            .O(N__87904),
            .I(N__87601));
    InMux I__21030 (
            .O(N__87903),
            .I(N__87596));
    InMux I__21029 (
            .O(N__87902),
            .I(N__87596));
    LocalMux I__21028 (
            .O(N__87897),
            .I(N__87591));
    LocalMux I__21027 (
            .O(N__87892),
            .I(N__87586));
    LocalMux I__21026 (
            .O(N__87887),
            .I(N__87586));
    InMux I__21025 (
            .O(N__87886),
            .I(N__87583));
    Span4Mux_h I__21024 (
            .O(N__87883),
            .I(N__87569));
    Span4Mux_v I__21023 (
            .O(N__87880),
            .I(N__87569));
    Span4Mux_v I__21022 (
            .O(N__87871),
            .I(N__87569));
    Span4Mux_h I__21021 (
            .O(N__87862),
            .I(N__87562));
    Span4Mux_v I__21020 (
            .O(N__87847),
            .I(N__87562));
    LocalMux I__21019 (
            .O(N__87844),
            .I(N__87562));
    Span4Mux_v I__21018 (
            .O(N__87841),
            .I(N__87553));
    Span4Mux_h I__21017 (
            .O(N__87836),
            .I(N__87553));
    LocalMux I__21016 (
            .O(N__87833),
            .I(N__87553));
    LocalMux I__21015 (
            .O(N__87830),
            .I(N__87553));
    Span4Mux_h I__21014 (
            .O(N__87823),
            .I(N__87544));
    LocalMux I__21013 (
            .O(N__87820),
            .I(N__87544));
    LocalMux I__21012 (
            .O(N__87815),
            .I(N__87544));
    LocalMux I__21011 (
            .O(N__87810),
            .I(N__87544));
    Span4Mux_v I__21010 (
            .O(N__87805),
            .I(N__87537));
    Span4Mux_h I__21009 (
            .O(N__87800),
            .I(N__87537));
    LocalMux I__21008 (
            .O(N__87797),
            .I(N__87537));
    InMux I__21007 (
            .O(N__87794),
            .I(N__87534));
    InMux I__21006 (
            .O(N__87793),
            .I(N__87531));
    CascadeMux I__21005 (
            .O(N__87792),
            .I(N__87524));
    CascadeMux I__21004 (
            .O(N__87791),
            .I(N__87521));
    Span4Mux_h I__21003 (
            .O(N__87784),
            .I(N__87512));
    Span4Mux_v I__21002 (
            .O(N__87781),
            .I(N__87512));
    LocalMux I__21001 (
            .O(N__87776),
            .I(N__87512));
    LocalMux I__21000 (
            .O(N__87771),
            .I(N__87512));
    LocalMux I__20999 (
            .O(N__87768),
            .I(N__87507));
    LocalMux I__20998 (
            .O(N__87763),
            .I(N__87507));
    LocalMux I__20997 (
            .O(N__87760),
            .I(N__87502));
    LocalMux I__20996 (
            .O(N__87757),
            .I(N__87502));
    InMux I__20995 (
            .O(N__87756),
            .I(N__87497));
    InMux I__20994 (
            .O(N__87755),
            .I(N__87497));
    InMux I__20993 (
            .O(N__87754),
            .I(N__87492));
    InMux I__20992 (
            .O(N__87753),
            .I(N__87492));
    InMux I__20991 (
            .O(N__87752),
            .I(N__87489));
    CascadeMux I__20990 (
            .O(N__87751),
            .I(N__87486));
    LocalMux I__20989 (
            .O(N__87742),
            .I(N__87481));
    LocalMux I__20988 (
            .O(N__87737),
            .I(N__87481));
    InMux I__20987 (
            .O(N__87736),
            .I(N__87476));
    InMux I__20986 (
            .O(N__87735),
            .I(N__87476));
    InMux I__20985 (
            .O(N__87734),
            .I(N__87473));
    CascadeMux I__20984 (
            .O(N__87733),
            .I(N__87469));
    Span4Mux_v I__20983 (
            .O(N__87730),
            .I(N__87460));
    LocalMux I__20982 (
            .O(N__87727),
            .I(N__87460));
    InMux I__20981 (
            .O(N__87726),
            .I(N__87457));
    LocalMux I__20980 (
            .O(N__87723),
            .I(N__87452));
    LocalMux I__20979 (
            .O(N__87718),
            .I(N__87452));
    InMux I__20978 (
            .O(N__87717),
            .I(N__87447));
    InMux I__20977 (
            .O(N__87716),
            .I(N__87447));
    InMux I__20976 (
            .O(N__87715),
            .I(N__87441));
    InMux I__20975 (
            .O(N__87714),
            .I(N__87436));
    InMux I__20974 (
            .O(N__87713),
            .I(N__87436));
    CascadeMux I__20973 (
            .O(N__87712),
            .I(N__87433));
    Span4Mux_v I__20972 (
            .O(N__87709),
            .I(N__87412));
    Span4Mux_h I__20971 (
            .O(N__87702),
            .I(N__87412));
    LocalMux I__20970 (
            .O(N__87699),
            .I(N__87412));
    LocalMux I__20969 (
            .O(N__87694),
            .I(N__87412));
    LocalMux I__20968 (
            .O(N__87689),
            .I(N__87407));
    LocalMux I__20967 (
            .O(N__87684),
            .I(N__87407));
    LocalMux I__20966 (
            .O(N__87679),
            .I(N__87404));
    InMux I__20965 (
            .O(N__87678),
            .I(N__87397));
    InMux I__20964 (
            .O(N__87677),
            .I(N__87397));
    InMux I__20963 (
            .O(N__87676),
            .I(N__87397));
    LocalMux I__20962 (
            .O(N__87667),
            .I(N__87389));
    InMux I__20961 (
            .O(N__87666),
            .I(N__87384));
    InMux I__20960 (
            .O(N__87665),
            .I(N__87384));
    InMux I__20959 (
            .O(N__87664),
            .I(N__87379));
    InMux I__20958 (
            .O(N__87663),
            .I(N__87379));
    InMux I__20957 (
            .O(N__87662),
            .I(N__87374));
    InMux I__20956 (
            .O(N__87661),
            .I(N__87374));
    Span4Mux_v I__20955 (
            .O(N__87658),
            .I(N__87369));
    Span4Mux_v I__20954 (
            .O(N__87651),
            .I(N__87369));
    InMux I__20953 (
            .O(N__87650),
            .I(N__87362));
    InMux I__20952 (
            .O(N__87649),
            .I(N__87362));
    InMux I__20951 (
            .O(N__87648),
            .I(N__87362));
    InMux I__20950 (
            .O(N__87647),
            .I(N__87357));
    InMux I__20949 (
            .O(N__87646),
            .I(N__87357));
    LocalMux I__20948 (
            .O(N__87643),
            .I(N__87351));
    Span4Mux_h I__20947 (
            .O(N__87634),
            .I(N__87344));
    Span4Mux_v I__20946 (
            .O(N__87627),
            .I(N__87344));
    Span4Mux_v I__20945 (
            .O(N__87620),
            .I(N__87344));
    Span4Mux_h I__20944 (
            .O(N__87615),
            .I(N__87337));
    Span4Mux_h I__20943 (
            .O(N__87610),
            .I(N__87337));
    LocalMux I__20942 (
            .O(N__87607),
            .I(N__87337));
    Span4Mux_v I__20941 (
            .O(N__87604),
            .I(N__87327));
    Span4Mux_v I__20940 (
            .O(N__87601),
            .I(N__87327));
    LocalMux I__20939 (
            .O(N__87596),
            .I(N__87327));
    InMux I__20938 (
            .O(N__87595),
            .I(N__87322));
    InMux I__20937 (
            .O(N__87594),
            .I(N__87322));
    Span4Mux_v I__20936 (
            .O(N__87591),
            .I(N__87315));
    Span4Mux_v I__20935 (
            .O(N__87586),
            .I(N__87315));
    LocalMux I__20934 (
            .O(N__87583),
            .I(N__87315));
    InMux I__20933 (
            .O(N__87582),
            .I(N__87306));
    InMux I__20932 (
            .O(N__87581),
            .I(N__87306));
    InMux I__20931 (
            .O(N__87580),
            .I(N__87306));
    InMux I__20930 (
            .O(N__87579),
            .I(N__87306));
    InMux I__20929 (
            .O(N__87578),
            .I(N__87303));
    InMux I__20928 (
            .O(N__87577),
            .I(N__87291));
    InMux I__20927 (
            .O(N__87576),
            .I(N__87291));
    Span4Mux_h I__20926 (
            .O(N__87569),
            .I(N__87276));
    Span4Mux_v I__20925 (
            .O(N__87562),
            .I(N__87276));
    Span4Mux_v I__20924 (
            .O(N__87553),
            .I(N__87276));
    Span4Mux_h I__20923 (
            .O(N__87544),
            .I(N__87276));
    Span4Mux_h I__20922 (
            .O(N__87537),
            .I(N__87276));
    LocalMux I__20921 (
            .O(N__87534),
            .I(N__87276));
    LocalMux I__20920 (
            .O(N__87531),
            .I(N__87276));
    InMux I__20919 (
            .O(N__87530),
            .I(N__87269));
    InMux I__20918 (
            .O(N__87529),
            .I(N__87269));
    InMux I__20917 (
            .O(N__87528),
            .I(N__87269));
    InMux I__20916 (
            .O(N__87527),
            .I(N__87266));
    InMux I__20915 (
            .O(N__87524),
            .I(N__87263));
    InMux I__20914 (
            .O(N__87521),
            .I(N__87260));
    Span4Mux_v I__20913 (
            .O(N__87512),
            .I(N__87246));
    Span4Mux_v I__20912 (
            .O(N__87507),
            .I(N__87246));
    Span4Mux_v I__20911 (
            .O(N__87502),
            .I(N__87246));
    LocalMux I__20910 (
            .O(N__87497),
            .I(N__87246));
    LocalMux I__20909 (
            .O(N__87492),
            .I(N__87246));
    LocalMux I__20908 (
            .O(N__87489),
            .I(N__87246));
    InMux I__20907 (
            .O(N__87486),
            .I(N__87243));
    Span4Mux_v I__20906 (
            .O(N__87481),
            .I(N__87238));
    LocalMux I__20905 (
            .O(N__87476),
            .I(N__87238));
    LocalMux I__20904 (
            .O(N__87473),
            .I(N__87235));
    InMux I__20903 (
            .O(N__87472),
            .I(N__87230));
    InMux I__20902 (
            .O(N__87469),
            .I(N__87230));
    CascadeMux I__20901 (
            .O(N__87468),
            .I(N__87227));
    CascadeMux I__20900 (
            .O(N__87467),
            .I(N__87224));
    InMux I__20899 (
            .O(N__87466),
            .I(N__87218));
    InMux I__20898 (
            .O(N__87465),
            .I(N__87218));
    Span4Mux_v I__20897 (
            .O(N__87460),
            .I(N__87211));
    LocalMux I__20896 (
            .O(N__87457),
            .I(N__87211));
    Span4Mux_h I__20895 (
            .O(N__87452),
            .I(N__87206));
    LocalMux I__20894 (
            .O(N__87447),
            .I(N__87206));
    InMux I__20893 (
            .O(N__87446),
            .I(N__87199));
    InMux I__20892 (
            .O(N__87445),
            .I(N__87199));
    InMux I__20891 (
            .O(N__87444),
            .I(N__87199));
    LocalMux I__20890 (
            .O(N__87441),
            .I(N__87194));
    LocalMux I__20889 (
            .O(N__87436),
            .I(N__87194));
    InMux I__20888 (
            .O(N__87433),
            .I(N__87189));
    InMux I__20887 (
            .O(N__87432),
            .I(N__87189));
    InMux I__20886 (
            .O(N__87431),
            .I(N__87186));
    InMux I__20885 (
            .O(N__87430),
            .I(N__87179));
    InMux I__20884 (
            .O(N__87429),
            .I(N__87179));
    InMux I__20883 (
            .O(N__87428),
            .I(N__87179));
    InMux I__20882 (
            .O(N__87427),
            .I(N__87170));
    InMux I__20881 (
            .O(N__87426),
            .I(N__87170));
    InMux I__20880 (
            .O(N__87425),
            .I(N__87165));
    InMux I__20879 (
            .O(N__87424),
            .I(N__87165));
    InMux I__20878 (
            .O(N__87423),
            .I(N__87158));
    InMux I__20877 (
            .O(N__87422),
            .I(N__87158));
    InMux I__20876 (
            .O(N__87421),
            .I(N__87158));
    Span4Mux_h I__20875 (
            .O(N__87412),
            .I(N__87149));
    Span4Mux_v I__20874 (
            .O(N__87407),
            .I(N__87149));
    Span4Mux_v I__20873 (
            .O(N__87404),
            .I(N__87149));
    LocalMux I__20872 (
            .O(N__87397),
            .I(N__87149));
    InMux I__20871 (
            .O(N__87396),
            .I(N__87144));
    InMux I__20870 (
            .O(N__87395),
            .I(N__87144));
    InMux I__20869 (
            .O(N__87394),
            .I(N__87139));
    InMux I__20868 (
            .O(N__87393),
            .I(N__87139));
    InMux I__20867 (
            .O(N__87392),
            .I(N__87136));
    Span4Mux_v I__20866 (
            .O(N__87389),
            .I(N__87131));
    LocalMux I__20865 (
            .O(N__87384),
            .I(N__87131));
    LocalMux I__20864 (
            .O(N__87379),
            .I(N__87120));
    LocalMux I__20863 (
            .O(N__87374),
            .I(N__87120));
    Span4Mux_h I__20862 (
            .O(N__87369),
            .I(N__87120));
    LocalMux I__20861 (
            .O(N__87362),
            .I(N__87120));
    LocalMux I__20860 (
            .O(N__87357),
            .I(N__87120));
    InMux I__20859 (
            .O(N__87356),
            .I(N__87117));
    InMux I__20858 (
            .O(N__87355),
            .I(N__87114));
    CascadeMux I__20857 (
            .O(N__87354),
            .I(N__87111));
    Span4Mux_v I__20856 (
            .O(N__87351),
            .I(N__87108));
    Span4Mux_h I__20855 (
            .O(N__87344),
            .I(N__87103));
    Span4Mux_h I__20854 (
            .O(N__87337),
            .I(N__87103));
    InMux I__20853 (
            .O(N__87336),
            .I(N__87098));
    InMux I__20852 (
            .O(N__87335),
            .I(N__87098));
    InMux I__20851 (
            .O(N__87334),
            .I(N__87095));
    Span4Mux_v I__20850 (
            .O(N__87327),
            .I(N__87092));
    LocalMux I__20849 (
            .O(N__87322),
            .I(N__87089));
    Span4Mux_v I__20848 (
            .O(N__87315),
            .I(N__87082));
    LocalMux I__20847 (
            .O(N__87306),
            .I(N__87082));
    LocalMux I__20846 (
            .O(N__87303),
            .I(N__87082));
    InMux I__20845 (
            .O(N__87302),
            .I(N__87077));
    InMux I__20844 (
            .O(N__87301),
            .I(N__87077));
    InMux I__20843 (
            .O(N__87300),
            .I(N__87070));
    InMux I__20842 (
            .O(N__87299),
            .I(N__87070));
    InMux I__20841 (
            .O(N__87298),
            .I(N__87070));
    InMux I__20840 (
            .O(N__87297),
            .I(N__87067));
    CascadeMux I__20839 (
            .O(N__87296),
            .I(N__87064));
    LocalMux I__20838 (
            .O(N__87291),
            .I(N__87056));
    Span4Mux_h I__20837 (
            .O(N__87276),
            .I(N__87056));
    LocalMux I__20836 (
            .O(N__87269),
            .I(N__87056));
    LocalMux I__20835 (
            .O(N__87266),
            .I(N__87053));
    LocalMux I__20834 (
            .O(N__87263),
            .I(N__87048));
    LocalMux I__20833 (
            .O(N__87260),
            .I(N__87048));
    InMux I__20832 (
            .O(N__87259),
            .I(N__87045));
    Span4Mux_v I__20831 (
            .O(N__87246),
            .I(N__87042));
    LocalMux I__20830 (
            .O(N__87243),
            .I(N__87039));
    Span4Mux_h I__20829 (
            .O(N__87238),
            .I(N__87032));
    Span4Mux_v I__20828 (
            .O(N__87235),
            .I(N__87032));
    LocalMux I__20827 (
            .O(N__87230),
            .I(N__87032));
    InMux I__20826 (
            .O(N__87227),
            .I(N__87027));
    InMux I__20825 (
            .O(N__87224),
            .I(N__87027));
    InMux I__20824 (
            .O(N__87223),
            .I(N__87024));
    LocalMux I__20823 (
            .O(N__87218),
            .I(N__87021));
    InMux I__20822 (
            .O(N__87217),
            .I(N__87016));
    InMux I__20821 (
            .O(N__87216),
            .I(N__87016));
    Span4Mux_v I__20820 (
            .O(N__87211),
            .I(N__87008));
    Span4Mux_v I__20819 (
            .O(N__87206),
            .I(N__87008));
    LocalMux I__20818 (
            .O(N__87199),
            .I(N__87008));
    Span4Mux_v I__20817 (
            .O(N__87194),
            .I(N__87001));
    LocalMux I__20816 (
            .O(N__87189),
            .I(N__87001));
    LocalMux I__20815 (
            .O(N__87186),
            .I(N__87001));
    LocalMux I__20814 (
            .O(N__87179),
            .I(N__86998));
    InMux I__20813 (
            .O(N__87178),
            .I(N__86993));
    InMux I__20812 (
            .O(N__87177),
            .I(N__86993));
    InMux I__20811 (
            .O(N__87176),
            .I(N__86990));
    CascadeMux I__20810 (
            .O(N__87175),
            .I(N__86985));
    LocalMux I__20809 (
            .O(N__87170),
            .I(N__86979));
    LocalMux I__20808 (
            .O(N__87165),
            .I(N__86974));
    LocalMux I__20807 (
            .O(N__87158),
            .I(N__86974));
    Sp12to4 I__20806 (
            .O(N__87149),
            .I(N__86965));
    LocalMux I__20805 (
            .O(N__87144),
            .I(N__86965));
    LocalMux I__20804 (
            .O(N__87139),
            .I(N__86965));
    LocalMux I__20803 (
            .O(N__87136),
            .I(N__86965));
    Span4Mux_h I__20802 (
            .O(N__87131),
            .I(N__86956));
    Span4Mux_v I__20801 (
            .O(N__87120),
            .I(N__86956));
    LocalMux I__20800 (
            .O(N__87117),
            .I(N__86956));
    LocalMux I__20799 (
            .O(N__87114),
            .I(N__86956));
    InMux I__20798 (
            .O(N__87111),
            .I(N__86953));
    Span4Mux_v I__20797 (
            .O(N__87108),
            .I(N__86950));
    Span4Mux_v I__20796 (
            .O(N__87103),
            .I(N__86945));
    LocalMux I__20795 (
            .O(N__87098),
            .I(N__86945));
    LocalMux I__20794 (
            .O(N__87095),
            .I(N__86942));
    Span4Mux_h I__20793 (
            .O(N__87092),
            .I(N__86929));
    Span4Mux_h I__20792 (
            .O(N__87089),
            .I(N__86929));
    Span4Mux_v I__20791 (
            .O(N__87082),
            .I(N__86929));
    LocalMux I__20790 (
            .O(N__87077),
            .I(N__86929));
    LocalMux I__20789 (
            .O(N__87070),
            .I(N__86929));
    LocalMux I__20788 (
            .O(N__87067),
            .I(N__86929));
    InMux I__20787 (
            .O(N__87064),
            .I(N__86926));
    InMux I__20786 (
            .O(N__87063),
            .I(N__86923));
    Span4Mux_v I__20785 (
            .O(N__87056),
            .I(N__86916));
    Span4Mux_v I__20784 (
            .O(N__87053),
            .I(N__86909));
    Span4Mux_v I__20783 (
            .O(N__87048),
            .I(N__86909));
    LocalMux I__20782 (
            .O(N__87045),
            .I(N__86909));
    Span4Mux_v I__20781 (
            .O(N__87042),
            .I(N__86898));
    Span4Mux_v I__20780 (
            .O(N__87039),
            .I(N__86898));
    Span4Mux_h I__20779 (
            .O(N__87032),
            .I(N__86898));
    LocalMux I__20778 (
            .O(N__87027),
            .I(N__86898));
    LocalMux I__20777 (
            .O(N__87024),
            .I(N__86898));
    Span4Mux_v I__20776 (
            .O(N__87021),
            .I(N__86893));
    LocalMux I__20775 (
            .O(N__87016),
            .I(N__86893));
    InMux I__20774 (
            .O(N__87015),
            .I(N__86890));
    Span4Mux_h I__20773 (
            .O(N__87008),
            .I(N__86879));
    Span4Mux_v I__20772 (
            .O(N__87001),
            .I(N__86879));
    Span4Mux_v I__20771 (
            .O(N__86998),
            .I(N__86879));
    LocalMux I__20770 (
            .O(N__86993),
            .I(N__86879));
    LocalMux I__20769 (
            .O(N__86990),
            .I(N__86879));
    InMux I__20768 (
            .O(N__86989),
            .I(N__86872));
    InMux I__20767 (
            .O(N__86988),
            .I(N__86872));
    InMux I__20766 (
            .O(N__86985),
            .I(N__86872));
    InMux I__20765 (
            .O(N__86984),
            .I(N__86867));
    InMux I__20764 (
            .O(N__86983),
            .I(N__86867));
    CascadeMux I__20763 (
            .O(N__86982),
            .I(N__86863));
    Span4Mux_v I__20762 (
            .O(N__86979),
            .I(N__86855));
    Span12Mux_h I__20761 (
            .O(N__86974),
            .I(N__86846));
    Span12Mux_v I__20760 (
            .O(N__86965),
            .I(N__86846));
    Sp12to4 I__20759 (
            .O(N__86956),
            .I(N__86846));
    LocalMux I__20758 (
            .O(N__86953),
            .I(N__86846));
    Span4Mux_v I__20757 (
            .O(N__86950),
            .I(N__86841));
    Span4Mux_v I__20756 (
            .O(N__86945),
            .I(N__86841));
    Span4Mux_h I__20755 (
            .O(N__86942),
            .I(N__86832));
    Span4Mux_h I__20754 (
            .O(N__86929),
            .I(N__86832));
    LocalMux I__20753 (
            .O(N__86926),
            .I(N__86832));
    LocalMux I__20752 (
            .O(N__86923),
            .I(N__86832));
    InMux I__20751 (
            .O(N__86922),
            .I(N__86827));
    InMux I__20750 (
            .O(N__86921),
            .I(N__86827));
    InMux I__20749 (
            .O(N__86920),
            .I(N__86822));
    InMux I__20748 (
            .O(N__86919),
            .I(N__86822));
    Span4Mux_v I__20747 (
            .O(N__86916),
            .I(N__86811));
    Span4Mux_v I__20746 (
            .O(N__86909),
            .I(N__86811));
    Span4Mux_v I__20745 (
            .O(N__86898),
            .I(N__86811));
    Span4Mux_v I__20744 (
            .O(N__86893),
            .I(N__86811));
    LocalMux I__20743 (
            .O(N__86890),
            .I(N__86811));
    Span4Mux_h I__20742 (
            .O(N__86879),
            .I(N__86804));
    LocalMux I__20741 (
            .O(N__86872),
            .I(N__86804));
    LocalMux I__20740 (
            .O(N__86867),
            .I(N__86804));
    InMux I__20739 (
            .O(N__86866),
            .I(N__86801));
    InMux I__20738 (
            .O(N__86863),
            .I(N__86798));
    InMux I__20737 (
            .O(N__86862),
            .I(N__86795));
    InMux I__20736 (
            .O(N__86861),
            .I(N__86792));
    InMux I__20735 (
            .O(N__86860),
            .I(N__86785));
    InMux I__20734 (
            .O(N__86859),
            .I(N__86785));
    InMux I__20733 (
            .O(N__86858),
            .I(N__86785));
    Odrv4 I__20732 (
            .O(N__86855),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    Odrv12 I__20731 (
            .O(N__86846),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    Odrv4 I__20730 (
            .O(N__86841),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    Odrv4 I__20729 (
            .O(N__86832),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    LocalMux I__20728 (
            .O(N__86827),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    LocalMux I__20727 (
            .O(N__86822),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    Odrv4 I__20726 (
            .O(N__86811),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    Odrv4 I__20725 (
            .O(N__86804),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    LocalMux I__20724 (
            .O(N__86801),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    LocalMux I__20723 (
            .O(N__86798),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    LocalMux I__20722 (
            .O(N__86795),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    LocalMux I__20721 (
            .O(N__86792),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    LocalMux I__20720 (
            .O(N__86785),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ));
    InMux I__20719 (
            .O(N__86758),
            .I(N__86755));
    LocalMux I__20718 (
            .O(N__86755),
            .I(N__86752));
    Span12Mux_v I__20717 (
            .O(N__86752),
            .I(N__86749));
    Odrv12 I__20716 (
            .O(N__86749),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11725 ));
    InMux I__20715 (
            .O(N__86746),
            .I(\timing_controller_inst.n10614 ));
    InMux I__20714 (
            .O(N__86743),
            .I(N__86740));
    LocalMux I__20713 (
            .O(N__86740),
            .I(N__86737));
    Span4Mux_v I__20712 (
            .O(N__86737),
            .I(N__86733));
    CascadeMux I__20711 (
            .O(N__86736),
            .I(N__86730));
    Span4Mux_h I__20710 (
            .O(N__86733),
            .I(N__86727));
    InMux I__20709 (
            .O(N__86730),
            .I(N__86724));
    Odrv4 I__20708 (
            .O(N__86727),
            .I(\timing_controller_inst.state_timeout_counter_28 ));
    LocalMux I__20707 (
            .O(N__86724),
            .I(\timing_controller_inst.state_timeout_counter_28 ));
    InMux I__20706 (
            .O(N__86719),
            .I(\timing_controller_inst.n10615 ));
    InMux I__20705 (
            .O(N__86716),
            .I(N__86713));
    LocalMux I__20704 (
            .O(N__86713),
            .I(N__86710));
    Span4Mux_h I__20703 (
            .O(N__86710),
            .I(N__86706));
    InMux I__20702 (
            .O(N__86709),
            .I(N__86703));
    Odrv4 I__20701 (
            .O(N__86706),
            .I(\timing_controller_inst.state_timeout_counter_29 ));
    LocalMux I__20700 (
            .O(N__86703),
            .I(\timing_controller_inst.state_timeout_counter_29 ));
    InMux I__20699 (
            .O(N__86698),
            .I(\timing_controller_inst.n10616 ));
    CascadeMux I__20698 (
            .O(N__86695),
            .I(N__86692));
    InMux I__20697 (
            .O(N__86692),
            .I(N__86689));
    LocalMux I__20696 (
            .O(N__86689),
            .I(N__86685));
    CascadeMux I__20695 (
            .O(N__86688),
            .I(N__86682));
    Span4Mux_v I__20694 (
            .O(N__86685),
            .I(N__86679));
    InMux I__20693 (
            .O(N__86682),
            .I(N__86676));
    Odrv4 I__20692 (
            .O(N__86679),
            .I(\timing_controller_inst.state_timeout_counter_30 ));
    LocalMux I__20691 (
            .O(N__86676),
            .I(\timing_controller_inst.state_timeout_counter_30 ));
    InMux I__20690 (
            .O(N__86671),
            .I(\timing_controller_inst.n10617 ));
    IoInMux I__20689 (
            .O(N__86668),
            .I(N__86665));
    LocalMux I__20688 (
            .O(N__86665),
            .I(N__86652));
    IoInMux I__20687 (
            .O(N__86664),
            .I(N__86649));
    IoInMux I__20686 (
            .O(N__86663),
            .I(N__86646));
    CascadeMux I__20685 (
            .O(N__86662),
            .I(N__86642));
    CascadeMux I__20684 (
            .O(N__86661),
            .I(N__86639));
    CascadeMux I__20683 (
            .O(N__86660),
            .I(N__86636));
    CascadeMux I__20682 (
            .O(N__86659),
            .I(N__86633));
    CascadeMux I__20681 (
            .O(N__86658),
            .I(N__86630));
    CascadeMux I__20680 (
            .O(N__86657),
            .I(N__86627));
    CascadeMux I__20679 (
            .O(N__86656),
            .I(N__86624));
    CascadeMux I__20678 (
            .O(N__86655),
            .I(N__86621));
    IoSpan4Mux I__20677 (
            .O(N__86652),
            .I(N__86618));
    LocalMux I__20676 (
            .O(N__86649),
            .I(N__86615));
    LocalMux I__20675 (
            .O(N__86646),
            .I(N__86612));
    InMux I__20674 (
            .O(N__86645),
            .I(N__86607));
    InMux I__20673 (
            .O(N__86642),
            .I(N__86607));
    InMux I__20672 (
            .O(N__86639),
            .I(N__86600));
    InMux I__20671 (
            .O(N__86636),
            .I(N__86600));
    InMux I__20670 (
            .O(N__86633),
            .I(N__86600));
    InMux I__20669 (
            .O(N__86630),
            .I(N__86591));
    InMux I__20668 (
            .O(N__86627),
            .I(N__86591));
    InMux I__20667 (
            .O(N__86624),
            .I(N__86591));
    InMux I__20666 (
            .O(N__86621),
            .I(N__86591));
    Span4Mux_s1_h I__20665 (
            .O(N__86618),
            .I(N__86579));
    Span4Mux_s1_h I__20664 (
            .O(N__86615),
            .I(N__86576));
    Span4Mux_s2_v I__20663 (
            .O(N__86612),
            .I(N__86568));
    LocalMux I__20662 (
            .O(N__86607),
            .I(N__86565));
    LocalMux I__20661 (
            .O(N__86600),
            .I(N__86560));
    LocalMux I__20660 (
            .O(N__86591),
            .I(N__86560));
    CascadeMux I__20659 (
            .O(N__86590),
            .I(N__86556));
    CascadeMux I__20658 (
            .O(N__86589),
            .I(N__86546));
    CascadeMux I__20657 (
            .O(N__86588),
            .I(N__86536));
    CascadeMux I__20656 (
            .O(N__86587),
            .I(N__86533));
    CascadeMux I__20655 (
            .O(N__86586),
            .I(N__86525));
    CascadeMux I__20654 (
            .O(N__86585),
            .I(N__86522));
    CascadeMux I__20653 (
            .O(N__86584),
            .I(N__86518));
    CascadeMux I__20652 (
            .O(N__86583),
            .I(N__86514));
    CascadeMux I__20651 (
            .O(N__86582),
            .I(N__86510));
    Sp12to4 I__20650 (
            .O(N__86579),
            .I(N__86501));
    Sp12to4 I__20649 (
            .O(N__86576),
            .I(N__86501));
    CascadeMux I__20648 (
            .O(N__86575),
            .I(N__86497));
    CascadeMux I__20647 (
            .O(N__86574),
            .I(N__86493));
    CascadeMux I__20646 (
            .O(N__86573),
            .I(N__86489));
    CascadeMux I__20645 (
            .O(N__86572),
            .I(N__86485));
    CascadeMux I__20644 (
            .O(N__86571),
            .I(N__86481));
    Span4Mux_v I__20643 (
            .O(N__86568),
            .I(N__86478));
    Span4Mux_v I__20642 (
            .O(N__86565),
            .I(N__86473));
    Span4Mux_v I__20641 (
            .O(N__86560),
            .I(N__86473));
    InMux I__20640 (
            .O(N__86559),
            .I(N__86470));
    InMux I__20639 (
            .O(N__86556),
            .I(N__86467));
    InMux I__20638 (
            .O(N__86555),
            .I(N__86460));
    InMux I__20637 (
            .O(N__86554),
            .I(N__86460));
    InMux I__20636 (
            .O(N__86553),
            .I(N__86460));
    InMux I__20635 (
            .O(N__86552),
            .I(N__86449));
    InMux I__20634 (
            .O(N__86551),
            .I(N__86449));
    InMux I__20633 (
            .O(N__86550),
            .I(N__86449));
    InMux I__20632 (
            .O(N__86549),
            .I(N__86449));
    InMux I__20631 (
            .O(N__86546),
            .I(N__86449));
    InMux I__20630 (
            .O(N__86545),
            .I(N__86442));
    InMux I__20629 (
            .O(N__86544),
            .I(N__86442));
    InMux I__20628 (
            .O(N__86543),
            .I(N__86442));
    InMux I__20627 (
            .O(N__86542),
            .I(N__86431));
    InMux I__20626 (
            .O(N__86541),
            .I(N__86431));
    InMux I__20625 (
            .O(N__86540),
            .I(N__86431));
    InMux I__20624 (
            .O(N__86539),
            .I(N__86431));
    InMux I__20623 (
            .O(N__86536),
            .I(N__86431));
    InMux I__20622 (
            .O(N__86533),
            .I(N__86416));
    InMux I__20621 (
            .O(N__86532),
            .I(N__86416));
    InMux I__20620 (
            .O(N__86531),
            .I(N__86416));
    InMux I__20619 (
            .O(N__86530),
            .I(N__86416));
    InMux I__20618 (
            .O(N__86529),
            .I(N__86409));
    InMux I__20617 (
            .O(N__86528),
            .I(N__86409));
    InMux I__20616 (
            .O(N__86525),
            .I(N__86409));
    InMux I__20615 (
            .O(N__86522),
            .I(N__86394));
    InMux I__20614 (
            .O(N__86521),
            .I(N__86394));
    InMux I__20613 (
            .O(N__86518),
            .I(N__86394));
    InMux I__20612 (
            .O(N__86517),
            .I(N__86394));
    InMux I__20611 (
            .O(N__86514),
            .I(N__86394));
    InMux I__20610 (
            .O(N__86513),
            .I(N__86394));
    InMux I__20609 (
            .O(N__86510),
            .I(N__86394));
    CascadeMux I__20608 (
            .O(N__86509),
            .I(N__86391));
    CascadeMux I__20607 (
            .O(N__86508),
            .I(N__86386));
    CascadeMux I__20606 (
            .O(N__86507),
            .I(N__86382));
    CascadeMux I__20605 (
            .O(N__86506),
            .I(N__86378));
    Span12Mux_v I__20604 (
            .O(N__86501),
            .I(N__86357));
    InMux I__20603 (
            .O(N__86500),
            .I(N__86350));
    InMux I__20602 (
            .O(N__86497),
            .I(N__86350));
    InMux I__20601 (
            .O(N__86496),
            .I(N__86350));
    InMux I__20600 (
            .O(N__86493),
            .I(N__86335));
    InMux I__20599 (
            .O(N__86492),
            .I(N__86335));
    InMux I__20598 (
            .O(N__86489),
            .I(N__86335));
    InMux I__20597 (
            .O(N__86488),
            .I(N__86335));
    InMux I__20596 (
            .O(N__86485),
            .I(N__86335));
    InMux I__20595 (
            .O(N__86484),
            .I(N__86335));
    InMux I__20594 (
            .O(N__86481),
            .I(N__86335));
    Span4Mux_v I__20593 (
            .O(N__86478),
            .I(N__86318));
    Span4Mux_h I__20592 (
            .O(N__86473),
            .I(N__86318));
    LocalMux I__20591 (
            .O(N__86470),
            .I(N__86318));
    LocalMux I__20590 (
            .O(N__86467),
            .I(N__86318));
    LocalMux I__20589 (
            .O(N__86460),
            .I(N__86318));
    LocalMux I__20588 (
            .O(N__86449),
            .I(N__86318));
    LocalMux I__20587 (
            .O(N__86442),
            .I(N__86318));
    LocalMux I__20586 (
            .O(N__86431),
            .I(N__86318));
    CascadeMux I__20585 (
            .O(N__86430),
            .I(N__86314));
    CascadeMux I__20584 (
            .O(N__86429),
            .I(N__86310));
    CascadeMux I__20583 (
            .O(N__86428),
            .I(N__86306));
    CascadeMux I__20582 (
            .O(N__86427),
            .I(N__86302));
    CascadeMux I__20581 (
            .O(N__86426),
            .I(N__86299));
    CascadeMux I__20580 (
            .O(N__86425),
            .I(N__86296));
    LocalMux I__20579 (
            .O(N__86416),
            .I(N__86288));
    LocalMux I__20578 (
            .O(N__86409),
            .I(N__86288));
    LocalMux I__20577 (
            .O(N__86394),
            .I(N__86288));
    InMux I__20576 (
            .O(N__86391),
            .I(N__86283));
    InMux I__20575 (
            .O(N__86390),
            .I(N__86283));
    InMux I__20574 (
            .O(N__86389),
            .I(N__86270));
    InMux I__20573 (
            .O(N__86386),
            .I(N__86270));
    InMux I__20572 (
            .O(N__86385),
            .I(N__86270));
    InMux I__20571 (
            .O(N__86382),
            .I(N__86270));
    InMux I__20570 (
            .O(N__86381),
            .I(N__86270));
    InMux I__20569 (
            .O(N__86378),
            .I(N__86270));
    CascadeMux I__20568 (
            .O(N__86377),
            .I(N__86267));
    CascadeMux I__20567 (
            .O(N__86376),
            .I(N__86264));
    CascadeMux I__20566 (
            .O(N__86375),
            .I(N__86261));
    CascadeMux I__20565 (
            .O(N__86374),
            .I(N__86258));
    CascadeMux I__20564 (
            .O(N__86373),
            .I(N__86255));
    CascadeMux I__20563 (
            .O(N__86372),
            .I(N__86251));
    CascadeMux I__20562 (
            .O(N__86371),
            .I(N__86248));
    CascadeMux I__20561 (
            .O(N__86370),
            .I(N__86245));
    CascadeMux I__20560 (
            .O(N__86369),
            .I(N__86242));
    CascadeMux I__20559 (
            .O(N__86368),
            .I(N__86239));
    CascadeMux I__20558 (
            .O(N__86367),
            .I(N__86236));
    CascadeMux I__20557 (
            .O(N__86366),
            .I(N__86233));
    CascadeMux I__20556 (
            .O(N__86365),
            .I(N__86230));
    CascadeMux I__20555 (
            .O(N__86364),
            .I(N__86227));
    CascadeMux I__20554 (
            .O(N__86363),
            .I(N__86224));
    CascadeMux I__20553 (
            .O(N__86362),
            .I(N__86220));
    CascadeMux I__20552 (
            .O(N__86361),
            .I(N__86216));
    CascadeMux I__20551 (
            .O(N__86360),
            .I(N__86211));
    Span12Mux_h I__20550 (
            .O(N__86357),
            .I(N__86208));
    LocalMux I__20549 (
            .O(N__86350),
            .I(N__86203));
    LocalMux I__20548 (
            .O(N__86335),
            .I(N__86203));
    Span4Mux_v I__20547 (
            .O(N__86318),
            .I(N__86200));
    InMux I__20546 (
            .O(N__86317),
            .I(N__86183));
    InMux I__20545 (
            .O(N__86314),
            .I(N__86183));
    InMux I__20544 (
            .O(N__86313),
            .I(N__86183));
    InMux I__20543 (
            .O(N__86310),
            .I(N__86183));
    InMux I__20542 (
            .O(N__86309),
            .I(N__86183));
    InMux I__20541 (
            .O(N__86306),
            .I(N__86183));
    InMux I__20540 (
            .O(N__86305),
            .I(N__86183));
    InMux I__20539 (
            .O(N__86302),
            .I(N__86183));
    InMux I__20538 (
            .O(N__86299),
            .I(N__86180));
    InMux I__20537 (
            .O(N__86296),
            .I(N__86175));
    InMux I__20536 (
            .O(N__86295),
            .I(N__86175));
    Span4Mux_h I__20535 (
            .O(N__86288),
            .I(N__86172));
    LocalMux I__20534 (
            .O(N__86283),
            .I(N__86167));
    LocalMux I__20533 (
            .O(N__86270),
            .I(N__86167));
    InMux I__20532 (
            .O(N__86267),
            .I(N__86160));
    InMux I__20531 (
            .O(N__86264),
            .I(N__86160));
    InMux I__20530 (
            .O(N__86261),
            .I(N__86160));
    InMux I__20529 (
            .O(N__86258),
            .I(N__86149));
    InMux I__20528 (
            .O(N__86255),
            .I(N__86149));
    InMux I__20527 (
            .O(N__86254),
            .I(N__86149));
    InMux I__20526 (
            .O(N__86251),
            .I(N__86149));
    InMux I__20525 (
            .O(N__86248),
            .I(N__86149));
    InMux I__20524 (
            .O(N__86245),
            .I(N__86140));
    InMux I__20523 (
            .O(N__86242),
            .I(N__86140));
    InMux I__20522 (
            .O(N__86239),
            .I(N__86140));
    InMux I__20521 (
            .O(N__86236),
            .I(N__86140));
    InMux I__20520 (
            .O(N__86233),
            .I(N__86131));
    InMux I__20519 (
            .O(N__86230),
            .I(N__86131));
    InMux I__20518 (
            .O(N__86227),
            .I(N__86131));
    InMux I__20517 (
            .O(N__86224),
            .I(N__86131));
    InMux I__20516 (
            .O(N__86223),
            .I(N__86116));
    InMux I__20515 (
            .O(N__86220),
            .I(N__86116));
    InMux I__20514 (
            .O(N__86219),
            .I(N__86116));
    InMux I__20513 (
            .O(N__86216),
            .I(N__86116));
    InMux I__20512 (
            .O(N__86215),
            .I(N__86116));
    InMux I__20511 (
            .O(N__86214),
            .I(N__86116));
    InMux I__20510 (
            .O(N__86211),
            .I(N__86116));
    Span12Mux_h I__20509 (
            .O(N__86208),
            .I(N__86113));
    Span12Mux_v I__20508 (
            .O(N__86203),
            .I(N__86102));
    Sp12to4 I__20507 (
            .O(N__86200),
            .I(N__86102));
    LocalMux I__20506 (
            .O(N__86183),
            .I(N__86102));
    LocalMux I__20505 (
            .O(N__86180),
            .I(N__86102));
    LocalMux I__20504 (
            .O(N__86175),
            .I(N__86102));
    Span4Mux_h I__20503 (
            .O(N__86172),
            .I(N__86089));
    Span4Mux_v I__20502 (
            .O(N__86167),
            .I(N__86089));
    LocalMux I__20501 (
            .O(N__86160),
            .I(N__86089));
    LocalMux I__20500 (
            .O(N__86149),
            .I(N__86089));
    LocalMux I__20499 (
            .O(N__86140),
            .I(N__86089));
    LocalMux I__20498 (
            .O(N__86131),
            .I(N__86089));
    LocalMux I__20497 (
            .O(N__86116),
            .I(N__86086));
    Odrv12 I__20496 (
            .O(N__86113),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__20495 (
            .O(N__86102),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__20494 (
            .O(N__86089),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__20493 (
            .O(N__86086),
            .I(CONSTANT_ONE_NET));
    InMux I__20492 (
            .O(N__86077),
            .I(\timing_controller_inst.n10618 ));
    InMux I__20491 (
            .O(N__86074),
            .I(N__86071));
    LocalMux I__20490 (
            .O(N__86071),
            .I(N__86068));
    Span4Mux_v I__20489 (
            .O(N__86068),
            .I(N__86064));
    InMux I__20488 (
            .O(N__86067),
            .I(N__86061));
    Odrv4 I__20487 (
            .O(N__86064),
            .I(\timing_controller_inst.state_timeout_counter_31 ));
    LocalMux I__20486 (
            .O(N__86061),
            .I(\timing_controller_inst.state_timeout_counter_31 ));
    CEMux I__20485 (
            .O(N__86056),
            .I(N__86051));
    CEMux I__20484 (
            .O(N__86055),
            .I(N__86048));
    CEMux I__20483 (
            .O(N__86054),
            .I(N__86045));
    LocalMux I__20482 (
            .O(N__86051),
            .I(N__86040));
    LocalMux I__20481 (
            .O(N__86048),
            .I(N__86032));
    LocalMux I__20480 (
            .O(N__86045),
            .I(N__86032));
    CEMux I__20479 (
            .O(N__86044),
            .I(N__86029));
    CEMux I__20478 (
            .O(N__86043),
            .I(N__86026));
    Span4Mux_v I__20477 (
            .O(N__86040),
            .I(N__86023));
    CEMux I__20476 (
            .O(N__86039),
            .I(N__86020));
    CEMux I__20475 (
            .O(N__86038),
            .I(N__86017));
    CEMux I__20474 (
            .O(N__86037),
            .I(N__86014));
    Span4Mux_v I__20473 (
            .O(N__86032),
            .I(N__86011));
    LocalMux I__20472 (
            .O(N__86029),
            .I(N__86002));
    LocalMux I__20471 (
            .O(N__86026),
            .I(N__86002));
    Span4Mux_v I__20470 (
            .O(N__86023),
            .I(N__86002));
    LocalMux I__20469 (
            .O(N__86020),
            .I(N__86002));
    LocalMux I__20468 (
            .O(N__86017),
            .I(N__85997));
    LocalMux I__20467 (
            .O(N__86014),
            .I(N__85997));
    Span4Mux_h I__20466 (
            .O(N__86011),
            .I(N__85992));
    Span4Mux_v I__20465 (
            .O(N__86002),
            .I(N__85992));
    Span4Mux_h I__20464 (
            .O(N__85997),
            .I(N__85989));
    Odrv4 I__20463 (
            .O(N__85992),
            .I(\timing_controller_inst.n4301 ));
    Odrv4 I__20462 (
            .O(N__85989),
            .I(\timing_controller_inst.n4301 ));
    SRMux I__20461 (
            .O(N__85984),
            .I(N__85978));
    SRMux I__20460 (
            .O(N__85983),
            .I(N__85975));
    SRMux I__20459 (
            .O(N__85982),
            .I(N__85972));
    SRMux I__20458 (
            .O(N__85981),
            .I(N__85969));
    LocalMux I__20457 (
            .O(N__85978),
            .I(N__85966));
    LocalMux I__20456 (
            .O(N__85975),
            .I(N__85961));
    LocalMux I__20455 (
            .O(N__85972),
            .I(N__85961));
    LocalMux I__20454 (
            .O(N__85969),
            .I(N__85958));
    Span4Mux_v I__20453 (
            .O(N__85966),
            .I(N__85955));
    Span4Mux_v I__20452 (
            .O(N__85961),
            .I(N__85952));
    Span4Mux_h I__20451 (
            .O(N__85958),
            .I(N__85949));
    Odrv4 I__20450 (
            .O(N__85955),
            .I(\timing_controller_inst.n4589 ));
    Odrv4 I__20449 (
            .O(N__85952),
            .I(\timing_controller_inst.n4589 ));
    Odrv4 I__20448 (
            .O(N__85949),
            .I(\timing_controller_inst.n4589 ));
    InMux I__20447 (
            .O(N__85942),
            .I(N__85939));
    LocalMux I__20446 (
            .O(N__85939),
            .I(N__85936));
    Span12Mux_h I__20445 (
            .O(N__85936),
            .I(N__85932));
    InMux I__20444 (
            .O(N__85935),
            .I(N__85929));
    Odrv12 I__20443 (
            .O(N__85932),
            .I(REG_mem_43_8));
    LocalMux I__20442 (
            .O(N__85929),
            .I(REG_mem_43_8));
    InMux I__20441 (
            .O(N__85924),
            .I(N__85921));
    LocalMux I__20440 (
            .O(N__85921),
            .I(N__85918));
    Span4Mux_v I__20439 (
            .O(N__85918),
            .I(N__85914));
    InMux I__20438 (
            .O(N__85917),
            .I(N__85911));
    Span4Mux_h I__20437 (
            .O(N__85914),
            .I(N__85906));
    LocalMux I__20436 (
            .O(N__85911),
            .I(N__85906));
    Odrv4 I__20435 (
            .O(N__85906),
            .I(REG_mem_42_8));
    InMux I__20434 (
            .O(N__85903),
            .I(N__85900));
    LocalMux I__20433 (
            .O(N__85900),
            .I(N__85897));
    Span4Mux_v I__20432 (
            .O(N__85897),
            .I(N__85894));
    Sp12to4 I__20431 (
            .O(N__85894),
            .I(N__85890));
    InMux I__20430 (
            .O(N__85893),
            .I(N__85887));
    Odrv12 I__20429 (
            .O(N__85890),
            .I(REG_mem_40_8));
    LocalMux I__20428 (
            .O(N__85887),
            .I(REG_mem_40_8));
    CascadeMux I__20427 (
            .O(N__85882),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13724_cascade_ ));
    InMux I__20426 (
            .O(N__85879),
            .I(N__85876));
    LocalMux I__20425 (
            .O(N__85876),
            .I(N__85873));
    Span12Mux_s7_h I__20424 (
            .O(N__85873),
            .I(N__85869));
    InMux I__20423 (
            .O(N__85872),
            .I(N__85866));
    Odrv12 I__20422 (
            .O(N__85869),
            .I(REG_mem_41_8));
    LocalMux I__20421 (
            .O(N__85866),
            .I(REG_mem_41_8));
    InMux I__20420 (
            .O(N__85861),
            .I(N__85858));
    LocalMux I__20419 (
            .O(N__85858),
            .I(N__85839));
    InMux I__20418 (
            .O(N__85857),
            .I(N__85834));
    InMux I__20417 (
            .O(N__85856),
            .I(N__85834));
    InMux I__20416 (
            .O(N__85855),
            .I(N__85831));
    InMux I__20415 (
            .O(N__85854),
            .I(N__85828));
    InMux I__20414 (
            .O(N__85853),
            .I(N__85797));
    InMux I__20413 (
            .O(N__85852),
            .I(N__85797));
    InMux I__20412 (
            .O(N__85851),
            .I(N__85797));
    InMux I__20411 (
            .O(N__85850),
            .I(N__85788));
    InMux I__20410 (
            .O(N__85849),
            .I(N__85788));
    InMux I__20409 (
            .O(N__85848),
            .I(N__85788));
    InMux I__20408 (
            .O(N__85847),
            .I(N__85788));
    InMux I__20407 (
            .O(N__85846),
            .I(N__85785));
    InMux I__20406 (
            .O(N__85845),
            .I(N__85778));
    InMux I__20405 (
            .O(N__85844),
            .I(N__85778));
    InMux I__20404 (
            .O(N__85843),
            .I(N__85778));
    InMux I__20403 (
            .O(N__85842),
            .I(N__85775));
    Span4Mux_v I__20402 (
            .O(N__85839),
            .I(N__85766));
    LocalMux I__20401 (
            .O(N__85834),
            .I(N__85766));
    LocalMux I__20400 (
            .O(N__85831),
            .I(N__85766));
    LocalMux I__20399 (
            .O(N__85828),
            .I(N__85766));
    InMux I__20398 (
            .O(N__85827),
            .I(N__85761));
    InMux I__20397 (
            .O(N__85826),
            .I(N__85761));
    InMux I__20396 (
            .O(N__85825),
            .I(N__85758));
    InMux I__20395 (
            .O(N__85824),
            .I(N__85755));
    InMux I__20394 (
            .O(N__85823),
            .I(N__85749));
    InMux I__20393 (
            .O(N__85822),
            .I(N__85749));
    InMux I__20392 (
            .O(N__85821),
            .I(N__85745));
    CascadeMux I__20391 (
            .O(N__85820),
            .I(N__85742));
    CascadeMux I__20390 (
            .O(N__85819),
            .I(N__85739));
    InMux I__20389 (
            .O(N__85818),
            .I(N__85736));
    InMux I__20388 (
            .O(N__85817),
            .I(N__85729));
    InMux I__20387 (
            .O(N__85816),
            .I(N__85729));
    InMux I__20386 (
            .O(N__85815),
            .I(N__85724));
    InMux I__20385 (
            .O(N__85814),
            .I(N__85724));
    InMux I__20384 (
            .O(N__85813),
            .I(N__85718));
    InMux I__20383 (
            .O(N__85812),
            .I(N__85711));
    InMux I__20382 (
            .O(N__85811),
            .I(N__85711));
    InMux I__20381 (
            .O(N__85810),
            .I(N__85711));
    InMux I__20380 (
            .O(N__85809),
            .I(N__85708));
    InMux I__20379 (
            .O(N__85808),
            .I(N__85705));
    InMux I__20378 (
            .O(N__85807),
            .I(N__85696));
    InMux I__20377 (
            .O(N__85806),
            .I(N__85696));
    InMux I__20376 (
            .O(N__85805),
            .I(N__85696));
    InMux I__20375 (
            .O(N__85804),
            .I(N__85696));
    LocalMux I__20374 (
            .O(N__85797),
            .I(N__85693));
    LocalMux I__20373 (
            .O(N__85788),
            .I(N__85688));
    LocalMux I__20372 (
            .O(N__85785),
            .I(N__85688));
    LocalMux I__20371 (
            .O(N__85778),
            .I(N__85679));
    LocalMux I__20370 (
            .O(N__85775),
            .I(N__85679));
    Span4Mux_v I__20369 (
            .O(N__85766),
            .I(N__85679));
    LocalMux I__20368 (
            .O(N__85761),
            .I(N__85679));
    LocalMux I__20367 (
            .O(N__85758),
            .I(N__85676));
    LocalMux I__20366 (
            .O(N__85755),
            .I(N__85673));
    InMux I__20365 (
            .O(N__85754),
            .I(N__85670));
    LocalMux I__20364 (
            .O(N__85749),
            .I(N__85667));
    InMux I__20363 (
            .O(N__85748),
            .I(N__85664));
    LocalMux I__20362 (
            .O(N__85745),
            .I(N__85649));
    InMux I__20361 (
            .O(N__85742),
            .I(N__85644));
    InMux I__20360 (
            .O(N__85739),
            .I(N__85644));
    LocalMux I__20359 (
            .O(N__85736),
            .I(N__85641));
    InMux I__20358 (
            .O(N__85735),
            .I(N__85636));
    InMux I__20357 (
            .O(N__85734),
            .I(N__85636));
    LocalMux I__20356 (
            .O(N__85729),
            .I(N__85618));
    LocalMux I__20355 (
            .O(N__85724),
            .I(N__85615));
    InMux I__20354 (
            .O(N__85723),
            .I(N__85610));
    InMux I__20353 (
            .O(N__85722),
            .I(N__85610));
    InMux I__20352 (
            .O(N__85721),
            .I(N__85607));
    LocalMux I__20351 (
            .O(N__85718),
            .I(N__85600));
    LocalMux I__20350 (
            .O(N__85711),
            .I(N__85600));
    LocalMux I__20349 (
            .O(N__85708),
            .I(N__85600));
    LocalMux I__20348 (
            .O(N__85705),
            .I(N__85597));
    LocalMux I__20347 (
            .O(N__85696),
            .I(N__85594));
    Span4Mux_v I__20346 (
            .O(N__85693),
            .I(N__85577));
    Span4Mux_v I__20345 (
            .O(N__85688),
            .I(N__85577));
    Span4Mux_h I__20344 (
            .O(N__85679),
            .I(N__85577));
    Span4Mux_v I__20343 (
            .O(N__85676),
            .I(N__85577));
    Span4Mux_h I__20342 (
            .O(N__85673),
            .I(N__85577));
    LocalMux I__20341 (
            .O(N__85670),
            .I(N__85577));
    Span4Mux_v I__20340 (
            .O(N__85667),
            .I(N__85577));
    LocalMux I__20339 (
            .O(N__85664),
            .I(N__85577));
    InMux I__20338 (
            .O(N__85663),
            .I(N__85572));
    InMux I__20337 (
            .O(N__85662),
            .I(N__85572));
    InMux I__20336 (
            .O(N__85661),
            .I(N__85569));
    InMux I__20335 (
            .O(N__85660),
            .I(N__85560));
    InMux I__20334 (
            .O(N__85659),
            .I(N__85557));
    InMux I__20333 (
            .O(N__85658),
            .I(N__85552));
    InMux I__20332 (
            .O(N__85657),
            .I(N__85552));
    InMux I__20331 (
            .O(N__85656),
            .I(N__85541));
    InMux I__20330 (
            .O(N__85655),
            .I(N__85541));
    InMux I__20329 (
            .O(N__85654),
            .I(N__85541));
    InMux I__20328 (
            .O(N__85653),
            .I(N__85541));
    InMux I__20327 (
            .O(N__85652),
            .I(N__85541));
    Span4Mux_v I__20326 (
            .O(N__85649),
            .I(N__85537));
    LocalMux I__20325 (
            .O(N__85644),
            .I(N__85534));
    Span4Mux_v I__20324 (
            .O(N__85641),
            .I(N__85529));
    LocalMux I__20323 (
            .O(N__85636),
            .I(N__85529));
    InMux I__20322 (
            .O(N__85635),
            .I(N__85524));
    InMux I__20321 (
            .O(N__85634),
            .I(N__85524));
    InMux I__20320 (
            .O(N__85633),
            .I(N__85516));
    InMux I__20319 (
            .O(N__85632),
            .I(N__85516));
    InMux I__20318 (
            .O(N__85631),
            .I(N__85512));
    InMux I__20317 (
            .O(N__85630),
            .I(N__85505));
    InMux I__20316 (
            .O(N__85629),
            .I(N__85505));
    InMux I__20315 (
            .O(N__85628),
            .I(N__85505));
    InMux I__20314 (
            .O(N__85627),
            .I(N__85499));
    InMux I__20313 (
            .O(N__85626),
            .I(N__85496));
    InMux I__20312 (
            .O(N__85625),
            .I(N__85493));
    InMux I__20311 (
            .O(N__85624),
            .I(N__85488));
    InMux I__20310 (
            .O(N__85623),
            .I(N__85488));
    CascadeMux I__20309 (
            .O(N__85622),
            .I(N__85485));
    CascadeMux I__20308 (
            .O(N__85621),
            .I(N__85482));
    Span4Mux_h I__20307 (
            .O(N__85618),
            .I(N__85473));
    Span4Mux_v I__20306 (
            .O(N__85615),
            .I(N__85473));
    LocalMux I__20305 (
            .O(N__85610),
            .I(N__85473));
    LocalMux I__20304 (
            .O(N__85607),
            .I(N__85470));
    Span4Mux_h I__20303 (
            .O(N__85600),
            .I(N__85457));
    Span4Mux_v I__20302 (
            .O(N__85597),
            .I(N__85457));
    Span4Mux_v I__20301 (
            .O(N__85594),
            .I(N__85457));
    Span4Mux_h I__20300 (
            .O(N__85577),
            .I(N__85457));
    LocalMux I__20299 (
            .O(N__85572),
            .I(N__85457));
    LocalMux I__20298 (
            .O(N__85569),
            .I(N__85457));
    CascadeMux I__20297 (
            .O(N__85568),
            .I(N__85453));
    InMux I__20296 (
            .O(N__85567),
            .I(N__85450));
    InMux I__20295 (
            .O(N__85566),
            .I(N__85441));
    InMux I__20294 (
            .O(N__85565),
            .I(N__85441));
    InMux I__20293 (
            .O(N__85564),
            .I(N__85441));
    InMux I__20292 (
            .O(N__85563),
            .I(N__85441));
    LocalMux I__20291 (
            .O(N__85560),
            .I(N__85432));
    LocalMux I__20290 (
            .O(N__85557),
            .I(N__85432));
    LocalMux I__20289 (
            .O(N__85552),
            .I(N__85426));
    LocalMux I__20288 (
            .O(N__85541),
            .I(N__85426));
    InMux I__20287 (
            .O(N__85540),
            .I(N__85423));
    Span4Mux_h I__20286 (
            .O(N__85537),
            .I(N__85414));
    Span4Mux_v I__20285 (
            .O(N__85534),
            .I(N__85414));
    Span4Mux_v I__20284 (
            .O(N__85529),
            .I(N__85414));
    LocalMux I__20283 (
            .O(N__85524),
            .I(N__85414));
    InMux I__20282 (
            .O(N__85523),
            .I(N__85407));
    InMux I__20281 (
            .O(N__85522),
            .I(N__85407));
    InMux I__20280 (
            .O(N__85521),
            .I(N__85407));
    LocalMux I__20279 (
            .O(N__85516),
            .I(N__85403));
    InMux I__20278 (
            .O(N__85515),
            .I(N__85400));
    LocalMux I__20277 (
            .O(N__85512),
            .I(N__85395));
    LocalMux I__20276 (
            .O(N__85505),
            .I(N__85395));
    InMux I__20275 (
            .O(N__85504),
            .I(N__85392));
    InMux I__20274 (
            .O(N__85503),
            .I(N__85382));
    InMux I__20273 (
            .O(N__85502),
            .I(N__85382));
    LocalMux I__20272 (
            .O(N__85499),
            .I(N__85378));
    LocalMux I__20271 (
            .O(N__85496),
            .I(N__85375));
    LocalMux I__20270 (
            .O(N__85493),
            .I(N__85370));
    LocalMux I__20269 (
            .O(N__85488),
            .I(N__85370));
    InMux I__20268 (
            .O(N__85485),
            .I(N__85365));
    InMux I__20267 (
            .O(N__85482),
            .I(N__85365));
    InMux I__20266 (
            .O(N__85481),
            .I(N__85360));
    InMux I__20265 (
            .O(N__85480),
            .I(N__85360));
    Span4Mux_h I__20264 (
            .O(N__85473),
            .I(N__85353));
    Span4Mux_h I__20263 (
            .O(N__85470),
            .I(N__85353));
    Span4Mux_v I__20262 (
            .O(N__85457),
            .I(N__85353));
    InMux I__20261 (
            .O(N__85456),
            .I(N__85349));
    InMux I__20260 (
            .O(N__85453),
            .I(N__85345));
    LocalMux I__20259 (
            .O(N__85450),
            .I(N__85338));
    LocalMux I__20258 (
            .O(N__85441),
            .I(N__85338));
    InMux I__20257 (
            .O(N__85440),
            .I(N__85335));
    InMux I__20256 (
            .O(N__85439),
            .I(N__85330));
    InMux I__20255 (
            .O(N__85438),
            .I(N__85330));
    CascadeMux I__20254 (
            .O(N__85437),
            .I(N__85326));
    Span4Mux_v I__20253 (
            .O(N__85432),
            .I(N__85319));
    InMux I__20252 (
            .O(N__85431),
            .I(N__85316));
    Span4Mux_v I__20251 (
            .O(N__85426),
            .I(N__85311));
    LocalMux I__20250 (
            .O(N__85423),
            .I(N__85311));
    Span4Mux_h I__20249 (
            .O(N__85414),
            .I(N__85306));
    LocalMux I__20248 (
            .O(N__85407),
            .I(N__85306));
    InMux I__20247 (
            .O(N__85406),
            .I(N__85303));
    Span4Mux_v I__20246 (
            .O(N__85403),
            .I(N__85297));
    LocalMux I__20245 (
            .O(N__85400),
            .I(N__85297));
    Span4Mux_v I__20244 (
            .O(N__85395),
            .I(N__85292));
    LocalMux I__20243 (
            .O(N__85392),
            .I(N__85292));
    InMux I__20242 (
            .O(N__85391),
            .I(N__85287));
    InMux I__20241 (
            .O(N__85390),
            .I(N__85287));
    InMux I__20240 (
            .O(N__85389),
            .I(N__85284));
    InMux I__20239 (
            .O(N__85388),
            .I(N__85281));
    InMux I__20238 (
            .O(N__85387),
            .I(N__85276));
    LocalMux I__20237 (
            .O(N__85382),
            .I(N__85273));
    CascadeMux I__20236 (
            .O(N__85381),
            .I(N__85270));
    Span4Mux_v I__20235 (
            .O(N__85378),
            .I(N__85266));
    Span4Mux_v I__20234 (
            .O(N__85375),
            .I(N__85263));
    Span4Mux_v I__20233 (
            .O(N__85370),
            .I(N__85254));
    LocalMux I__20232 (
            .O(N__85365),
            .I(N__85254));
    LocalMux I__20231 (
            .O(N__85360),
            .I(N__85254));
    Span4Mux_v I__20230 (
            .O(N__85353),
            .I(N__85251));
    InMux I__20229 (
            .O(N__85352),
            .I(N__85248));
    LocalMux I__20228 (
            .O(N__85349),
            .I(N__85245));
    InMux I__20227 (
            .O(N__85348),
            .I(N__85242));
    LocalMux I__20226 (
            .O(N__85345),
            .I(N__85238));
    InMux I__20225 (
            .O(N__85344),
            .I(N__85235));
    InMux I__20224 (
            .O(N__85343),
            .I(N__85232));
    Span4Mux_v I__20223 (
            .O(N__85338),
            .I(N__85219));
    LocalMux I__20222 (
            .O(N__85335),
            .I(N__85219));
    LocalMux I__20221 (
            .O(N__85330),
            .I(N__85219));
    InMux I__20220 (
            .O(N__85329),
            .I(N__85214));
    InMux I__20219 (
            .O(N__85326),
            .I(N__85214));
    InMux I__20218 (
            .O(N__85325),
            .I(N__85211));
    InMux I__20217 (
            .O(N__85324),
            .I(N__85206));
    InMux I__20216 (
            .O(N__85323),
            .I(N__85206));
    InMux I__20215 (
            .O(N__85322),
            .I(N__85203));
    Span4Mux_h I__20214 (
            .O(N__85319),
            .I(N__85196));
    LocalMux I__20213 (
            .O(N__85316),
            .I(N__85196));
    Span4Mux_v I__20212 (
            .O(N__85311),
            .I(N__85189));
    Span4Mux_h I__20211 (
            .O(N__85306),
            .I(N__85189));
    LocalMux I__20210 (
            .O(N__85303),
            .I(N__85189));
    CascadeMux I__20209 (
            .O(N__85302),
            .I(N__85186));
    Span4Mux_v I__20208 (
            .O(N__85297),
            .I(N__85181));
    Span4Mux_v I__20207 (
            .O(N__85292),
            .I(N__85181));
    LocalMux I__20206 (
            .O(N__85287),
            .I(N__85174));
    LocalMux I__20205 (
            .O(N__85284),
            .I(N__85174));
    LocalMux I__20204 (
            .O(N__85281),
            .I(N__85174));
    InMux I__20203 (
            .O(N__85280),
            .I(N__85171));
    InMux I__20202 (
            .O(N__85279),
            .I(N__85161));
    LocalMux I__20201 (
            .O(N__85276),
            .I(N__85156));
    Span4Mux_v I__20200 (
            .O(N__85273),
            .I(N__85156));
    InMux I__20199 (
            .O(N__85270),
            .I(N__85151));
    InMux I__20198 (
            .O(N__85269),
            .I(N__85151));
    Span4Mux_v I__20197 (
            .O(N__85266),
            .I(N__85146));
    Span4Mux_v I__20196 (
            .O(N__85263),
            .I(N__85146));
    InMux I__20195 (
            .O(N__85262),
            .I(N__85141));
    InMux I__20194 (
            .O(N__85261),
            .I(N__85141));
    Span4Mux_h I__20193 (
            .O(N__85254),
            .I(N__85134));
    Span4Mux_h I__20192 (
            .O(N__85251),
            .I(N__85134));
    LocalMux I__20191 (
            .O(N__85248),
            .I(N__85134));
    Span4Mux_v I__20190 (
            .O(N__85245),
            .I(N__85129));
    LocalMux I__20189 (
            .O(N__85242),
            .I(N__85129));
    InMux I__20188 (
            .O(N__85241),
            .I(N__85126));
    Span4Mux_v I__20187 (
            .O(N__85238),
            .I(N__85119));
    LocalMux I__20186 (
            .O(N__85235),
            .I(N__85119));
    LocalMux I__20185 (
            .O(N__85232),
            .I(N__85119));
    InMux I__20184 (
            .O(N__85231),
            .I(N__85116));
    InMux I__20183 (
            .O(N__85230),
            .I(N__85111));
    InMux I__20182 (
            .O(N__85229),
            .I(N__85111));
    InMux I__20181 (
            .O(N__85228),
            .I(N__85103));
    InMux I__20180 (
            .O(N__85227),
            .I(N__85103));
    InMux I__20179 (
            .O(N__85226),
            .I(N__85103));
    Span4Mux_v I__20178 (
            .O(N__85219),
            .I(N__85090));
    LocalMux I__20177 (
            .O(N__85214),
            .I(N__85090));
    LocalMux I__20176 (
            .O(N__85211),
            .I(N__85090));
    LocalMux I__20175 (
            .O(N__85206),
            .I(N__85090));
    LocalMux I__20174 (
            .O(N__85203),
            .I(N__85090));
    InMux I__20173 (
            .O(N__85202),
            .I(N__85085));
    InMux I__20172 (
            .O(N__85201),
            .I(N__85085));
    Span4Mux_v I__20171 (
            .O(N__85196),
            .I(N__85082));
    Span4Mux_h I__20170 (
            .O(N__85189),
            .I(N__85079));
    InMux I__20169 (
            .O(N__85186),
            .I(N__85076));
    Span4Mux_h I__20168 (
            .O(N__85181),
            .I(N__85068));
    Span4Mux_v I__20167 (
            .O(N__85174),
            .I(N__85068));
    LocalMux I__20166 (
            .O(N__85171),
            .I(N__85068));
    InMux I__20165 (
            .O(N__85170),
            .I(N__85065));
    InMux I__20164 (
            .O(N__85169),
            .I(N__85056));
    InMux I__20163 (
            .O(N__85168),
            .I(N__85056));
    InMux I__20162 (
            .O(N__85167),
            .I(N__85056));
    InMux I__20161 (
            .O(N__85166),
            .I(N__85056));
    CascadeMux I__20160 (
            .O(N__85165),
            .I(N__85053));
    CascadeMux I__20159 (
            .O(N__85164),
            .I(N__85047));
    LocalMux I__20158 (
            .O(N__85161),
            .I(N__85044));
    Sp12to4 I__20157 (
            .O(N__85156),
            .I(N__85035));
    LocalMux I__20156 (
            .O(N__85151),
            .I(N__85035));
    Sp12to4 I__20155 (
            .O(N__85146),
            .I(N__85035));
    LocalMux I__20154 (
            .O(N__85141),
            .I(N__85035));
    Span4Mux_h I__20153 (
            .O(N__85134),
            .I(N__85032));
    Span4Mux_v I__20152 (
            .O(N__85129),
            .I(N__85027));
    LocalMux I__20151 (
            .O(N__85126),
            .I(N__85027));
    Span4Mux_v I__20150 (
            .O(N__85119),
            .I(N__85022));
    LocalMux I__20149 (
            .O(N__85116),
            .I(N__85022));
    LocalMux I__20148 (
            .O(N__85111),
            .I(N__85019));
    InMux I__20147 (
            .O(N__85110),
            .I(N__85016));
    LocalMux I__20146 (
            .O(N__85103),
            .I(N__85013));
    InMux I__20145 (
            .O(N__85102),
            .I(N__85010));
    InMux I__20144 (
            .O(N__85101),
            .I(N__85007));
    Span4Mux_v I__20143 (
            .O(N__85090),
            .I(N__85002));
    LocalMux I__20142 (
            .O(N__85085),
            .I(N__84999));
    Span4Mux_v I__20141 (
            .O(N__85082),
            .I(N__84996));
    Span4Mux_v I__20140 (
            .O(N__85079),
            .I(N__84991));
    LocalMux I__20139 (
            .O(N__85076),
            .I(N__84991));
    InMux I__20138 (
            .O(N__85075),
            .I(N__84988));
    Span4Mux_v I__20137 (
            .O(N__85068),
            .I(N__84981));
    LocalMux I__20136 (
            .O(N__85065),
            .I(N__84981));
    LocalMux I__20135 (
            .O(N__85056),
            .I(N__84981));
    InMux I__20134 (
            .O(N__85053),
            .I(N__84976));
    InMux I__20133 (
            .O(N__85052),
            .I(N__84976));
    InMux I__20132 (
            .O(N__85051),
            .I(N__84973));
    InMux I__20131 (
            .O(N__85050),
            .I(N__84968));
    InMux I__20130 (
            .O(N__85047),
            .I(N__84968));
    Span12Mux_v I__20129 (
            .O(N__85044),
            .I(N__84962));
    Span12Mux_h I__20128 (
            .O(N__85035),
            .I(N__84959));
    Span4Mux_v I__20127 (
            .O(N__85032),
            .I(N__84956));
    Span4Mux_v I__20126 (
            .O(N__85027),
            .I(N__84941));
    Span4Mux_h I__20125 (
            .O(N__85022),
            .I(N__84941));
    Span4Mux_h I__20124 (
            .O(N__85019),
            .I(N__84941));
    LocalMux I__20123 (
            .O(N__85016),
            .I(N__84941));
    Span4Mux_v I__20122 (
            .O(N__85013),
            .I(N__84941));
    LocalMux I__20121 (
            .O(N__85010),
            .I(N__84941));
    LocalMux I__20120 (
            .O(N__85007),
            .I(N__84941));
    InMux I__20119 (
            .O(N__85006),
            .I(N__84938));
    CascadeMux I__20118 (
            .O(N__85005),
            .I(N__84935));
    Span4Mux_v I__20117 (
            .O(N__85002),
            .I(N__84929));
    Span4Mux_v I__20116 (
            .O(N__84999),
            .I(N__84929));
    Span4Mux_v I__20115 (
            .O(N__84996),
            .I(N__84924));
    Span4Mux_h I__20114 (
            .O(N__84991),
            .I(N__84924));
    LocalMux I__20113 (
            .O(N__84988),
            .I(N__84921));
    Span4Mux_v I__20112 (
            .O(N__84981),
            .I(N__84912));
    LocalMux I__20111 (
            .O(N__84976),
            .I(N__84912));
    LocalMux I__20110 (
            .O(N__84973),
            .I(N__84912));
    LocalMux I__20109 (
            .O(N__84968),
            .I(N__84912));
    InMux I__20108 (
            .O(N__84967),
            .I(N__84909));
    CascadeMux I__20107 (
            .O(N__84966),
            .I(N__84905));
    CascadeMux I__20106 (
            .O(N__84965),
            .I(N__84902));
    Span12Mux_v I__20105 (
            .O(N__84962),
            .I(N__84899));
    Span12Mux_v I__20104 (
            .O(N__84959),
            .I(N__84896));
    Span4Mux_h I__20103 (
            .O(N__84956),
            .I(N__84889));
    Span4Mux_h I__20102 (
            .O(N__84941),
            .I(N__84889));
    LocalMux I__20101 (
            .O(N__84938),
            .I(N__84889));
    InMux I__20100 (
            .O(N__84935),
            .I(N__84886));
    InMux I__20099 (
            .O(N__84934),
            .I(N__84883));
    Span4Mux_h I__20098 (
            .O(N__84929),
            .I(N__84872));
    Span4Mux_v I__20097 (
            .O(N__84924),
            .I(N__84872));
    Span4Mux_v I__20096 (
            .O(N__84921),
            .I(N__84872));
    Span4Mux_v I__20095 (
            .O(N__84912),
            .I(N__84872));
    LocalMux I__20094 (
            .O(N__84909),
            .I(N__84872));
    InMux I__20093 (
            .O(N__84908),
            .I(N__84867));
    InMux I__20092 (
            .O(N__84905),
            .I(N__84867));
    InMux I__20091 (
            .O(N__84902),
            .I(N__84864));
    Odrv12 I__20090 (
            .O(N__84899),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2 ));
    Odrv12 I__20089 (
            .O(N__84896),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2 ));
    Odrv4 I__20088 (
            .O(N__84889),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2 ));
    LocalMux I__20087 (
            .O(N__84886),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2 ));
    LocalMux I__20086 (
            .O(N__84883),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2 ));
    Odrv4 I__20085 (
            .O(N__84872),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2 ));
    LocalMux I__20084 (
            .O(N__84867),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2 ));
    LocalMux I__20083 (
            .O(N__84864),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2 ));
    CascadeMux I__20082 (
            .O(N__84847),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11811_cascade_ ));
    InMux I__20081 (
            .O(N__84844),
            .I(N__84841));
    LocalMux I__20080 (
            .O(N__84841),
            .I(N__84838));
    Span4Mux_v I__20079 (
            .O(N__84838),
            .I(N__84834));
    InMux I__20078 (
            .O(N__84837),
            .I(N__84831));
    Sp12to4 I__20077 (
            .O(N__84834),
            .I(N__84828));
    LocalMux I__20076 (
            .O(N__84831),
            .I(N__84825));
    Odrv12 I__20075 (
            .O(N__84828),
            .I(REG_mem_47_8));
    Odrv4 I__20074 (
            .O(N__84825),
            .I(REG_mem_47_8));
    InMux I__20073 (
            .O(N__84820),
            .I(\timing_controller_inst.n10606 ));
    InMux I__20072 (
            .O(N__84817),
            .I(N__84814));
    LocalMux I__20071 (
            .O(N__84814),
            .I(N__84810));
    InMux I__20070 (
            .O(N__84813),
            .I(N__84807));
    Span4Mux_h I__20069 (
            .O(N__84810),
            .I(N__84804));
    LocalMux I__20068 (
            .O(N__84807),
            .I(N__84801));
    Odrv4 I__20067 (
            .O(N__84804),
            .I(\timing_controller_inst.state_timeout_counter_20 ));
    Odrv12 I__20066 (
            .O(N__84801),
            .I(\timing_controller_inst.state_timeout_counter_20 ));
    InMux I__20065 (
            .O(N__84796),
            .I(N__84793));
    LocalMux I__20064 (
            .O(N__84793),
            .I(N__84790));
    Span4Mux_v I__20063 (
            .O(N__84790),
            .I(N__84787));
    Span4Mux_h I__20062 (
            .O(N__84787),
            .I(N__84784));
    Odrv4 I__20061 (
            .O(N__84784),
            .I(\timing_controller_inst.n12542 ));
    InMux I__20060 (
            .O(N__84781),
            .I(\timing_controller_inst.n10607 ));
    InMux I__20059 (
            .O(N__84778),
            .I(N__84775));
    LocalMux I__20058 (
            .O(N__84775),
            .I(N__84771));
    InMux I__20057 (
            .O(N__84774),
            .I(N__84768));
    Odrv4 I__20056 (
            .O(N__84771),
            .I(\timing_controller_inst.state_timeout_counter_21 ));
    LocalMux I__20055 (
            .O(N__84768),
            .I(\timing_controller_inst.state_timeout_counter_21 ));
    InMux I__20054 (
            .O(N__84763),
            .I(\timing_controller_inst.n10608 ));
    InMux I__20053 (
            .O(N__84760),
            .I(N__84756));
    InMux I__20052 (
            .O(N__84759),
            .I(N__84753));
    LocalMux I__20051 (
            .O(N__84756),
            .I(\timing_controller_inst.state_timeout_counter_22 ));
    LocalMux I__20050 (
            .O(N__84753),
            .I(\timing_controller_inst.state_timeout_counter_22 ));
    InMux I__20049 (
            .O(N__84748),
            .I(N__84745));
    LocalMux I__20048 (
            .O(N__84745),
            .I(\timing_controller_inst.n12541 ));
    InMux I__20047 (
            .O(N__84742),
            .I(\timing_controller_inst.n10609 ));
    InMux I__20046 (
            .O(N__84739),
            .I(N__84736));
    LocalMux I__20045 (
            .O(N__84736),
            .I(N__84733));
    Span4Mux_v I__20044 (
            .O(N__84733),
            .I(N__84729));
    InMux I__20043 (
            .O(N__84732),
            .I(N__84726));
    Odrv4 I__20042 (
            .O(N__84729),
            .I(\timing_controller_inst.state_timeout_counter_23 ));
    LocalMux I__20041 (
            .O(N__84726),
            .I(\timing_controller_inst.state_timeout_counter_23 ));
    InMux I__20040 (
            .O(N__84721),
            .I(N__84718));
    LocalMux I__20039 (
            .O(N__84718),
            .I(\timing_controller_inst.n12540 ));
    InMux I__20038 (
            .O(N__84715),
            .I(\timing_controller_inst.n10610 ));
    InMux I__20037 (
            .O(N__84712),
            .I(N__84709));
    LocalMux I__20036 (
            .O(N__84709),
            .I(N__84706));
    Span4Mux_v I__20035 (
            .O(N__84706),
            .I(N__84702));
    InMux I__20034 (
            .O(N__84705),
            .I(N__84699));
    Span4Mux_h I__20033 (
            .O(N__84702),
            .I(N__84691));
    LocalMux I__20032 (
            .O(N__84699),
            .I(N__84688));
    InMux I__20031 (
            .O(N__84698),
            .I(N__84683));
    InMux I__20030 (
            .O(N__84697),
            .I(N__84683));
    InMux I__20029 (
            .O(N__84696),
            .I(N__84676));
    InMux I__20028 (
            .O(N__84695),
            .I(N__84676));
    InMux I__20027 (
            .O(N__84694),
            .I(N__84676));
    Span4Mux_h I__20026 (
            .O(N__84691),
            .I(N__84664));
    Span4Mux_v I__20025 (
            .O(N__84688),
            .I(N__84657));
    LocalMux I__20024 (
            .O(N__84683),
            .I(N__84657));
    LocalMux I__20023 (
            .O(N__84676),
            .I(N__84657));
    InMux I__20022 (
            .O(N__84675),
            .I(N__84650));
    InMux I__20021 (
            .O(N__84674),
            .I(N__84650));
    InMux I__20020 (
            .O(N__84673),
            .I(N__84650));
    InMux I__20019 (
            .O(N__84672),
            .I(N__84645));
    InMux I__20018 (
            .O(N__84671),
            .I(N__84645));
    InMux I__20017 (
            .O(N__84670),
            .I(N__84642));
    InMux I__20016 (
            .O(N__84669),
            .I(N__84637));
    InMux I__20015 (
            .O(N__84668),
            .I(N__84637));
    InMux I__20014 (
            .O(N__84667),
            .I(N__84634));
    Odrv4 I__20013 (
            .O(N__84664),
            .I(n1616));
    Odrv4 I__20012 (
            .O(N__84657),
            .I(n1616));
    LocalMux I__20011 (
            .O(N__84650),
            .I(n1616));
    LocalMux I__20010 (
            .O(N__84645),
            .I(n1616));
    LocalMux I__20009 (
            .O(N__84642),
            .I(n1616));
    LocalMux I__20008 (
            .O(N__84637),
            .I(n1616));
    LocalMux I__20007 (
            .O(N__84634),
            .I(n1616));
    InMux I__20006 (
            .O(N__84619),
            .I(N__84615));
    InMux I__20005 (
            .O(N__84618),
            .I(N__84612));
    LocalMux I__20004 (
            .O(N__84615),
            .I(\timing_controller_inst.state_timeout_counter_24 ));
    LocalMux I__20003 (
            .O(N__84612),
            .I(\timing_controller_inst.state_timeout_counter_24 ));
    InMux I__20002 (
            .O(N__84607),
            .I(N__84604));
    LocalMux I__20001 (
            .O(N__84604),
            .I(\timing_controller_inst.n12539 ));
    InMux I__20000 (
            .O(N__84601),
            .I(bfn_23_16_0_));
    InMux I__19999 (
            .O(N__84598),
            .I(N__84594));
    InMux I__19998 (
            .O(N__84597),
            .I(N__84591));
    LocalMux I__19997 (
            .O(N__84594),
            .I(\timing_controller_inst.state_timeout_counter_25 ));
    LocalMux I__19996 (
            .O(N__84591),
            .I(\timing_controller_inst.state_timeout_counter_25 ));
    InMux I__19995 (
            .O(N__84586),
            .I(\timing_controller_inst.n10612 ));
    CascadeMux I__19994 (
            .O(N__84583),
            .I(N__84579));
    InMux I__19993 (
            .O(N__84582),
            .I(N__84576));
    InMux I__19992 (
            .O(N__84579),
            .I(N__84573));
    LocalMux I__19991 (
            .O(N__84576),
            .I(\timing_controller_inst.state_timeout_counter_26 ));
    LocalMux I__19990 (
            .O(N__84573),
            .I(\timing_controller_inst.state_timeout_counter_26 ));
    InMux I__19989 (
            .O(N__84568),
            .I(\timing_controller_inst.n10613 ));
    InMux I__19988 (
            .O(N__84565),
            .I(N__84562));
    LocalMux I__19987 (
            .O(N__84562),
            .I(N__84559));
    Span4Mux_h I__19986 (
            .O(N__84559),
            .I(N__84555));
    InMux I__19985 (
            .O(N__84558),
            .I(N__84552));
    Odrv4 I__19984 (
            .O(N__84555),
            .I(\timing_controller_inst.state_timeout_counter_27 ));
    LocalMux I__19983 (
            .O(N__84552),
            .I(\timing_controller_inst.state_timeout_counter_27 ));
    InMux I__19982 (
            .O(N__84547),
            .I(\timing_controller_inst.n10598 ));
    InMux I__19981 (
            .O(N__84544),
            .I(N__84540));
    InMux I__19980 (
            .O(N__84543),
            .I(N__84537));
    LocalMux I__19979 (
            .O(N__84540),
            .I(N__84532));
    LocalMux I__19978 (
            .O(N__84537),
            .I(N__84532));
    Span4Mux_v I__19977 (
            .O(N__84532),
            .I(N__84529));
    Odrv4 I__19976 (
            .O(N__84529),
            .I(\timing_controller_inst.state_timeout_counter_12 ));
    InMux I__19975 (
            .O(N__84526),
            .I(N__84523));
    LocalMux I__19974 (
            .O(N__84523),
            .I(N__84520));
    Span4Mux_h I__19973 (
            .O(N__84520),
            .I(N__84517));
    Odrv4 I__19972 (
            .O(N__84517),
            .I(\timing_controller_inst.n12549 ));
    InMux I__19971 (
            .O(N__84514),
            .I(\timing_controller_inst.n10599 ));
    CascadeMux I__19970 (
            .O(N__84511),
            .I(N__84508));
    InMux I__19969 (
            .O(N__84508),
            .I(N__84505));
    LocalMux I__19968 (
            .O(N__84505),
            .I(N__84502));
    Span4Mux_v I__19967 (
            .O(N__84502),
            .I(N__84498));
    InMux I__19966 (
            .O(N__84501),
            .I(N__84495));
    Odrv4 I__19965 (
            .O(N__84498),
            .I(\timing_controller_inst.state_timeout_counter_13 ));
    LocalMux I__19964 (
            .O(N__84495),
            .I(\timing_controller_inst.state_timeout_counter_13 ));
    InMux I__19963 (
            .O(N__84490),
            .I(\timing_controller_inst.n10600 ));
    InMux I__19962 (
            .O(N__84487),
            .I(N__84484));
    LocalMux I__19961 (
            .O(N__84484),
            .I(N__84481));
    Span4Mux_v I__19960 (
            .O(N__84481),
            .I(N__84477));
    InMux I__19959 (
            .O(N__84480),
            .I(N__84474));
    Odrv4 I__19958 (
            .O(N__84477),
            .I(\timing_controller_inst.state_timeout_counter_14 ));
    LocalMux I__19957 (
            .O(N__84474),
            .I(\timing_controller_inst.state_timeout_counter_14 ));
    InMux I__19956 (
            .O(N__84469),
            .I(N__84466));
    LocalMux I__19955 (
            .O(N__84466),
            .I(N__84463));
    Span4Mux_v I__19954 (
            .O(N__84463),
            .I(N__84460));
    Odrv4 I__19953 (
            .O(N__84460),
            .I(\timing_controller_inst.n12548 ));
    InMux I__19952 (
            .O(N__84457),
            .I(\timing_controller_inst.n10601 ));
    InMux I__19951 (
            .O(N__84454),
            .I(N__84450));
    CascadeMux I__19950 (
            .O(N__84453),
            .I(N__84447));
    LocalMux I__19949 (
            .O(N__84450),
            .I(N__84444));
    InMux I__19948 (
            .O(N__84447),
            .I(N__84441));
    Span4Mux_v I__19947 (
            .O(N__84444),
            .I(N__84438));
    LocalMux I__19946 (
            .O(N__84441),
            .I(N__84435));
    Odrv4 I__19945 (
            .O(N__84438),
            .I(\timing_controller_inst.state_timeout_counter_15 ));
    Odrv12 I__19944 (
            .O(N__84435),
            .I(\timing_controller_inst.state_timeout_counter_15 ));
    InMux I__19943 (
            .O(N__84430),
            .I(N__84427));
    LocalMux I__19942 (
            .O(N__84427),
            .I(N__84424));
    Span4Mux_v I__19941 (
            .O(N__84424),
            .I(N__84421));
    Odrv4 I__19940 (
            .O(N__84421),
            .I(\timing_controller_inst.n12547 ));
    InMux I__19939 (
            .O(N__84418),
            .I(\timing_controller_inst.n10602 ));
    CascadeMux I__19938 (
            .O(N__84415),
            .I(N__84412));
    InMux I__19937 (
            .O(N__84412),
            .I(N__84409));
    LocalMux I__19936 (
            .O(N__84409),
            .I(N__84406));
    Span4Mux_v I__19935 (
            .O(N__84406),
            .I(N__84402));
    InMux I__19934 (
            .O(N__84405),
            .I(N__84399));
    Odrv4 I__19933 (
            .O(N__84402),
            .I(\timing_controller_inst.state_timeout_counter_16 ));
    LocalMux I__19932 (
            .O(N__84399),
            .I(\timing_controller_inst.state_timeout_counter_16 ));
    InMux I__19931 (
            .O(N__84394),
            .I(bfn_23_15_0_));
    InMux I__19930 (
            .O(N__84391),
            .I(N__84387));
    InMux I__19929 (
            .O(N__84390),
            .I(N__84384));
    LocalMux I__19928 (
            .O(N__84387),
            .I(\timing_controller_inst.state_timeout_counter_17 ));
    LocalMux I__19927 (
            .O(N__84384),
            .I(\timing_controller_inst.state_timeout_counter_17 ));
    InMux I__19926 (
            .O(N__84379),
            .I(\timing_controller_inst.n10604 ));
    InMux I__19925 (
            .O(N__84376),
            .I(N__84373));
    LocalMux I__19924 (
            .O(N__84373),
            .I(N__84369));
    InMux I__19923 (
            .O(N__84372),
            .I(N__84366));
    Span4Mux_v I__19922 (
            .O(N__84369),
            .I(N__84363));
    LocalMux I__19921 (
            .O(N__84366),
            .I(N__84360));
    Odrv4 I__19920 (
            .O(N__84363),
            .I(\timing_controller_inst.state_timeout_counter_18 ));
    Odrv4 I__19919 (
            .O(N__84360),
            .I(\timing_controller_inst.state_timeout_counter_18 ));
    InMux I__19918 (
            .O(N__84355),
            .I(N__84352));
    LocalMux I__19917 (
            .O(N__84352),
            .I(N__84349));
    Span4Mux_v I__19916 (
            .O(N__84349),
            .I(N__84346));
    Odrv4 I__19915 (
            .O(N__84346),
            .I(\timing_controller_inst.n12545 ));
    InMux I__19914 (
            .O(N__84343),
            .I(\timing_controller_inst.n10605 ));
    CascadeMux I__19913 (
            .O(N__84340),
            .I(N__84336));
    CascadeMux I__19912 (
            .O(N__84339),
            .I(N__84333));
    InMux I__19911 (
            .O(N__84336),
            .I(N__84330));
    InMux I__19910 (
            .O(N__84333),
            .I(N__84327));
    LocalMux I__19909 (
            .O(N__84330),
            .I(N__84322));
    LocalMux I__19908 (
            .O(N__84327),
            .I(N__84322));
    Span4Mux_v I__19907 (
            .O(N__84322),
            .I(N__84319));
    Odrv4 I__19906 (
            .O(N__84319),
            .I(\timing_controller_inst.state_timeout_counter_19 ));
    InMux I__19905 (
            .O(N__84316),
            .I(N__84313));
    LocalMux I__19904 (
            .O(N__84313),
            .I(N__84310));
    Span12Mux_h I__19903 (
            .O(N__84310),
            .I(N__84307));
    Odrv12 I__19902 (
            .O(N__84307),
            .I(\timing_controller_inst.n12544 ));
    InMux I__19901 (
            .O(N__84304),
            .I(\timing_controller_inst.n10590 ));
    InMux I__19900 (
            .O(N__84301),
            .I(N__84298));
    LocalMux I__19899 (
            .O(N__84298),
            .I(N__84294));
    InMux I__19898 (
            .O(N__84297),
            .I(N__84291));
    Odrv4 I__19897 (
            .O(N__84294),
            .I(\timing_controller_inst.state_timeout_counter_4 ));
    LocalMux I__19896 (
            .O(N__84291),
            .I(\timing_controller_inst.state_timeout_counter_4 ));
    InMux I__19895 (
            .O(N__84286),
            .I(N__84283));
    LocalMux I__19894 (
            .O(N__84283),
            .I(N__84280));
    Odrv4 I__19893 (
            .O(N__84280),
            .I(\timing_controller_inst.n12604 ));
    InMux I__19892 (
            .O(N__84277),
            .I(\timing_controller_inst.n10591 ));
    InMux I__19891 (
            .O(N__84274),
            .I(N__84271));
    LocalMux I__19890 (
            .O(N__84271),
            .I(\timing_controller_inst.n11347 ));
    CascadeMux I__19889 (
            .O(N__84268),
            .I(N__84265));
    InMux I__19888 (
            .O(N__84265),
            .I(N__84261));
    InMux I__19887 (
            .O(N__84264),
            .I(N__84258));
    LocalMux I__19886 (
            .O(N__84261),
            .I(\timing_controller_inst.state_timeout_counter_5 ));
    LocalMux I__19885 (
            .O(N__84258),
            .I(\timing_controller_inst.state_timeout_counter_5 ));
    InMux I__19884 (
            .O(N__84253),
            .I(N__84250));
    LocalMux I__19883 (
            .O(N__84250),
            .I(\timing_controller_inst.n12555 ));
    InMux I__19882 (
            .O(N__84247),
            .I(\timing_controller_inst.n10592 ));
    InMux I__19881 (
            .O(N__84244),
            .I(N__84240));
    InMux I__19880 (
            .O(N__84243),
            .I(N__84237));
    LocalMux I__19879 (
            .O(N__84240),
            .I(\timing_controller_inst.state_timeout_counter_6 ));
    LocalMux I__19878 (
            .O(N__84237),
            .I(\timing_controller_inst.state_timeout_counter_6 ));
    InMux I__19877 (
            .O(N__84232),
            .I(\timing_controller_inst.n10593 ));
    InMux I__19876 (
            .O(N__84229),
            .I(N__84225));
    CascadeMux I__19875 (
            .O(N__84228),
            .I(N__84222));
    LocalMux I__19874 (
            .O(N__84225),
            .I(N__84219));
    InMux I__19873 (
            .O(N__84222),
            .I(N__84216));
    Odrv12 I__19872 (
            .O(N__84219),
            .I(\timing_controller_inst.state_timeout_counter_7 ));
    LocalMux I__19871 (
            .O(N__84216),
            .I(\timing_controller_inst.state_timeout_counter_7 ));
    InMux I__19870 (
            .O(N__84211),
            .I(\timing_controller_inst.n10594 ));
    InMux I__19869 (
            .O(N__84208),
            .I(N__84205));
    LocalMux I__19868 (
            .O(N__84205),
            .I(N__84201));
    InMux I__19867 (
            .O(N__84204),
            .I(N__84198));
    Odrv4 I__19866 (
            .O(N__84201),
            .I(\timing_controller_inst.state_timeout_counter_8 ));
    LocalMux I__19865 (
            .O(N__84198),
            .I(\timing_controller_inst.state_timeout_counter_8 ));
    InMux I__19864 (
            .O(N__84193),
            .I(bfn_23_14_0_));
    InMux I__19863 (
            .O(N__84190),
            .I(N__84186));
    InMux I__19862 (
            .O(N__84189),
            .I(N__84183));
    LocalMux I__19861 (
            .O(N__84186),
            .I(\timing_controller_inst.state_timeout_counter_9 ));
    LocalMux I__19860 (
            .O(N__84183),
            .I(\timing_controller_inst.state_timeout_counter_9 ));
    InMux I__19859 (
            .O(N__84178),
            .I(N__84175));
    LocalMux I__19858 (
            .O(N__84175),
            .I(\timing_controller_inst.n12551 ));
    InMux I__19857 (
            .O(N__84172),
            .I(\timing_controller_inst.n10596 ));
    InMux I__19856 (
            .O(N__84169),
            .I(N__84165));
    InMux I__19855 (
            .O(N__84168),
            .I(N__84162));
    LocalMux I__19854 (
            .O(N__84165),
            .I(N__84159));
    LocalMux I__19853 (
            .O(N__84162),
            .I(\timing_controller_inst.state_timeout_counter_10 ));
    Odrv4 I__19852 (
            .O(N__84159),
            .I(\timing_controller_inst.state_timeout_counter_10 ));
    InMux I__19851 (
            .O(N__84154),
            .I(N__84151));
    LocalMux I__19850 (
            .O(N__84151),
            .I(\timing_controller_inst.n12550 ));
    InMux I__19849 (
            .O(N__84148),
            .I(\timing_controller_inst.n10597 ));
    InMux I__19848 (
            .O(N__84145),
            .I(N__84142));
    LocalMux I__19847 (
            .O(N__84142),
            .I(N__84138));
    InMux I__19846 (
            .O(N__84141),
            .I(N__84135));
    Odrv4 I__19845 (
            .O(N__84138),
            .I(\timing_controller_inst.state_timeout_counter_11 ));
    LocalMux I__19844 (
            .O(N__84135),
            .I(\timing_controller_inst.state_timeout_counter_11 ));
    InMux I__19843 (
            .O(N__84130),
            .I(N__84127));
    LocalMux I__19842 (
            .O(N__84127),
            .I(\timing_controller_inst.n7592 ));
    InMux I__19841 (
            .O(N__84124),
            .I(N__84121));
    LocalMux I__19840 (
            .O(N__84121),
            .I(N__84118));
    Odrv12 I__19839 (
            .O(N__84118),
            .I(\timing_controller_inst.n7 ));
    InMux I__19838 (
            .O(N__84115),
            .I(N__84102));
    InMux I__19837 (
            .O(N__84114),
            .I(N__84102));
    InMux I__19836 (
            .O(N__84113),
            .I(N__84102));
    InMux I__19835 (
            .O(N__84112),
            .I(N__84102));
    CascadeMux I__19834 (
            .O(N__84111),
            .I(N__84099));
    LocalMux I__19833 (
            .O(N__84102),
            .I(N__84096));
    InMux I__19832 (
            .O(N__84099),
            .I(N__84090));
    Span4Mux_v I__19831 (
            .O(N__84096),
            .I(N__84083));
    InMux I__19830 (
            .O(N__84095),
            .I(N__84076));
    InMux I__19829 (
            .O(N__84094),
            .I(N__84076));
    InMux I__19828 (
            .O(N__84093),
            .I(N__84076));
    LocalMux I__19827 (
            .O(N__84090),
            .I(N__84067));
    InMux I__19826 (
            .O(N__84089),
            .I(N__84058));
    InMux I__19825 (
            .O(N__84088),
            .I(N__84058));
    InMux I__19824 (
            .O(N__84087),
            .I(N__84058));
    InMux I__19823 (
            .O(N__84086),
            .I(N__84058));
    Span4Mux_h I__19822 (
            .O(N__84083),
            .I(N__84053));
    LocalMux I__19821 (
            .O(N__84076),
            .I(N__84053));
    InMux I__19820 (
            .O(N__84075),
            .I(N__84044));
    InMux I__19819 (
            .O(N__84074),
            .I(N__84044));
    InMux I__19818 (
            .O(N__84073),
            .I(N__84044));
    InMux I__19817 (
            .O(N__84072),
            .I(N__84044));
    InMux I__19816 (
            .O(N__84071),
            .I(N__84039));
    InMux I__19815 (
            .O(N__84070),
            .I(N__84039));
    Odrv4 I__19814 (
            .O(N__84067),
            .I(state_3));
    LocalMux I__19813 (
            .O(N__84058),
            .I(state_3));
    Odrv4 I__19812 (
            .O(N__84053),
            .I(state_3));
    LocalMux I__19811 (
            .O(N__84044),
            .I(state_3));
    LocalMux I__19810 (
            .O(N__84039),
            .I(state_3));
    CascadeMux I__19809 (
            .O(N__84028),
            .I(N__84023));
    CascadeMux I__19808 (
            .O(N__84027),
            .I(N__84019));
    InMux I__19807 (
            .O(N__84026),
            .I(N__84005));
    InMux I__19806 (
            .O(N__84023),
            .I(N__84005));
    InMux I__19805 (
            .O(N__84022),
            .I(N__84005));
    InMux I__19804 (
            .O(N__84019),
            .I(N__84005));
    InMux I__19803 (
            .O(N__84018),
            .I(N__84005));
    CascadeMux I__19802 (
            .O(N__84017),
            .I(N__83999));
    CascadeMux I__19801 (
            .O(N__84016),
            .I(N__83992));
    LocalMux I__19800 (
            .O(N__84005),
            .I(N__83988));
    InMux I__19799 (
            .O(N__84004),
            .I(N__83985));
    InMux I__19798 (
            .O(N__84003),
            .I(N__83974));
    InMux I__19797 (
            .O(N__84002),
            .I(N__83974));
    InMux I__19796 (
            .O(N__83999),
            .I(N__83974));
    InMux I__19795 (
            .O(N__83998),
            .I(N__83974));
    InMux I__19794 (
            .O(N__83997),
            .I(N__83974));
    InMux I__19793 (
            .O(N__83996),
            .I(N__83967));
    InMux I__19792 (
            .O(N__83995),
            .I(N__83967));
    InMux I__19791 (
            .O(N__83992),
            .I(N__83967));
    CascadeMux I__19790 (
            .O(N__83991),
            .I(N__83961));
    Span12Mux_v I__19789 (
            .O(N__83988),
            .I(N__83950));
    LocalMux I__19788 (
            .O(N__83985),
            .I(N__83950));
    LocalMux I__19787 (
            .O(N__83974),
            .I(N__83950));
    LocalMux I__19786 (
            .O(N__83967),
            .I(N__83950));
    InMux I__19785 (
            .O(N__83966),
            .I(N__83947));
    InMux I__19784 (
            .O(N__83965),
            .I(N__83938));
    InMux I__19783 (
            .O(N__83964),
            .I(N__83938));
    InMux I__19782 (
            .O(N__83961),
            .I(N__83938));
    InMux I__19781 (
            .O(N__83960),
            .I(N__83938));
    InMux I__19780 (
            .O(N__83959),
            .I(N__83935));
    Odrv12 I__19779 (
            .O(N__83950),
            .I(state_0));
    LocalMux I__19778 (
            .O(N__83947),
            .I(state_0));
    LocalMux I__19777 (
            .O(N__83938),
            .I(state_0));
    LocalMux I__19776 (
            .O(N__83935),
            .I(state_0));
    CEMux I__19775 (
            .O(N__83926),
            .I(N__83923));
    LocalMux I__19774 (
            .O(N__83923),
            .I(N__83920));
    Span4Mux_h I__19773 (
            .O(N__83920),
            .I(N__83917));
    Odrv4 I__19772 (
            .O(N__83917),
            .I(\timing_controller_inst.n11377 ));
    SRMux I__19771 (
            .O(N__83914),
            .I(N__83910));
    InMux I__19770 (
            .O(N__83913),
            .I(N__83901));
    LocalMux I__19769 (
            .O(N__83910),
            .I(N__83898));
    InMux I__19768 (
            .O(N__83909),
            .I(N__83885));
    InMux I__19767 (
            .O(N__83908),
            .I(N__83885));
    InMux I__19766 (
            .O(N__83907),
            .I(N__83885));
    InMux I__19765 (
            .O(N__83906),
            .I(N__83885));
    InMux I__19764 (
            .O(N__83905),
            .I(N__83885));
    InMux I__19763 (
            .O(N__83904),
            .I(N__83885));
    LocalMux I__19762 (
            .O(N__83901),
            .I(r_SM_Main_2));
    Odrv4 I__19761 (
            .O(N__83898),
            .I(r_SM_Main_2));
    LocalMux I__19760 (
            .O(N__83885),
            .I(r_SM_Main_2));
    IoInMux I__19759 (
            .O(N__83878),
            .I(N__83875));
    LocalMux I__19758 (
            .O(N__83875),
            .I(N__83872));
    Span12Mux_s5_h I__19757 (
            .O(N__83872),
            .I(N__83869));
    Span12Mux_v I__19756 (
            .O(N__83869),
            .I(N__83866));
    Odrv12 I__19755 (
            .O(N__83866),
            .I(GB_BUFFER_DEBUG_6_c_c_THRU_CO));
    IoInMux I__19754 (
            .O(N__83863),
            .I(N__83860));
    LocalMux I__19753 (
            .O(N__83860),
            .I(N__83857));
    IoSpan4Mux I__19752 (
            .O(N__83857),
            .I(N__83854));
    Span4Mux_s3_h I__19751 (
            .O(N__83854),
            .I(N__83851));
    Odrv4 I__19750 (
            .O(N__83851),
            .I(GB_BUFFER_SLM_CLK_c_THRU_CO));
    InMux I__19749 (
            .O(N__83848),
            .I(N__83844));
    InMux I__19748 (
            .O(N__83847),
            .I(N__83841));
    LocalMux I__19747 (
            .O(N__83844),
            .I(N__83838));
    LocalMux I__19746 (
            .O(N__83841),
            .I(N__83835));
    Odrv4 I__19745 (
            .O(N__83838),
            .I(\timing_controller_inst.state_timeout_counter_0 ));
    Odrv12 I__19744 (
            .O(N__83835),
            .I(\timing_controller_inst.state_timeout_counter_0 ));
    InMux I__19743 (
            .O(N__83830),
            .I(N__83827));
    LocalMux I__19742 (
            .O(N__83827),
            .I(N__83824));
    Span4Mux_v I__19741 (
            .O(N__83824),
            .I(N__83821));
    Odrv4 I__19740 (
            .O(N__83821),
            .I(\timing_controller_inst.n12532 ));
    InMux I__19739 (
            .O(N__83818),
            .I(bfn_23_13_0_));
    CascadeMux I__19738 (
            .O(N__83815),
            .I(N__83812));
    InMux I__19737 (
            .O(N__83812),
            .I(N__83808));
    CascadeMux I__19736 (
            .O(N__83811),
            .I(N__83805));
    LocalMux I__19735 (
            .O(N__83808),
            .I(N__83802));
    InMux I__19734 (
            .O(N__83805),
            .I(N__83799));
    Odrv12 I__19733 (
            .O(N__83802),
            .I(\timing_controller_inst.state_timeout_counter_1 ));
    LocalMux I__19732 (
            .O(N__83799),
            .I(\timing_controller_inst.state_timeout_counter_1 ));
    InMux I__19731 (
            .O(N__83794),
            .I(N__83791));
    LocalMux I__19730 (
            .O(N__83791),
            .I(\timing_controller_inst.n12554 ));
    InMux I__19729 (
            .O(N__83788),
            .I(\timing_controller_inst.n10588 ));
    InMux I__19728 (
            .O(N__83785),
            .I(N__83779));
    InMux I__19727 (
            .O(N__83784),
            .I(N__83779));
    LocalMux I__19726 (
            .O(N__83779),
            .I(N__83776));
    Span4Mux_v I__19725 (
            .O(N__83776),
            .I(N__83773));
    Sp12to4 I__19724 (
            .O(N__83773),
            .I(N__83770));
    Odrv12 I__19723 (
            .O(N__83770),
            .I(n7383));
    CascadeMux I__19722 (
            .O(N__83767),
            .I(N__83764));
    InMux I__19721 (
            .O(N__83764),
            .I(N__83761));
    LocalMux I__19720 (
            .O(N__83761),
            .I(N__83758));
    Span4Mux_v I__19719 (
            .O(N__83758),
            .I(N__83754));
    InMux I__19718 (
            .O(N__83757),
            .I(N__83751));
    Odrv4 I__19717 (
            .O(N__83754),
            .I(\timing_controller_inst.state_timeout_counter_2 ));
    LocalMux I__19716 (
            .O(N__83751),
            .I(\timing_controller_inst.state_timeout_counter_2 ));
    InMux I__19715 (
            .O(N__83746),
            .I(N__83743));
    LocalMux I__19714 (
            .O(N__83743),
            .I(\timing_controller_inst.n12553 ));
    InMux I__19713 (
            .O(N__83740),
            .I(\timing_controller_inst.n10589 ));
    InMux I__19712 (
            .O(N__83737),
            .I(N__83734));
    LocalMux I__19711 (
            .O(N__83734),
            .I(N__83730));
    CascadeMux I__19710 (
            .O(N__83733),
            .I(N__83727));
    Span4Mux_v I__19709 (
            .O(N__83730),
            .I(N__83724));
    InMux I__19708 (
            .O(N__83727),
            .I(N__83721));
    Odrv4 I__19707 (
            .O(N__83724),
            .I(\timing_controller_inst.state_timeout_counter_3 ));
    LocalMux I__19706 (
            .O(N__83721),
            .I(\timing_controller_inst.state_timeout_counter_3 ));
    InMux I__19705 (
            .O(N__83716),
            .I(N__83713));
    LocalMux I__19704 (
            .O(N__83713),
            .I(\timing_controller_inst.n12552 ));
    SRMux I__19703 (
            .O(N__83710),
            .I(N__83707));
    LocalMux I__19702 (
            .O(N__83707),
            .I(N__83704));
    Span4Mux_h I__19701 (
            .O(N__83704),
            .I(N__83701));
    Odrv4 I__19700 (
            .O(N__83701),
            .I(\pc_tx.n4468 ));
    CascadeMux I__19699 (
            .O(N__83698),
            .I(\pc_tx.n4_cascade_ ));
    InMux I__19698 (
            .O(N__83695),
            .I(N__83692));
    LocalMux I__19697 (
            .O(N__83692),
            .I(\pc_tx.n8 ));
    InMux I__19696 (
            .O(N__83689),
            .I(N__83686));
    LocalMux I__19695 (
            .O(N__83686),
            .I(\pc_tx.n7 ));
    InMux I__19694 (
            .O(N__83683),
            .I(N__83680));
    LocalMux I__19693 (
            .O(N__83680),
            .I(\pc_tx.n2813 ));
    CascadeMux I__19692 (
            .O(N__83677),
            .I(r_SM_Main_2_N_808_1_cascade_));
    InMux I__19691 (
            .O(N__83674),
            .I(N__83667));
    CascadeMux I__19690 (
            .O(N__83673),
            .I(N__83664));
    CascadeMux I__19689 (
            .O(N__83672),
            .I(N__83661));
    CascadeMux I__19688 (
            .O(N__83671),
            .I(N__83658));
    CascadeMux I__19687 (
            .O(N__83670),
            .I(N__83654));
    LocalMux I__19686 (
            .O(N__83667),
            .I(N__83648));
    InMux I__19685 (
            .O(N__83664),
            .I(N__83643));
    InMux I__19684 (
            .O(N__83661),
            .I(N__83643));
    InMux I__19683 (
            .O(N__83658),
            .I(N__83634));
    InMux I__19682 (
            .O(N__83657),
            .I(N__83634));
    InMux I__19681 (
            .O(N__83654),
            .I(N__83634));
    InMux I__19680 (
            .O(N__83653),
            .I(N__83634));
    InMux I__19679 (
            .O(N__83652),
            .I(N__83631));
    InMux I__19678 (
            .O(N__83651),
            .I(N__83628));
    Odrv4 I__19677 (
            .O(N__83648),
            .I(r_SM_Main_0));
    LocalMux I__19676 (
            .O(N__83643),
            .I(r_SM_Main_0));
    LocalMux I__19675 (
            .O(N__83634),
            .I(r_SM_Main_0));
    LocalMux I__19674 (
            .O(N__83631),
            .I(r_SM_Main_0));
    LocalMux I__19673 (
            .O(N__83628),
            .I(r_SM_Main_0));
    InMux I__19672 (
            .O(N__83617),
            .I(N__83614));
    LocalMux I__19671 (
            .O(N__83614),
            .I(N__83610));
    InMux I__19670 (
            .O(N__83613),
            .I(N__83607));
    Span4Mux_v I__19669 (
            .O(N__83610),
            .I(N__83593));
    LocalMux I__19668 (
            .O(N__83607),
            .I(N__83593));
    InMux I__19667 (
            .O(N__83606),
            .I(N__83590));
    InMux I__19666 (
            .O(N__83605),
            .I(N__83575));
    InMux I__19665 (
            .O(N__83604),
            .I(N__83575));
    InMux I__19664 (
            .O(N__83603),
            .I(N__83575));
    InMux I__19663 (
            .O(N__83602),
            .I(N__83575));
    InMux I__19662 (
            .O(N__83601),
            .I(N__83575));
    InMux I__19661 (
            .O(N__83600),
            .I(N__83575));
    InMux I__19660 (
            .O(N__83599),
            .I(N__83575));
    InMux I__19659 (
            .O(N__83598),
            .I(N__83572));
    Odrv4 I__19658 (
            .O(N__83593),
            .I(r_SM_Main_1));
    LocalMux I__19657 (
            .O(N__83590),
            .I(r_SM_Main_1));
    LocalMux I__19656 (
            .O(N__83575),
            .I(r_SM_Main_1));
    LocalMux I__19655 (
            .O(N__83572),
            .I(r_SM_Main_1));
    CascadeMux I__19654 (
            .O(N__83563),
            .I(N__83557));
    InMux I__19653 (
            .O(N__83562),
            .I(N__83546));
    InMux I__19652 (
            .O(N__83561),
            .I(N__83546));
    InMux I__19651 (
            .O(N__83560),
            .I(N__83546));
    InMux I__19650 (
            .O(N__83557),
            .I(N__83546));
    InMux I__19649 (
            .O(N__83556),
            .I(N__83541));
    InMux I__19648 (
            .O(N__83555),
            .I(N__83541));
    LocalMux I__19647 (
            .O(N__83546),
            .I(r_SM_Main_2_N_808_1));
    LocalMux I__19646 (
            .O(N__83541),
            .I(r_SM_Main_2_N_808_1));
    CascadeMux I__19645 (
            .O(N__83536),
            .I(N__83533));
    InMux I__19644 (
            .O(N__83533),
            .I(N__83527));
    InMux I__19643 (
            .O(N__83532),
            .I(N__83527));
    LocalMux I__19642 (
            .O(N__83527),
            .I(\pc_tx.r_SM_Main_2_N_805_0 ));
    InMux I__19641 (
            .O(N__83524),
            .I(N__83521));
    LocalMux I__19640 (
            .O(N__83521),
            .I(N__83518));
    Span4Mux_h I__19639 (
            .O(N__83518),
            .I(N__83511));
    InMux I__19638 (
            .O(N__83517),
            .I(N__83506));
    InMux I__19637 (
            .O(N__83516),
            .I(N__83506));
    InMux I__19636 (
            .O(N__83515),
            .I(N__83503));
    InMux I__19635 (
            .O(N__83514),
            .I(N__83500));
    Odrv4 I__19634 (
            .O(N__83511),
            .I(\pc_tx.r_Bit_Index_1 ));
    LocalMux I__19633 (
            .O(N__83506),
            .I(\pc_tx.r_Bit_Index_1 ));
    LocalMux I__19632 (
            .O(N__83503),
            .I(\pc_tx.r_Bit_Index_1 ));
    LocalMux I__19631 (
            .O(N__83500),
            .I(\pc_tx.r_Bit_Index_1 ));
    InMux I__19630 (
            .O(N__83491),
            .I(N__83485));
    InMux I__19629 (
            .O(N__83490),
            .I(N__83485));
    LocalMux I__19628 (
            .O(N__83485),
            .I(N__83481));
    CascadeMux I__19627 (
            .O(N__83484),
            .I(N__83478));
    Span4Mux_h I__19626 (
            .O(N__83481),
            .I(N__83473));
    InMux I__19625 (
            .O(N__83478),
            .I(N__83468));
    InMux I__19624 (
            .O(N__83477),
            .I(N__83468));
    InMux I__19623 (
            .O(N__83476),
            .I(N__83465));
    Odrv4 I__19622 (
            .O(N__83473),
            .I(\pc_tx.r_Bit_Index_2 ));
    LocalMux I__19621 (
            .O(N__83468),
            .I(\pc_tx.r_Bit_Index_2 ));
    LocalMux I__19620 (
            .O(N__83465),
            .I(\pc_tx.r_Bit_Index_2 ));
    InMux I__19619 (
            .O(N__83458),
            .I(N__83450));
    InMux I__19618 (
            .O(N__83457),
            .I(N__83450));
    InMux I__19617 (
            .O(N__83456),
            .I(N__83441));
    InMux I__19616 (
            .O(N__83455),
            .I(N__83441));
    LocalMux I__19615 (
            .O(N__83450),
            .I(N__83438));
    InMux I__19614 (
            .O(N__83449),
            .I(N__83429));
    InMux I__19613 (
            .O(N__83448),
            .I(N__83429));
    InMux I__19612 (
            .O(N__83447),
            .I(N__83429));
    InMux I__19611 (
            .O(N__83446),
            .I(N__83429));
    LocalMux I__19610 (
            .O(N__83441),
            .I(N__83425));
    Span4Mux_v I__19609 (
            .O(N__83438),
            .I(N__83420));
    LocalMux I__19608 (
            .O(N__83429),
            .I(N__83420));
    CascadeMux I__19607 (
            .O(N__83428),
            .I(N__83417));
    Span4Mux_h I__19606 (
            .O(N__83425),
            .I(N__83412));
    Span4Mux_h I__19605 (
            .O(N__83420),
            .I(N__83412));
    InMux I__19604 (
            .O(N__83417),
            .I(N__83409));
    Odrv4 I__19603 (
            .O(N__83412),
            .I(r_Bit_Index_0));
    LocalMux I__19602 (
            .O(N__83409),
            .I(r_Bit_Index_0));
    InMux I__19601 (
            .O(N__83404),
            .I(N__83401));
    LocalMux I__19600 (
            .O(N__83401),
            .I(N__83398));
    Span4Mux_h I__19599 (
            .O(N__83398),
            .I(N__83395));
    Span4Mux_v I__19598 (
            .O(N__83395),
            .I(N__83392));
    Odrv4 I__19597 (
            .O(N__83392),
            .I(n11319));
    InMux I__19596 (
            .O(N__83389),
            .I(N__83371));
    InMux I__19595 (
            .O(N__83388),
            .I(N__83362));
    InMux I__19594 (
            .O(N__83387),
            .I(N__83362));
    InMux I__19593 (
            .O(N__83386),
            .I(N__83362));
    InMux I__19592 (
            .O(N__83385),
            .I(N__83362));
    CascadeMux I__19591 (
            .O(N__83384),
            .I(N__83358));
    CascadeMux I__19590 (
            .O(N__83383),
            .I(N__83354));
    InMux I__19589 (
            .O(N__83382),
            .I(N__83345));
    InMux I__19588 (
            .O(N__83381),
            .I(N__83345));
    InMux I__19587 (
            .O(N__83380),
            .I(N__83345));
    InMux I__19586 (
            .O(N__83379),
            .I(N__83345));
    InMux I__19585 (
            .O(N__83378),
            .I(N__83336));
    InMux I__19584 (
            .O(N__83377),
            .I(N__83332));
    InMux I__19583 (
            .O(N__83376),
            .I(N__83329));
    InMux I__19582 (
            .O(N__83375),
            .I(N__83325));
    InMux I__19581 (
            .O(N__83374),
            .I(N__83322));
    LocalMux I__19580 (
            .O(N__83371),
            .I(N__83317));
    LocalMux I__19579 (
            .O(N__83362),
            .I(N__83317));
    InMux I__19578 (
            .O(N__83361),
            .I(N__83314));
    InMux I__19577 (
            .O(N__83358),
            .I(N__83308));
    InMux I__19576 (
            .O(N__83357),
            .I(N__83305));
    InMux I__19575 (
            .O(N__83354),
            .I(N__83302));
    LocalMux I__19574 (
            .O(N__83345),
            .I(N__83299));
    InMux I__19573 (
            .O(N__83344),
            .I(N__83295));
    InMux I__19572 (
            .O(N__83343),
            .I(N__83292));
    InMux I__19571 (
            .O(N__83342),
            .I(N__83287));
    InMux I__19570 (
            .O(N__83341),
            .I(N__83284));
    InMux I__19569 (
            .O(N__83340),
            .I(N__83281));
    InMux I__19568 (
            .O(N__83339),
            .I(N__83278));
    LocalMux I__19567 (
            .O(N__83336),
            .I(N__83275));
    InMux I__19566 (
            .O(N__83335),
            .I(N__83272));
    LocalMux I__19565 (
            .O(N__83332),
            .I(N__83267));
    LocalMux I__19564 (
            .O(N__83329),
            .I(N__83267));
    InMux I__19563 (
            .O(N__83328),
            .I(N__83264));
    LocalMux I__19562 (
            .O(N__83325),
            .I(N__83261));
    LocalMux I__19561 (
            .O(N__83322),
            .I(N__83258));
    Span4Mux_v I__19560 (
            .O(N__83317),
            .I(N__83255));
    LocalMux I__19559 (
            .O(N__83314),
            .I(N__83252));
    InMux I__19558 (
            .O(N__83313),
            .I(N__83247));
    InMux I__19557 (
            .O(N__83312),
            .I(N__83247));
    InMux I__19556 (
            .O(N__83311),
            .I(N__83244));
    LocalMux I__19555 (
            .O(N__83308),
            .I(N__83241));
    LocalMux I__19554 (
            .O(N__83305),
            .I(N__83234));
    LocalMux I__19553 (
            .O(N__83302),
            .I(N__83234));
    Span4Mux_h I__19552 (
            .O(N__83299),
            .I(N__83234));
    InMux I__19551 (
            .O(N__83298),
            .I(N__83231));
    LocalMux I__19550 (
            .O(N__83295),
            .I(N__83228));
    LocalMux I__19549 (
            .O(N__83292),
            .I(N__83225));
    InMux I__19548 (
            .O(N__83291),
            .I(N__83222));
    InMux I__19547 (
            .O(N__83290),
            .I(N__83219));
    LocalMux I__19546 (
            .O(N__83287),
            .I(N__83216));
    LocalMux I__19545 (
            .O(N__83284),
            .I(N__83209));
    LocalMux I__19544 (
            .O(N__83281),
            .I(N__83209));
    LocalMux I__19543 (
            .O(N__83278),
            .I(N__83209));
    Span4Mux_v I__19542 (
            .O(N__83275),
            .I(N__83206));
    LocalMux I__19541 (
            .O(N__83272),
            .I(N__83201));
    Span4Mux_v I__19540 (
            .O(N__83267),
            .I(N__83201));
    LocalMux I__19539 (
            .O(N__83264),
            .I(N__83198));
    Span4Mux_v I__19538 (
            .O(N__83261),
            .I(N__83191));
    Span4Mux_v I__19537 (
            .O(N__83258),
            .I(N__83191));
    Span4Mux_h I__19536 (
            .O(N__83255),
            .I(N__83191));
    Span4Mux_h I__19535 (
            .O(N__83252),
            .I(N__83180));
    LocalMux I__19534 (
            .O(N__83247),
            .I(N__83180));
    LocalMux I__19533 (
            .O(N__83244),
            .I(N__83180));
    Span4Mux_h I__19532 (
            .O(N__83241),
            .I(N__83180));
    Span4Mux_h I__19531 (
            .O(N__83234),
            .I(N__83180));
    LocalMux I__19530 (
            .O(N__83231),
            .I(N__83177));
    Span4Mux_h I__19529 (
            .O(N__83228),
            .I(N__83174));
    Span4Mux_v I__19528 (
            .O(N__83225),
            .I(N__83171));
    LocalMux I__19527 (
            .O(N__83222),
            .I(N__83158));
    LocalMux I__19526 (
            .O(N__83219),
            .I(N__83158));
    Span12Mux_s7_h I__19525 (
            .O(N__83216),
            .I(N__83158));
    Span12Mux_v I__19524 (
            .O(N__83209),
            .I(N__83158));
    Sp12to4 I__19523 (
            .O(N__83206),
            .I(N__83158));
    Sp12to4 I__19522 (
            .O(N__83201),
            .I(N__83158));
    Span4Mux_v I__19521 (
            .O(N__83198),
            .I(N__83153));
    Span4Mux_h I__19520 (
            .O(N__83191),
            .I(N__83153));
    Span4Mux_v I__19519 (
            .O(N__83180),
            .I(N__83150));
    Odrv12 I__19518 (
            .O(N__83177),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n44 ));
    Odrv4 I__19517 (
            .O(N__83174),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n44 ));
    Odrv4 I__19516 (
            .O(N__83171),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n44 ));
    Odrv12 I__19515 (
            .O(N__83158),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n44 ));
    Odrv4 I__19514 (
            .O(N__83153),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n44 ));
    Odrv4 I__19513 (
            .O(N__83150),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n44 ));
    InMux I__19512 (
            .O(N__83137),
            .I(N__83131));
    InMux I__19511 (
            .O(N__83136),
            .I(N__83131));
    LocalMux I__19510 (
            .O(N__83131),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_8 ));
    CascadeMux I__19509 (
            .O(N__83128),
            .I(N__83125));
    InMux I__19508 (
            .O(N__83125),
            .I(N__83122));
    LocalMux I__19507 (
            .O(N__83122),
            .I(N__83118));
    CascadeMux I__19506 (
            .O(N__83121),
            .I(N__83115));
    Span4Mux_h I__19505 (
            .O(N__83118),
            .I(N__83112));
    InMux I__19504 (
            .O(N__83115),
            .I(N__83109));
    Odrv4 I__19503 (
            .O(N__83112),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_8 ));
    LocalMux I__19502 (
            .O(N__83109),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_8 ));
    CascadeMux I__19501 (
            .O(N__83104),
            .I(N__83100));
    InMux I__19500 (
            .O(N__83103),
            .I(N__83097));
    InMux I__19499 (
            .O(N__83100),
            .I(N__83094));
    LocalMux I__19498 (
            .O(N__83097),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_8 ));
    LocalMux I__19497 (
            .O(N__83094),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_8 ));
    CascadeMux I__19496 (
            .O(N__83089),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13070_cascade_ ));
    CascadeMux I__19495 (
            .O(N__83086),
            .I(N__83083));
    InMux I__19494 (
            .O(N__83083),
            .I(N__83080));
    LocalMux I__19493 (
            .O(N__83080),
            .I(N__83077));
    Span4Mux_h I__19492 (
            .O(N__83077),
            .I(N__83073));
    InMux I__19491 (
            .O(N__83076),
            .I(N__83070));
    Odrv4 I__19490 (
            .O(N__83073),
            .I(REG_mem_6_8));
    LocalMux I__19489 (
            .O(N__83070),
            .I(REG_mem_6_8));
    InMux I__19488 (
            .O(N__83065),
            .I(N__83062));
    LocalMux I__19487 (
            .O(N__83062),
            .I(N__83058));
    InMux I__19486 (
            .O(N__83061),
            .I(N__83055));
    Odrv12 I__19485 (
            .O(N__83058),
            .I(REG_mem_7_8));
    LocalMux I__19484 (
            .O(N__83055),
            .I(REG_mem_7_8));
    CascadeMux I__19483 (
            .O(N__83050),
            .I(N__83047));
    InMux I__19482 (
            .O(N__83047),
            .I(N__83044));
    LocalMux I__19481 (
            .O(N__83044),
            .I(N__83041));
    Span4Mux_v I__19480 (
            .O(N__83041),
            .I(N__83038));
    Odrv4 I__19479 (
            .O(N__83038),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12824 ));
    InMux I__19478 (
            .O(N__83035),
            .I(N__83032));
    LocalMux I__19477 (
            .O(N__83032),
            .I(N__83029));
    Span4Mux_v I__19476 (
            .O(N__83029),
            .I(N__83026));
    Span4Mux_h I__19475 (
            .O(N__83026),
            .I(N__83023));
    Odrv4 I__19474 (
            .O(N__83023),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14246 ));
    CascadeMux I__19473 (
            .O(N__83020),
            .I(N__83017));
    InMux I__19472 (
            .O(N__83017),
            .I(N__83014));
    LocalMux I__19471 (
            .O(N__83014),
            .I(N__83011));
    Span4Mux_v I__19470 (
            .O(N__83011),
            .I(N__83008));
    Sp12to4 I__19469 (
            .O(N__83008),
            .I(N__83004));
    InMux I__19468 (
            .O(N__83007),
            .I(N__83001));
    Odrv12 I__19467 (
            .O(N__83004),
            .I(REG_mem_9_8));
    LocalMux I__19466 (
            .O(N__83001),
            .I(REG_mem_9_8));
    InMux I__19465 (
            .O(N__82996),
            .I(N__82993));
    LocalMux I__19464 (
            .O(N__82993),
            .I(N__82990));
    Span4Mux_h I__19463 (
            .O(N__82990),
            .I(N__82987));
    Span4Mux_h I__19462 (
            .O(N__82987),
            .I(N__82983));
    InMux I__19461 (
            .O(N__82986),
            .I(N__82980));
    Odrv4 I__19460 (
            .O(N__82983),
            .I(REG_mem_8_8));
    LocalMux I__19459 (
            .O(N__82980),
            .I(REG_mem_8_8));
    CascadeMux I__19458 (
            .O(N__82975),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11646_cascade_ ));
    InMux I__19457 (
            .O(N__82972),
            .I(N__82969));
    LocalMux I__19456 (
            .O(N__82969),
            .I(N__82966));
    Span4Mux_v I__19455 (
            .O(N__82966),
            .I(N__82963));
    Sp12to4 I__19454 (
            .O(N__82963),
            .I(N__82960));
    Span12Mux_h I__19453 (
            .O(N__82960),
            .I(N__82957));
    Odrv12 I__19452 (
            .O(N__82957),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11667 ));
    InMux I__19451 (
            .O(N__82954),
            .I(N__82946));
    InMux I__19450 (
            .O(N__82953),
            .I(N__82941));
    InMux I__19449 (
            .O(N__82952),
            .I(N__82941));
    InMux I__19448 (
            .O(N__82951),
            .I(N__82936));
    InMux I__19447 (
            .O(N__82950),
            .I(N__82931));
    InMux I__19446 (
            .O(N__82949),
            .I(N__82928));
    LocalMux I__19445 (
            .O(N__82946),
            .I(N__82922));
    LocalMux I__19444 (
            .O(N__82941),
            .I(N__82916));
    InMux I__19443 (
            .O(N__82940),
            .I(N__82911));
    InMux I__19442 (
            .O(N__82939),
            .I(N__82911));
    LocalMux I__19441 (
            .O(N__82936),
            .I(N__82905));
    InMux I__19440 (
            .O(N__82935),
            .I(N__82899));
    InMux I__19439 (
            .O(N__82934),
            .I(N__82899));
    LocalMux I__19438 (
            .O(N__82931),
            .I(N__82894));
    LocalMux I__19437 (
            .O(N__82928),
            .I(N__82891));
    InMux I__19436 (
            .O(N__82927),
            .I(N__82888));
    InMux I__19435 (
            .O(N__82926),
            .I(N__82882));
    InMux I__19434 (
            .O(N__82925),
            .I(N__82879));
    Span4Mux_v I__19433 (
            .O(N__82922),
            .I(N__82876));
    InMux I__19432 (
            .O(N__82921),
            .I(N__82873));
    InMux I__19431 (
            .O(N__82920),
            .I(N__82864));
    InMux I__19430 (
            .O(N__82919),
            .I(N__82864));
    Span4Mux_v I__19429 (
            .O(N__82916),
            .I(N__82859));
    LocalMux I__19428 (
            .O(N__82911),
            .I(N__82859));
    InMux I__19427 (
            .O(N__82910),
            .I(N__82856));
    InMux I__19426 (
            .O(N__82909),
            .I(N__82853));
    InMux I__19425 (
            .O(N__82908),
            .I(N__82850));
    Span4Mux_h I__19424 (
            .O(N__82905),
            .I(N__82847));
    InMux I__19423 (
            .O(N__82904),
            .I(N__82844));
    LocalMux I__19422 (
            .O(N__82899),
            .I(N__82841));
    InMux I__19421 (
            .O(N__82898),
            .I(N__82838));
    InMux I__19420 (
            .O(N__82897),
            .I(N__82835));
    Span4Mux_h I__19419 (
            .O(N__82894),
            .I(N__82832));
    Span4Mux_v I__19418 (
            .O(N__82891),
            .I(N__82827));
    LocalMux I__19417 (
            .O(N__82888),
            .I(N__82827));
    InMux I__19416 (
            .O(N__82887),
            .I(N__82824));
    InMux I__19415 (
            .O(N__82886),
            .I(N__82821));
    InMux I__19414 (
            .O(N__82885),
            .I(N__82818));
    LocalMux I__19413 (
            .O(N__82882),
            .I(N__82812));
    LocalMux I__19412 (
            .O(N__82879),
            .I(N__82812));
    Span4Mux_h I__19411 (
            .O(N__82876),
            .I(N__82807));
    LocalMux I__19410 (
            .O(N__82873),
            .I(N__82807));
    InMux I__19409 (
            .O(N__82872),
            .I(N__82798));
    InMux I__19408 (
            .O(N__82871),
            .I(N__82798));
    InMux I__19407 (
            .O(N__82870),
            .I(N__82798));
    InMux I__19406 (
            .O(N__82869),
            .I(N__82798));
    LocalMux I__19405 (
            .O(N__82864),
            .I(N__82795));
    Span4Mux_h I__19404 (
            .O(N__82859),
            .I(N__82788));
    LocalMux I__19403 (
            .O(N__82856),
            .I(N__82788));
    LocalMux I__19402 (
            .O(N__82853),
            .I(N__82788));
    LocalMux I__19401 (
            .O(N__82850),
            .I(N__82785));
    Span4Mux_h I__19400 (
            .O(N__82847),
            .I(N__82780));
    LocalMux I__19399 (
            .O(N__82844),
            .I(N__82780));
    Span4Mux_v I__19398 (
            .O(N__82841),
            .I(N__82777));
    LocalMux I__19397 (
            .O(N__82838),
            .I(N__82774));
    LocalMux I__19396 (
            .O(N__82835),
            .I(N__82771));
    Span4Mux_h I__19395 (
            .O(N__82832),
            .I(N__82760));
    Span4Mux_v I__19394 (
            .O(N__82827),
            .I(N__82760));
    LocalMux I__19393 (
            .O(N__82824),
            .I(N__82760));
    LocalMux I__19392 (
            .O(N__82821),
            .I(N__82760));
    LocalMux I__19391 (
            .O(N__82818),
            .I(N__82760));
    InMux I__19390 (
            .O(N__82817),
            .I(N__82757));
    Span12Mux_h I__19389 (
            .O(N__82812),
            .I(N__82753));
    Span4Mux_h I__19388 (
            .O(N__82807),
            .I(N__82750));
    LocalMux I__19387 (
            .O(N__82798),
            .I(N__82747));
    Span4Mux_v I__19386 (
            .O(N__82795),
            .I(N__82744));
    Span4Mux_v I__19385 (
            .O(N__82788),
            .I(N__82739));
    Span4Mux_v I__19384 (
            .O(N__82785),
            .I(N__82739));
    Span4Mux_h I__19383 (
            .O(N__82780),
            .I(N__82736));
    Span4Mux_h I__19382 (
            .O(N__82777),
            .I(N__82725));
    Span4Mux_v I__19381 (
            .O(N__82774),
            .I(N__82725));
    Span4Mux_v I__19380 (
            .O(N__82771),
            .I(N__82725));
    Span4Mux_v I__19379 (
            .O(N__82760),
            .I(N__82725));
    LocalMux I__19378 (
            .O(N__82757),
            .I(N__82725));
    InMux I__19377 (
            .O(N__82756),
            .I(N__82722));
    Odrv12 I__19376 (
            .O(N__82753),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616 ));
    Odrv4 I__19375 (
            .O(N__82750),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616 ));
    Odrv12 I__19374 (
            .O(N__82747),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616 ));
    Odrv4 I__19373 (
            .O(N__82744),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616 ));
    Odrv4 I__19372 (
            .O(N__82739),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616 ));
    Odrv4 I__19371 (
            .O(N__82736),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616 ));
    Odrv4 I__19370 (
            .O(N__82725),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616 ));
    LocalMux I__19369 (
            .O(N__82722),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616 ));
    InMux I__19368 (
            .O(N__82705),
            .I(N__82701));
    InMux I__19367 (
            .O(N__82704),
            .I(N__82698));
    LocalMux I__19366 (
            .O(N__82701),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_8 ));
    LocalMux I__19365 (
            .O(N__82698),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_8 ));
    InMux I__19364 (
            .O(N__82693),
            .I(N__82690));
    LocalMux I__19363 (
            .O(N__82690),
            .I(N__82687));
    Span4Mux_h I__19362 (
            .O(N__82687),
            .I(N__82683));
    CEMux I__19361 (
            .O(N__82686),
            .I(N__82680));
    Odrv4 I__19360 (
            .O(N__82683),
            .I(n4133));
    LocalMux I__19359 (
            .O(N__82680),
            .I(n4133));
    InMux I__19358 (
            .O(N__82675),
            .I(N__82672));
    LocalMux I__19357 (
            .O(N__82672),
            .I(n8));
    InMux I__19356 (
            .O(N__82669),
            .I(n10686));
    InMux I__19355 (
            .O(N__82666),
            .I(N__82663));
    LocalMux I__19354 (
            .O(N__82663),
            .I(n7_adj_1200));
    InMux I__19353 (
            .O(N__82660),
            .I(n10687));
    InMux I__19352 (
            .O(N__82657),
            .I(N__82654));
    LocalMux I__19351 (
            .O(N__82654),
            .I(n6));
    InMux I__19350 (
            .O(N__82651),
            .I(n10688));
    InMux I__19349 (
            .O(N__82648),
            .I(N__82645));
    LocalMux I__19348 (
            .O(N__82645),
            .I(n5_adj_1201));
    InMux I__19347 (
            .O(N__82642),
            .I(n10689));
    InMux I__19346 (
            .O(N__82639),
            .I(N__82636));
    LocalMux I__19345 (
            .O(N__82636),
            .I(n4_adj_1202));
    InMux I__19344 (
            .O(N__82633),
            .I(n10690));
    InMux I__19343 (
            .O(N__82630),
            .I(N__82627));
    LocalMux I__19342 (
            .O(N__82627),
            .I(n3));
    InMux I__19341 (
            .O(N__82624),
            .I(n10691));
    InMux I__19340 (
            .O(N__82621),
            .I(N__82618));
    LocalMux I__19339 (
            .O(N__82618),
            .I(n2_adj_1203));
    InMux I__19338 (
            .O(N__82615),
            .I(n10692));
    InMux I__19337 (
            .O(N__82612),
            .I(bfn_23_8_0_));
    IoInMux I__19336 (
            .O(N__82609),
            .I(N__82606));
    LocalMux I__19335 (
            .O(N__82606),
            .I(N__82603));
    Span4Mux_s2_h I__19334 (
            .O(N__82603),
            .I(N__82600));
    Span4Mux_v I__19333 (
            .O(N__82600),
            .I(N__82597));
    Span4Mux_v I__19332 (
            .O(N__82597),
            .I(N__82593));
    InMux I__19331 (
            .O(N__82596),
            .I(N__82590));
    Odrv4 I__19330 (
            .O(N__82593),
            .I(DEBUG_0_c_24));
    LocalMux I__19329 (
            .O(N__82590),
            .I(DEBUG_0_c_24));
    InMux I__19328 (
            .O(N__82585),
            .I(N__82582));
    LocalMux I__19327 (
            .O(N__82582),
            .I(n17_adj_1195));
    InMux I__19326 (
            .O(N__82579),
            .I(bfn_23_6_0_));
    InMux I__19325 (
            .O(N__82576),
            .I(N__82573));
    LocalMux I__19324 (
            .O(N__82573),
            .I(n16_adj_1196));
    InMux I__19323 (
            .O(N__82570),
            .I(n10678));
    InMux I__19322 (
            .O(N__82567),
            .I(N__82564));
    LocalMux I__19321 (
            .O(N__82564),
            .I(n15_adj_1197));
    InMux I__19320 (
            .O(N__82561),
            .I(n10679));
    InMux I__19319 (
            .O(N__82558),
            .I(N__82555));
    LocalMux I__19318 (
            .O(N__82555),
            .I(n14_adj_1198));
    InMux I__19317 (
            .O(N__82552),
            .I(n10680));
    InMux I__19316 (
            .O(N__82549),
            .I(N__82546));
    LocalMux I__19315 (
            .O(N__82546),
            .I(n13));
    InMux I__19314 (
            .O(N__82543),
            .I(n10681));
    InMux I__19313 (
            .O(N__82540),
            .I(N__82537));
    LocalMux I__19312 (
            .O(N__82537),
            .I(n12));
    InMux I__19311 (
            .O(N__82534),
            .I(n10682));
    InMux I__19310 (
            .O(N__82531),
            .I(N__82528));
    LocalMux I__19309 (
            .O(N__82528),
            .I(n11));
    InMux I__19308 (
            .O(N__82525),
            .I(n10683));
    InMux I__19307 (
            .O(N__82522),
            .I(N__82519));
    LocalMux I__19306 (
            .O(N__82519),
            .I(n10_adj_1199));
    InMux I__19305 (
            .O(N__82516),
            .I(n10684));
    InMux I__19304 (
            .O(N__82513),
            .I(N__82510));
    LocalMux I__19303 (
            .O(N__82510),
            .I(n9));
    InMux I__19302 (
            .O(N__82507),
            .I(bfn_23_7_0_));
    InMux I__19301 (
            .O(N__82504),
            .I(N__82501));
    LocalMux I__19300 (
            .O(N__82501),
            .I(n25_adj_1187));
    InMux I__19299 (
            .O(N__82498),
            .I(bfn_23_5_0_));
    InMux I__19298 (
            .O(N__82495),
            .I(N__82492));
    LocalMux I__19297 (
            .O(N__82492),
            .I(n24_adj_1188));
    InMux I__19296 (
            .O(N__82489),
            .I(n10670));
    InMux I__19295 (
            .O(N__82486),
            .I(N__82483));
    LocalMux I__19294 (
            .O(N__82483),
            .I(n23_adj_1189));
    InMux I__19293 (
            .O(N__82480),
            .I(n10671));
    InMux I__19292 (
            .O(N__82477),
            .I(N__82474));
    LocalMux I__19291 (
            .O(N__82474),
            .I(n22_adj_1190));
    InMux I__19290 (
            .O(N__82471),
            .I(n10672));
    InMux I__19289 (
            .O(N__82468),
            .I(N__82465));
    LocalMux I__19288 (
            .O(N__82465),
            .I(n21_adj_1191));
    InMux I__19287 (
            .O(N__82462),
            .I(n10673));
    InMux I__19286 (
            .O(N__82459),
            .I(N__82456));
    LocalMux I__19285 (
            .O(N__82456),
            .I(n20_adj_1192));
    InMux I__19284 (
            .O(N__82453),
            .I(n10674));
    InMux I__19283 (
            .O(N__82450),
            .I(N__82447));
    LocalMux I__19282 (
            .O(N__82447),
            .I(n19_adj_1193));
    InMux I__19281 (
            .O(N__82444),
            .I(n10675));
    InMux I__19280 (
            .O(N__82441),
            .I(N__82438));
    LocalMux I__19279 (
            .O(N__82438),
            .I(n18_adj_1194));
    InMux I__19278 (
            .O(N__82435),
            .I(n10676));
    CascadeMux I__19277 (
            .O(N__82432),
            .I(\timing_controller_inst.n1730_cascade_ ));
    CascadeMux I__19276 (
            .O(N__82429),
            .I(\timing_controller_inst.n1745_cascade_ ));
    CascadeMux I__19275 (
            .O(N__82426),
            .I(N__82421));
    CascadeMux I__19274 (
            .O(N__82425),
            .I(N__82417));
    CascadeMux I__19273 (
            .O(N__82424),
            .I(N__82414));
    InMux I__19272 (
            .O(N__82421),
            .I(N__82406));
    InMux I__19271 (
            .O(N__82420),
            .I(N__82406));
    InMux I__19270 (
            .O(N__82417),
            .I(N__82399));
    InMux I__19269 (
            .O(N__82414),
            .I(N__82399));
    InMux I__19268 (
            .O(N__82413),
            .I(N__82399));
    CascadeMux I__19267 (
            .O(N__82412),
            .I(N__82394));
    CascadeMux I__19266 (
            .O(N__82411),
            .I(N__82391));
    LocalMux I__19265 (
            .O(N__82406),
            .I(N__82386));
    LocalMux I__19264 (
            .O(N__82399),
            .I(N__82383));
    InMux I__19263 (
            .O(N__82398),
            .I(N__82378));
    InMux I__19262 (
            .O(N__82397),
            .I(N__82378));
    InMux I__19261 (
            .O(N__82394),
            .I(N__82369));
    InMux I__19260 (
            .O(N__82391),
            .I(N__82369));
    InMux I__19259 (
            .O(N__82390),
            .I(N__82369));
    InMux I__19258 (
            .O(N__82389),
            .I(N__82369));
    Span4Mux_h I__19257 (
            .O(N__82386),
            .I(N__82361));
    Span4Mux_v I__19256 (
            .O(N__82383),
            .I(N__82358));
    LocalMux I__19255 (
            .O(N__82378),
            .I(N__82355));
    LocalMux I__19254 (
            .O(N__82369),
            .I(N__82352));
    InMux I__19253 (
            .O(N__82368),
            .I(N__82345));
    InMux I__19252 (
            .O(N__82367),
            .I(N__82345));
    InMux I__19251 (
            .O(N__82366),
            .I(N__82345));
    InMux I__19250 (
            .O(N__82365),
            .I(N__82342));
    InMux I__19249 (
            .O(N__82364),
            .I(N__82339));
    Odrv4 I__19248 (
            .O(N__82361),
            .I(n1721));
    Odrv4 I__19247 (
            .O(N__82358),
            .I(n1721));
    Odrv12 I__19246 (
            .O(N__82355),
            .I(n1721));
    Odrv4 I__19245 (
            .O(N__82352),
            .I(n1721));
    LocalMux I__19244 (
            .O(N__82345),
            .I(n1721));
    LocalMux I__19243 (
            .O(N__82342),
            .I(n1721));
    LocalMux I__19242 (
            .O(N__82339),
            .I(n1721));
    CascadeMux I__19241 (
            .O(N__82324),
            .I(N__82307));
    CascadeMux I__19240 (
            .O(N__82323),
            .I(N__82304));
    CascadeMux I__19239 (
            .O(N__82322),
            .I(N__82301));
    CascadeMux I__19238 (
            .O(N__82321),
            .I(N__82298));
    CascadeMux I__19237 (
            .O(N__82320),
            .I(N__82294));
    InMux I__19236 (
            .O(N__82319),
            .I(N__82276));
    InMux I__19235 (
            .O(N__82318),
            .I(N__82276));
    InMux I__19234 (
            .O(N__82317),
            .I(N__82276));
    InMux I__19233 (
            .O(N__82316),
            .I(N__82276));
    InMux I__19232 (
            .O(N__82315),
            .I(N__82276));
    InMux I__19231 (
            .O(N__82314),
            .I(N__82276));
    InMux I__19230 (
            .O(N__82313),
            .I(N__82276));
    InMux I__19229 (
            .O(N__82312),
            .I(N__82269));
    InMux I__19228 (
            .O(N__82311),
            .I(N__82269));
    InMux I__19227 (
            .O(N__82310),
            .I(N__82269));
    InMux I__19226 (
            .O(N__82307),
            .I(N__82260));
    InMux I__19225 (
            .O(N__82304),
            .I(N__82260));
    InMux I__19224 (
            .O(N__82301),
            .I(N__82260));
    InMux I__19223 (
            .O(N__82298),
            .I(N__82260));
    InMux I__19222 (
            .O(N__82297),
            .I(N__82253));
    InMux I__19221 (
            .O(N__82294),
            .I(N__82253));
    InMux I__19220 (
            .O(N__82293),
            .I(N__82253));
    InMux I__19219 (
            .O(N__82292),
            .I(N__82248));
    InMux I__19218 (
            .O(N__82291),
            .I(N__82248));
    LocalMux I__19217 (
            .O(N__82276),
            .I(N__82234));
    LocalMux I__19216 (
            .O(N__82269),
            .I(N__82227));
    LocalMux I__19215 (
            .O(N__82260),
            .I(N__82227));
    LocalMux I__19214 (
            .O(N__82253),
            .I(N__82227));
    LocalMux I__19213 (
            .O(N__82248),
            .I(N__82224));
    InMux I__19212 (
            .O(N__82247),
            .I(N__82219));
    InMux I__19211 (
            .O(N__82246),
            .I(N__82219));
    InMux I__19210 (
            .O(N__82245),
            .I(N__82214));
    InMux I__19209 (
            .O(N__82244),
            .I(N__82214));
    CascadeMux I__19208 (
            .O(N__82243),
            .I(N__82210));
    CascadeMux I__19207 (
            .O(N__82242),
            .I(N__82207));
    CascadeMux I__19206 (
            .O(N__82241),
            .I(N__82203));
    CascadeMux I__19205 (
            .O(N__82240),
            .I(N__82200));
    CascadeMux I__19204 (
            .O(N__82239),
            .I(N__82197));
    CascadeMux I__19203 (
            .O(N__82238),
            .I(N__82181));
    CascadeMux I__19202 (
            .O(N__82237),
            .I(N__82178));
    Span4Mux_v I__19201 (
            .O(N__82234),
            .I(N__82171));
    Span4Mux_v I__19200 (
            .O(N__82227),
            .I(N__82162));
    Span4Mux_v I__19199 (
            .O(N__82224),
            .I(N__82162));
    LocalMux I__19198 (
            .O(N__82219),
            .I(N__82162));
    LocalMux I__19197 (
            .O(N__82214),
            .I(N__82162));
    InMux I__19196 (
            .O(N__82213),
            .I(N__82155));
    InMux I__19195 (
            .O(N__82210),
            .I(N__82155));
    InMux I__19194 (
            .O(N__82207),
            .I(N__82155));
    InMux I__19193 (
            .O(N__82206),
            .I(N__82146));
    InMux I__19192 (
            .O(N__82203),
            .I(N__82146));
    InMux I__19191 (
            .O(N__82200),
            .I(N__82146));
    InMux I__19190 (
            .O(N__82197),
            .I(N__82146));
    InMux I__19189 (
            .O(N__82196),
            .I(N__82131));
    InMux I__19188 (
            .O(N__82195),
            .I(N__82131));
    InMux I__19187 (
            .O(N__82194),
            .I(N__82131));
    InMux I__19186 (
            .O(N__82193),
            .I(N__82131));
    InMux I__19185 (
            .O(N__82192),
            .I(N__82131));
    InMux I__19184 (
            .O(N__82191),
            .I(N__82131));
    InMux I__19183 (
            .O(N__82190),
            .I(N__82131));
    InMux I__19182 (
            .O(N__82189),
            .I(N__82118));
    InMux I__19181 (
            .O(N__82188),
            .I(N__82118));
    InMux I__19180 (
            .O(N__82187),
            .I(N__82118));
    InMux I__19179 (
            .O(N__82186),
            .I(N__82118));
    InMux I__19178 (
            .O(N__82185),
            .I(N__82118));
    InMux I__19177 (
            .O(N__82184),
            .I(N__82118));
    InMux I__19176 (
            .O(N__82181),
            .I(N__82115));
    InMux I__19175 (
            .O(N__82178),
            .I(N__82104));
    InMux I__19174 (
            .O(N__82177),
            .I(N__82104));
    InMux I__19173 (
            .O(N__82176),
            .I(N__82104));
    InMux I__19172 (
            .O(N__82175),
            .I(N__82104));
    InMux I__19171 (
            .O(N__82174),
            .I(N__82104));
    Odrv4 I__19170 (
            .O(N__82171),
            .I(state_1));
    Odrv4 I__19169 (
            .O(N__82162),
            .I(state_1));
    LocalMux I__19168 (
            .O(N__82155),
            .I(state_1));
    LocalMux I__19167 (
            .O(N__82146),
            .I(state_1));
    LocalMux I__19166 (
            .O(N__82131),
            .I(state_1));
    LocalMux I__19165 (
            .O(N__82118),
            .I(state_1));
    LocalMux I__19164 (
            .O(N__82115),
            .I(state_1));
    LocalMux I__19163 (
            .O(N__82104),
            .I(state_1));
    InMux I__19162 (
            .O(N__82087),
            .I(N__82066));
    InMux I__19161 (
            .O(N__82086),
            .I(N__82066));
    InMux I__19160 (
            .O(N__82085),
            .I(N__82066));
    InMux I__19159 (
            .O(N__82084),
            .I(N__82066));
    InMux I__19158 (
            .O(N__82083),
            .I(N__82066));
    InMux I__19157 (
            .O(N__82082),
            .I(N__82066));
    InMux I__19156 (
            .O(N__82081),
            .I(N__82066));
    LocalMux I__19155 (
            .O(N__82066),
            .I(N__82063));
    Sp12to4 I__19154 (
            .O(N__82063),
            .I(N__82052));
    InMux I__19153 (
            .O(N__82062),
            .I(N__82049));
    InMux I__19152 (
            .O(N__82061),
            .I(N__82042));
    InMux I__19151 (
            .O(N__82060),
            .I(N__82042));
    InMux I__19150 (
            .O(N__82059),
            .I(N__82042));
    InMux I__19149 (
            .O(N__82058),
            .I(N__82033));
    InMux I__19148 (
            .O(N__82057),
            .I(N__82033));
    InMux I__19147 (
            .O(N__82056),
            .I(N__82033));
    InMux I__19146 (
            .O(N__82055),
            .I(N__82033));
    Span12Mux_v I__19145 (
            .O(N__82052),
            .I(N__82028));
    LocalMux I__19144 (
            .O(N__82049),
            .I(N__82023));
    LocalMux I__19143 (
            .O(N__82042),
            .I(N__82023));
    LocalMux I__19142 (
            .O(N__82033),
            .I(N__82020));
    InMux I__19141 (
            .O(N__82032),
            .I(N__82015));
    InMux I__19140 (
            .O(N__82031),
            .I(N__82015));
    Odrv12 I__19139 (
            .O(N__82028),
            .I(\timing_controller_inst.n1793 ));
    Odrv4 I__19138 (
            .O(N__82023),
            .I(\timing_controller_inst.n1793 ));
    Odrv12 I__19137 (
            .O(N__82020),
            .I(\timing_controller_inst.n1793 ));
    LocalMux I__19136 (
            .O(N__82015),
            .I(\timing_controller_inst.n1793 ));
    CascadeMux I__19135 (
            .O(N__82006),
            .I(\timing_controller_inst.n1744_cascade_ ));
    InMux I__19134 (
            .O(N__82003),
            .I(N__81982));
    InMux I__19133 (
            .O(N__82002),
            .I(N__81982));
    InMux I__19132 (
            .O(N__82001),
            .I(N__81982));
    InMux I__19131 (
            .O(N__82000),
            .I(N__81982));
    InMux I__19130 (
            .O(N__81999),
            .I(N__81982));
    InMux I__19129 (
            .O(N__81998),
            .I(N__81982));
    InMux I__19128 (
            .O(N__81997),
            .I(N__81982));
    LocalMux I__19127 (
            .O(N__81982),
            .I(N__81973));
    InMux I__19126 (
            .O(N__81981),
            .I(N__81966));
    InMux I__19125 (
            .O(N__81980),
            .I(N__81966));
    InMux I__19124 (
            .O(N__81979),
            .I(N__81966));
    InMux I__19123 (
            .O(N__81978),
            .I(N__81963));
    InMux I__19122 (
            .O(N__81977),
            .I(N__81958));
    InMux I__19121 (
            .O(N__81976),
            .I(N__81958));
    Span4Mux_v I__19120 (
            .O(N__81973),
            .I(N__81955));
    LocalMux I__19119 (
            .O(N__81966),
            .I(N__81952));
    LocalMux I__19118 (
            .O(N__81963),
            .I(N__81947));
    LocalMux I__19117 (
            .O(N__81958),
            .I(N__81947));
    Odrv4 I__19116 (
            .O(N__81955),
            .I(\timing_controller_inst.n11368 ));
    Odrv12 I__19115 (
            .O(N__81952),
            .I(\timing_controller_inst.n11368 ));
    Odrv4 I__19114 (
            .O(N__81947),
            .I(\timing_controller_inst.n11368 ));
    InMux I__19113 (
            .O(N__81940),
            .I(N__81937));
    LocalMux I__19112 (
            .O(N__81937),
            .I(\timing_controller_inst.n52 ));
    CascadeMux I__19111 (
            .O(N__81934),
            .I(\timing_controller_inst.n38_cascade_ ));
    InMux I__19110 (
            .O(N__81931),
            .I(N__81928));
    LocalMux I__19109 (
            .O(N__81928),
            .I(N__81925));
    Odrv4 I__19108 (
            .O(N__81925),
            .I(\timing_controller_inst.n58 ));
    SRMux I__19107 (
            .O(N__81922),
            .I(N__81919));
    LocalMux I__19106 (
            .O(N__81919),
            .I(\timing_controller_inst.n4586 ));
    InMux I__19105 (
            .O(N__81916),
            .I(N__81913));
    LocalMux I__19104 (
            .O(N__81913),
            .I(N__81905));
    InMux I__19103 (
            .O(N__81912),
            .I(N__81896));
    InMux I__19102 (
            .O(N__81911),
            .I(N__81896));
    InMux I__19101 (
            .O(N__81910),
            .I(N__81896));
    InMux I__19100 (
            .O(N__81909),
            .I(N__81896));
    CascadeMux I__19099 (
            .O(N__81908),
            .I(N__81893));
    Span4Mux_v I__19098 (
            .O(N__81905),
            .I(N__81876));
    LocalMux I__19097 (
            .O(N__81896),
            .I(N__81876));
    InMux I__19096 (
            .O(N__81893),
            .I(N__81867));
    InMux I__19095 (
            .O(N__81892),
            .I(N__81867));
    InMux I__19094 (
            .O(N__81891),
            .I(N__81867));
    InMux I__19093 (
            .O(N__81890),
            .I(N__81867));
    InMux I__19092 (
            .O(N__81889),
            .I(N__81860));
    InMux I__19091 (
            .O(N__81888),
            .I(N__81860));
    InMux I__19090 (
            .O(N__81887),
            .I(N__81860));
    InMux I__19089 (
            .O(N__81886),
            .I(N__81847));
    InMux I__19088 (
            .O(N__81885),
            .I(N__81847));
    InMux I__19087 (
            .O(N__81884),
            .I(N__81847));
    InMux I__19086 (
            .O(N__81883),
            .I(N__81847));
    InMux I__19085 (
            .O(N__81882),
            .I(N__81847));
    InMux I__19084 (
            .O(N__81881),
            .I(N__81847));
    Odrv4 I__19083 (
            .O(N__81876),
            .I(state_2));
    LocalMux I__19082 (
            .O(N__81867),
            .I(state_2));
    LocalMux I__19081 (
            .O(N__81860),
            .I(state_2));
    LocalMux I__19080 (
            .O(N__81847),
            .I(state_2));
    CascadeMux I__19079 (
            .O(N__81838),
            .I(N__81834));
    CascadeMux I__19078 (
            .O(N__81837),
            .I(N__81830));
    InMux I__19077 (
            .O(N__81834),
            .I(N__81823));
    InMux I__19076 (
            .O(N__81833),
            .I(N__81823));
    InMux I__19075 (
            .O(N__81830),
            .I(N__81823));
    LocalMux I__19074 (
            .O(N__81823),
            .I(n3929));
    InMux I__19073 (
            .O(N__81820),
            .I(N__81817));
    LocalMux I__19072 (
            .O(N__81817),
            .I(N__81814));
    Odrv12 I__19071 (
            .O(N__81814),
            .I(\timing_controller_inst.n54 ));
    CascadeMux I__19070 (
            .O(N__81811),
            .I(\timing_controller_inst.n1751_cascade_ ));
    CascadeMux I__19069 (
            .O(N__81808),
            .I(\timing_controller_inst.n1732_cascade_ ));
    InMux I__19068 (
            .O(N__81805),
            .I(N__81802));
    LocalMux I__19067 (
            .O(N__81802),
            .I(N__81799));
    Odrv4 I__19066 (
            .O(N__81799),
            .I(\timing_controller_inst.n1731 ));
    InMux I__19065 (
            .O(N__81796),
            .I(N__81793));
    LocalMux I__19064 (
            .O(N__81793),
            .I(\timing_controller_inst.n1875 ));
    InMux I__19063 (
            .O(N__81790),
            .I(N__81784));
    InMux I__19062 (
            .O(N__81789),
            .I(N__81784));
    LocalMux I__19061 (
            .O(N__81784),
            .I(N__81781));
    Odrv12 I__19060 (
            .O(N__81781),
            .I(n7566));
    InMux I__19059 (
            .O(N__81778),
            .I(N__81764));
    InMux I__19058 (
            .O(N__81777),
            .I(N__81764));
    InMux I__19057 (
            .O(N__81776),
            .I(N__81764));
    InMux I__19056 (
            .O(N__81775),
            .I(N__81764));
    CascadeMux I__19055 (
            .O(N__81774),
            .I(N__81761));
    CascadeMux I__19054 (
            .O(N__81773),
            .I(N__81757));
    LocalMux I__19053 (
            .O(N__81764),
            .I(N__81751));
    InMux I__19052 (
            .O(N__81761),
            .I(N__81746));
    InMux I__19051 (
            .O(N__81760),
            .I(N__81746));
    InMux I__19050 (
            .O(N__81757),
            .I(N__81743));
    InMux I__19049 (
            .O(N__81756),
            .I(N__81740));
    CascadeMux I__19048 (
            .O(N__81755),
            .I(N__81735));
    CascadeMux I__19047 (
            .O(N__81754),
            .I(N__81732));
    Span4Mux_h I__19046 (
            .O(N__81751),
            .I(N__81727));
    LocalMux I__19045 (
            .O(N__81746),
            .I(N__81727));
    LocalMux I__19044 (
            .O(N__81743),
            .I(N__81722));
    LocalMux I__19043 (
            .O(N__81740),
            .I(N__81722));
    InMux I__19042 (
            .O(N__81739),
            .I(N__81713));
    InMux I__19041 (
            .O(N__81738),
            .I(N__81713));
    InMux I__19040 (
            .O(N__81735),
            .I(N__81713));
    InMux I__19039 (
            .O(N__81732),
            .I(N__81713));
    Span4Mux_v I__19038 (
            .O(N__81727),
            .I(N__81710));
    Span4Mux_v I__19037 (
            .O(N__81722),
            .I(N__81707));
    LocalMux I__19036 (
            .O(N__81713),
            .I(N__81704));
    Odrv4 I__19035 (
            .O(N__81710),
            .I(n63));
    Odrv4 I__19034 (
            .O(N__81707),
            .I(n63));
    Odrv12 I__19033 (
            .O(N__81704),
            .I(n63));
    InMux I__19032 (
            .O(N__81697),
            .I(N__81694));
    LocalMux I__19031 (
            .O(N__81694),
            .I(N__81691));
    Span4Mux_v I__19030 (
            .O(N__81691),
            .I(N__81688));
    Odrv4 I__19029 (
            .O(N__81688),
            .I(n1876));
    CascadeMux I__19028 (
            .O(N__81685),
            .I(n1721_cascade_));
    CascadeMux I__19027 (
            .O(N__81682),
            .I(\timing_controller_inst.n11347_cascade_ ));
    InMux I__19026 (
            .O(N__81679),
            .I(N__81667));
    InMux I__19025 (
            .O(N__81678),
            .I(N__81667));
    InMux I__19024 (
            .O(N__81677),
            .I(N__81660));
    InMux I__19023 (
            .O(N__81676),
            .I(N__81660));
    InMux I__19022 (
            .O(N__81675),
            .I(N__81660));
    InMux I__19021 (
            .O(N__81674),
            .I(N__81653));
    InMux I__19020 (
            .O(N__81673),
            .I(N__81653));
    InMux I__19019 (
            .O(N__81672),
            .I(N__81653));
    LocalMux I__19018 (
            .O(N__81667),
            .I(N__81650));
    LocalMux I__19017 (
            .O(N__81660),
            .I(N__81647));
    LocalMux I__19016 (
            .O(N__81653),
            .I(N__81644));
    Span4Mux_v I__19015 (
            .O(N__81650),
            .I(N__81641));
    Span4Mux_h I__19014 (
            .O(N__81647),
            .I(N__81636));
    Span4Mux_h I__19013 (
            .O(N__81644),
            .I(N__81636));
    Odrv4 I__19012 (
            .O(N__81641),
            .I(n3710));
    Odrv4 I__19011 (
            .O(N__81636),
            .I(n3710));
    InMux I__19010 (
            .O(N__81631),
            .I(N__81622));
    InMux I__19009 (
            .O(N__81630),
            .I(N__81622));
    InMux I__19008 (
            .O(N__81629),
            .I(N__81622));
    LocalMux I__19007 (
            .O(N__81622),
            .I(N__81619));
    Span4Mux_h I__19006 (
            .O(N__81619),
            .I(N__81615));
    CascadeMux I__19005 (
            .O(N__81618),
            .I(N__81612));
    Span4Mux_v I__19004 (
            .O(N__81615),
            .I(N__81609));
    InMux I__19003 (
            .O(N__81612),
            .I(N__81606));
    Odrv4 I__19002 (
            .O(N__81609),
            .I(r_SM_Main_2_N_811_0));
    LocalMux I__19001 (
            .O(N__81606),
            .I(r_SM_Main_2_N_811_0));
    InMux I__19000 (
            .O(N__81601),
            .I(N__81598));
    LocalMux I__18999 (
            .O(N__81598),
            .I(N__81595));
    Span4Mux_v I__18998 (
            .O(N__81595),
            .I(N__81592));
    Odrv4 I__18997 (
            .O(N__81592),
            .I(\timing_controller_inst.n50 ));
    IoInMux I__18996 (
            .O(N__81589),
            .I(N__81586));
    LocalMux I__18995 (
            .O(N__81586),
            .I(N__81583));
    Span4Mux_s2_h I__18994 (
            .O(N__81583),
            .I(N__81580));
    Span4Mux_h I__18993 (
            .O(N__81580),
            .I(N__81577));
    Odrv4 I__18992 (
            .O(N__81577),
            .I(UPDATE_c_3));
    SRMux I__18991 (
            .O(N__81574),
            .I(N__81571));
    LocalMux I__18990 (
            .O(N__81571),
            .I(N__81568));
    Odrv4 I__18989 (
            .O(N__81568),
            .I(\timing_controller_inst.n5 ));
    CascadeMux I__18988 (
            .O(N__81565),
            .I(n7495_cascade_));
    InMux I__18987 (
            .O(N__81562),
            .I(N__81559));
    LocalMux I__18986 (
            .O(N__81559),
            .I(N__81556));
    Odrv12 I__18985 (
            .O(N__81556),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11874 ));
    InMux I__18984 (
            .O(N__81553),
            .I(N__81550));
    LocalMux I__18983 (
            .O(N__81550),
            .I(N__81547));
    Odrv4 I__18982 (
            .O(N__81547),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11862 ));
    InMux I__18981 (
            .O(N__81544),
            .I(N__81541));
    LocalMux I__18980 (
            .O(N__81541),
            .I(N__81538));
    Odrv12 I__18979 (
            .O(N__81538),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11853 ));
    CascadeMux I__18978 (
            .O(N__81535),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13082_cascade_ ));
    InMux I__18977 (
            .O(N__81532),
            .I(N__81529));
    LocalMux I__18976 (
            .O(N__81529),
            .I(N__81526));
    Span4Mux_h I__18975 (
            .O(N__81526),
            .I(N__81523));
    Span4Mux_h I__18974 (
            .O(N__81523),
            .I(N__81520));
    Odrv4 I__18973 (
            .O(N__81520),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11841 ));
    CascadeMux I__18972 (
            .O(N__81517),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11913_cascade_ ));
    InMux I__18971 (
            .O(N__81514),
            .I(N__81507));
    InMux I__18970 (
            .O(N__81513),
            .I(N__81504));
    InMux I__18969 (
            .O(N__81512),
            .I(N__81499));
    InMux I__18968 (
            .O(N__81511),
            .I(N__81499));
    InMux I__18967 (
            .O(N__81510),
            .I(N__81496));
    LocalMux I__18966 (
            .O(N__81507),
            .I(N__81492));
    LocalMux I__18965 (
            .O(N__81504),
            .I(N__81489));
    LocalMux I__18964 (
            .O(N__81499),
            .I(N__81486));
    LocalMux I__18963 (
            .O(N__81496),
            .I(N__81483));
    InMux I__18962 (
            .O(N__81495),
            .I(N__81475));
    Span4Mux_h I__18961 (
            .O(N__81492),
            .I(N__81457));
    Span4Mux_h I__18960 (
            .O(N__81489),
            .I(N__81457));
    Span4Mux_v I__18959 (
            .O(N__81486),
            .I(N__81457));
    Span4Mux_v I__18958 (
            .O(N__81483),
            .I(N__81457));
    InMux I__18957 (
            .O(N__81482),
            .I(N__81454));
    InMux I__18956 (
            .O(N__81481),
            .I(N__81451));
    InMux I__18955 (
            .O(N__81480),
            .I(N__81443));
    InMux I__18954 (
            .O(N__81479),
            .I(N__81443));
    InMux I__18953 (
            .O(N__81478),
            .I(N__81434));
    LocalMux I__18952 (
            .O(N__81475),
            .I(N__81430));
    InMux I__18951 (
            .O(N__81474),
            .I(N__81425));
    InMux I__18950 (
            .O(N__81473),
            .I(N__81425));
    InMux I__18949 (
            .O(N__81472),
            .I(N__81422));
    InMux I__18948 (
            .O(N__81471),
            .I(N__81417));
    InMux I__18947 (
            .O(N__81470),
            .I(N__81417));
    InMux I__18946 (
            .O(N__81469),
            .I(N__81413));
    InMux I__18945 (
            .O(N__81468),
            .I(N__81410));
    InMux I__18944 (
            .O(N__81467),
            .I(N__81405));
    InMux I__18943 (
            .O(N__81466),
            .I(N__81405));
    Span4Mux_h I__18942 (
            .O(N__81457),
            .I(N__81400));
    LocalMux I__18941 (
            .O(N__81454),
            .I(N__81400));
    LocalMux I__18940 (
            .O(N__81451),
            .I(N__81396));
    InMux I__18939 (
            .O(N__81450),
            .I(N__81393));
    InMux I__18938 (
            .O(N__81449),
            .I(N__81388));
    InMux I__18937 (
            .O(N__81448),
            .I(N__81388));
    LocalMux I__18936 (
            .O(N__81443),
            .I(N__81385));
    InMux I__18935 (
            .O(N__81442),
            .I(N__81382));
    InMux I__18934 (
            .O(N__81441),
            .I(N__81377));
    InMux I__18933 (
            .O(N__81440),
            .I(N__81377));
    InMux I__18932 (
            .O(N__81439),
            .I(N__81374));
    InMux I__18931 (
            .O(N__81438),
            .I(N__81369));
    InMux I__18930 (
            .O(N__81437),
            .I(N__81369));
    LocalMux I__18929 (
            .O(N__81434),
            .I(N__81366));
    InMux I__18928 (
            .O(N__81433),
            .I(N__81363));
    Span4Mux_v I__18927 (
            .O(N__81430),
            .I(N__81358));
    LocalMux I__18926 (
            .O(N__81425),
            .I(N__81358));
    LocalMux I__18925 (
            .O(N__81422),
            .I(N__81355));
    LocalMux I__18924 (
            .O(N__81417),
            .I(N__81352));
    InMux I__18923 (
            .O(N__81416),
            .I(N__81349));
    LocalMux I__18922 (
            .O(N__81413),
            .I(N__81343));
    LocalMux I__18921 (
            .O(N__81410),
            .I(N__81343));
    LocalMux I__18920 (
            .O(N__81405),
            .I(N__81340));
    Span4Mux_h I__18919 (
            .O(N__81400),
            .I(N__81337));
    CascadeMux I__18918 (
            .O(N__81399),
            .I(N__81334));
    Span4Mux_v I__18917 (
            .O(N__81396),
            .I(N__81329));
    LocalMux I__18916 (
            .O(N__81393),
            .I(N__81329));
    LocalMux I__18915 (
            .O(N__81388),
            .I(N__81326));
    Span4Mux_h I__18914 (
            .O(N__81385),
            .I(N__81321));
    LocalMux I__18913 (
            .O(N__81382),
            .I(N__81321));
    LocalMux I__18912 (
            .O(N__81377),
            .I(N__81314));
    LocalMux I__18911 (
            .O(N__81374),
            .I(N__81314));
    LocalMux I__18910 (
            .O(N__81369),
            .I(N__81314));
    Span4Mux_v I__18909 (
            .O(N__81366),
            .I(N__81309));
    LocalMux I__18908 (
            .O(N__81363),
            .I(N__81309));
    Span4Mux_v I__18907 (
            .O(N__81358),
            .I(N__81306));
    Span4Mux_v I__18906 (
            .O(N__81355),
            .I(N__81302));
    Span4Mux_v I__18905 (
            .O(N__81352),
            .I(N__81297));
    LocalMux I__18904 (
            .O(N__81349),
            .I(N__81297));
    InMux I__18903 (
            .O(N__81348),
            .I(N__81294));
    Span4Mux_v I__18902 (
            .O(N__81343),
            .I(N__81290));
    Span4Mux_h I__18901 (
            .O(N__81340),
            .I(N__81283));
    Span4Mux_v I__18900 (
            .O(N__81337),
            .I(N__81283));
    InMux I__18899 (
            .O(N__81334),
            .I(N__81280));
    Span4Mux_v I__18898 (
            .O(N__81329),
            .I(N__81277));
    Span4Mux_v I__18897 (
            .O(N__81326),
            .I(N__81274));
    Span4Mux_v I__18896 (
            .O(N__81321),
            .I(N__81270));
    Span4Mux_v I__18895 (
            .O(N__81314),
            .I(N__81265));
    Span4Mux_h I__18894 (
            .O(N__81309),
            .I(N__81265));
    Span4Mux_v I__18893 (
            .O(N__81306),
            .I(N__81262));
    InMux I__18892 (
            .O(N__81305),
            .I(N__81259));
    Span4Mux_h I__18891 (
            .O(N__81302),
            .I(N__81252));
    Span4Mux_h I__18890 (
            .O(N__81297),
            .I(N__81252));
    LocalMux I__18889 (
            .O(N__81294),
            .I(N__81252));
    CascadeMux I__18888 (
            .O(N__81293),
            .I(N__81249));
    Span4Mux_v I__18887 (
            .O(N__81290),
            .I(N__81246));
    InMux I__18886 (
            .O(N__81289),
            .I(N__81240));
    InMux I__18885 (
            .O(N__81288),
            .I(N__81240));
    Span4Mux_v I__18884 (
            .O(N__81283),
            .I(N__81234));
    LocalMux I__18883 (
            .O(N__81280),
            .I(N__81234));
    Span4Mux_v I__18882 (
            .O(N__81277),
            .I(N__81230));
    Span4Mux_v I__18881 (
            .O(N__81274),
            .I(N__81227));
    InMux I__18880 (
            .O(N__81273),
            .I(N__81224));
    Span4Mux_h I__18879 (
            .O(N__81270),
            .I(N__81219));
    Span4Mux_v I__18878 (
            .O(N__81265),
            .I(N__81219));
    Span4Mux_h I__18877 (
            .O(N__81262),
            .I(N__81214));
    LocalMux I__18876 (
            .O(N__81259),
            .I(N__81214));
    Span4Mux_v I__18875 (
            .O(N__81252),
            .I(N__81211));
    InMux I__18874 (
            .O(N__81249),
            .I(N__81208));
    Span4Mux_h I__18873 (
            .O(N__81246),
            .I(N__81205));
    InMux I__18872 (
            .O(N__81245),
            .I(N__81202));
    LocalMux I__18871 (
            .O(N__81240),
            .I(N__81199));
    InMux I__18870 (
            .O(N__81239),
            .I(N__81196));
    Span4Mux_h I__18869 (
            .O(N__81234),
            .I(N__81192));
    CascadeMux I__18868 (
            .O(N__81233),
            .I(N__81188));
    Sp12to4 I__18867 (
            .O(N__81230),
            .I(N__81179));
    Sp12to4 I__18866 (
            .O(N__81227),
            .I(N__81179));
    LocalMux I__18865 (
            .O(N__81224),
            .I(N__81179));
    Span4Mux_v I__18864 (
            .O(N__81219),
            .I(N__81174));
    Span4Mux_h I__18863 (
            .O(N__81214),
            .I(N__81174));
    Span4Mux_h I__18862 (
            .O(N__81211),
            .I(N__81169));
    LocalMux I__18861 (
            .O(N__81208),
            .I(N__81169));
    Span4Mux_v I__18860 (
            .O(N__81205),
            .I(N__81164));
    LocalMux I__18859 (
            .O(N__81202),
            .I(N__81164));
    Span12Mux_v I__18858 (
            .O(N__81199),
            .I(N__81159));
    LocalMux I__18857 (
            .O(N__81196),
            .I(N__81159));
    InMux I__18856 (
            .O(N__81195),
            .I(N__81156));
    Span4Mux_v I__18855 (
            .O(N__81192),
            .I(N__81153));
    InMux I__18854 (
            .O(N__81191),
            .I(N__81146));
    InMux I__18853 (
            .O(N__81188),
            .I(N__81146));
    InMux I__18852 (
            .O(N__81187),
            .I(N__81146));
    CascadeMux I__18851 (
            .O(N__81186),
            .I(N__81143));
    Span12Mux_h I__18850 (
            .O(N__81179),
            .I(N__81140));
    Span4Mux_v I__18849 (
            .O(N__81174),
            .I(N__81135));
    Span4Mux_h I__18848 (
            .O(N__81169),
            .I(N__81135));
    Span4Mux_v I__18847 (
            .O(N__81164),
            .I(N__81132));
    Span12Mux_v I__18846 (
            .O(N__81159),
            .I(N__81127));
    LocalMux I__18845 (
            .O(N__81156),
            .I(N__81127));
    Span4Mux_h I__18844 (
            .O(N__81153),
            .I(N__81122));
    LocalMux I__18843 (
            .O(N__81146),
            .I(N__81122));
    InMux I__18842 (
            .O(N__81143),
            .I(N__81119));
    Odrv12 I__18841 (
            .O(N__81140),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4 ));
    Odrv4 I__18840 (
            .O(N__81135),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4 ));
    Odrv4 I__18839 (
            .O(N__81132),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4 ));
    Odrv12 I__18838 (
            .O(N__81127),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4 ));
    Odrv4 I__18837 (
            .O(N__81122),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4 ));
    LocalMux I__18836 (
            .O(N__81119),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4 ));
    InMux I__18835 (
            .O(N__81106),
            .I(N__81103));
    LocalMux I__18834 (
            .O(N__81103),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11898 ));
    InMux I__18833 (
            .O(N__81100),
            .I(N__81094));
    InMux I__18832 (
            .O(N__81099),
            .I(N__81094));
    LocalMux I__18831 (
            .O(N__81094),
            .I(N__81088));
    InMux I__18830 (
            .O(N__81093),
            .I(N__81083));
    InMux I__18829 (
            .O(N__81092),
            .I(N__81078));
    InMux I__18828 (
            .O(N__81091),
            .I(N__81078));
    Span4Mux_h I__18827 (
            .O(N__81088),
            .I(N__81075));
    InMux I__18826 (
            .O(N__81087),
            .I(N__81070));
    InMux I__18825 (
            .O(N__81086),
            .I(N__81070));
    LocalMux I__18824 (
            .O(N__81083),
            .I(N__81067));
    LocalMux I__18823 (
            .O(N__81078),
            .I(N__81064));
    Span4Mux_v I__18822 (
            .O(N__81075),
            .I(N__81057));
    LocalMux I__18821 (
            .O(N__81070),
            .I(N__81057));
    Span4Mux_v I__18820 (
            .O(N__81067),
            .I(N__81046));
    Span4Mux_h I__18819 (
            .O(N__81064),
            .I(N__81043));
    InMux I__18818 (
            .O(N__81063),
            .I(N__81038));
    InMux I__18817 (
            .O(N__81062),
            .I(N__81038));
    Span4Mux_v I__18816 (
            .O(N__81057),
            .I(N__81034));
    InMux I__18815 (
            .O(N__81056),
            .I(N__81017));
    InMux I__18814 (
            .O(N__81055),
            .I(N__81017));
    InMux I__18813 (
            .O(N__81054),
            .I(N__81017));
    InMux I__18812 (
            .O(N__81053),
            .I(N__81017));
    InMux I__18811 (
            .O(N__81052),
            .I(N__81017));
    InMux I__18810 (
            .O(N__81051),
            .I(N__81017));
    InMux I__18809 (
            .O(N__81050),
            .I(N__81017));
    InMux I__18808 (
            .O(N__81049),
            .I(N__81017));
    Span4Mux_v I__18807 (
            .O(N__81046),
            .I(N__81012));
    Span4Mux_h I__18806 (
            .O(N__81043),
            .I(N__81007));
    LocalMux I__18805 (
            .O(N__81038),
            .I(N__81007));
    InMux I__18804 (
            .O(N__81037),
            .I(N__81004));
    Span4Mux_h I__18803 (
            .O(N__81034),
            .I(N__80999));
    LocalMux I__18802 (
            .O(N__81017),
            .I(N__80999));
    InMux I__18801 (
            .O(N__81016),
            .I(N__80994));
    InMux I__18800 (
            .O(N__81015),
            .I(N__80994));
    Span4Mux_v I__18799 (
            .O(N__81012),
            .I(N__80989));
    Span4Mux_h I__18798 (
            .O(N__81007),
            .I(N__80986));
    LocalMux I__18797 (
            .O(N__81004),
            .I(N__80983));
    Span4Mux_h I__18796 (
            .O(N__80999),
            .I(N__80980));
    LocalMux I__18795 (
            .O(N__80994),
            .I(N__80977));
    InMux I__18794 (
            .O(N__80993),
            .I(N__80972));
    InMux I__18793 (
            .O(N__80992),
            .I(N__80972));
    Span4Mux_v I__18792 (
            .O(N__80989),
            .I(N__80969));
    Span4Mux_v I__18791 (
            .O(N__80986),
            .I(N__80966));
    Span4Mux_v I__18790 (
            .O(N__80983),
            .I(N__80963));
    Span4Mux_h I__18789 (
            .O(N__80980),
            .I(N__80958));
    Span4Mux_h I__18788 (
            .O(N__80977),
            .I(N__80958));
    LocalMux I__18787 (
            .O(N__80972),
            .I(N__80955));
    Sp12to4 I__18786 (
            .O(N__80969),
            .I(N__80946));
    Span4Mux_v I__18785 (
            .O(N__80966),
            .I(N__80941));
    Span4Mux_h I__18784 (
            .O(N__80963),
            .I(N__80941));
    Span4Mux_v I__18783 (
            .O(N__80958),
            .I(N__80938));
    Span4Mux_v I__18782 (
            .O(N__80955),
            .I(N__80935));
    InMux I__18781 (
            .O(N__80954),
            .I(N__80932));
    InMux I__18780 (
            .O(N__80953),
            .I(N__80927));
    InMux I__18779 (
            .O(N__80952),
            .I(N__80927));
    InMux I__18778 (
            .O(N__80951),
            .I(N__80920));
    InMux I__18777 (
            .O(N__80950),
            .I(N__80920));
    InMux I__18776 (
            .O(N__80949),
            .I(N__80920));
    Odrv12 I__18775 (
            .O(N__80946),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_5 ));
    Odrv4 I__18774 (
            .O(N__80941),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_5 ));
    Odrv4 I__18773 (
            .O(N__80938),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_5 ));
    Odrv4 I__18772 (
            .O(N__80935),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_5 ));
    LocalMux I__18771 (
            .O(N__80932),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_5 ));
    LocalMux I__18770 (
            .O(N__80927),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_5 ));
    LocalMux I__18769 (
            .O(N__80920),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_5 ));
    CascadeMux I__18768 (
            .O(N__80905),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13058_cascade_ ));
    CascadeMux I__18767 (
            .O(N__80902),
            .I(N__80899));
    InMux I__18766 (
            .O(N__80899),
            .I(N__80896));
    LocalMux I__18765 (
            .O(N__80896),
            .I(N__80893));
    Span4Mux_v I__18764 (
            .O(N__80893),
            .I(N__80890));
    Span4Mux_h I__18763 (
            .O(N__80890),
            .I(N__80887));
    Span4Mux_v I__18762 (
            .O(N__80887),
            .I(N__80884));
    Odrv4 I__18761 (
            .O(N__80884),
            .I(REG_out_raw_8));
    CEMux I__18760 (
            .O(N__80881),
            .I(N__80877));
    CEMux I__18759 (
            .O(N__80880),
            .I(N__80873));
    LocalMux I__18758 (
            .O(N__80877),
            .I(N__80868));
    CEMux I__18757 (
            .O(N__80876),
            .I(N__80863));
    LocalMux I__18756 (
            .O(N__80873),
            .I(N__80858));
    CEMux I__18755 (
            .O(N__80872),
            .I(N__80855));
    CEMux I__18754 (
            .O(N__80871),
            .I(N__80851));
    Span4Mux_v I__18753 (
            .O(N__80868),
            .I(N__80848));
    CEMux I__18752 (
            .O(N__80867),
            .I(N__80845));
    InMux I__18751 (
            .O(N__80866),
            .I(N__80842));
    LocalMux I__18750 (
            .O(N__80863),
            .I(N__80839));
    CEMux I__18749 (
            .O(N__80862),
            .I(N__80836));
    InMux I__18748 (
            .O(N__80861),
            .I(N__80832));
    Span4Mux_v I__18747 (
            .O(N__80858),
            .I(N__80823));
    LocalMux I__18746 (
            .O(N__80855),
            .I(N__80820));
    CEMux I__18745 (
            .O(N__80854),
            .I(N__80817));
    LocalMux I__18744 (
            .O(N__80851),
            .I(N__80813));
    Span4Mux_v I__18743 (
            .O(N__80848),
            .I(N__80810));
    LocalMux I__18742 (
            .O(N__80845),
            .I(N__80807));
    LocalMux I__18741 (
            .O(N__80842),
            .I(N__80804));
    Span4Mux_h I__18740 (
            .O(N__80839),
            .I(N__80799));
    LocalMux I__18739 (
            .O(N__80836),
            .I(N__80799));
    CEMux I__18738 (
            .O(N__80835),
            .I(N__80796));
    LocalMux I__18737 (
            .O(N__80832),
            .I(N__80793));
    InMux I__18736 (
            .O(N__80831),
            .I(N__80790));
    InMux I__18735 (
            .O(N__80830),
            .I(N__80779));
    InMux I__18734 (
            .O(N__80829),
            .I(N__80779));
    InMux I__18733 (
            .O(N__80828),
            .I(N__80779));
    InMux I__18732 (
            .O(N__80827),
            .I(N__80779));
    InMux I__18731 (
            .O(N__80826),
            .I(N__80779));
    Span4Mux_h I__18730 (
            .O(N__80823),
            .I(N__80774));
    Span4Mux_v I__18729 (
            .O(N__80820),
            .I(N__80774));
    LocalMux I__18728 (
            .O(N__80817),
            .I(N__80771));
    CEMux I__18727 (
            .O(N__80816),
            .I(N__80768));
    Sp12to4 I__18726 (
            .O(N__80813),
            .I(N__80765));
    Span4Mux_v I__18725 (
            .O(N__80810),
            .I(N__80762));
    Span4Mux_v I__18724 (
            .O(N__80807),
            .I(N__80759));
    Span4Mux_v I__18723 (
            .O(N__80804),
            .I(N__80756));
    Span4Mux_v I__18722 (
            .O(N__80799),
            .I(N__80753));
    LocalMux I__18721 (
            .O(N__80796),
            .I(N__80750));
    Span4Mux_h I__18720 (
            .O(N__80793),
            .I(N__80743));
    LocalMux I__18719 (
            .O(N__80790),
            .I(N__80743));
    LocalMux I__18718 (
            .O(N__80779),
            .I(N__80743));
    Span4Mux_h I__18717 (
            .O(N__80774),
            .I(N__80736));
    Span4Mux_h I__18716 (
            .O(N__80771),
            .I(N__80736));
    LocalMux I__18715 (
            .O(N__80768),
            .I(N__80736));
    Span12Mux_v I__18714 (
            .O(N__80765),
            .I(N__80725));
    Span4Mux_h I__18713 (
            .O(N__80762),
            .I(N__80720));
    Span4Mux_h I__18712 (
            .O(N__80759),
            .I(N__80720));
    Span4Mux_h I__18711 (
            .O(N__80756),
            .I(N__80717));
    Span4Mux_h I__18710 (
            .O(N__80753),
            .I(N__80714));
    Span4Mux_v I__18709 (
            .O(N__80750),
            .I(N__80707));
    Span4Mux_v I__18708 (
            .O(N__80743),
            .I(N__80707));
    Span4Mux_v I__18707 (
            .O(N__80736),
            .I(N__80707));
    InMux I__18706 (
            .O(N__80735),
            .I(N__80698));
    InMux I__18705 (
            .O(N__80734),
            .I(N__80698));
    InMux I__18704 (
            .O(N__80733),
            .I(N__80698));
    InMux I__18703 (
            .O(N__80732),
            .I(N__80698));
    InMux I__18702 (
            .O(N__80731),
            .I(N__80693));
    InMux I__18701 (
            .O(N__80730),
            .I(N__80693));
    InMux I__18700 (
            .O(N__80729),
            .I(N__80690));
    InMux I__18699 (
            .O(N__80728),
            .I(N__80687));
    Odrv12 I__18698 (
            .O(N__80725),
            .I(t_rd_fifo_en_w));
    Odrv4 I__18697 (
            .O(N__80720),
            .I(t_rd_fifo_en_w));
    Odrv4 I__18696 (
            .O(N__80717),
            .I(t_rd_fifo_en_w));
    Odrv4 I__18695 (
            .O(N__80714),
            .I(t_rd_fifo_en_w));
    Odrv4 I__18694 (
            .O(N__80707),
            .I(t_rd_fifo_en_w));
    LocalMux I__18693 (
            .O(N__80698),
            .I(t_rd_fifo_en_w));
    LocalMux I__18692 (
            .O(N__80693),
            .I(t_rd_fifo_en_w));
    LocalMux I__18691 (
            .O(N__80690),
            .I(t_rd_fifo_en_w));
    LocalMux I__18690 (
            .O(N__80687),
            .I(t_rd_fifo_en_w));
    CascadeMux I__18689 (
            .O(N__80668),
            .I(n11339_cascade_));
    InMux I__18688 (
            .O(N__80665),
            .I(N__80662));
    LocalMux I__18687 (
            .O(N__80662),
            .I(N__80658));
    InMux I__18686 (
            .O(N__80661),
            .I(N__80655));
    Span4Mux_v I__18685 (
            .O(N__80658),
            .I(N__80650));
    LocalMux I__18684 (
            .O(N__80655),
            .I(N__80650));
    Span4Mux_v I__18683 (
            .O(N__80650),
            .I(N__80646));
    InMux I__18682 (
            .O(N__80649),
            .I(N__80643));
    Odrv4 I__18681 (
            .O(N__80646),
            .I(tx_uart_active_flag));
    LocalMux I__18680 (
            .O(N__80643),
            .I(tx_uart_active_flag));
    CascadeMux I__18679 (
            .O(N__80638),
            .I(N__80634));
    InMux I__18678 (
            .O(N__80637),
            .I(N__80631));
    InMux I__18677 (
            .O(N__80634),
            .I(N__80628));
    LocalMux I__18676 (
            .O(N__80631),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_8 ));
    LocalMux I__18675 (
            .O(N__80628),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_8 ));
    CascadeMux I__18674 (
            .O(N__80623),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13928_cascade_ ));
    CascadeMux I__18673 (
            .O(N__80620),
            .I(N__80616));
    InMux I__18672 (
            .O(N__80619),
            .I(N__80611));
    InMux I__18671 (
            .O(N__80616),
            .I(N__80611));
    LocalMux I__18670 (
            .O(N__80611),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_8 ));
    InMux I__18669 (
            .O(N__80608),
            .I(N__80595));
    InMux I__18668 (
            .O(N__80607),
            .I(N__80591));
    InMux I__18667 (
            .O(N__80606),
            .I(N__80586));
    InMux I__18666 (
            .O(N__80605),
            .I(N__80586));
    InMux I__18665 (
            .O(N__80604),
            .I(N__80583));
    InMux I__18664 (
            .O(N__80603),
            .I(N__80578));
    InMux I__18663 (
            .O(N__80602),
            .I(N__80572));
    InMux I__18662 (
            .O(N__80601),
            .I(N__80566));
    InMux I__18661 (
            .O(N__80600),
            .I(N__80563));
    InMux I__18660 (
            .O(N__80599),
            .I(N__80560));
    InMux I__18659 (
            .O(N__80598),
            .I(N__80557));
    LocalMux I__18658 (
            .O(N__80595),
            .I(N__80551));
    InMux I__18657 (
            .O(N__80594),
            .I(N__80548));
    LocalMux I__18656 (
            .O(N__80591),
            .I(N__80544));
    LocalMux I__18655 (
            .O(N__80586),
            .I(N__80539));
    LocalMux I__18654 (
            .O(N__80583),
            .I(N__80539));
    InMux I__18653 (
            .O(N__80582),
            .I(N__80534));
    InMux I__18652 (
            .O(N__80581),
            .I(N__80534));
    LocalMux I__18651 (
            .O(N__80578),
            .I(N__80531));
    InMux I__18650 (
            .O(N__80577),
            .I(N__80528));
    InMux I__18649 (
            .O(N__80576),
            .I(N__80522));
    InMux I__18648 (
            .O(N__80575),
            .I(N__80519));
    LocalMux I__18647 (
            .O(N__80572),
            .I(N__80516));
    InMux I__18646 (
            .O(N__80571),
            .I(N__80513));
    CascadeMux I__18645 (
            .O(N__80570),
            .I(N__80509));
    InMux I__18644 (
            .O(N__80569),
            .I(N__80504));
    LocalMux I__18643 (
            .O(N__80566),
            .I(N__80499));
    LocalMux I__18642 (
            .O(N__80563),
            .I(N__80499));
    LocalMux I__18641 (
            .O(N__80560),
            .I(N__80494));
    LocalMux I__18640 (
            .O(N__80557),
            .I(N__80494));
    InMux I__18639 (
            .O(N__80556),
            .I(N__80491));
    InMux I__18638 (
            .O(N__80555),
            .I(N__80486));
    InMux I__18637 (
            .O(N__80554),
            .I(N__80486));
    Span4Mux_h I__18636 (
            .O(N__80551),
            .I(N__80483));
    LocalMux I__18635 (
            .O(N__80548),
            .I(N__80480));
    InMux I__18634 (
            .O(N__80547),
            .I(N__80477));
    Span4Mux_v I__18633 (
            .O(N__80544),
            .I(N__80472));
    Span4Mux_h I__18632 (
            .O(N__80539),
            .I(N__80472));
    LocalMux I__18631 (
            .O(N__80534),
            .I(N__80464));
    Span4Mux_v I__18630 (
            .O(N__80531),
            .I(N__80464));
    LocalMux I__18629 (
            .O(N__80528),
            .I(N__80464));
    InMux I__18628 (
            .O(N__80527),
            .I(N__80457));
    InMux I__18627 (
            .O(N__80526),
            .I(N__80457));
    InMux I__18626 (
            .O(N__80525),
            .I(N__80457));
    LocalMux I__18625 (
            .O(N__80522),
            .I(N__80454));
    LocalMux I__18624 (
            .O(N__80519),
            .I(N__80451));
    Span4Mux_v I__18623 (
            .O(N__80516),
            .I(N__80446));
    LocalMux I__18622 (
            .O(N__80513),
            .I(N__80446));
    InMux I__18621 (
            .O(N__80512),
            .I(N__80440));
    InMux I__18620 (
            .O(N__80509),
            .I(N__80440));
    InMux I__18619 (
            .O(N__80508),
            .I(N__80437));
    InMux I__18618 (
            .O(N__80507),
            .I(N__80434));
    LocalMux I__18617 (
            .O(N__80504),
            .I(N__80431));
    Span4Mux_v I__18616 (
            .O(N__80499),
            .I(N__80426));
    Span4Mux_v I__18615 (
            .O(N__80494),
            .I(N__80426));
    LocalMux I__18614 (
            .O(N__80491),
            .I(N__80417));
    LocalMux I__18613 (
            .O(N__80486),
            .I(N__80417));
    Span4Mux_v I__18612 (
            .O(N__80483),
            .I(N__80417));
    Span4Mux_h I__18611 (
            .O(N__80480),
            .I(N__80417));
    LocalMux I__18610 (
            .O(N__80477),
            .I(N__80412));
    Span4Mux_h I__18609 (
            .O(N__80472),
            .I(N__80412));
    InMux I__18608 (
            .O(N__80471),
            .I(N__80409));
    Span4Mux_h I__18607 (
            .O(N__80464),
            .I(N__80406));
    LocalMux I__18606 (
            .O(N__80457),
            .I(N__80403));
    Span12Mux_h I__18605 (
            .O(N__80454),
            .I(N__80398));
    Span12Mux_v I__18604 (
            .O(N__80451),
            .I(N__80398));
    Sp12to4 I__18603 (
            .O(N__80446),
            .I(N__80395));
    InMux I__18602 (
            .O(N__80445),
            .I(N__80392));
    LocalMux I__18601 (
            .O(N__80440),
            .I(N__80389));
    LocalMux I__18600 (
            .O(N__80437),
            .I(N__80382));
    LocalMux I__18599 (
            .O(N__80434),
            .I(N__80382));
    Span4Mux_h I__18598 (
            .O(N__80431),
            .I(N__80382));
    Span4Mux_h I__18597 (
            .O(N__80426),
            .I(N__80377));
    Span4Mux_v I__18596 (
            .O(N__80417),
            .I(N__80377));
    Span4Mux_h I__18595 (
            .O(N__80412),
            .I(N__80374));
    LocalMux I__18594 (
            .O(N__80409),
            .I(N__80365));
    Sp12to4 I__18593 (
            .O(N__80406),
            .I(N__80365));
    Span12Mux_s7_v I__18592 (
            .O(N__80403),
            .I(N__80365));
    Span12Mux_h I__18591 (
            .O(N__80398),
            .I(N__80365));
    Span12Mux_v I__18590 (
            .O(N__80395),
            .I(N__80362));
    LocalMux I__18589 (
            .O(N__80392),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n42 ));
    Odrv12 I__18588 (
            .O(N__80389),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n42 ));
    Odrv4 I__18587 (
            .O(N__80382),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n42 ));
    Odrv4 I__18586 (
            .O(N__80377),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n42 ));
    Odrv4 I__18585 (
            .O(N__80374),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n42 ));
    Odrv12 I__18584 (
            .O(N__80365),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n42 ));
    Odrv12 I__18583 (
            .O(N__80362),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n42 ));
    CascadeMux I__18582 (
            .O(N__80347),
            .I(N__80343));
    InMux I__18581 (
            .O(N__80346),
            .I(N__80338));
    InMux I__18580 (
            .O(N__80343),
            .I(N__80338));
    LocalMux I__18579 (
            .O(N__80338),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_8 ));
    CascadeMux I__18578 (
            .O(N__80335),
            .I(N__80331));
    InMux I__18577 (
            .O(N__80334),
            .I(N__80326));
    InMux I__18576 (
            .O(N__80331),
            .I(N__80326));
    LocalMux I__18575 (
            .O(N__80326),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_8 ));
    InMux I__18574 (
            .O(N__80323),
            .I(N__80314));
    InMux I__18573 (
            .O(N__80322),
            .I(N__80303));
    InMux I__18572 (
            .O(N__80321),
            .I(N__80303));
    InMux I__18571 (
            .O(N__80320),
            .I(N__80303));
    InMux I__18570 (
            .O(N__80319),
            .I(N__80294));
    InMux I__18569 (
            .O(N__80318),
            .I(N__80290));
    InMux I__18568 (
            .O(N__80317),
            .I(N__80284));
    LocalMux I__18567 (
            .O(N__80314),
            .I(N__80280));
    InMux I__18566 (
            .O(N__80313),
            .I(N__80277));
    InMux I__18565 (
            .O(N__80312),
            .I(N__80274));
    InMux I__18564 (
            .O(N__80311),
            .I(N__80269));
    InMux I__18563 (
            .O(N__80310),
            .I(N__80269));
    LocalMux I__18562 (
            .O(N__80303),
            .I(N__80263));
    InMux I__18561 (
            .O(N__80302),
            .I(N__80260));
    InMux I__18560 (
            .O(N__80301),
            .I(N__80255));
    InMux I__18559 (
            .O(N__80300),
            .I(N__80255));
    InMux I__18558 (
            .O(N__80299),
            .I(N__80252));
    InMux I__18557 (
            .O(N__80298),
            .I(N__80249));
    InMux I__18556 (
            .O(N__80297),
            .I(N__80245));
    LocalMux I__18555 (
            .O(N__80294),
            .I(N__80242));
    InMux I__18554 (
            .O(N__80293),
            .I(N__80239));
    LocalMux I__18553 (
            .O(N__80290),
            .I(N__80236));
    InMux I__18552 (
            .O(N__80289),
            .I(N__80233));
    InMux I__18551 (
            .O(N__80288),
            .I(N__80227));
    InMux I__18550 (
            .O(N__80287),
            .I(N__80227));
    LocalMux I__18549 (
            .O(N__80284),
            .I(N__80224));
    InMux I__18548 (
            .O(N__80283),
            .I(N__80221));
    Span4Mux_v I__18547 (
            .O(N__80280),
            .I(N__80216));
    LocalMux I__18546 (
            .O(N__80277),
            .I(N__80216));
    LocalMux I__18545 (
            .O(N__80274),
            .I(N__80210));
    LocalMux I__18544 (
            .O(N__80269),
            .I(N__80210));
    InMux I__18543 (
            .O(N__80268),
            .I(N__80207));
    InMux I__18542 (
            .O(N__80267),
            .I(N__80202));
    InMux I__18541 (
            .O(N__80266),
            .I(N__80202));
    Span4Mux_h I__18540 (
            .O(N__80263),
            .I(N__80198));
    LocalMux I__18539 (
            .O(N__80260),
            .I(N__80195));
    LocalMux I__18538 (
            .O(N__80255),
            .I(N__80192));
    LocalMux I__18537 (
            .O(N__80252),
            .I(N__80189));
    LocalMux I__18536 (
            .O(N__80249),
            .I(N__80186));
    InMux I__18535 (
            .O(N__80248),
            .I(N__80183));
    LocalMux I__18534 (
            .O(N__80245),
            .I(N__80176));
    Span4Mux_v I__18533 (
            .O(N__80242),
            .I(N__80176));
    LocalMux I__18532 (
            .O(N__80239),
            .I(N__80176));
    Span4Mux_h I__18531 (
            .O(N__80236),
            .I(N__80171));
    LocalMux I__18530 (
            .O(N__80233),
            .I(N__80171));
    InMux I__18529 (
            .O(N__80232),
            .I(N__80168));
    LocalMux I__18528 (
            .O(N__80227),
            .I(N__80162));
    Span4Mux_v I__18527 (
            .O(N__80224),
            .I(N__80157));
    LocalMux I__18526 (
            .O(N__80221),
            .I(N__80157));
    Span4Mux_v I__18525 (
            .O(N__80216),
            .I(N__80154));
    InMux I__18524 (
            .O(N__80215),
            .I(N__80151));
    Span4Mux_v I__18523 (
            .O(N__80210),
            .I(N__80148));
    LocalMux I__18522 (
            .O(N__80207),
            .I(N__80145));
    LocalMux I__18521 (
            .O(N__80202),
            .I(N__80142));
    InMux I__18520 (
            .O(N__80201),
            .I(N__80139));
    Span4Mux_h I__18519 (
            .O(N__80198),
            .I(N__80134));
    Span4Mux_v I__18518 (
            .O(N__80195),
            .I(N__80134));
    Span4Mux_h I__18517 (
            .O(N__80192),
            .I(N__80131));
    Span4Mux_v I__18516 (
            .O(N__80189),
            .I(N__80124));
    Span4Mux_h I__18515 (
            .O(N__80186),
            .I(N__80124));
    LocalMux I__18514 (
            .O(N__80183),
            .I(N__80124));
    Span4Mux_h I__18513 (
            .O(N__80176),
            .I(N__80121));
    Span4Mux_h I__18512 (
            .O(N__80171),
            .I(N__80116));
    LocalMux I__18511 (
            .O(N__80168),
            .I(N__80116));
    InMux I__18510 (
            .O(N__80167),
            .I(N__80113));
    InMux I__18509 (
            .O(N__80166),
            .I(N__80108));
    InMux I__18508 (
            .O(N__80165),
            .I(N__80108));
    Span4Mux_v I__18507 (
            .O(N__80162),
            .I(N__80105));
    Span4Mux_v I__18506 (
            .O(N__80157),
            .I(N__80102));
    Span4Mux_h I__18505 (
            .O(N__80154),
            .I(N__80097));
    LocalMux I__18504 (
            .O(N__80151),
            .I(N__80097));
    Span4Mux_h I__18503 (
            .O(N__80148),
            .I(N__80090));
    Span4Mux_v I__18502 (
            .O(N__80145),
            .I(N__80090));
    Span4Mux_v I__18501 (
            .O(N__80142),
            .I(N__80090));
    LocalMux I__18500 (
            .O(N__80139),
            .I(N__80087));
    Span4Mux_v I__18499 (
            .O(N__80134),
            .I(N__80084));
    Span4Mux_h I__18498 (
            .O(N__80131),
            .I(N__80079));
    Span4Mux_v I__18497 (
            .O(N__80124),
            .I(N__80079));
    Span4Mux_v I__18496 (
            .O(N__80121),
            .I(N__80074));
    Span4Mux_h I__18495 (
            .O(N__80116),
            .I(N__80074));
    LocalMux I__18494 (
            .O(N__80113),
            .I(N__80071));
    LocalMux I__18493 (
            .O(N__80108),
            .I(N__80068));
    Span4Mux_v I__18492 (
            .O(N__80105),
            .I(N__80061));
    Span4Mux_h I__18491 (
            .O(N__80102),
            .I(N__80061));
    Span4Mux_h I__18490 (
            .O(N__80097),
            .I(N__80061));
    Span4Mux_h I__18489 (
            .O(N__80090),
            .I(N__80056));
    Span4Mux_v I__18488 (
            .O(N__80087),
            .I(N__80056));
    Odrv4 I__18487 (
            .O(N__80084),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n40 ));
    Odrv4 I__18486 (
            .O(N__80079),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n40 ));
    Odrv4 I__18485 (
            .O(N__80074),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n40 ));
    Odrv12 I__18484 (
            .O(N__80071),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n40 ));
    Odrv12 I__18483 (
            .O(N__80068),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n40 ));
    Odrv4 I__18482 (
            .O(N__80061),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n40 ));
    Odrv4 I__18481 (
            .O(N__80056),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n40 ));
    InMux I__18480 (
            .O(N__80041),
            .I(N__80038));
    LocalMux I__18479 (
            .O(N__80038),
            .I(N__80035));
    Odrv4 I__18478 (
            .O(N__80035),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11718 ));
    InMux I__18477 (
            .O(N__80032),
            .I(N__80029));
    LocalMux I__18476 (
            .O(N__80029),
            .I(N__80026));
    Odrv12 I__18475 (
            .O(N__80026),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11709 ));
    CascadeMux I__18474 (
            .O(N__80023),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13136_cascade_ ));
    InMux I__18473 (
            .O(N__80020),
            .I(N__80017));
    LocalMux I__18472 (
            .O(N__80017),
            .I(N__80014));
    Span4Mux_v I__18471 (
            .O(N__80014),
            .I(N__80011));
    Odrv4 I__18470 (
            .O(N__80011),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11691 ));
    CascadeMux I__18469 (
            .O(N__80008),
            .I(N__80004));
    InMux I__18468 (
            .O(N__80007),
            .I(N__79999));
    InMux I__18467 (
            .O(N__80004),
            .I(N__79999));
    LocalMux I__18466 (
            .O(N__79999),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_6 ));
    InMux I__18465 (
            .O(N__79996),
            .I(N__79991));
    InMux I__18464 (
            .O(N__79995),
            .I(N__79986));
    InMux I__18463 (
            .O(N__79994),
            .I(N__79983));
    LocalMux I__18462 (
            .O(N__79991),
            .I(N__79978));
    InMux I__18461 (
            .O(N__79990),
            .I(N__79975));
    InMux I__18460 (
            .O(N__79989),
            .I(N__79971));
    LocalMux I__18459 (
            .O(N__79986),
            .I(N__79964));
    LocalMux I__18458 (
            .O(N__79983),
            .I(N__79961));
    InMux I__18457 (
            .O(N__79982),
            .I(N__79958));
    InMux I__18456 (
            .O(N__79981),
            .I(N__79955));
    Span4Mux_h I__18455 (
            .O(N__79978),
            .I(N__79950));
    LocalMux I__18454 (
            .O(N__79975),
            .I(N__79950));
    InMux I__18453 (
            .O(N__79974),
            .I(N__79947));
    LocalMux I__18452 (
            .O(N__79971),
            .I(N__79943));
    InMux I__18451 (
            .O(N__79970),
            .I(N__79940));
    InMux I__18450 (
            .O(N__79969),
            .I(N__79937));
    InMux I__18449 (
            .O(N__79968),
            .I(N__79932));
    InMux I__18448 (
            .O(N__79967),
            .I(N__79929));
    Span4Mux_h I__18447 (
            .O(N__79964),
            .I(N__79926));
    Span4Mux_v I__18446 (
            .O(N__79961),
            .I(N__79923));
    LocalMux I__18445 (
            .O(N__79958),
            .I(N__79920));
    LocalMux I__18444 (
            .O(N__79955),
            .I(N__79917));
    Span4Mux_v I__18443 (
            .O(N__79950),
            .I(N__79912));
    LocalMux I__18442 (
            .O(N__79947),
            .I(N__79912));
    InMux I__18441 (
            .O(N__79946),
            .I(N__79908));
    Span4Mux_h I__18440 (
            .O(N__79943),
            .I(N__79905));
    LocalMux I__18439 (
            .O(N__79940),
            .I(N__79900));
    LocalMux I__18438 (
            .O(N__79937),
            .I(N__79900));
    InMux I__18437 (
            .O(N__79936),
            .I(N__79897));
    InMux I__18436 (
            .O(N__79935),
            .I(N__79894));
    LocalMux I__18435 (
            .O(N__79932),
            .I(N__79891));
    LocalMux I__18434 (
            .O(N__79929),
            .I(N__79888));
    Span4Mux_v I__18433 (
            .O(N__79926),
            .I(N__79885));
    Sp12to4 I__18432 (
            .O(N__79923),
            .I(N__79882));
    Span4Mux_v I__18431 (
            .O(N__79920),
            .I(N__79879));
    Span4Mux_v I__18430 (
            .O(N__79917),
            .I(N__79874));
    Span4Mux_v I__18429 (
            .O(N__79912),
            .I(N__79874));
    InMux I__18428 (
            .O(N__79911),
            .I(N__79871));
    LocalMux I__18427 (
            .O(N__79908),
            .I(N__79866));
    Span4Mux_h I__18426 (
            .O(N__79905),
            .I(N__79866));
    Sp12to4 I__18425 (
            .O(N__79900),
            .I(N__79855));
    LocalMux I__18424 (
            .O(N__79897),
            .I(N__79855));
    LocalMux I__18423 (
            .O(N__79894),
            .I(N__79855));
    Span12Mux_v I__18422 (
            .O(N__79891),
            .I(N__79855));
    Span12Mux_v I__18421 (
            .O(N__79888),
            .I(N__79855));
    Span4Mux_h I__18420 (
            .O(N__79885),
            .I(N__79852));
    Span12Mux_h I__18419 (
            .O(N__79882),
            .I(N__79845));
    Sp12to4 I__18418 (
            .O(N__79879),
            .I(N__79845));
    Sp12to4 I__18417 (
            .O(N__79874),
            .I(N__79845));
    LocalMux I__18416 (
            .O(N__79871),
            .I(n7_adj_1183));
    Odrv4 I__18415 (
            .O(N__79866),
            .I(n7_adj_1183));
    Odrv12 I__18414 (
            .O(N__79855),
            .I(n7_adj_1183));
    Odrv4 I__18413 (
            .O(N__79852),
            .I(n7_adj_1183));
    Odrv12 I__18412 (
            .O(N__79845),
            .I(n7_adj_1183));
    InMux I__18411 (
            .O(N__79834),
            .I(N__79828));
    InMux I__18410 (
            .O(N__79833),
            .I(N__79828));
    LocalMux I__18409 (
            .O(N__79828),
            .I(REG_mem_58_8));
    CascadeMux I__18408 (
            .O(N__79825),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13448_cascade_ ));
    CascadeMux I__18407 (
            .O(N__79822),
            .I(N__79818));
    InMux I__18406 (
            .O(N__79821),
            .I(N__79813));
    InMux I__18405 (
            .O(N__79818),
            .I(N__79813));
    LocalMux I__18404 (
            .O(N__79813),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_8 ));
    CascadeMux I__18403 (
            .O(N__79810),
            .I(N__79806));
    InMux I__18402 (
            .O(N__79809),
            .I(N__79801));
    InMux I__18401 (
            .O(N__79806),
            .I(N__79801));
    LocalMux I__18400 (
            .O(N__79801),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_8 ));
    CascadeMux I__18399 (
            .O(N__79798),
            .I(N__79789));
    InMux I__18398 (
            .O(N__79797),
            .I(N__79780));
    InMux I__18397 (
            .O(N__79796),
            .I(N__79780));
    InMux I__18396 (
            .O(N__79795),
            .I(N__79777));
    InMux I__18395 (
            .O(N__79794),
            .I(N__79772));
    InMux I__18394 (
            .O(N__79793),
            .I(N__79772));
    InMux I__18393 (
            .O(N__79792),
            .I(N__79767));
    InMux I__18392 (
            .O(N__79789),
            .I(N__79764));
    InMux I__18391 (
            .O(N__79788),
            .I(N__79761));
    InMux I__18390 (
            .O(N__79787),
            .I(N__79756));
    InMux I__18389 (
            .O(N__79786),
            .I(N__79751));
    InMux I__18388 (
            .O(N__79785),
            .I(N__79747));
    LocalMux I__18387 (
            .O(N__79780),
            .I(N__79736));
    LocalMux I__18386 (
            .O(N__79777),
            .I(N__79733));
    LocalMux I__18385 (
            .O(N__79772),
            .I(N__79730));
    InMux I__18384 (
            .O(N__79771),
            .I(N__79725));
    InMux I__18383 (
            .O(N__79770),
            .I(N__79725));
    LocalMux I__18382 (
            .O(N__79767),
            .I(N__79720));
    LocalMux I__18381 (
            .O(N__79764),
            .I(N__79720));
    LocalMux I__18380 (
            .O(N__79761),
            .I(N__79717));
    InMux I__18379 (
            .O(N__79760),
            .I(N__79714));
    InMux I__18378 (
            .O(N__79759),
            .I(N__79711));
    LocalMux I__18377 (
            .O(N__79756),
            .I(N__79708));
    InMux I__18376 (
            .O(N__79755),
            .I(N__79703));
    InMux I__18375 (
            .O(N__79754),
            .I(N__79703));
    LocalMux I__18374 (
            .O(N__79751),
            .I(N__79699));
    InMux I__18373 (
            .O(N__79750),
            .I(N__79696));
    LocalMux I__18372 (
            .O(N__79747),
            .I(N__79693));
    InMux I__18371 (
            .O(N__79746),
            .I(N__79690));
    InMux I__18370 (
            .O(N__79745),
            .I(N__79687));
    InMux I__18369 (
            .O(N__79744),
            .I(N__79684));
    InMux I__18368 (
            .O(N__79743),
            .I(N__79681));
    InMux I__18367 (
            .O(N__79742),
            .I(N__79678));
    InMux I__18366 (
            .O(N__79741),
            .I(N__79675));
    InMux I__18365 (
            .O(N__79740),
            .I(N__79670));
    InMux I__18364 (
            .O(N__79739),
            .I(N__79670));
    Span4Mux_v I__18363 (
            .O(N__79736),
            .I(N__79665));
    Span4Mux_h I__18362 (
            .O(N__79733),
            .I(N__79665));
    Span4Mux_v I__18361 (
            .O(N__79730),
            .I(N__79662));
    LocalMux I__18360 (
            .O(N__79725),
            .I(N__79655));
    Span4Mux_v I__18359 (
            .O(N__79720),
            .I(N__79652));
    Span4Mux_v I__18358 (
            .O(N__79717),
            .I(N__79649));
    LocalMux I__18357 (
            .O(N__79714),
            .I(N__79646));
    LocalMux I__18356 (
            .O(N__79711),
            .I(N__79643));
    Span4Mux_v I__18355 (
            .O(N__79708),
            .I(N__79638));
    LocalMux I__18354 (
            .O(N__79703),
            .I(N__79638));
    InMux I__18353 (
            .O(N__79702),
            .I(N__79634));
    Span4Mux_v I__18352 (
            .O(N__79699),
            .I(N__79631));
    LocalMux I__18351 (
            .O(N__79696),
            .I(N__79628));
    Span4Mux_v I__18350 (
            .O(N__79693),
            .I(N__79625));
    LocalMux I__18349 (
            .O(N__79690),
            .I(N__79622));
    LocalMux I__18348 (
            .O(N__79687),
            .I(N__79619));
    LocalMux I__18347 (
            .O(N__79684),
            .I(N__79616));
    LocalMux I__18346 (
            .O(N__79681),
            .I(N__79613));
    LocalMux I__18345 (
            .O(N__79678),
            .I(N__79608));
    LocalMux I__18344 (
            .O(N__79675),
            .I(N__79608));
    LocalMux I__18343 (
            .O(N__79670),
            .I(N__79605));
    Span4Mux_h I__18342 (
            .O(N__79665),
            .I(N__79602));
    Sp12to4 I__18341 (
            .O(N__79662),
            .I(N__79599));
    InMux I__18340 (
            .O(N__79661),
            .I(N__79596));
    InMux I__18339 (
            .O(N__79660),
            .I(N__79593));
    InMux I__18338 (
            .O(N__79659),
            .I(N__79590));
    InMux I__18337 (
            .O(N__79658),
            .I(N__79587));
    Span4Mux_v I__18336 (
            .O(N__79655),
            .I(N__79584));
    Span4Mux_h I__18335 (
            .O(N__79652),
            .I(N__79579));
    Span4Mux_v I__18334 (
            .O(N__79649),
            .I(N__79579));
    Sp12to4 I__18333 (
            .O(N__79646),
            .I(N__79576));
    Span4Mux_v I__18332 (
            .O(N__79643),
            .I(N__79571));
    Span4Mux_v I__18331 (
            .O(N__79638),
            .I(N__79571));
    InMux I__18330 (
            .O(N__79637),
            .I(N__79568));
    LocalMux I__18329 (
            .O(N__79634),
            .I(N__79565));
    Span4Mux_h I__18328 (
            .O(N__79631),
            .I(N__79560));
    Span4Mux_v I__18327 (
            .O(N__79628),
            .I(N__79560));
    Span4Mux_h I__18326 (
            .O(N__79625),
            .I(N__79557));
    Span4Mux_h I__18325 (
            .O(N__79622),
            .I(N__79554));
    Span4Mux_h I__18324 (
            .O(N__79619),
            .I(N__79549));
    Span4Mux_h I__18323 (
            .O(N__79616),
            .I(N__79549));
    Span4Mux_v I__18322 (
            .O(N__79613),
            .I(N__79542));
    Span4Mux_h I__18321 (
            .O(N__79608),
            .I(N__79542));
    Span4Mux_v I__18320 (
            .O(N__79605),
            .I(N__79542));
    Sp12to4 I__18319 (
            .O(N__79602),
            .I(N__79535));
    Span12Mux_h I__18318 (
            .O(N__79599),
            .I(N__79535));
    LocalMux I__18317 (
            .O(N__79596),
            .I(N__79535));
    LocalMux I__18316 (
            .O(N__79593),
            .I(N__79520));
    LocalMux I__18315 (
            .O(N__79590),
            .I(N__79520));
    LocalMux I__18314 (
            .O(N__79587),
            .I(N__79520));
    Sp12to4 I__18313 (
            .O(N__79584),
            .I(N__79520));
    Sp12to4 I__18312 (
            .O(N__79579),
            .I(N__79520));
    Span12Mux_v I__18311 (
            .O(N__79576),
            .I(N__79520));
    Sp12to4 I__18310 (
            .O(N__79571),
            .I(N__79520));
    LocalMux I__18309 (
            .O(N__79568),
            .I(N__79515));
    Span4Mux_v I__18308 (
            .O(N__79565),
            .I(N__79515));
    Span4Mux_h I__18307 (
            .O(N__79560),
            .I(N__79510));
    Span4Mux_h I__18306 (
            .O(N__79557),
            .I(N__79510));
    Span4Mux_v I__18305 (
            .O(N__79554),
            .I(N__79503));
    Span4Mux_h I__18304 (
            .O(N__79549),
            .I(N__79503));
    Span4Mux_h I__18303 (
            .O(N__79542),
            .I(N__79503));
    Span12Mux_s11_v I__18302 (
            .O(N__79535),
            .I(N__79498));
    Span12Mux_h I__18301 (
            .O(N__79520),
            .I(N__79498));
    Odrv4 I__18300 (
            .O(N__79515),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n59 ));
    Odrv4 I__18299 (
            .O(N__79510),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n59 ));
    Odrv4 I__18298 (
            .O(N__79503),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n59 ));
    Odrv12 I__18297 (
            .O(N__79498),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n59 ));
    CascadeMux I__18296 (
            .O(N__79489),
            .I(N__79485));
    CascadeMux I__18295 (
            .O(N__79488),
            .I(N__79482));
    InMux I__18294 (
            .O(N__79485),
            .I(N__79477));
    InMux I__18293 (
            .O(N__79482),
            .I(N__79477));
    LocalMux I__18292 (
            .O(N__79477),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_8 ));
    InMux I__18291 (
            .O(N__79474),
            .I(N__79470));
    CascadeMux I__18290 (
            .O(N__79473),
            .I(N__79467));
    LocalMux I__18289 (
            .O(N__79470),
            .I(N__79464));
    InMux I__18288 (
            .O(N__79467),
            .I(N__79461));
    Odrv12 I__18287 (
            .O(N__79464),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_8 ));
    LocalMux I__18286 (
            .O(N__79461),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_8 ));
    CascadeMux I__18285 (
            .O(N__79456),
            .I(N__79453));
    InMux I__18284 (
            .O(N__79453),
            .I(N__79450));
    LocalMux I__18283 (
            .O(N__79450),
            .I(N__79447));
    Span4Mux_v I__18282 (
            .O(N__79447),
            .I(N__79444));
    Odrv4 I__18281 (
            .O(N__79444),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14042 ));
    CascadeMux I__18280 (
            .O(N__79441),
            .I(N__79437));
    InMux I__18279 (
            .O(N__79440),
            .I(N__79432));
    InMux I__18278 (
            .O(N__79437),
            .I(N__79432));
    LocalMux I__18277 (
            .O(N__79432),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_8 ));
    CascadeMux I__18276 (
            .O(N__79429),
            .I(N__79425));
    InMux I__18275 (
            .O(N__79428),
            .I(N__79422));
    InMux I__18274 (
            .O(N__79425),
            .I(N__79419));
    LocalMux I__18273 (
            .O(N__79422),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_6 ));
    LocalMux I__18272 (
            .O(N__79419),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_6 ));
    CascadeMux I__18271 (
            .O(N__79414),
            .I(N__79410));
    InMux I__18270 (
            .O(N__79413),
            .I(N__79405));
    InMux I__18269 (
            .O(N__79410),
            .I(N__79405));
    LocalMux I__18268 (
            .O(N__79405),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_6 ));
    CascadeMux I__18267 (
            .O(N__79402),
            .I(N__79398));
    InMux I__18266 (
            .O(N__79401),
            .I(N__79395));
    InMux I__18265 (
            .O(N__79398),
            .I(N__79392));
    LocalMux I__18264 (
            .O(N__79395),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_6 ));
    LocalMux I__18263 (
            .O(N__79392),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_6 ));
    InMux I__18262 (
            .O(N__79387),
            .I(N__79384));
    LocalMux I__18261 (
            .O(N__79384),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11789 ));
    InMux I__18260 (
            .O(N__79381),
            .I(N__79378));
    LocalMux I__18259 (
            .O(N__79378),
            .I(N__79375));
    Odrv12 I__18258 (
            .O(N__79375),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11788 ));
    CascadeMux I__18257 (
            .O(N__79372),
            .I(N__79368));
    InMux I__18256 (
            .O(N__79371),
            .I(N__79365));
    InMux I__18255 (
            .O(N__79368),
            .I(N__79362));
    LocalMux I__18254 (
            .O(N__79365),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_6 ));
    LocalMux I__18253 (
            .O(N__79362),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_6 ));
    InMux I__18252 (
            .O(N__79357),
            .I(N__79354));
    LocalMux I__18251 (
            .O(N__79354),
            .I(N__79351));
    Odrv12 I__18250 (
            .O(N__79351),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11785 ));
    InMux I__18249 (
            .O(N__79348),
            .I(N__79345));
    LocalMux I__18248 (
            .O(N__79345),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13526 ));
    CascadeMux I__18247 (
            .O(N__79342),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11786_cascade_ ));
    InMux I__18246 (
            .O(N__79339),
            .I(N__79336));
    LocalMux I__18245 (
            .O(N__79336),
            .I(N__79333));
    Odrv4 I__18244 (
            .O(N__79333),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13529 ));
    InMux I__18243 (
            .O(N__79330),
            .I(N__79326));
    InMux I__18242 (
            .O(N__79329),
            .I(N__79323));
    LocalMux I__18241 (
            .O(N__79326),
            .I(REG_mem_7_6));
    LocalMux I__18240 (
            .O(N__79323),
            .I(REG_mem_7_6));
    CascadeMux I__18239 (
            .O(N__79318),
            .I(N__79314));
    InMux I__18238 (
            .O(N__79317),
            .I(N__79309));
    InMux I__18237 (
            .O(N__79314),
            .I(N__79309));
    LocalMux I__18236 (
            .O(N__79309),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_6 ));
    InMux I__18235 (
            .O(N__79306),
            .I(N__79303));
    LocalMux I__18234 (
            .O(N__79303),
            .I(N__79300));
    Odrv12 I__18233 (
            .O(N__79300),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13007 ));
    InMux I__18232 (
            .O(N__79297),
            .I(N__79294));
    LocalMux I__18231 (
            .O(N__79294),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14342 ));
    InMux I__18230 (
            .O(N__79291),
            .I(N__79288));
    LocalMux I__18229 (
            .O(N__79288),
            .I(N__79285));
    Span12Mux_s8_h I__18228 (
            .O(N__79285),
            .I(N__79282));
    Odrv12 I__18227 (
            .O(N__79282),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12315 ));
    InMux I__18226 (
            .O(N__79279),
            .I(N__79276));
    LocalMux I__18225 (
            .O(N__79276),
            .I(N__79273));
    Odrv4 I__18224 (
            .O(N__79273),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11844 ));
    InMux I__18223 (
            .O(N__79270),
            .I(N__79267));
    LocalMux I__18222 (
            .O(N__79267),
            .I(N__79264));
    Span4Mux_h I__18221 (
            .O(N__79264),
            .I(N__79261));
    Span4Mux_h I__18220 (
            .O(N__79261),
            .I(N__79258));
    Odrv4 I__18219 (
            .O(N__79258),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11838 ));
    CascadeMux I__18218 (
            .O(N__79255),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13370_cascade_ ));
    CascadeMux I__18217 (
            .O(N__79252),
            .I(N__79249));
    InMux I__18216 (
            .O(N__79249),
            .I(N__79246));
    LocalMux I__18215 (
            .O(N__79246),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13373 ));
    InMux I__18214 (
            .O(N__79243),
            .I(N__79240));
    LocalMux I__18213 (
            .O(N__79240),
            .I(N__79237));
    Span4Mux_v I__18212 (
            .O(N__79237),
            .I(N__79234));
    Odrv4 I__18211 (
            .O(N__79234),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13775 ));
    InMux I__18210 (
            .O(N__79231),
            .I(N__79228));
    LocalMux I__18209 (
            .O(N__79228),
            .I(N__79225));
    Odrv4 I__18208 (
            .O(N__79225),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13781 ));
    CascadeMux I__18207 (
            .O(N__79222),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12002_cascade_ ));
    CascadeMux I__18206 (
            .O(N__79219),
            .I(N__79216));
    InMux I__18205 (
            .O(N__79216),
            .I(N__79213));
    LocalMux I__18204 (
            .O(N__79213),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12003 ));
    InMux I__18203 (
            .O(N__79210),
            .I(N__79207));
    LocalMux I__18202 (
            .O(N__79207),
            .I(N__79203));
    CascadeMux I__18201 (
            .O(N__79206),
            .I(N__79200));
    Span4Mux_v I__18200 (
            .O(N__79203),
            .I(N__79197));
    InMux I__18199 (
            .O(N__79200),
            .I(N__79194));
    Odrv4 I__18198 (
            .O(N__79197),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_6 ));
    LocalMux I__18197 (
            .O(N__79194),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_6 ));
    CascadeMux I__18196 (
            .O(N__79189),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13568_cascade_ ));
    InMux I__18195 (
            .O(N__79186),
            .I(N__79183));
    LocalMux I__18194 (
            .O(N__79183),
            .I(N__79179));
    CascadeMux I__18193 (
            .O(N__79182),
            .I(N__79176));
    Span4Mux_v I__18192 (
            .O(N__79179),
            .I(N__79173));
    InMux I__18191 (
            .O(N__79176),
            .I(N__79170));
    Odrv4 I__18190 (
            .O(N__79173),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_6 ));
    LocalMux I__18189 (
            .O(N__79170),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_6 ));
    InMux I__18188 (
            .O(N__79165),
            .I(N__79162));
    LocalMux I__18187 (
            .O(N__79162),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11835 ));
    InMux I__18186 (
            .O(N__79159),
            .I(N__79156));
    LocalMux I__18185 (
            .O(N__79156),
            .I(N__79153));
    Span4Mux_h I__18184 (
            .O(N__79153),
            .I(N__79149));
    InMux I__18183 (
            .O(N__79152),
            .I(N__79146));
    Odrv4 I__18182 (
            .O(N__79149),
            .I(REG_mem_6_6));
    LocalMux I__18181 (
            .O(N__79146),
            .I(REG_mem_6_6));
    InMux I__18180 (
            .O(N__79141),
            .I(N__79138));
    LocalMux I__18179 (
            .O(N__79138),
            .I(N__79135));
    Span4Mux_v I__18178 (
            .O(N__79135),
            .I(N__79131));
    InMux I__18177 (
            .O(N__79134),
            .I(N__79128));
    Odrv4 I__18176 (
            .O(N__79131),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_1 ));
    LocalMux I__18175 (
            .O(N__79128),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_1 ));
    InMux I__18174 (
            .O(N__79123),
            .I(N__79119));
    InMux I__18173 (
            .O(N__79122),
            .I(N__79116));
    LocalMux I__18172 (
            .O(N__79119),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1 ));
    LocalMux I__18171 (
            .O(N__79116),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1 ));
    InMux I__18170 (
            .O(N__79111),
            .I(N__79108));
    LocalMux I__18169 (
            .O(N__79108),
            .I(N__79104));
    CascadeMux I__18168 (
            .O(N__79107),
            .I(N__79101));
    Span4Mux_v I__18167 (
            .O(N__79104),
            .I(N__79098));
    InMux I__18166 (
            .O(N__79101),
            .I(N__79095));
    Odrv4 I__18165 (
            .O(N__79098),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_1 ));
    LocalMux I__18164 (
            .O(N__79095),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_1 ));
    CascadeMux I__18163 (
            .O(N__79090),
            .I(\tx_fifo.lscc_fifo_inst.n13538_cascade_ ));
    InMux I__18162 (
            .O(N__79087),
            .I(N__79083));
    InMux I__18161 (
            .O(N__79086),
            .I(N__79080));
    LocalMux I__18160 (
            .O(N__79083),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1 ));
    LocalMux I__18159 (
            .O(N__79080),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1 ));
    InMux I__18158 (
            .O(N__79075),
            .I(N__79072));
    LocalMux I__18157 (
            .O(N__79072),
            .I(mem_LUT_data_raw_r_1));
    InMux I__18156 (
            .O(N__79069),
            .I(N__79066));
    LocalMux I__18155 (
            .O(N__79066),
            .I(N__79063));
    Span4Mux_v I__18154 (
            .O(N__79063),
            .I(N__79059));
    InMux I__18153 (
            .O(N__79062),
            .I(N__79056));
    Odrv4 I__18152 (
            .O(N__79059),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_7 ));
    LocalMux I__18151 (
            .O(N__79056),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_7 ));
    CascadeMux I__18150 (
            .O(N__79051),
            .I(N__79048));
    InMux I__18149 (
            .O(N__79048),
            .I(N__79045));
    LocalMux I__18148 (
            .O(N__79045),
            .I(N__79041));
    CascadeMux I__18147 (
            .O(N__79044),
            .I(N__79038));
    Span4Mux_v I__18146 (
            .O(N__79041),
            .I(N__79035));
    InMux I__18145 (
            .O(N__79038),
            .I(N__79032));
    Odrv4 I__18144 (
            .O(N__79035),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7 ));
    LocalMux I__18143 (
            .O(N__79032),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7 ));
    CascadeMux I__18142 (
            .O(N__79027),
            .I(N__79021));
    CascadeMux I__18141 (
            .O(N__79026),
            .I(N__79018));
    CascadeMux I__18140 (
            .O(N__79025),
            .I(N__79015));
    CascadeMux I__18139 (
            .O(N__79024),
            .I(N__79011));
    InMux I__18138 (
            .O(N__79021),
            .I(N__79005));
    InMux I__18137 (
            .O(N__79018),
            .I(N__79000));
    InMux I__18136 (
            .O(N__79015),
            .I(N__79000));
    InMux I__18135 (
            .O(N__79014),
            .I(N__78997));
    InMux I__18134 (
            .O(N__79011),
            .I(N__78994));
    InMux I__18133 (
            .O(N__79010),
            .I(N__78989));
    InMux I__18132 (
            .O(N__79009),
            .I(N__78989));
    CascadeMux I__18131 (
            .O(N__79008),
            .I(N__78985));
    LocalMux I__18130 (
            .O(N__79005),
            .I(N__78981));
    LocalMux I__18129 (
            .O(N__79000),
            .I(N__78978));
    LocalMux I__18128 (
            .O(N__78997),
            .I(N__78973));
    LocalMux I__18127 (
            .O(N__78994),
            .I(N__78973));
    LocalMux I__18126 (
            .O(N__78989),
            .I(N__78970));
    InMux I__18125 (
            .O(N__78988),
            .I(N__78967));
    InMux I__18124 (
            .O(N__78985),
            .I(N__78964));
    CascadeMux I__18123 (
            .O(N__78984),
            .I(N__78957));
    Span4Mux_v I__18122 (
            .O(N__78981),
            .I(N__78951));
    Span4Mux_h I__18121 (
            .O(N__78978),
            .I(N__78951));
    Span4Mux_h I__18120 (
            .O(N__78973),
            .I(N__78942));
    Span4Mux_h I__18119 (
            .O(N__78970),
            .I(N__78942));
    LocalMux I__18118 (
            .O(N__78967),
            .I(N__78942));
    LocalMux I__18117 (
            .O(N__78964),
            .I(N__78942));
    InMux I__18116 (
            .O(N__78963),
            .I(N__78937));
    InMux I__18115 (
            .O(N__78962),
            .I(N__78937));
    InMux I__18114 (
            .O(N__78961),
            .I(N__78934));
    InMux I__18113 (
            .O(N__78960),
            .I(N__78931));
    InMux I__18112 (
            .O(N__78957),
            .I(N__78928));
    InMux I__18111 (
            .O(N__78956),
            .I(N__78925));
    Odrv4 I__18110 (
            .O(N__78951),
            .I(rd_addr_r_0));
    Odrv4 I__18109 (
            .O(N__78942),
            .I(rd_addr_r_0));
    LocalMux I__18108 (
            .O(N__78937),
            .I(rd_addr_r_0));
    LocalMux I__18107 (
            .O(N__78934),
            .I(rd_addr_r_0));
    LocalMux I__18106 (
            .O(N__78931),
            .I(rd_addr_r_0));
    LocalMux I__18105 (
            .O(N__78928),
            .I(rd_addr_r_0));
    LocalMux I__18104 (
            .O(N__78925),
            .I(rd_addr_r_0));
    InMux I__18103 (
            .O(N__78910),
            .I(N__78907));
    LocalMux I__18102 (
            .O(N__78907),
            .I(N__78904));
    Odrv4 I__18101 (
            .O(N__78904),
            .I(\tx_fifo.lscc_fifo_inst.n14234 ));
    InMux I__18100 (
            .O(N__78901),
            .I(N__78898));
    LocalMux I__18099 (
            .O(N__78898),
            .I(\tx_fifo.lscc_fifo_inst.n13556 ));
    CascadeMux I__18098 (
            .O(N__78895),
            .I(N__78892));
    InMux I__18097 (
            .O(N__78892),
            .I(N__78888));
    CascadeMux I__18096 (
            .O(N__78891),
            .I(N__78885));
    LocalMux I__18095 (
            .O(N__78888),
            .I(N__78882));
    InMux I__18094 (
            .O(N__78885),
            .I(N__78879));
    Odrv4 I__18093 (
            .O(N__78882),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_3 ));
    LocalMux I__18092 (
            .O(N__78879),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_3 ));
    InMux I__18091 (
            .O(N__78874),
            .I(N__78870));
    InMux I__18090 (
            .O(N__78873),
            .I(N__78867));
    LocalMux I__18089 (
            .O(N__78870),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3 ));
    LocalMux I__18088 (
            .O(N__78867),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3 ));
    InMux I__18087 (
            .O(N__78862),
            .I(N__78859));
    LocalMux I__18086 (
            .O(N__78859),
            .I(N__78856));
    Span4Mux_v I__18085 (
            .O(N__78856),
            .I(N__78853));
    Odrv4 I__18084 (
            .O(N__78853),
            .I(mem_LUT_data_raw_r_3));
    InMux I__18083 (
            .O(N__78850),
            .I(N__78846));
    CascadeMux I__18082 (
            .O(N__78849),
            .I(N__78843));
    LocalMux I__18081 (
            .O(N__78846),
            .I(N__78840));
    InMux I__18080 (
            .O(N__78843),
            .I(N__78837));
    Odrv4 I__18079 (
            .O(N__78840),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0 ));
    LocalMux I__18078 (
            .O(N__78837),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0 ));
    InMux I__18077 (
            .O(N__78832),
            .I(N__78829));
    LocalMux I__18076 (
            .O(N__78829),
            .I(N__78826));
    Span4Mux_h I__18075 (
            .O(N__78826),
            .I(N__78823));
    Odrv4 I__18074 (
            .O(N__78823),
            .I(\tx_fifo.lscc_fifo_inst.n13496 ));
    CascadeMux I__18073 (
            .O(N__78820),
            .I(N__78817));
    InMux I__18072 (
            .O(N__78817),
            .I(N__78814));
    LocalMux I__18071 (
            .O(N__78814),
            .I(N__78811));
    Span4Mux_v I__18070 (
            .O(N__78811),
            .I(N__78807));
    InMux I__18069 (
            .O(N__78810),
            .I(N__78804));
    Odrv4 I__18068 (
            .O(N__78807),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_0 ));
    LocalMux I__18067 (
            .O(N__78804),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_0 ));
    CascadeMux I__18066 (
            .O(N__78799),
            .I(N__78788));
    InMux I__18065 (
            .O(N__78798),
            .I(N__78781));
    InMux I__18064 (
            .O(N__78797),
            .I(N__78781));
    InMux I__18063 (
            .O(N__78796),
            .I(N__78781));
    InMux I__18062 (
            .O(N__78795),
            .I(N__78778));
    InMux I__18061 (
            .O(N__78794),
            .I(N__78775));
    InMux I__18060 (
            .O(N__78793),
            .I(N__78761));
    InMux I__18059 (
            .O(N__78792),
            .I(N__78761));
    InMux I__18058 (
            .O(N__78791),
            .I(N__78761));
    InMux I__18057 (
            .O(N__78788),
            .I(N__78758));
    LocalMux I__18056 (
            .O(N__78781),
            .I(N__78753));
    LocalMux I__18055 (
            .O(N__78778),
            .I(N__78753));
    LocalMux I__18054 (
            .O(N__78775),
            .I(N__78750));
    InMux I__18053 (
            .O(N__78774),
            .I(N__78747));
    InMux I__18052 (
            .O(N__78773),
            .I(N__78734));
    InMux I__18051 (
            .O(N__78772),
            .I(N__78734));
    InMux I__18050 (
            .O(N__78771),
            .I(N__78734));
    InMux I__18049 (
            .O(N__78770),
            .I(N__78734));
    InMux I__18048 (
            .O(N__78769),
            .I(N__78734));
    InMux I__18047 (
            .O(N__78768),
            .I(N__78734));
    LocalMux I__18046 (
            .O(N__78761),
            .I(N__78728));
    LocalMux I__18045 (
            .O(N__78758),
            .I(N__78725));
    Span4Mux_v I__18044 (
            .O(N__78753),
            .I(N__78716));
    Span4Mux_h I__18043 (
            .O(N__78750),
            .I(N__78716));
    LocalMux I__18042 (
            .O(N__78747),
            .I(N__78716));
    LocalMux I__18041 (
            .O(N__78734),
            .I(N__78716));
    InMux I__18040 (
            .O(N__78733),
            .I(N__78713));
    InMux I__18039 (
            .O(N__78732),
            .I(N__78710));
    CascadeMux I__18038 (
            .O(N__78731),
            .I(N__78706));
    Span4Mux_h I__18037 (
            .O(N__78728),
            .I(N__78701));
    Span4Mux_v I__18036 (
            .O(N__78725),
            .I(N__78696));
    Span4Mux_v I__18035 (
            .O(N__78716),
            .I(N__78696));
    LocalMux I__18034 (
            .O(N__78713),
            .I(N__78693));
    LocalMux I__18033 (
            .O(N__78710),
            .I(N__78690));
    InMux I__18032 (
            .O(N__78709),
            .I(N__78683));
    InMux I__18031 (
            .O(N__78706),
            .I(N__78683));
    InMux I__18030 (
            .O(N__78705),
            .I(N__78683));
    InMux I__18029 (
            .O(N__78704),
            .I(N__78680));
    Odrv4 I__18028 (
            .O(N__78701),
            .I(rd_addr_r_1));
    Odrv4 I__18027 (
            .O(N__78696),
            .I(rd_addr_r_1));
    Odrv12 I__18026 (
            .O(N__78693),
            .I(rd_addr_r_1));
    Odrv4 I__18025 (
            .O(N__78690),
            .I(rd_addr_r_1));
    LocalMux I__18024 (
            .O(N__78683),
            .I(rd_addr_r_1));
    LocalMux I__18023 (
            .O(N__78680),
            .I(rd_addr_r_1));
    InMux I__18022 (
            .O(N__78667),
            .I(N__78664));
    LocalMux I__18021 (
            .O(N__78664),
            .I(N__78661));
    Odrv4 I__18020 (
            .O(N__78661),
            .I(mem_LUT_data_raw_r_0));
    CEMux I__18019 (
            .O(N__78658),
            .I(N__78651));
    InMux I__18018 (
            .O(N__78657),
            .I(N__78648));
    CEMux I__18017 (
            .O(N__78656),
            .I(N__78645));
    CEMux I__18016 (
            .O(N__78655),
            .I(N__78642));
    CEMux I__18015 (
            .O(N__78654),
            .I(N__78639));
    LocalMux I__18014 (
            .O(N__78651),
            .I(N__78636));
    LocalMux I__18013 (
            .O(N__78648),
            .I(N__78630));
    LocalMux I__18012 (
            .O(N__78645),
            .I(N__78630));
    LocalMux I__18011 (
            .O(N__78642),
            .I(N__78625));
    LocalMux I__18010 (
            .O(N__78639),
            .I(N__78625));
    Span4Mux_v I__18009 (
            .O(N__78636),
            .I(N__78622));
    CEMux I__18008 (
            .O(N__78635),
            .I(N__78619));
    Span4Mux_v I__18007 (
            .O(N__78630),
            .I(N__78616));
    Span4Mux_v I__18006 (
            .O(N__78625),
            .I(N__78613));
    Sp12to4 I__18005 (
            .O(N__78622),
            .I(N__78608));
    LocalMux I__18004 (
            .O(N__78619),
            .I(N__78608));
    Odrv4 I__18003 (
            .O(N__78616),
            .I(rd_fifo_en_w));
    Odrv4 I__18002 (
            .O(N__78613),
            .I(rd_fifo_en_w));
    Odrv12 I__18001 (
            .O(N__78608),
            .I(rd_fifo_en_w));
    InMux I__18000 (
            .O(N__78601),
            .I(N__78598));
    LocalMux I__17999 (
            .O(N__78598),
            .I(N__78595));
    Span4Mux_v I__17998 (
            .O(N__78595),
            .I(N__78592));
    Odrv4 I__17997 (
            .O(N__78592),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13649 ));
    CascadeMux I__17996 (
            .O(N__78589),
            .I(N__78586));
    InMux I__17995 (
            .O(N__78586),
            .I(N__78583));
    LocalMux I__17994 (
            .O(N__78583),
            .I(N__78580));
    Odrv4 I__17993 (
            .O(N__78580),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13946 ));
    InMux I__17992 (
            .O(N__78577),
            .I(N__78574));
    LocalMux I__17991 (
            .O(N__78574),
            .I(N__78571));
    Odrv12 I__17990 (
            .O(N__78571),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13661 ));
    InMux I__17989 (
            .O(N__78568),
            .I(N__78565));
    LocalMux I__17988 (
            .O(N__78565),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13949 ));
    InMux I__17987 (
            .O(N__78562),
            .I(N__78559));
    LocalMux I__17986 (
            .O(N__78559),
            .I(N__78556));
    Span4Mux_v I__17985 (
            .O(N__78556),
            .I(N__78553));
    Sp12to4 I__17984 (
            .O(N__78553),
            .I(N__78550));
    Span12Mux_v I__17983 (
            .O(N__78550),
            .I(N__78547));
    Odrv12 I__17982 (
            .O(N__78547),
            .I(REG_out_raw_6));
    InMux I__17981 (
            .O(N__78544),
            .I(N__78538));
    InMux I__17980 (
            .O(N__78543),
            .I(N__78538));
    LocalMux I__17979 (
            .O(N__78538),
            .I(fifo_temp_output_0));
    InMux I__17978 (
            .O(N__78535),
            .I(N__78532));
    LocalMux I__17977 (
            .O(N__78532),
            .I(N__78528));
    InMux I__17976 (
            .O(N__78531),
            .I(N__78525));
    Odrv4 I__17975 (
            .O(N__78528),
            .I(r_Tx_Data_0));
    LocalMux I__17974 (
            .O(N__78525),
            .I(r_Tx_Data_0));
    InMux I__17973 (
            .O(N__78520),
            .I(N__78516));
    InMux I__17972 (
            .O(N__78519),
            .I(N__78513));
    LocalMux I__17971 (
            .O(N__78516),
            .I(fifo_temp_output_1));
    LocalMux I__17970 (
            .O(N__78513),
            .I(fifo_temp_output_1));
    InMux I__17969 (
            .O(N__78508),
            .I(N__78505));
    LocalMux I__17968 (
            .O(N__78505),
            .I(N__78501));
    InMux I__17967 (
            .O(N__78504),
            .I(N__78498));
    Odrv4 I__17966 (
            .O(N__78501),
            .I(r_Tx_Data_1));
    LocalMux I__17965 (
            .O(N__78498),
            .I(r_Tx_Data_1));
    InMux I__17964 (
            .O(N__78493),
            .I(N__78490));
    LocalMux I__17963 (
            .O(N__78490),
            .I(N__78487));
    Span4Mux_v I__17962 (
            .O(N__78487),
            .I(N__78484));
    Odrv4 I__17961 (
            .O(N__78484),
            .I(mem_LUT_data_raw_r_2));
    InMux I__17960 (
            .O(N__78481),
            .I(N__78477));
    InMux I__17959 (
            .O(N__78480),
            .I(N__78474));
    LocalMux I__17958 (
            .O(N__78477),
            .I(fifo_temp_output_2));
    LocalMux I__17957 (
            .O(N__78474),
            .I(fifo_temp_output_2));
    InMux I__17956 (
            .O(N__78469),
            .I(N__78466));
    LocalMux I__17955 (
            .O(N__78466),
            .I(N__78462));
    InMux I__17954 (
            .O(N__78465),
            .I(N__78459));
    Odrv12 I__17953 (
            .O(N__78462),
            .I(r_Tx_Data_2));
    LocalMux I__17952 (
            .O(N__78459),
            .I(r_Tx_Data_2));
    InMux I__17951 (
            .O(N__78454),
            .I(N__78436));
    InMux I__17950 (
            .O(N__78453),
            .I(N__78436));
    InMux I__17949 (
            .O(N__78452),
            .I(N__78436));
    InMux I__17948 (
            .O(N__78451),
            .I(N__78436));
    InMux I__17947 (
            .O(N__78450),
            .I(N__78436));
    InMux I__17946 (
            .O(N__78449),
            .I(N__78428));
    InMux I__17945 (
            .O(N__78448),
            .I(N__78428));
    InMux I__17944 (
            .O(N__78447),
            .I(N__78428));
    LocalMux I__17943 (
            .O(N__78436),
            .I(N__78421));
    InMux I__17942 (
            .O(N__78435),
            .I(N__78418));
    LocalMux I__17941 (
            .O(N__78428),
            .I(N__78415));
    InMux I__17940 (
            .O(N__78427),
            .I(N__78408));
    InMux I__17939 (
            .O(N__78426),
            .I(N__78408));
    InMux I__17938 (
            .O(N__78425),
            .I(N__78403));
    SRMux I__17937 (
            .O(N__78424),
            .I(N__78403));
    Span4Mux_v I__17936 (
            .O(N__78421),
            .I(N__78398));
    LocalMux I__17935 (
            .O(N__78418),
            .I(N__78398));
    Span4Mux_v I__17934 (
            .O(N__78415),
            .I(N__78395));
    InMux I__17933 (
            .O(N__78414),
            .I(N__78390));
    InMux I__17932 (
            .O(N__78413),
            .I(N__78390));
    LocalMux I__17931 (
            .O(N__78408),
            .I(N__78382));
    LocalMux I__17930 (
            .O(N__78403),
            .I(N__78382));
    Span4Mux_h I__17929 (
            .O(N__78398),
            .I(N__78379));
    Span4Mux_v I__17928 (
            .O(N__78395),
            .I(N__78374));
    LocalMux I__17927 (
            .O(N__78390),
            .I(N__78374));
    InMux I__17926 (
            .O(N__78389),
            .I(N__78369));
    InMux I__17925 (
            .O(N__78388),
            .I(N__78369));
    CascadeMux I__17924 (
            .O(N__78387),
            .I(N__78366));
    Span4Mux_v I__17923 (
            .O(N__78382),
            .I(N__78362));
    Span4Mux_v I__17922 (
            .O(N__78379),
            .I(N__78357));
    Span4Mux_h I__17921 (
            .O(N__78374),
            .I(N__78357));
    LocalMux I__17920 (
            .O(N__78369),
            .I(N__78354));
    InMux I__17919 (
            .O(N__78366),
            .I(N__78351));
    InMux I__17918 (
            .O(N__78365),
            .I(N__78348));
    Odrv4 I__17917 (
            .O(N__78362),
            .I(reset_all_w));
    Odrv4 I__17916 (
            .O(N__78357),
            .I(reset_all_w));
    Odrv12 I__17915 (
            .O(N__78354),
            .I(reset_all_w));
    LocalMux I__17914 (
            .O(N__78351),
            .I(reset_all_w));
    LocalMux I__17913 (
            .O(N__78348),
            .I(reset_all_w));
    CascadeMux I__17912 (
            .O(N__78337),
            .I(N__78328));
    CascadeMux I__17911 (
            .O(N__78336),
            .I(N__78325));
    CascadeMux I__17910 (
            .O(N__78335),
            .I(N__78322));
    CascadeMux I__17909 (
            .O(N__78334),
            .I(N__78319));
    CascadeMux I__17908 (
            .O(N__78333),
            .I(N__78315));
    CascadeMux I__17907 (
            .O(N__78332),
            .I(N__78312));
    CascadeMux I__17906 (
            .O(N__78331),
            .I(N__78309));
    InMux I__17905 (
            .O(N__78328),
            .I(N__78300));
    InMux I__17904 (
            .O(N__78325),
            .I(N__78300));
    InMux I__17903 (
            .O(N__78322),
            .I(N__78300));
    InMux I__17902 (
            .O(N__78319),
            .I(N__78300));
    CascadeMux I__17901 (
            .O(N__78318),
            .I(N__78297));
    InMux I__17900 (
            .O(N__78315),
            .I(N__78290));
    InMux I__17899 (
            .O(N__78312),
            .I(N__78290));
    InMux I__17898 (
            .O(N__78309),
            .I(N__78290));
    LocalMux I__17897 (
            .O(N__78300),
            .I(N__78287));
    InMux I__17896 (
            .O(N__78297),
            .I(N__78284));
    LocalMux I__17895 (
            .O(N__78290),
            .I(N__78281));
    Span4Mux_h I__17894 (
            .O(N__78287),
            .I(N__78276));
    LocalMux I__17893 (
            .O(N__78284),
            .I(N__78276));
    Odrv12 I__17892 (
            .O(N__78281),
            .I(n4249));
    Odrv4 I__17891 (
            .O(N__78276),
            .I(n4249));
    InMux I__17890 (
            .O(N__78271),
            .I(N__78267));
    InMux I__17889 (
            .O(N__78270),
            .I(N__78264));
    LocalMux I__17888 (
            .O(N__78267),
            .I(fifo_temp_output_3));
    LocalMux I__17887 (
            .O(N__78264),
            .I(fifo_temp_output_3));
    InMux I__17886 (
            .O(N__78259),
            .I(N__78256));
    LocalMux I__17885 (
            .O(N__78256),
            .I(\timing_controller_inst.n55 ));
    InMux I__17884 (
            .O(N__78253),
            .I(N__78250));
    LocalMux I__17883 (
            .O(N__78250),
            .I(\timing_controller_inst.n56 ));
    CascadeMux I__17882 (
            .O(N__78247),
            .I(N__78244));
    InMux I__17881 (
            .O(N__78244),
            .I(N__78241));
    LocalMux I__17880 (
            .O(N__78241),
            .I(\timing_controller_inst.n53 ));
    InMux I__17879 (
            .O(N__78238),
            .I(N__78235));
    LocalMux I__17878 (
            .O(N__78235),
            .I(\timing_controller_inst.n1740 ));
    InMux I__17877 (
            .O(N__78232),
            .I(N__78229));
    LocalMux I__17876 (
            .O(N__78229),
            .I(\timing_controller_inst.n1742 ));
    InMux I__17875 (
            .O(N__78226),
            .I(N__78223));
    LocalMux I__17874 (
            .O(N__78223),
            .I(\timing_controller_inst.n1739 ));
    InMux I__17873 (
            .O(N__78220),
            .I(N__78217));
    LocalMux I__17872 (
            .O(N__78217),
            .I(\timing_controller_inst.n1736 ));
    InMux I__17871 (
            .O(N__78214),
            .I(N__78211));
    LocalMux I__17870 (
            .O(N__78211),
            .I(\timing_controller_inst.n1754 ));
    CascadeMux I__17869 (
            .O(N__78208),
            .I(N__78205));
    InMux I__17868 (
            .O(N__78205),
            .I(N__78202));
    LocalMux I__17867 (
            .O(N__78202),
            .I(N__78199));
    Span4Mux_h I__17866 (
            .O(N__78199),
            .I(N__78196));
    Odrv4 I__17865 (
            .O(N__78196),
            .I(\timing_controller_inst.n1735 ));
    CascadeMux I__17864 (
            .O(N__78193),
            .I(N__78190));
    InMux I__17863 (
            .O(N__78190),
            .I(N__78187));
    LocalMux I__17862 (
            .O(N__78187),
            .I(N__78184));
    Span4Mux_h I__17861 (
            .O(N__78184),
            .I(N__78181));
    Odrv4 I__17860 (
            .O(N__78181),
            .I(\timing_controller_inst.n1734 ));
    InMux I__17859 (
            .O(N__78178),
            .I(N__78175));
    LocalMux I__17858 (
            .O(N__78175),
            .I(N__78172));
    Span4Mux_v I__17857 (
            .O(N__78172),
            .I(N__78169));
    Span4Mux_h I__17856 (
            .O(N__78169),
            .I(N__78165));
    InMux I__17855 (
            .O(N__78168),
            .I(N__78162));
    Odrv4 I__17854 (
            .O(N__78165),
            .I(r_Tx_Data_7));
    LocalMux I__17853 (
            .O(N__78162),
            .I(r_Tx_Data_7));
    InMux I__17852 (
            .O(N__78157),
            .I(N__78154));
    LocalMux I__17851 (
            .O(N__78154),
            .I(N__78150));
    InMux I__17850 (
            .O(N__78153),
            .I(N__78147));
    Odrv4 I__17849 (
            .O(N__78150),
            .I(r_Tx_Data_6));
    LocalMux I__17848 (
            .O(N__78147),
            .I(r_Tx_Data_6));
    InMux I__17847 (
            .O(N__78142),
            .I(N__78139));
    LocalMux I__17846 (
            .O(N__78139),
            .I(\pc_tx.n12140 ));
    InMux I__17845 (
            .O(N__78136),
            .I(N__78133));
    LocalMux I__17844 (
            .O(N__78133),
            .I(N__78130));
    Span4Mux_v I__17843 (
            .O(N__78130),
            .I(N__78123));
    InMux I__17842 (
            .O(N__78129),
            .I(N__78120));
    InMux I__17841 (
            .O(N__78128),
            .I(N__78115));
    InMux I__17840 (
            .O(N__78127),
            .I(N__78115));
    InMux I__17839 (
            .O(N__78126),
            .I(N__78112));
    Odrv4 I__17838 (
            .O(N__78123),
            .I(\bluejay_data_inst.n710 ));
    LocalMux I__17837 (
            .O(N__78120),
            .I(\bluejay_data_inst.n710 ));
    LocalMux I__17836 (
            .O(N__78115),
            .I(\bluejay_data_inst.n710 ));
    LocalMux I__17835 (
            .O(N__78112),
            .I(\bluejay_data_inst.n710 ));
    InMux I__17834 (
            .O(N__78103),
            .I(N__78100));
    LocalMux I__17833 (
            .O(N__78100),
            .I(N__78097));
    Span4Mux_v I__17832 (
            .O(N__78097),
            .I(N__78091));
    InMux I__17831 (
            .O(N__78096),
            .I(N__78084));
    InMux I__17830 (
            .O(N__78095),
            .I(N__78084));
    InMux I__17829 (
            .O(N__78094),
            .I(N__78084));
    Odrv4 I__17828 (
            .O(N__78091),
            .I(n718));
    LocalMux I__17827 (
            .O(N__78084),
            .I(n718));
    InMux I__17826 (
            .O(N__78079),
            .I(N__78076));
    LocalMux I__17825 (
            .O(N__78076),
            .I(N__78073));
    Span4Mux_v I__17824 (
            .O(N__78073),
            .I(N__78070));
    Span4Mux_h I__17823 (
            .O(N__78070),
            .I(N__78065));
    InMux I__17822 (
            .O(N__78069),
            .I(N__78060));
    InMux I__17821 (
            .O(N__78068),
            .I(N__78060));
    Odrv4 I__17820 (
            .O(N__78065),
            .I(\bluejay_data_inst.n715 ));
    LocalMux I__17819 (
            .O(N__78060),
            .I(\bluejay_data_inst.n715 ));
    InMux I__17818 (
            .O(N__78055),
            .I(N__78051));
    InMux I__17817 (
            .O(N__78054),
            .I(N__78048));
    LocalMux I__17816 (
            .O(N__78051),
            .I(N__78041));
    LocalMux I__17815 (
            .O(N__78048),
            .I(N__78041));
    InMux I__17814 (
            .O(N__78047),
            .I(N__78038));
    InMux I__17813 (
            .O(N__78046),
            .I(N__78035));
    Span4Mux_v I__17812 (
            .O(N__78041),
            .I(N__78027));
    LocalMux I__17811 (
            .O(N__78038),
            .I(N__78027));
    LocalMux I__17810 (
            .O(N__78035),
            .I(N__78024));
    InMux I__17809 (
            .O(N__78034),
            .I(N__78021));
    InMux I__17808 (
            .O(N__78033),
            .I(N__78016));
    InMux I__17807 (
            .O(N__78032),
            .I(N__78016));
    Span4Mux_h I__17806 (
            .O(N__78027),
            .I(N__78013));
    Span4Mux_v I__17805 (
            .O(N__78024),
            .I(N__78010));
    LocalMux I__17804 (
            .O(N__78021),
            .I(N__78005));
    LocalMux I__17803 (
            .O(N__78016),
            .I(N__78005));
    Odrv4 I__17802 (
            .O(N__78013),
            .I(\bluejay_data_inst.n1137 ));
    Odrv4 I__17801 (
            .O(N__78010),
            .I(\bluejay_data_inst.n1137 ));
    Odrv12 I__17800 (
            .O(N__78005),
            .I(\bluejay_data_inst.n1137 ));
    CascadeMux I__17799 (
            .O(N__77998),
            .I(N__77995));
    InMux I__17798 (
            .O(N__77995),
            .I(N__77992));
    LocalMux I__17797 (
            .O(N__77992),
            .I(n4_adj_1182));
    InMux I__17796 (
            .O(N__77989),
            .I(N__77986));
    LocalMux I__17795 (
            .O(N__77986),
            .I(n3514));
    CascadeMux I__17794 (
            .O(N__77983),
            .I(n4_adj_1182_cascade_));
    InMux I__17793 (
            .O(N__77980),
            .I(N__77977));
    LocalMux I__17792 (
            .O(N__77977),
            .I(n12601));
    InMux I__17791 (
            .O(N__77974),
            .I(N__77970));
    InMux I__17790 (
            .O(N__77973),
            .I(N__77965));
    LocalMux I__17789 (
            .O(N__77970),
            .I(N__77961));
    InMux I__17788 (
            .O(N__77969),
            .I(N__77958));
    CascadeMux I__17787 (
            .O(N__77968),
            .I(N__77952));
    LocalMux I__17786 (
            .O(N__77965),
            .I(N__77947));
    InMux I__17785 (
            .O(N__77964),
            .I(N__77944));
    Span4Mux_v I__17784 (
            .O(N__77961),
            .I(N__77938));
    LocalMux I__17783 (
            .O(N__77958),
            .I(N__77938));
    InMux I__17782 (
            .O(N__77957),
            .I(N__77931));
    InMux I__17781 (
            .O(N__77956),
            .I(N__77927));
    InMux I__17780 (
            .O(N__77955),
            .I(N__77924));
    InMux I__17779 (
            .O(N__77952),
            .I(N__77920));
    InMux I__17778 (
            .O(N__77951),
            .I(N__77917));
    InMux I__17777 (
            .O(N__77950),
            .I(N__77914));
    Span4Mux_v I__17776 (
            .O(N__77947),
            .I(N__77911));
    LocalMux I__17775 (
            .O(N__77944),
            .I(N__77908));
    InMux I__17774 (
            .O(N__77943),
            .I(N__77905));
    Span4Mux_h I__17773 (
            .O(N__77938),
            .I(N__77901));
    InMux I__17772 (
            .O(N__77937),
            .I(N__77898));
    InMux I__17771 (
            .O(N__77936),
            .I(N__77894));
    InMux I__17770 (
            .O(N__77935),
            .I(N__77886));
    InMux I__17769 (
            .O(N__77934),
            .I(N__77883));
    LocalMux I__17768 (
            .O(N__77931),
            .I(N__77880));
    InMux I__17767 (
            .O(N__77930),
            .I(N__77877));
    LocalMux I__17766 (
            .O(N__77927),
            .I(N__77872));
    LocalMux I__17765 (
            .O(N__77924),
            .I(N__77872));
    InMux I__17764 (
            .O(N__77923),
            .I(N__77869));
    LocalMux I__17763 (
            .O(N__77920),
            .I(N__77862));
    LocalMux I__17762 (
            .O(N__77917),
            .I(N__77862));
    LocalMux I__17761 (
            .O(N__77914),
            .I(N__77862));
    Span4Mux_h I__17760 (
            .O(N__77911),
            .I(N__77857));
    Span4Mux_h I__17759 (
            .O(N__77908),
            .I(N__77857));
    LocalMux I__17758 (
            .O(N__77905),
            .I(N__77854));
    InMux I__17757 (
            .O(N__77904),
            .I(N__77851));
    Span4Mux_v I__17756 (
            .O(N__77901),
            .I(N__77845));
    LocalMux I__17755 (
            .O(N__77898),
            .I(N__77845));
    InMux I__17754 (
            .O(N__77897),
            .I(N__77842));
    LocalMux I__17753 (
            .O(N__77894),
            .I(N__77837));
    InMux I__17752 (
            .O(N__77893),
            .I(N__77834));
    InMux I__17751 (
            .O(N__77892),
            .I(N__77827));
    InMux I__17750 (
            .O(N__77891),
            .I(N__77827));
    InMux I__17749 (
            .O(N__77890),
            .I(N__77822));
    InMux I__17748 (
            .O(N__77889),
            .I(N__77822));
    LocalMux I__17747 (
            .O(N__77886),
            .I(N__77819));
    LocalMux I__17746 (
            .O(N__77883),
            .I(N__77812));
    Span4Mux_h I__17745 (
            .O(N__77880),
            .I(N__77812));
    LocalMux I__17744 (
            .O(N__77877),
            .I(N__77812));
    Span4Mux_v I__17743 (
            .O(N__77872),
            .I(N__77809));
    LocalMux I__17742 (
            .O(N__77869),
            .I(N__77806));
    Span4Mux_v I__17741 (
            .O(N__77862),
            .I(N__77801));
    Span4Mux_h I__17740 (
            .O(N__77857),
            .I(N__77801));
    Span4Mux_h I__17739 (
            .O(N__77854),
            .I(N__77796));
    LocalMux I__17738 (
            .O(N__77851),
            .I(N__77796));
    InMux I__17737 (
            .O(N__77850),
            .I(N__77793));
    Span4Mux_h I__17736 (
            .O(N__77845),
            .I(N__77790));
    LocalMux I__17735 (
            .O(N__77842),
            .I(N__77787));
    InMux I__17734 (
            .O(N__77841),
            .I(N__77784));
    InMux I__17733 (
            .O(N__77840),
            .I(N__77780));
    Span4Mux_v I__17732 (
            .O(N__77837),
            .I(N__77777));
    LocalMux I__17731 (
            .O(N__77834),
            .I(N__77774));
    InMux I__17730 (
            .O(N__77833),
            .I(N__77771));
    InMux I__17729 (
            .O(N__77832),
            .I(N__77768));
    LocalMux I__17728 (
            .O(N__77827),
            .I(N__77765));
    LocalMux I__17727 (
            .O(N__77822),
            .I(N__77762));
    Span4Mux_v I__17726 (
            .O(N__77819),
            .I(N__77759));
    Span4Mux_v I__17725 (
            .O(N__77812),
            .I(N__77753));
    Span4Mux_h I__17724 (
            .O(N__77809),
            .I(N__77753));
    Span4Mux_v I__17723 (
            .O(N__77806),
            .I(N__77750));
    Span4Mux_v I__17722 (
            .O(N__77801),
            .I(N__77745));
    Span4Mux_v I__17721 (
            .O(N__77796),
            .I(N__77745));
    LocalMux I__17720 (
            .O(N__77793),
            .I(N__77741));
    Span4Mux_v I__17719 (
            .O(N__77790),
            .I(N__77736));
    Span4Mux_h I__17718 (
            .O(N__77787),
            .I(N__77736));
    LocalMux I__17717 (
            .O(N__77784),
            .I(N__77733));
    InMux I__17716 (
            .O(N__77783),
            .I(N__77730));
    LocalMux I__17715 (
            .O(N__77780),
            .I(N__77721));
    Span4Mux_h I__17714 (
            .O(N__77777),
            .I(N__77721));
    Span4Mux_v I__17713 (
            .O(N__77774),
            .I(N__77721));
    LocalMux I__17712 (
            .O(N__77771),
            .I(N__77721));
    LocalMux I__17711 (
            .O(N__77768),
            .I(N__77716));
    Span4Mux_h I__17710 (
            .O(N__77765),
            .I(N__77716));
    Span4Mux_h I__17709 (
            .O(N__77762),
            .I(N__77711));
    Span4Mux_v I__17708 (
            .O(N__77759),
            .I(N__77711));
    InMux I__17707 (
            .O(N__77758),
            .I(N__77708));
    Sp12to4 I__17706 (
            .O(N__77753),
            .I(N__77703));
    Sp12to4 I__17705 (
            .O(N__77750),
            .I(N__77703));
    Sp12to4 I__17704 (
            .O(N__77745),
            .I(N__77700));
    InMux I__17703 (
            .O(N__77744),
            .I(N__77697));
    Span4Mux_h I__17702 (
            .O(N__77741),
            .I(N__77692));
    Span4Mux_h I__17701 (
            .O(N__77736),
            .I(N__77692));
    Span4Mux_h I__17700 (
            .O(N__77733),
            .I(N__77689));
    LocalMux I__17699 (
            .O(N__77730),
            .I(N__77686));
    Span4Mux_h I__17698 (
            .O(N__77721),
            .I(N__77679));
    Span4Mux_v I__17697 (
            .O(N__77716),
            .I(N__77679));
    Span4Mux_v I__17696 (
            .O(N__77711),
            .I(N__77679));
    LocalMux I__17695 (
            .O(N__77708),
            .I(N__77672));
    Span12Mux_h I__17694 (
            .O(N__77703),
            .I(N__77672));
    Span12Mux_h I__17693 (
            .O(N__77700),
            .I(N__77672));
    LocalMux I__17692 (
            .O(N__77697),
            .I(N__77667));
    Span4Mux_v I__17691 (
            .O(N__77692),
            .I(N__77667));
    Odrv4 I__17690 (
            .O(N__77689),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n65 ));
    Odrv12 I__17689 (
            .O(N__77686),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n65 ));
    Odrv4 I__17688 (
            .O(N__77679),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n65 ));
    Odrv12 I__17687 (
            .O(N__77672),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n65 ));
    Odrv4 I__17686 (
            .O(N__77667),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n65 ));
    InMux I__17685 (
            .O(N__77656),
            .I(N__77653));
    LocalMux I__17684 (
            .O(N__77653),
            .I(N__77649));
    CascadeMux I__17683 (
            .O(N__77652),
            .I(N__77646));
    Sp12to4 I__17682 (
            .O(N__77649),
            .I(N__77643));
    InMux I__17681 (
            .O(N__77646),
            .I(N__77640));
    Odrv12 I__17680 (
            .O(N__77643),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_6 ));
    LocalMux I__17679 (
            .O(N__77640),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_6 ));
    InMux I__17678 (
            .O(N__77635),
            .I(N__77632));
    LocalMux I__17677 (
            .O(N__77632),
            .I(N__77629));
    Span4Mux_v I__17676 (
            .O(N__77629),
            .I(N__77625));
    InMux I__17675 (
            .O(N__77628),
            .I(N__77622));
    Odrv4 I__17674 (
            .O(N__77625),
            .I(REG_mem_5_8));
    LocalMux I__17673 (
            .O(N__77622),
            .I(REG_mem_5_8));
    InMux I__17672 (
            .O(N__77617),
            .I(N__77614));
    LocalMux I__17671 (
            .O(N__77614),
            .I(N__77611));
    Span4Mux_v I__17670 (
            .O(N__77611),
            .I(N__77608));
    Span4Mux_v I__17669 (
            .O(N__77608),
            .I(N__77604));
    InMux I__17668 (
            .O(N__77607),
            .I(N__77601));
    Odrv4 I__17667 (
            .O(N__77604),
            .I(REG_mem_4_8));
    LocalMux I__17666 (
            .O(N__77601),
            .I(REG_mem_4_8));
    CascadeMux I__17665 (
            .O(N__77596),
            .I(\pc_tx.n12133_cascade_ ));
    CascadeMux I__17664 (
            .O(N__77593),
            .I(\pc_tx.o_Tx_Serial_N_840_cascade_ ));
    IoInMux I__17663 (
            .O(N__77590),
            .I(N__77587));
    LocalMux I__17662 (
            .O(N__77587),
            .I(N__77584));
    IoSpan4Mux I__17661 (
            .O(N__77584),
            .I(N__77581));
    Span4Mux_s2_h I__17660 (
            .O(N__77581),
            .I(N__77578));
    Sp12to4 I__17659 (
            .O(N__77578),
            .I(N__77575));
    Span12Mux_v I__17658 (
            .O(N__77575),
            .I(N__77572));
    Odrv12 I__17657 (
            .O(N__77572),
            .I(UART_TX_c));
    InMux I__17656 (
            .O(N__77569),
            .I(N__77566));
    LocalMux I__17655 (
            .O(N__77566),
            .I(N__77563));
    Span4Mux_v I__17654 (
            .O(N__77563),
            .I(N__77559));
    InMux I__17653 (
            .O(N__77562),
            .I(N__77556));
    Odrv4 I__17652 (
            .O(N__77559),
            .I(r_Tx_Data_3));
    LocalMux I__17651 (
            .O(N__77556),
            .I(r_Tx_Data_3));
    InMux I__17650 (
            .O(N__77551),
            .I(N__77548));
    LocalMux I__17649 (
            .O(N__77548),
            .I(\pc_tx.n12134 ));
    InMux I__17648 (
            .O(N__77545),
            .I(N__77542));
    LocalMux I__17647 (
            .O(N__77542),
            .I(N__77539));
    Span4Mux_v I__17646 (
            .O(N__77539),
            .I(N__77535));
    InMux I__17645 (
            .O(N__77538),
            .I(N__77532));
    Odrv4 I__17644 (
            .O(N__77535),
            .I(r_Tx_Data_5));
    LocalMux I__17643 (
            .O(N__77532),
            .I(r_Tx_Data_5));
    InMux I__17642 (
            .O(N__77527),
            .I(N__77524));
    LocalMux I__17641 (
            .O(N__77524),
            .I(N__77520));
    InMux I__17640 (
            .O(N__77523),
            .I(N__77517));
    Odrv4 I__17639 (
            .O(N__77520),
            .I(r_Tx_Data_4));
    LocalMux I__17638 (
            .O(N__77517),
            .I(r_Tx_Data_4));
    CascadeMux I__17637 (
            .O(N__77512),
            .I(\pc_tx.n12139_cascade_ ));
    InMux I__17636 (
            .O(N__77509),
            .I(N__77506));
    LocalMux I__17635 (
            .O(N__77506),
            .I(\pc_tx.n13790 ));
    CascadeMux I__17634 (
            .O(N__77503),
            .I(N__77499));
    InMux I__17633 (
            .O(N__77502),
            .I(N__77494));
    InMux I__17632 (
            .O(N__77499),
            .I(N__77494));
    LocalMux I__17631 (
            .O(N__77494),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_4 ));
    CascadeMux I__17630 (
            .O(N__77491),
            .I(N__77487));
    InMux I__17629 (
            .O(N__77490),
            .I(N__77482));
    InMux I__17628 (
            .O(N__77487),
            .I(N__77482));
    LocalMux I__17627 (
            .O(N__77482),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_4 ));
    CascadeMux I__17626 (
            .O(N__77479),
            .I(N__77476));
    InMux I__17625 (
            .O(N__77476),
            .I(N__77468));
    InMux I__17624 (
            .O(N__77475),
            .I(N__77459));
    InMux I__17623 (
            .O(N__77474),
            .I(N__77459));
    InMux I__17622 (
            .O(N__77473),
            .I(N__77452));
    InMux I__17621 (
            .O(N__77472),
            .I(N__77444));
    InMux I__17620 (
            .O(N__77471),
            .I(N__77444));
    LocalMux I__17619 (
            .O(N__77468),
            .I(N__77435));
    InMux I__17618 (
            .O(N__77467),
            .I(N__77432));
    CascadeMux I__17617 (
            .O(N__77466),
            .I(N__77429));
    InMux I__17616 (
            .O(N__77465),
            .I(N__77426));
    InMux I__17615 (
            .O(N__77464),
            .I(N__77423));
    LocalMux I__17614 (
            .O(N__77459),
            .I(N__77420));
    InMux I__17613 (
            .O(N__77458),
            .I(N__77413));
    InMux I__17612 (
            .O(N__77457),
            .I(N__77410));
    InMux I__17611 (
            .O(N__77456),
            .I(N__77405));
    InMux I__17610 (
            .O(N__77455),
            .I(N__77405));
    LocalMux I__17609 (
            .O(N__77452),
            .I(N__77402));
    InMux I__17608 (
            .O(N__77451),
            .I(N__77395));
    InMux I__17607 (
            .O(N__77450),
            .I(N__77395));
    InMux I__17606 (
            .O(N__77449),
            .I(N__77395));
    LocalMux I__17605 (
            .O(N__77444),
            .I(N__77392));
    InMux I__17604 (
            .O(N__77443),
            .I(N__77384));
    InMux I__17603 (
            .O(N__77442),
            .I(N__77379));
    InMux I__17602 (
            .O(N__77441),
            .I(N__77379));
    InMux I__17601 (
            .O(N__77440),
            .I(N__77372));
    InMux I__17600 (
            .O(N__77439),
            .I(N__77372));
    InMux I__17599 (
            .O(N__77438),
            .I(N__77372));
    Span4Mux_h I__17598 (
            .O(N__77435),
            .I(N__77367));
    LocalMux I__17597 (
            .O(N__77432),
            .I(N__77367));
    InMux I__17596 (
            .O(N__77429),
            .I(N__77364));
    LocalMux I__17595 (
            .O(N__77426),
            .I(N__77361));
    LocalMux I__17594 (
            .O(N__77423),
            .I(N__77356));
    Span4Mux_h I__17593 (
            .O(N__77420),
            .I(N__77356));
    InMux I__17592 (
            .O(N__77419),
            .I(N__77353));
    InMux I__17591 (
            .O(N__77418),
            .I(N__77350));
    InMux I__17590 (
            .O(N__77417),
            .I(N__77345));
    InMux I__17589 (
            .O(N__77416),
            .I(N__77345));
    LocalMux I__17588 (
            .O(N__77413),
            .I(N__77338));
    LocalMux I__17587 (
            .O(N__77410),
            .I(N__77338));
    LocalMux I__17586 (
            .O(N__77405),
            .I(N__77338));
    Sp12to4 I__17585 (
            .O(N__77402),
            .I(N__77335));
    LocalMux I__17584 (
            .O(N__77395),
            .I(N__77330));
    Span4Mux_v I__17583 (
            .O(N__77392),
            .I(N__77330));
    InMux I__17582 (
            .O(N__77391),
            .I(N__77327));
    InMux I__17581 (
            .O(N__77390),
            .I(N__77324));
    InMux I__17580 (
            .O(N__77389),
            .I(N__77317));
    InMux I__17579 (
            .O(N__77388),
            .I(N__77317));
    InMux I__17578 (
            .O(N__77387),
            .I(N__77317));
    LocalMux I__17577 (
            .O(N__77384),
            .I(N__77312));
    LocalMux I__17576 (
            .O(N__77379),
            .I(N__77312));
    LocalMux I__17575 (
            .O(N__77372),
            .I(N__77309));
    Span4Mux_v I__17574 (
            .O(N__77367),
            .I(N__77306));
    LocalMux I__17573 (
            .O(N__77364),
            .I(N__77299));
    Span4Mux_h I__17572 (
            .O(N__77361),
            .I(N__77299));
    Span4Mux_h I__17571 (
            .O(N__77356),
            .I(N__77299));
    LocalMux I__17570 (
            .O(N__77353),
            .I(N__77286));
    LocalMux I__17569 (
            .O(N__77350),
            .I(N__77286));
    LocalMux I__17568 (
            .O(N__77345),
            .I(N__77286));
    Span12Mux_v I__17567 (
            .O(N__77338),
            .I(N__77286));
    Span12Mux_v I__17566 (
            .O(N__77335),
            .I(N__77286));
    Sp12to4 I__17565 (
            .O(N__77330),
            .I(N__77286));
    LocalMux I__17564 (
            .O(N__77327),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n45 ));
    LocalMux I__17563 (
            .O(N__77324),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n45 ));
    LocalMux I__17562 (
            .O(N__77317),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n45 ));
    Odrv12 I__17561 (
            .O(N__77312),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n45 ));
    Odrv4 I__17560 (
            .O(N__77309),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n45 ));
    Odrv4 I__17559 (
            .O(N__77306),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n45 ));
    Odrv4 I__17558 (
            .O(N__77299),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n45 ));
    Odrv12 I__17557 (
            .O(N__77286),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n45 ));
    InMux I__17556 (
            .O(N__77269),
            .I(N__77266));
    LocalMux I__17555 (
            .O(N__77266),
            .I(N__77262));
    CascadeMux I__17554 (
            .O(N__77265),
            .I(N__77259));
    Span4Mux_h I__17553 (
            .O(N__77262),
            .I(N__77256));
    InMux I__17552 (
            .O(N__77259),
            .I(N__77253));
    Odrv4 I__17551 (
            .O(N__77256),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_4 ));
    LocalMux I__17550 (
            .O(N__77253),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_4 ));
    InMux I__17549 (
            .O(N__77248),
            .I(N__77241));
    InMux I__17548 (
            .O(N__77247),
            .I(N__77237));
    InMux I__17547 (
            .O(N__77246),
            .I(N__77233));
    InMux I__17546 (
            .O(N__77245),
            .I(N__77226));
    InMux I__17545 (
            .O(N__77244),
            .I(N__77223));
    LocalMux I__17544 (
            .O(N__77241),
            .I(N__77220));
    InMux I__17543 (
            .O(N__77240),
            .I(N__77217));
    LocalMux I__17542 (
            .O(N__77237),
            .I(N__77214));
    InMux I__17541 (
            .O(N__77236),
            .I(N__77211));
    LocalMux I__17540 (
            .O(N__77233),
            .I(N__77206));
    InMux I__17539 (
            .O(N__77232),
            .I(N__77203));
    InMux I__17538 (
            .O(N__77231),
            .I(N__77199));
    InMux I__17537 (
            .O(N__77230),
            .I(N__77196));
    InMux I__17536 (
            .O(N__77229),
            .I(N__77193));
    LocalMux I__17535 (
            .O(N__77226),
            .I(N__77187));
    LocalMux I__17534 (
            .O(N__77223),
            .I(N__77187));
    Span4Mux_v I__17533 (
            .O(N__77220),
            .I(N__77184));
    LocalMux I__17532 (
            .O(N__77217),
            .I(N__77181));
    Span4Mux_v I__17531 (
            .O(N__77214),
            .I(N__77178));
    LocalMux I__17530 (
            .O(N__77211),
            .I(N__77175));
    InMux I__17529 (
            .O(N__77210),
            .I(N__77172));
    InMux I__17528 (
            .O(N__77209),
            .I(N__77169));
    Span4Mux_h I__17527 (
            .O(N__77206),
            .I(N__77166));
    LocalMux I__17526 (
            .O(N__77203),
            .I(N__77163));
    InMux I__17525 (
            .O(N__77202),
            .I(N__77160));
    LocalMux I__17524 (
            .O(N__77199),
            .I(N__77157));
    LocalMux I__17523 (
            .O(N__77196),
            .I(N__77154));
    LocalMux I__17522 (
            .O(N__77193),
            .I(N__77151));
    InMux I__17521 (
            .O(N__77192),
            .I(N__77148));
    Span4Mux_h I__17520 (
            .O(N__77187),
            .I(N__77145));
    Span4Mux_h I__17519 (
            .O(N__77184),
            .I(N__77140));
    Span4Mux_v I__17518 (
            .O(N__77181),
            .I(N__77140));
    Span4Mux_v I__17517 (
            .O(N__77178),
            .I(N__77135));
    Span4Mux_v I__17516 (
            .O(N__77175),
            .I(N__77135));
    LocalMux I__17515 (
            .O(N__77172),
            .I(N__77132));
    LocalMux I__17514 (
            .O(N__77169),
            .I(N__77129));
    Span4Mux_h I__17513 (
            .O(N__77166),
            .I(N__77122));
    Span4Mux_v I__17512 (
            .O(N__77163),
            .I(N__77122));
    LocalMux I__17511 (
            .O(N__77160),
            .I(N__77122));
    Span4Mux_v I__17510 (
            .O(N__77157),
            .I(N__77119));
    Span4Mux_v I__17509 (
            .O(N__77154),
            .I(N__77116));
    Span4Mux_v I__17508 (
            .O(N__77151),
            .I(N__77113));
    LocalMux I__17507 (
            .O(N__77148),
            .I(N__77110));
    Span4Mux_h I__17506 (
            .O(N__77145),
            .I(N__77101));
    Span4Mux_v I__17505 (
            .O(N__77140),
            .I(N__77101));
    Span4Mux_h I__17504 (
            .O(N__77135),
            .I(N__77101));
    Span4Mux_v I__17503 (
            .O(N__77132),
            .I(N__77101));
    Span4Mux_v I__17502 (
            .O(N__77129),
            .I(N__77096));
    Span4Mux_h I__17501 (
            .O(N__77122),
            .I(N__77096));
    Span4Mux_v I__17500 (
            .O(N__77119),
            .I(N__77087));
    Span4Mux_h I__17499 (
            .O(N__77116),
            .I(N__77087));
    Span4Mux_v I__17498 (
            .O(N__77113),
            .I(N__77087));
    Span4Mux_v I__17497 (
            .O(N__77110),
            .I(N__77087));
    Odrv4 I__17496 (
            .O(N__77101),
            .I(n10));
    Odrv4 I__17495 (
            .O(N__77096),
            .I(n10));
    Odrv4 I__17494 (
            .O(N__77087),
            .I(n10));
    InMux I__17493 (
            .O(N__77080),
            .I(N__77074));
    InMux I__17492 (
            .O(N__77079),
            .I(N__77074));
    LocalMux I__17491 (
            .O(N__77074),
            .I(REG_mem_55_8));
    CascadeMux I__17490 (
            .O(N__77071),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13460_cascade_ ));
    InMux I__17489 (
            .O(N__77068),
            .I(N__77064));
    InMux I__17488 (
            .O(N__77067),
            .I(N__77061));
    LocalMux I__17487 (
            .O(N__77064),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_8 ));
    LocalMux I__17486 (
            .O(N__77061),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_8 ));
    InMux I__17485 (
            .O(N__77056),
            .I(N__77050));
    InMux I__17484 (
            .O(N__77055),
            .I(N__77050));
    LocalMux I__17483 (
            .O(N__77050),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_8 ));
    InMux I__17482 (
            .O(N__77047),
            .I(N__77042));
    InMux I__17481 (
            .O(N__77046),
            .I(N__77032));
    InMux I__17480 (
            .O(N__77045),
            .I(N__77029));
    LocalMux I__17479 (
            .O(N__77042),
            .I(N__77026));
    InMux I__17478 (
            .O(N__77041),
            .I(N__77023));
    InMux I__17477 (
            .O(N__77040),
            .I(N__77016));
    InMux I__17476 (
            .O(N__77039),
            .I(N__77010));
    InMux I__17475 (
            .O(N__77038),
            .I(N__77007));
    InMux I__17474 (
            .O(N__77037),
            .I(N__77004));
    InMux I__17473 (
            .O(N__77036),
            .I(N__77000));
    InMux I__17472 (
            .O(N__77035),
            .I(N__76997));
    LocalMux I__17471 (
            .O(N__77032),
            .I(N__76992));
    LocalMux I__17470 (
            .O(N__77029),
            .I(N__76992));
    Span4Mux_v I__17469 (
            .O(N__77026),
            .I(N__76987));
    LocalMux I__17468 (
            .O(N__77023),
            .I(N__76987));
    InMux I__17467 (
            .O(N__77022),
            .I(N__76980));
    InMux I__17466 (
            .O(N__77021),
            .I(N__76980));
    InMux I__17465 (
            .O(N__77020),
            .I(N__76977));
    InMux I__17464 (
            .O(N__77019),
            .I(N__76972));
    LocalMux I__17463 (
            .O(N__77016),
            .I(N__76969));
    InMux I__17462 (
            .O(N__77015),
            .I(N__76966));
    InMux I__17461 (
            .O(N__77014),
            .I(N__76961));
    InMux I__17460 (
            .O(N__77013),
            .I(N__76961));
    LocalMux I__17459 (
            .O(N__77010),
            .I(N__76958));
    LocalMux I__17458 (
            .O(N__77007),
            .I(N__76955));
    LocalMux I__17457 (
            .O(N__77004),
            .I(N__76952));
    InMux I__17456 (
            .O(N__77003),
            .I(N__76949));
    LocalMux I__17455 (
            .O(N__77000),
            .I(N__76946));
    LocalMux I__17454 (
            .O(N__76997),
            .I(N__76940));
    Span4Mux_v I__17453 (
            .O(N__76992),
            .I(N__76937));
    Span4Mux_v I__17452 (
            .O(N__76987),
            .I(N__76934));
    InMux I__17451 (
            .O(N__76986),
            .I(N__76931));
    InMux I__17450 (
            .O(N__76985),
            .I(N__76928));
    LocalMux I__17449 (
            .O(N__76980),
            .I(N__76922));
    LocalMux I__17448 (
            .O(N__76977),
            .I(N__76922));
    InMux I__17447 (
            .O(N__76976),
            .I(N__76919));
    InMux I__17446 (
            .O(N__76975),
            .I(N__76912));
    LocalMux I__17445 (
            .O(N__76972),
            .I(N__76908));
    Span4Mux_v I__17444 (
            .O(N__76969),
            .I(N__76903));
    LocalMux I__17443 (
            .O(N__76966),
            .I(N__76903));
    LocalMux I__17442 (
            .O(N__76961),
            .I(N__76900));
    Span4Mux_h I__17441 (
            .O(N__76958),
            .I(N__76891));
    Span4Mux_h I__17440 (
            .O(N__76955),
            .I(N__76891));
    Span4Mux_v I__17439 (
            .O(N__76952),
            .I(N__76891));
    LocalMux I__17438 (
            .O(N__76949),
            .I(N__76891));
    Span4Mux_h I__17437 (
            .O(N__76946),
            .I(N__76888));
    InMux I__17436 (
            .O(N__76945),
            .I(N__76881));
    InMux I__17435 (
            .O(N__76944),
            .I(N__76881));
    InMux I__17434 (
            .O(N__76943),
            .I(N__76881));
    Span4Mux_v I__17433 (
            .O(N__76940),
            .I(N__76878));
    Span4Mux_v I__17432 (
            .O(N__76937),
            .I(N__76871));
    Span4Mux_h I__17431 (
            .O(N__76934),
            .I(N__76871));
    LocalMux I__17430 (
            .O(N__76931),
            .I(N__76871));
    LocalMux I__17429 (
            .O(N__76928),
            .I(N__76868));
    InMux I__17428 (
            .O(N__76927),
            .I(N__76865));
    Span4Mux_h I__17427 (
            .O(N__76922),
            .I(N__76862));
    LocalMux I__17426 (
            .O(N__76919),
            .I(N__76859));
    InMux I__17425 (
            .O(N__76918),
            .I(N__76854));
    InMux I__17424 (
            .O(N__76917),
            .I(N__76854));
    InMux I__17423 (
            .O(N__76916),
            .I(N__76851));
    InMux I__17422 (
            .O(N__76915),
            .I(N__76848));
    LocalMux I__17421 (
            .O(N__76912),
            .I(N__76845));
    InMux I__17420 (
            .O(N__76911),
            .I(N__76842));
    Span4Mux_v I__17419 (
            .O(N__76908),
            .I(N__76836));
    Span4Mux_h I__17418 (
            .O(N__76903),
            .I(N__76836));
    Span4Mux_h I__17417 (
            .O(N__76900),
            .I(N__76833));
    Span4Mux_h I__17416 (
            .O(N__76891),
            .I(N__76830));
    Span4Mux_h I__17415 (
            .O(N__76888),
            .I(N__76825));
    LocalMux I__17414 (
            .O(N__76881),
            .I(N__76825));
    Span4Mux_h I__17413 (
            .O(N__76878),
            .I(N__76816));
    Span4Mux_v I__17412 (
            .O(N__76871),
            .I(N__76816));
    Span4Mux_v I__17411 (
            .O(N__76868),
            .I(N__76816));
    LocalMux I__17410 (
            .O(N__76865),
            .I(N__76816));
    Span4Mux_h I__17409 (
            .O(N__76862),
            .I(N__76813));
    Span4Mux_v I__17408 (
            .O(N__76859),
            .I(N__76806));
    LocalMux I__17407 (
            .O(N__76854),
            .I(N__76806));
    LocalMux I__17406 (
            .O(N__76851),
            .I(N__76806));
    LocalMux I__17405 (
            .O(N__76848),
            .I(N__76803));
    Span4Mux_v I__17404 (
            .O(N__76845),
            .I(N__76798));
    LocalMux I__17403 (
            .O(N__76842),
            .I(N__76798));
    InMux I__17402 (
            .O(N__76841),
            .I(N__76795));
    Span4Mux_h I__17401 (
            .O(N__76836),
            .I(N__76788));
    Span4Mux_h I__17400 (
            .O(N__76833),
            .I(N__76788));
    Span4Mux_v I__17399 (
            .O(N__76830),
            .I(N__76788));
    Span4Mux_h I__17398 (
            .O(N__76825),
            .I(N__76783));
    Span4Mux_h I__17397 (
            .O(N__76816),
            .I(N__76783));
    Span4Mux_h I__17396 (
            .O(N__76813),
            .I(N__76778));
    Span4Mux_h I__17395 (
            .O(N__76806),
            .I(N__76778));
    Span4Mux_v I__17394 (
            .O(N__76803),
            .I(N__76771));
    Span4Mux_h I__17393 (
            .O(N__76798),
            .I(N__76771));
    LocalMux I__17392 (
            .O(N__76795),
            .I(N__76771));
    Odrv4 I__17391 (
            .O(N__76788),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n47 ));
    Odrv4 I__17390 (
            .O(N__76783),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n47 ));
    Odrv4 I__17389 (
            .O(N__76778),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n47 ));
    Odrv4 I__17388 (
            .O(N__76771),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n47 ));
    CascadeMux I__17387 (
            .O(N__76762),
            .I(N__76755));
    InMux I__17386 (
            .O(N__76761),
            .I(N__76746));
    InMux I__17385 (
            .O(N__76760),
            .I(N__76746));
    InMux I__17384 (
            .O(N__76759),
            .I(N__76740));
    InMux I__17383 (
            .O(N__76758),
            .I(N__76737));
    InMux I__17382 (
            .O(N__76755),
            .I(N__76726));
    InMux I__17381 (
            .O(N__76754),
            .I(N__76726));
    InMux I__17380 (
            .O(N__76753),
            .I(N__76726));
    CascadeMux I__17379 (
            .O(N__76752),
            .I(N__76723));
    InMux I__17378 (
            .O(N__76751),
            .I(N__76717));
    LocalMux I__17377 (
            .O(N__76746),
            .I(N__76699));
    InMux I__17376 (
            .O(N__76745),
            .I(N__76696));
    InMux I__17375 (
            .O(N__76744),
            .I(N__76692));
    InMux I__17374 (
            .O(N__76743),
            .I(N__76687));
    LocalMux I__17373 (
            .O(N__76740),
            .I(N__76682));
    LocalMux I__17372 (
            .O(N__76737),
            .I(N__76682));
    InMux I__17371 (
            .O(N__76736),
            .I(N__76673));
    InMux I__17370 (
            .O(N__76735),
            .I(N__76673));
    InMux I__17369 (
            .O(N__76734),
            .I(N__76673));
    InMux I__17368 (
            .O(N__76733),
            .I(N__76673));
    LocalMux I__17367 (
            .O(N__76726),
            .I(N__76670));
    InMux I__17366 (
            .O(N__76723),
            .I(N__76661));
    InMux I__17365 (
            .O(N__76722),
            .I(N__76661));
    InMux I__17364 (
            .O(N__76721),
            .I(N__76661));
    InMux I__17363 (
            .O(N__76720),
            .I(N__76661));
    LocalMux I__17362 (
            .O(N__76717),
            .I(N__76658));
    InMux I__17361 (
            .O(N__76716),
            .I(N__76647));
    InMux I__17360 (
            .O(N__76715),
            .I(N__76647));
    InMux I__17359 (
            .O(N__76714),
            .I(N__76647));
    InMux I__17358 (
            .O(N__76713),
            .I(N__76647));
    InMux I__17357 (
            .O(N__76712),
            .I(N__76647));
    InMux I__17356 (
            .O(N__76711),
            .I(N__76640));
    InMux I__17355 (
            .O(N__76710),
            .I(N__76640));
    InMux I__17354 (
            .O(N__76709),
            .I(N__76640));
    InMux I__17353 (
            .O(N__76708),
            .I(N__76630));
    InMux I__17352 (
            .O(N__76707),
            .I(N__76630));
    InMux I__17351 (
            .O(N__76706),
            .I(N__76623));
    InMux I__17350 (
            .O(N__76705),
            .I(N__76623));
    InMux I__17349 (
            .O(N__76704),
            .I(N__76623));
    InMux I__17348 (
            .O(N__76703),
            .I(N__76607));
    InMux I__17347 (
            .O(N__76702),
            .I(N__76597));
    Span4Mux_h I__17346 (
            .O(N__76699),
            .I(N__76592));
    LocalMux I__17345 (
            .O(N__76696),
            .I(N__76592));
    InMux I__17344 (
            .O(N__76695),
            .I(N__76589));
    LocalMux I__17343 (
            .O(N__76692),
            .I(N__76585));
    InMux I__17342 (
            .O(N__76691),
            .I(N__76580));
    InMux I__17341 (
            .O(N__76690),
            .I(N__76580));
    LocalMux I__17340 (
            .O(N__76687),
            .I(N__76575));
    Span4Mux_h I__17339 (
            .O(N__76682),
            .I(N__76575));
    LocalMux I__17338 (
            .O(N__76673),
            .I(N__76568));
    Span4Mux_h I__17337 (
            .O(N__76670),
            .I(N__76568));
    LocalMux I__17336 (
            .O(N__76661),
            .I(N__76568));
    Span4Mux_v I__17335 (
            .O(N__76658),
            .I(N__76565));
    LocalMux I__17334 (
            .O(N__76647),
            .I(N__76560));
    LocalMux I__17333 (
            .O(N__76640),
            .I(N__76560));
    InMux I__17332 (
            .O(N__76639),
            .I(N__76557));
    InMux I__17331 (
            .O(N__76638),
            .I(N__76552));
    InMux I__17330 (
            .O(N__76637),
            .I(N__76552));
    InMux I__17329 (
            .O(N__76636),
            .I(N__76547));
    InMux I__17328 (
            .O(N__76635),
            .I(N__76547));
    LocalMux I__17327 (
            .O(N__76630),
            .I(N__76544));
    LocalMux I__17326 (
            .O(N__76623),
            .I(N__76541));
    InMux I__17325 (
            .O(N__76622),
            .I(N__76538));
    InMux I__17324 (
            .O(N__76621),
            .I(N__76535));
    InMux I__17323 (
            .O(N__76620),
            .I(N__76532));
    InMux I__17322 (
            .O(N__76619),
            .I(N__76525));
    InMux I__17321 (
            .O(N__76618),
            .I(N__76525));
    InMux I__17320 (
            .O(N__76617),
            .I(N__76525));
    InMux I__17319 (
            .O(N__76616),
            .I(N__76514));
    InMux I__17318 (
            .O(N__76615),
            .I(N__76514));
    InMux I__17317 (
            .O(N__76614),
            .I(N__76514));
    InMux I__17316 (
            .O(N__76613),
            .I(N__76514));
    InMux I__17315 (
            .O(N__76612),
            .I(N__76514));
    InMux I__17314 (
            .O(N__76611),
            .I(N__76510));
    InMux I__17313 (
            .O(N__76610),
            .I(N__76507));
    LocalMux I__17312 (
            .O(N__76607),
            .I(N__76504));
    InMux I__17311 (
            .O(N__76606),
            .I(N__76499));
    InMux I__17310 (
            .O(N__76605),
            .I(N__76499));
    InMux I__17309 (
            .O(N__76604),
            .I(N__76488));
    InMux I__17308 (
            .O(N__76603),
            .I(N__76488));
    InMux I__17307 (
            .O(N__76602),
            .I(N__76488));
    InMux I__17306 (
            .O(N__76601),
            .I(N__76488));
    InMux I__17305 (
            .O(N__76600),
            .I(N__76488));
    LocalMux I__17304 (
            .O(N__76597),
            .I(N__76483));
    Span4Mux_v I__17303 (
            .O(N__76592),
            .I(N__76483));
    LocalMux I__17302 (
            .O(N__76589),
            .I(N__76480));
    InMux I__17301 (
            .O(N__76588),
            .I(N__76477));
    Span4Mux_v I__17300 (
            .O(N__76585),
            .I(N__76474));
    LocalMux I__17299 (
            .O(N__76580),
            .I(N__76463));
    Span4Mux_h I__17298 (
            .O(N__76575),
            .I(N__76463));
    Span4Mux_h I__17297 (
            .O(N__76568),
            .I(N__76463));
    Span4Mux_h I__17296 (
            .O(N__76565),
            .I(N__76463));
    Span4Mux_v I__17295 (
            .O(N__76560),
            .I(N__76463));
    LocalMux I__17294 (
            .O(N__76557),
            .I(N__76456));
    LocalMux I__17293 (
            .O(N__76552),
            .I(N__76456));
    LocalMux I__17292 (
            .O(N__76547),
            .I(N__76456));
    Span4Mux_v I__17291 (
            .O(N__76544),
            .I(N__76453));
    Span4Mux_v I__17290 (
            .O(N__76541),
            .I(N__76448));
    LocalMux I__17289 (
            .O(N__76538),
            .I(N__76448));
    LocalMux I__17288 (
            .O(N__76535),
            .I(N__76439));
    LocalMux I__17287 (
            .O(N__76532),
            .I(N__76439));
    LocalMux I__17286 (
            .O(N__76525),
            .I(N__76439));
    LocalMux I__17285 (
            .O(N__76514),
            .I(N__76439));
    InMux I__17284 (
            .O(N__76513),
            .I(N__76436));
    LocalMux I__17283 (
            .O(N__76510),
            .I(N__76431));
    LocalMux I__17282 (
            .O(N__76507),
            .I(N__76431));
    Span4Mux_v I__17281 (
            .O(N__76504),
            .I(N__76428));
    LocalMux I__17280 (
            .O(N__76499),
            .I(N__76421));
    LocalMux I__17279 (
            .O(N__76488),
            .I(N__76421));
    Span4Mux_h I__17278 (
            .O(N__76483),
            .I(N__76421));
    Sp12to4 I__17277 (
            .O(N__76480),
            .I(N__76418));
    LocalMux I__17276 (
            .O(N__76477),
            .I(N__76415));
    Span4Mux_h I__17275 (
            .O(N__76474),
            .I(N__76410));
    Span4Mux_v I__17274 (
            .O(N__76463),
            .I(N__76410));
    Span4Mux_v I__17273 (
            .O(N__76456),
            .I(N__76405));
    Span4Mux_h I__17272 (
            .O(N__76453),
            .I(N__76405));
    Span4Mux_v I__17271 (
            .O(N__76448),
            .I(N__76402));
    Span12Mux_v I__17270 (
            .O(N__76439),
            .I(N__76399));
    LocalMux I__17269 (
            .O(N__76436),
            .I(N__76390));
    Span4Mux_v I__17268 (
            .O(N__76431),
            .I(N__76390));
    Span4Mux_h I__17267 (
            .O(N__76428),
            .I(N__76390));
    Span4Mux_v I__17266 (
            .O(N__76421),
            .I(N__76390));
    Span12Mux_v I__17265 (
            .O(N__76418),
            .I(N__76387));
    Span4Mux_v I__17264 (
            .O(N__76415),
            .I(N__76382));
    Span4Mux_v I__17263 (
            .O(N__76410),
            .I(N__76382));
    Odrv4 I__17262 (
            .O(N__76405),
            .I(dc32_fifo_data_in_4));
    Odrv4 I__17261 (
            .O(N__76402),
            .I(dc32_fifo_data_in_4));
    Odrv12 I__17260 (
            .O(N__76399),
            .I(dc32_fifo_data_in_4));
    Odrv4 I__17259 (
            .O(N__76390),
            .I(dc32_fifo_data_in_4));
    Odrv12 I__17258 (
            .O(N__76387),
            .I(dc32_fifo_data_in_4));
    Odrv4 I__17257 (
            .O(N__76382),
            .I(dc32_fifo_data_in_4));
    CascadeMux I__17256 (
            .O(N__76369),
            .I(N__76365));
    InMux I__17255 (
            .O(N__76368),
            .I(N__76362));
    InMux I__17254 (
            .O(N__76365),
            .I(N__76359));
    LocalMux I__17253 (
            .O(N__76362),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_4 ));
    LocalMux I__17252 (
            .O(N__76359),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_4 ));
    InMux I__17251 (
            .O(N__76354),
            .I(N__76347));
    InMux I__17250 (
            .O(N__76353),
            .I(N__76341));
    InMux I__17249 (
            .O(N__76352),
            .I(N__76338));
    InMux I__17248 (
            .O(N__76351),
            .I(N__76326));
    InMux I__17247 (
            .O(N__76350),
            .I(N__76326));
    LocalMux I__17246 (
            .O(N__76347),
            .I(N__76320));
    InMux I__17245 (
            .O(N__76346),
            .I(N__76317));
    InMux I__17244 (
            .O(N__76345),
            .I(N__76314));
    InMux I__17243 (
            .O(N__76344),
            .I(N__76309));
    LocalMux I__17242 (
            .O(N__76341),
            .I(N__76301));
    LocalMux I__17241 (
            .O(N__76338),
            .I(N__76301));
    InMux I__17240 (
            .O(N__76337),
            .I(N__76298));
    InMux I__17239 (
            .O(N__76336),
            .I(N__76295));
    InMux I__17238 (
            .O(N__76335),
            .I(N__76292));
    InMux I__17237 (
            .O(N__76334),
            .I(N__76287));
    InMux I__17236 (
            .O(N__76333),
            .I(N__76287));
    InMux I__17235 (
            .O(N__76332),
            .I(N__76284));
    InMux I__17234 (
            .O(N__76331),
            .I(N__76280));
    LocalMux I__17233 (
            .O(N__76326),
            .I(N__76277));
    InMux I__17232 (
            .O(N__76325),
            .I(N__76274));
    InMux I__17231 (
            .O(N__76324),
            .I(N__76269));
    InMux I__17230 (
            .O(N__76323),
            .I(N__76269));
    Span4Mux_h I__17229 (
            .O(N__76320),
            .I(N__76261));
    LocalMux I__17228 (
            .O(N__76317),
            .I(N__76261));
    LocalMux I__17227 (
            .O(N__76314),
            .I(N__76261));
    InMux I__17226 (
            .O(N__76313),
            .I(N__76256));
    InMux I__17225 (
            .O(N__76312),
            .I(N__76256));
    LocalMux I__17224 (
            .O(N__76309),
            .I(N__76252));
    InMux I__17223 (
            .O(N__76308),
            .I(N__76249));
    InMux I__17222 (
            .O(N__76307),
            .I(N__76244));
    InMux I__17221 (
            .O(N__76306),
            .I(N__76244));
    Span4Mux_v I__17220 (
            .O(N__76301),
            .I(N__76241));
    LocalMux I__17219 (
            .O(N__76298),
            .I(N__76238));
    LocalMux I__17218 (
            .O(N__76295),
            .I(N__76232));
    LocalMux I__17217 (
            .O(N__76292),
            .I(N__76229));
    LocalMux I__17216 (
            .O(N__76287),
            .I(N__76226));
    LocalMux I__17215 (
            .O(N__76284),
            .I(N__76223));
    InMux I__17214 (
            .O(N__76283),
            .I(N__76220));
    LocalMux I__17213 (
            .O(N__76280),
            .I(N__76217));
    Span4Mux_h I__17212 (
            .O(N__76277),
            .I(N__76212));
    LocalMux I__17211 (
            .O(N__76274),
            .I(N__76212));
    LocalMux I__17210 (
            .O(N__76269),
            .I(N__76208));
    InMux I__17209 (
            .O(N__76268),
            .I(N__76205));
    Span4Mux_h I__17208 (
            .O(N__76261),
            .I(N__76202));
    LocalMux I__17207 (
            .O(N__76256),
            .I(N__76199));
    InMux I__17206 (
            .O(N__76255),
            .I(N__76196));
    Span4Mux_v I__17205 (
            .O(N__76252),
            .I(N__76192));
    LocalMux I__17204 (
            .O(N__76249),
            .I(N__76189));
    LocalMux I__17203 (
            .O(N__76244),
            .I(N__76186));
    Span4Mux_h I__17202 (
            .O(N__76241),
            .I(N__76181));
    Span4Mux_v I__17201 (
            .O(N__76238),
            .I(N__76181));
    InMux I__17200 (
            .O(N__76237),
            .I(N__76178));
    InMux I__17199 (
            .O(N__76236),
            .I(N__76175));
    InMux I__17198 (
            .O(N__76235),
            .I(N__76172));
    Span4Mux_h I__17197 (
            .O(N__76232),
            .I(N__76167));
    Span4Mux_v I__17196 (
            .O(N__76229),
            .I(N__76167));
    Span4Mux_v I__17195 (
            .O(N__76226),
            .I(N__76162));
    Span4Mux_h I__17194 (
            .O(N__76223),
            .I(N__76162));
    LocalMux I__17193 (
            .O(N__76220),
            .I(N__76159));
    Span4Mux_h I__17192 (
            .O(N__76217),
            .I(N__76156));
    Span4Mux_h I__17191 (
            .O(N__76212),
            .I(N__76153));
    InMux I__17190 (
            .O(N__76211),
            .I(N__76150));
    Span4Mux_h I__17189 (
            .O(N__76208),
            .I(N__76145));
    LocalMux I__17188 (
            .O(N__76205),
            .I(N__76145));
    Span4Mux_h I__17187 (
            .O(N__76202),
            .I(N__76138));
    Span4Mux_v I__17186 (
            .O(N__76199),
            .I(N__76138));
    LocalMux I__17185 (
            .O(N__76196),
            .I(N__76138));
    InMux I__17184 (
            .O(N__76195),
            .I(N__76135));
    Sp12to4 I__17183 (
            .O(N__76192),
            .I(N__76119));
    Span12Mux_s10_h I__17182 (
            .O(N__76189),
            .I(N__76119));
    Span12Mux_v I__17181 (
            .O(N__76186),
            .I(N__76119));
    Sp12to4 I__17180 (
            .O(N__76181),
            .I(N__76119));
    LocalMux I__17179 (
            .O(N__76178),
            .I(N__76119));
    LocalMux I__17178 (
            .O(N__76175),
            .I(N__76119));
    LocalMux I__17177 (
            .O(N__76172),
            .I(N__76119));
    Span4Mux_v I__17176 (
            .O(N__76167),
            .I(N__76112));
    Span4Mux_v I__17175 (
            .O(N__76162),
            .I(N__76112));
    Span4Mux_h I__17174 (
            .O(N__76159),
            .I(N__76112));
    Span4Mux_v I__17173 (
            .O(N__76156),
            .I(N__76105));
    Span4Mux_v I__17172 (
            .O(N__76153),
            .I(N__76105));
    LocalMux I__17171 (
            .O(N__76150),
            .I(N__76105));
    Span4Mux_v I__17170 (
            .O(N__76145),
            .I(N__76098));
    Span4Mux_v I__17169 (
            .O(N__76138),
            .I(N__76098));
    LocalMux I__17168 (
            .O(N__76135),
            .I(N__76098));
    InMux I__17167 (
            .O(N__76134),
            .I(N__76095));
    Odrv12 I__17166 (
            .O(N__76119),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n49 ));
    Odrv4 I__17165 (
            .O(N__76112),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n49 ));
    Odrv4 I__17164 (
            .O(N__76105),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n49 ));
    Odrv4 I__17163 (
            .O(N__76098),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n49 ));
    LocalMux I__17162 (
            .O(N__76095),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n49 ));
    CascadeMux I__17161 (
            .O(N__76084),
            .I(N__76080));
    CascadeMux I__17160 (
            .O(N__76083),
            .I(N__76077));
    InMux I__17159 (
            .O(N__76080),
            .I(N__76072));
    InMux I__17158 (
            .O(N__76077),
            .I(N__76072));
    LocalMux I__17157 (
            .O(N__76072),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_8 ));
    InMux I__17156 (
            .O(N__76069),
            .I(N__76066));
    LocalMux I__17155 (
            .O(N__76066),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14372 ));
    InMux I__17154 (
            .O(N__76063),
            .I(N__76060));
    LocalMux I__17153 (
            .O(N__76060),
            .I(N__76057));
    Span4Mux_h I__17152 (
            .O(N__76057),
            .I(N__76053));
    CascadeMux I__17151 (
            .O(N__76056),
            .I(N__76050));
    Span4Mux_h I__17150 (
            .O(N__76053),
            .I(N__76047));
    InMux I__17149 (
            .O(N__76050),
            .I(N__76044));
    Odrv4 I__17148 (
            .O(N__76047),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_6 ));
    LocalMux I__17147 (
            .O(N__76044),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_6 ));
    InMux I__17146 (
            .O(N__76039),
            .I(N__76036));
    LocalMux I__17145 (
            .O(N__76036),
            .I(N__76033));
    Odrv4 I__17144 (
            .O(N__76033),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12474 ));
    CascadeMux I__17143 (
            .O(N__76030),
            .I(N__76026));
    InMux I__17142 (
            .O(N__76029),
            .I(N__76021));
    InMux I__17141 (
            .O(N__76026),
            .I(N__76021));
    LocalMux I__17140 (
            .O(N__76021),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_2 ));
    CascadeMux I__17139 (
            .O(N__76018),
            .I(N__76014));
    CascadeMux I__17138 (
            .O(N__76017),
            .I(N__76011));
    InMux I__17137 (
            .O(N__76014),
            .I(N__76006));
    InMux I__17136 (
            .O(N__76011),
            .I(N__76006));
    LocalMux I__17135 (
            .O(N__76006),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_2 ));
    InMux I__17134 (
            .O(N__76003),
            .I(N__76000));
    LocalMux I__17133 (
            .O(N__76000),
            .I(N__75995));
    CascadeMux I__17132 (
            .O(N__75999),
            .I(N__75992));
    InMux I__17131 (
            .O(N__75998),
            .I(N__75989));
    Span4Mux_v I__17130 (
            .O(N__75995),
            .I(N__75983));
    InMux I__17129 (
            .O(N__75992),
            .I(N__75980));
    LocalMux I__17128 (
            .O(N__75989),
            .I(N__75977));
    InMux I__17127 (
            .O(N__75988),
            .I(N__75968));
    InMux I__17126 (
            .O(N__75987),
            .I(N__75951));
    InMux I__17125 (
            .O(N__75986),
            .I(N__75948));
    Span4Mux_h I__17124 (
            .O(N__75983),
            .I(N__75943));
    LocalMux I__17123 (
            .O(N__75980),
            .I(N__75943));
    Span4Mux_v I__17122 (
            .O(N__75977),
            .I(N__75916));
    InMux I__17121 (
            .O(N__75976),
            .I(N__75911));
    InMux I__17120 (
            .O(N__75975),
            .I(N__75911));
    InMux I__17119 (
            .O(N__75974),
            .I(N__75906));
    InMux I__17118 (
            .O(N__75973),
            .I(N__75906));
    InMux I__17117 (
            .O(N__75972),
            .I(N__75898));
    InMux I__17116 (
            .O(N__75971),
            .I(N__75898));
    LocalMux I__17115 (
            .O(N__75968),
            .I(N__75893));
    InMux I__17114 (
            .O(N__75967),
            .I(N__75888));
    InMux I__17113 (
            .O(N__75966),
            .I(N__75888));
    InMux I__17112 (
            .O(N__75965),
            .I(N__75885));
    InMux I__17111 (
            .O(N__75964),
            .I(N__75876));
    InMux I__17110 (
            .O(N__75963),
            .I(N__75876));
    InMux I__17109 (
            .O(N__75962),
            .I(N__75876));
    InMux I__17108 (
            .O(N__75961),
            .I(N__75876));
    CascadeMux I__17107 (
            .O(N__75960),
            .I(N__75872));
    CascadeMux I__17106 (
            .O(N__75959),
            .I(N__75869));
    CascadeMux I__17105 (
            .O(N__75958),
            .I(N__75866));
    InMux I__17104 (
            .O(N__75957),
            .I(N__75859));
    InMux I__17103 (
            .O(N__75956),
            .I(N__75859));
    InMux I__17102 (
            .O(N__75955),
            .I(N__75856));
    InMux I__17101 (
            .O(N__75954),
            .I(N__75853));
    LocalMux I__17100 (
            .O(N__75951),
            .I(N__75846));
    LocalMux I__17099 (
            .O(N__75948),
            .I(N__75846));
    Span4Mux_h I__17098 (
            .O(N__75943),
            .I(N__75846));
    InMux I__17097 (
            .O(N__75942),
            .I(N__75841));
    InMux I__17096 (
            .O(N__75941),
            .I(N__75841));
    InMux I__17095 (
            .O(N__75940),
            .I(N__75836));
    InMux I__17094 (
            .O(N__75939),
            .I(N__75836));
    InMux I__17093 (
            .O(N__75938),
            .I(N__75827));
    InMux I__17092 (
            .O(N__75937),
            .I(N__75827));
    InMux I__17091 (
            .O(N__75936),
            .I(N__75827));
    InMux I__17090 (
            .O(N__75935),
            .I(N__75827));
    InMux I__17089 (
            .O(N__75934),
            .I(N__75822));
    InMux I__17088 (
            .O(N__75933),
            .I(N__75822));
    InMux I__17087 (
            .O(N__75932),
            .I(N__75816));
    InMux I__17086 (
            .O(N__75931),
            .I(N__75807));
    InMux I__17085 (
            .O(N__75930),
            .I(N__75807));
    InMux I__17084 (
            .O(N__75929),
            .I(N__75807));
    InMux I__17083 (
            .O(N__75928),
            .I(N__75807));
    InMux I__17082 (
            .O(N__75927),
            .I(N__75791));
    InMux I__17081 (
            .O(N__75926),
            .I(N__75791));
    InMux I__17080 (
            .O(N__75925),
            .I(N__75791));
    InMux I__17079 (
            .O(N__75924),
            .I(N__75791));
    InMux I__17078 (
            .O(N__75923),
            .I(N__75791));
    InMux I__17077 (
            .O(N__75922),
            .I(N__75791));
    InMux I__17076 (
            .O(N__75921),
            .I(N__75786));
    InMux I__17075 (
            .O(N__75920),
            .I(N__75786));
    InMux I__17074 (
            .O(N__75919),
            .I(N__75783));
    Span4Mux_h I__17073 (
            .O(N__75916),
            .I(N__75778));
    LocalMux I__17072 (
            .O(N__75911),
            .I(N__75778));
    LocalMux I__17071 (
            .O(N__75906),
            .I(N__75775));
    InMux I__17070 (
            .O(N__75905),
            .I(N__75768));
    InMux I__17069 (
            .O(N__75904),
            .I(N__75768));
    InMux I__17068 (
            .O(N__75903),
            .I(N__75768));
    LocalMux I__17067 (
            .O(N__75898),
            .I(N__75765));
    InMux I__17066 (
            .O(N__75897),
            .I(N__75762));
    InMux I__17065 (
            .O(N__75896),
            .I(N__75759));
    Span4Mux_h I__17064 (
            .O(N__75893),
            .I(N__75750));
    LocalMux I__17063 (
            .O(N__75888),
            .I(N__75750));
    LocalMux I__17062 (
            .O(N__75885),
            .I(N__75750));
    LocalMux I__17061 (
            .O(N__75876),
            .I(N__75750));
    InMux I__17060 (
            .O(N__75875),
            .I(N__75739));
    InMux I__17059 (
            .O(N__75872),
            .I(N__75739));
    InMux I__17058 (
            .O(N__75869),
            .I(N__75739));
    InMux I__17057 (
            .O(N__75866),
            .I(N__75739));
    InMux I__17056 (
            .O(N__75865),
            .I(N__75739));
    InMux I__17055 (
            .O(N__75864),
            .I(N__75736));
    LocalMux I__17054 (
            .O(N__75859),
            .I(N__75733));
    LocalMux I__17053 (
            .O(N__75856),
            .I(N__75722));
    LocalMux I__17052 (
            .O(N__75853),
            .I(N__75722));
    Span4Mux_v I__17051 (
            .O(N__75846),
            .I(N__75722));
    LocalMux I__17050 (
            .O(N__75841),
            .I(N__75722));
    LocalMux I__17049 (
            .O(N__75836),
            .I(N__75722));
    LocalMux I__17048 (
            .O(N__75827),
            .I(N__75717));
    LocalMux I__17047 (
            .O(N__75822),
            .I(N__75717));
    InMux I__17046 (
            .O(N__75821),
            .I(N__75714));
    InMux I__17045 (
            .O(N__75820),
            .I(N__75711));
    InMux I__17044 (
            .O(N__75819),
            .I(N__75708));
    LocalMux I__17043 (
            .O(N__75816),
            .I(N__75705));
    LocalMux I__17042 (
            .O(N__75807),
            .I(N__75702));
    InMux I__17041 (
            .O(N__75806),
            .I(N__75699));
    InMux I__17040 (
            .O(N__75805),
            .I(N__75694));
    InMux I__17039 (
            .O(N__75804),
            .I(N__75694));
    LocalMux I__17038 (
            .O(N__75791),
            .I(N__75689));
    LocalMux I__17037 (
            .O(N__75786),
            .I(N__75689));
    LocalMux I__17036 (
            .O(N__75783),
            .I(N__75686));
    Sp12to4 I__17035 (
            .O(N__75778),
            .I(N__75681));
    Sp12to4 I__17034 (
            .O(N__75775),
            .I(N__75681));
    LocalMux I__17033 (
            .O(N__75768),
            .I(N__75674));
    Span4Mux_h I__17032 (
            .O(N__75765),
            .I(N__75674));
    LocalMux I__17031 (
            .O(N__75762),
            .I(N__75674));
    LocalMux I__17030 (
            .O(N__75759),
            .I(N__75667));
    Span4Mux_v I__17029 (
            .O(N__75750),
            .I(N__75667));
    LocalMux I__17028 (
            .O(N__75739),
            .I(N__75667));
    LocalMux I__17027 (
            .O(N__75736),
            .I(N__75660));
    Span4Mux_v I__17026 (
            .O(N__75733),
            .I(N__75660));
    Span4Mux_v I__17025 (
            .O(N__75722),
            .I(N__75660));
    Span4Mux_v I__17024 (
            .O(N__75717),
            .I(N__75657));
    LocalMux I__17023 (
            .O(N__75714),
            .I(N__75652));
    LocalMux I__17022 (
            .O(N__75711),
            .I(N__75652));
    LocalMux I__17021 (
            .O(N__75708),
            .I(N__75645));
    Span4Mux_h I__17020 (
            .O(N__75705),
            .I(N__75645));
    Span4Mux_h I__17019 (
            .O(N__75702),
            .I(N__75645));
    LocalMux I__17018 (
            .O(N__75699),
            .I(N__75638));
    LocalMux I__17017 (
            .O(N__75694),
            .I(N__75638));
    Span4Mux_v I__17016 (
            .O(N__75689),
            .I(N__75638));
    Span12Mux_h I__17015 (
            .O(N__75686),
            .I(N__75635));
    Span12Mux_v I__17014 (
            .O(N__75681),
            .I(N__75632));
    Span4Mux_v I__17013 (
            .O(N__75674),
            .I(N__75623));
    Span4Mux_v I__17012 (
            .O(N__75667),
            .I(N__75623));
    Span4Mux_h I__17011 (
            .O(N__75660),
            .I(N__75623));
    Span4Mux_v I__17010 (
            .O(N__75657),
            .I(N__75623));
    Odrv12 I__17009 (
            .O(N__75652),
            .I(dc32_fifo_data_in_2));
    Odrv4 I__17008 (
            .O(N__75645),
            .I(dc32_fifo_data_in_2));
    Odrv4 I__17007 (
            .O(N__75638),
            .I(dc32_fifo_data_in_2));
    Odrv12 I__17006 (
            .O(N__75635),
            .I(dc32_fifo_data_in_2));
    Odrv12 I__17005 (
            .O(N__75632),
            .I(dc32_fifo_data_in_2));
    Odrv4 I__17004 (
            .O(N__75623),
            .I(dc32_fifo_data_in_2));
    InMux I__17003 (
            .O(N__75610),
            .I(N__75607));
    LocalMux I__17002 (
            .O(N__75607),
            .I(N__75603));
    CascadeMux I__17001 (
            .O(N__75606),
            .I(N__75600));
    Span4Mux_h I__17000 (
            .O(N__75603),
            .I(N__75597));
    InMux I__16999 (
            .O(N__75600),
            .I(N__75594));
    Odrv4 I__16998 (
            .O(N__75597),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_2 ));
    LocalMux I__16997 (
            .O(N__75594),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_2 ));
    InMux I__16996 (
            .O(N__75589),
            .I(N__75585));
    InMux I__16995 (
            .O(N__75588),
            .I(N__75581));
    LocalMux I__16994 (
            .O(N__75585),
            .I(N__75573));
    InMux I__16993 (
            .O(N__75584),
            .I(N__75569));
    LocalMux I__16992 (
            .O(N__75581),
            .I(N__75563));
    InMux I__16991 (
            .O(N__75580),
            .I(N__75560));
    InMux I__16990 (
            .O(N__75579),
            .I(N__75555));
    InMux I__16989 (
            .O(N__75578),
            .I(N__75552));
    InMux I__16988 (
            .O(N__75577),
            .I(N__75549));
    InMux I__16987 (
            .O(N__75576),
            .I(N__75546));
    Span4Mux_v I__16986 (
            .O(N__75573),
            .I(N__75543));
    InMux I__16985 (
            .O(N__75572),
            .I(N__75540));
    LocalMux I__16984 (
            .O(N__75569),
            .I(N__75537));
    InMux I__16983 (
            .O(N__75568),
            .I(N__75534));
    InMux I__16982 (
            .O(N__75567),
            .I(N__75531));
    InMux I__16981 (
            .O(N__75566),
            .I(N__75528));
    Span4Mux_h I__16980 (
            .O(N__75563),
            .I(N__75523));
    LocalMux I__16979 (
            .O(N__75560),
            .I(N__75523));
    InMux I__16978 (
            .O(N__75559),
            .I(N__75520));
    InMux I__16977 (
            .O(N__75558),
            .I(N__75517));
    LocalMux I__16976 (
            .O(N__75555),
            .I(N__75514));
    LocalMux I__16975 (
            .O(N__75552),
            .I(N__75510));
    LocalMux I__16974 (
            .O(N__75549),
            .I(N__75507));
    LocalMux I__16973 (
            .O(N__75546),
            .I(N__75504));
    Span4Mux_h I__16972 (
            .O(N__75543),
            .I(N__75499));
    LocalMux I__16971 (
            .O(N__75540),
            .I(N__75499));
    Span4Mux_v I__16970 (
            .O(N__75537),
            .I(N__75494));
    LocalMux I__16969 (
            .O(N__75534),
            .I(N__75494));
    LocalMux I__16968 (
            .O(N__75531),
            .I(N__75491));
    LocalMux I__16967 (
            .O(N__75528),
            .I(N__75488));
    Span4Mux_h I__16966 (
            .O(N__75523),
            .I(N__75483));
    LocalMux I__16965 (
            .O(N__75520),
            .I(N__75483));
    LocalMux I__16964 (
            .O(N__75517),
            .I(N__75480));
    Span4Mux_h I__16963 (
            .O(N__75514),
            .I(N__75477));
    InMux I__16962 (
            .O(N__75513),
            .I(N__75474));
    Sp12to4 I__16961 (
            .O(N__75510),
            .I(N__75470));
    Span4Mux_h I__16960 (
            .O(N__75507),
            .I(N__75467));
    Span4Mux_h I__16959 (
            .O(N__75504),
            .I(N__75464));
    Span4Mux_h I__16958 (
            .O(N__75499),
            .I(N__75461));
    Span4Mux_v I__16957 (
            .O(N__75494),
            .I(N__75456));
    Span4Mux_h I__16956 (
            .O(N__75491),
            .I(N__75456));
    Span4Mux_h I__16955 (
            .O(N__75488),
            .I(N__75449));
    Span4Mux_h I__16954 (
            .O(N__75483),
            .I(N__75449));
    Span4Mux_v I__16953 (
            .O(N__75480),
            .I(N__75449));
    Span4Mux_v I__16952 (
            .O(N__75477),
            .I(N__75444));
    LocalMux I__16951 (
            .O(N__75474),
            .I(N__75444));
    InMux I__16950 (
            .O(N__75473),
            .I(N__75441));
    Odrv12 I__16949 (
            .O(N__75470),
            .I(n17));
    Odrv4 I__16948 (
            .O(N__75467),
            .I(n17));
    Odrv4 I__16947 (
            .O(N__75464),
            .I(n17));
    Odrv4 I__16946 (
            .O(N__75461),
            .I(n17));
    Odrv4 I__16945 (
            .O(N__75456),
            .I(n17));
    Odrv4 I__16944 (
            .O(N__75449),
            .I(n17));
    Odrv4 I__16943 (
            .O(N__75444),
            .I(n17));
    LocalMux I__16942 (
            .O(N__75441),
            .I(n17));
    InMux I__16941 (
            .O(N__75424),
            .I(N__75421));
    LocalMux I__16940 (
            .O(N__75421),
            .I(N__75417));
    InMux I__16939 (
            .O(N__75420),
            .I(N__75414));
    Odrv4 I__16938 (
            .O(N__75417),
            .I(REG_mem_48_6));
    LocalMux I__16937 (
            .O(N__75414),
            .I(REG_mem_48_6));
    InMux I__16936 (
            .O(N__75409),
            .I(N__75405));
    InMux I__16935 (
            .O(N__75408),
            .I(N__75402));
    LocalMux I__16934 (
            .O(N__75405),
            .I(REG_mem_44_6));
    LocalMux I__16933 (
            .O(N__75402),
            .I(REG_mem_44_6));
    CascadeMux I__16932 (
            .O(N__75397),
            .I(N__75394));
    InMux I__16931 (
            .O(N__75394),
            .I(N__75391));
    LocalMux I__16930 (
            .O(N__75391),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13388 ));
    InMux I__16929 (
            .O(N__75388),
            .I(N__75384));
    InMux I__16928 (
            .O(N__75387),
            .I(N__75381));
    LocalMux I__16927 (
            .O(N__75384),
            .I(REG_mem_45_6));
    LocalMux I__16926 (
            .O(N__75381),
            .I(REG_mem_45_6));
    InMux I__16925 (
            .O(N__75376),
            .I(N__75372));
    InMux I__16924 (
            .O(N__75375),
            .I(N__75369));
    LocalMux I__16923 (
            .O(N__75372),
            .I(N__75366));
    LocalMux I__16922 (
            .O(N__75369),
            .I(REG_mem_55_4));
    Odrv4 I__16921 (
            .O(N__75366),
            .I(REG_mem_55_4));
    CascadeMux I__16920 (
            .O(N__75361),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14216_cascade_ ));
    InMux I__16919 (
            .O(N__75358),
            .I(N__75355));
    LocalMux I__16918 (
            .O(N__75355),
            .I(N__75352));
    Odrv4 I__16917 (
            .O(N__75352),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12054 ));
    InMux I__16916 (
            .O(N__75349),
            .I(N__75345));
    InMux I__16915 (
            .O(N__75348),
            .I(N__75342));
    LocalMux I__16914 (
            .O(N__75345),
            .I(REG_mem_23_6));
    LocalMux I__16913 (
            .O(N__75342),
            .I(REG_mem_23_6));
    CascadeMux I__16912 (
            .O(N__75337),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13646_cascade_ ));
    CascadeMux I__16911 (
            .O(N__75334),
            .I(N__75331));
    InMux I__16910 (
            .O(N__75331),
            .I(N__75327));
    InMux I__16909 (
            .O(N__75330),
            .I(N__75324));
    LocalMux I__16908 (
            .O(N__75327),
            .I(N__75321));
    LocalMux I__16907 (
            .O(N__75324),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_6 ));
    Odrv4 I__16906 (
            .O(N__75321),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_6 ));
    CascadeMux I__16905 (
            .O(N__75316),
            .I(N__75312));
    InMux I__16904 (
            .O(N__75315),
            .I(N__75307));
    InMux I__16903 (
            .O(N__75312),
            .I(N__75307));
    LocalMux I__16902 (
            .O(N__75307),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_6 ));
    CascadeMux I__16901 (
            .O(N__75304),
            .I(N__75300));
    InMux I__16900 (
            .O(N__75303),
            .I(N__75295));
    InMux I__16899 (
            .O(N__75300),
            .I(N__75295));
    LocalMux I__16898 (
            .O(N__75295),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_6 ));
    CascadeMux I__16897 (
            .O(N__75292),
            .I(N__75288));
    InMux I__16896 (
            .O(N__75291),
            .I(N__75285));
    InMux I__16895 (
            .O(N__75288),
            .I(N__75282));
    LocalMux I__16894 (
            .O(N__75285),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_6 ));
    LocalMux I__16893 (
            .O(N__75282),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_6 ));
    CascadeMux I__16892 (
            .O(N__75277),
            .I(N__75273));
    InMux I__16891 (
            .O(N__75276),
            .I(N__75270));
    InMux I__16890 (
            .O(N__75273),
            .I(N__75267));
    LocalMux I__16889 (
            .O(N__75270),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_6 ));
    LocalMux I__16888 (
            .O(N__75267),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_6 ));
    InMux I__16887 (
            .O(N__75262),
            .I(N__75256));
    InMux I__16886 (
            .O(N__75261),
            .I(N__75256));
    LocalMux I__16885 (
            .O(N__75256),
            .I(REG_mem_58_2));
    CascadeMux I__16884 (
            .O(N__75253),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13730_cascade_ ));
    CascadeMux I__16883 (
            .O(N__75250),
            .I(N__75246));
    InMux I__16882 (
            .O(N__75249),
            .I(N__75243));
    InMux I__16881 (
            .O(N__75246),
            .I(N__75240));
    LocalMux I__16880 (
            .O(N__75243),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_2 ));
    LocalMux I__16879 (
            .O(N__75240),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_2 ));
    InMux I__16878 (
            .O(N__75235),
            .I(N__75232));
    LocalMux I__16877 (
            .O(N__75232),
            .I(N__75229));
    Span4Mux_h I__16876 (
            .O(N__75229),
            .I(N__75226));
    Odrv4 I__16875 (
            .O(N__75226),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13733 ));
    InMux I__16874 (
            .O(N__75223),
            .I(N__75219));
    InMux I__16873 (
            .O(N__75222),
            .I(N__75216));
    LocalMux I__16872 (
            .O(N__75219),
            .I(N__75213));
    LocalMux I__16871 (
            .O(N__75216),
            .I(N__75210));
    Odrv4 I__16870 (
            .O(N__75213),
            .I(REG_mem_40_6));
    Odrv4 I__16869 (
            .O(N__75210),
            .I(REG_mem_40_6));
    InMux I__16868 (
            .O(N__75205),
            .I(N__75202));
    LocalMux I__16867 (
            .O(N__75202),
            .I(N__75198));
    InMux I__16866 (
            .O(N__75201),
            .I(N__75195));
    Odrv4 I__16865 (
            .O(N__75198),
            .I(REG_mem_51_6));
    LocalMux I__16864 (
            .O(N__75195),
            .I(REG_mem_51_6));
    InMux I__16863 (
            .O(N__75190),
            .I(N__75186));
    InMux I__16862 (
            .O(N__75189),
            .I(N__75183));
    LocalMux I__16861 (
            .O(N__75186),
            .I(REG_mem_50_6));
    LocalMux I__16860 (
            .O(N__75183),
            .I(REG_mem_50_6));
    CascadeMux I__16859 (
            .O(N__75178),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12782_cascade_ ));
    InMux I__16858 (
            .O(N__75175),
            .I(N__75172));
    LocalMux I__16857 (
            .O(N__75172),
            .I(N__75169));
    Span4Mux_v I__16856 (
            .O(N__75169),
            .I(N__75165));
    InMux I__16855 (
            .O(N__75168),
            .I(N__75162));
    Span4Mux_h I__16854 (
            .O(N__75165),
            .I(N__75159));
    LocalMux I__16853 (
            .O(N__75162),
            .I(N__75156));
    Odrv4 I__16852 (
            .O(N__75159),
            .I(REG_mem_49_6));
    Odrv4 I__16851 (
            .O(N__75156),
            .I(REG_mem_49_6));
    InMux I__16850 (
            .O(N__75151),
            .I(N__75148));
    LocalMux I__16849 (
            .O(N__75148),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12785 ));
    InMux I__16848 (
            .O(N__75145),
            .I(N__75142));
    LocalMux I__16847 (
            .O(N__75142),
            .I(N__75138));
    CascadeMux I__16846 (
            .O(N__75141),
            .I(N__75135));
    Span4Mux_v I__16845 (
            .O(N__75138),
            .I(N__75132));
    InMux I__16844 (
            .O(N__75135),
            .I(N__75129));
    Odrv4 I__16843 (
            .O(N__75132),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_4 ));
    LocalMux I__16842 (
            .O(N__75129),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_4 ));
    CascadeMux I__16841 (
            .O(N__75124),
            .I(N__75121));
    InMux I__16840 (
            .O(N__75121),
            .I(N__75118));
    LocalMux I__16839 (
            .O(N__75118),
            .I(N__75114));
    CascadeMux I__16838 (
            .O(N__75117),
            .I(N__75111));
    Span12Mux_h I__16837 (
            .O(N__75114),
            .I(N__75108));
    InMux I__16836 (
            .O(N__75111),
            .I(N__75105));
    Odrv12 I__16835 (
            .O(N__75108),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_6 ));
    LocalMux I__16834 (
            .O(N__75105),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_6 ));
    CascadeMux I__16833 (
            .O(N__75100),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14390_cascade_ ));
    CascadeMux I__16832 (
            .O(N__75097),
            .I(N__75094));
    InMux I__16831 (
            .O(N__75094),
            .I(N__75091));
    LocalMux I__16830 (
            .O(N__75091),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12459 ));
    InMux I__16829 (
            .O(N__75088),
            .I(N__75085));
    LocalMux I__16828 (
            .O(N__75085),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11634 ));
    InMux I__16827 (
            .O(N__75082),
            .I(N__75079));
    LocalMux I__16826 (
            .O(N__75079),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13004 ));
    InMux I__16825 (
            .O(N__75076),
            .I(N__75070));
    InMux I__16824 (
            .O(N__75075),
            .I(N__75070));
    LocalMux I__16823 (
            .O(N__75070),
            .I(REG_mem_55_6));
    InMux I__16822 (
            .O(N__75067),
            .I(N__75061));
    InMux I__16821 (
            .O(N__75066),
            .I(N__75058));
    InMux I__16820 (
            .O(N__75065),
            .I(N__75055));
    InMux I__16819 (
            .O(N__75064),
            .I(N__75052));
    LocalMux I__16818 (
            .O(N__75061),
            .I(N__75045));
    LocalMux I__16817 (
            .O(N__75058),
            .I(N__75042));
    LocalMux I__16816 (
            .O(N__75055),
            .I(N__75036));
    LocalMux I__16815 (
            .O(N__75052),
            .I(N__75033));
    InMux I__16814 (
            .O(N__75051),
            .I(N__75030));
    InMux I__16813 (
            .O(N__75050),
            .I(N__75027));
    InMux I__16812 (
            .O(N__75049),
            .I(N__75024));
    InMux I__16811 (
            .O(N__75048),
            .I(N__75021));
    Span4Mux_v I__16810 (
            .O(N__75045),
            .I(N__75016));
    Span4Mux_h I__16809 (
            .O(N__75042),
            .I(N__75013));
    InMux I__16808 (
            .O(N__75041),
            .I(N__75009));
    InMux I__16807 (
            .O(N__75040),
            .I(N__75006));
    InMux I__16806 (
            .O(N__75039),
            .I(N__75003));
    Span4Mux_h I__16805 (
            .O(N__75036),
            .I(N__74999));
    Span4Mux_h I__16804 (
            .O(N__75033),
            .I(N__74992));
    LocalMux I__16803 (
            .O(N__75030),
            .I(N__74992));
    LocalMux I__16802 (
            .O(N__75027),
            .I(N__74992));
    LocalMux I__16801 (
            .O(N__75024),
            .I(N__74989));
    LocalMux I__16800 (
            .O(N__75021),
            .I(N__74986));
    InMux I__16799 (
            .O(N__75020),
            .I(N__74983));
    InMux I__16798 (
            .O(N__75019),
            .I(N__74980));
    Span4Mux_h I__16797 (
            .O(N__75016),
            .I(N__74975));
    Span4Mux_v I__16796 (
            .O(N__75013),
            .I(N__74975));
    InMux I__16795 (
            .O(N__75012),
            .I(N__74972));
    LocalMux I__16794 (
            .O(N__75009),
            .I(N__74965));
    LocalMux I__16793 (
            .O(N__75006),
            .I(N__74965));
    LocalMux I__16792 (
            .O(N__75003),
            .I(N__74965));
    InMux I__16791 (
            .O(N__75002),
            .I(N__74962));
    Span4Mux_v I__16790 (
            .O(N__74999),
            .I(N__74958));
    Span4Mux_v I__16789 (
            .O(N__74992),
            .I(N__74955));
    Span4Mux_h I__16788 (
            .O(N__74989),
            .I(N__74952));
    Span12Mux_h I__16787 (
            .O(N__74986),
            .I(N__74945));
    LocalMux I__16786 (
            .O(N__74983),
            .I(N__74945));
    LocalMux I__16785 (
            .O(N__74980),
            .I(N__74945));
    Sp12to4 I__16784 (
            .O(N__74975),
            .I(N__74936));
    LocalMux I__16783 (
            .O(N__74972),
            .I(N__74936));
    Span12Mux_v I__16782 (
            .O(N__74965),
            .I(N__74936));
    LocalMux I__16781 (
            .O(N__74962),
            .I(N__74936));
    InMux I__16780 (
            .O(N__74961),
            .I(N__74933));
    Odrv4 I__16779 (
            .O(N__74958),
            .I(n42));
    Odrv4 I__16778 (
            .O(N__74955),
            .I(n42));
    Odrv4 I__16777 (
            .O(N__74952),
            .I(n42));
    Odrv12 I__16776 (
            .O(N__74945),
            .I(n42));
    Odrv12 I__16775 (
            .O(N__74936),
            .I(n42));
    LocalMux I__16774 (
            .O(N__74933),
            .I(n42));
    InMux I__16773 (
            .O(N__74920),
            .I(N__74917));
    LocalMux I__16772 (
            .O(N__74917),
            .I(N__74914));
    Odrv4 I__16771 (
            .O(N__74914),
            .I(n11410));
    CascadeMux I__16770 (
            .O(N__74911),
            .I(n4_adj_1186_cascade_));
    InMux I__16769 (
            .O(N__74908),
            .I(N__74905));
    LocalMux I__16768 (
            .O(N__74905),
            .I(N__74902));
    Odrv4 I__16767 (
            .O(N__74902),
            .I(n24));
    InMux I__16766 (
            .O(N__74899),
            .I(N__74895));
    InMux I__16765 (
            .O(N__74898),
            .I(N__74888));
    LocalMux I__16764 (
            .O(N__74895),
            .I(N__74885));
    InMux I__16763 (
            .O(N__74894),
            .I(N__74876));
    InMux I__16762 (
            .O(N__74893),
            .I(N__74876));
    InMux I__16761 (
            .O(N__74892),
            .I(N__74876));
    InMux I__16760 (
            .O(N__74891),
            .I(N__74876));
    LocalMux I__16759 (
            .O(N__74888),
            .I(N__74870));
    Span4Mux_v I__16758 (
            .O(N__74885),
            .I(N__74865));
    LocalMux I__16757 (
            .O(N__74876),
            .I(N__74865));
    InMux I__16756 (
            .O(N__74875),
            .I(N__74862));
    InMux I__16755 (
            .O(N__74874),
            .I(N__74857));
    InMux I__16754 (
            .O(N__74873),
            .I(N__74857));
    Odrv12 I__16753 (
            .O(N__74870),
            .I(is_fifo_empty_flag));
    Odrv4 I__16752 (
            .O(N__74865),
            .I(is_fifo_empty_flag));
    LocalMux I__16751 (
            .O(N__74862),
            .I(is_fifo_empty_flag));
    LocalMux I__16750 (
            .O(N__74857),
            .I(is_fifo_empty_flag));
    InMux I__16749 (
            .O(N__74848),
            .I(N__74845));
    LocalMux I__16748 (
            .O(N__74845),
            .I(N__74842));
    Span12Mux_h I__16747 (
            .O(N__74842),
            .I(N__74838));
    InMux I__16746 (
            .O(N__74841),
            .I(N__74835));
    Odrv12 I__16745 (
            .O(N__74838),
            .I(REG_mem_12_6));
    LocalMux I__16744 (
            .O(N__74835),
            .I(REG_mem_12_6));
    CascadeMux I__16743 (
            .O(N__74830),
            .I(N__74827));
    InMux I__16742 (
            .O(N__74827),
            .I(N__74823));
    InMux I__16741 (
            .O(N__74826),
            .I(N__74820));
    LocalMux I__16740 (
            .O(N__74823),
            .I(REG_mem_13_6));
    LocalMux I__16739 (
            .O(N__74820),
            .I(REG_mem_13_6));
    CascadeMux I__16738 (
            .O(N__74815),
            .I(N__74812));
    InMux I__16737 (
            .O(N__74812),
            .I(N__74809));
    LocalMux I__16736 (
            .O(N__74809),
            .I(N__74806));
    Span4Mux_v I__16735 (
            .O(N__74806),
            .I(N__74803));
    Span4Mux_v I__16734 (
            .O(N__74803),
            .I(N__74799));
    InMux I__16733 (
            .O(N__74802),
            .I(N__74796));
    Odrv4 I__16732 (
            .O(N__74799),
            .I(REG_mem_15_6));
    LocalMux I__16731 (
            .O(N__74796),
            .I(REG_mem_15_6));
    InMux I__16730 (
            .O(N__74791),
            .I(N__74788));
    LocalMux I__16729 (
            .O(N__74788),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13772 ));
    CascadeMux I__16728 (
            .O(N__74785),
            .I(N__74781));
    InMux I__16727 (
            .O(N__74784),
            .I(N__74778));
    InMux I__16726 (
            .O(N__74781),
            .I(N__74775));
    LocalMux I__16725 (
            .O(N__74778),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_8 ));
    LocalMux I__16724 (
            .O(N__74775),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_8 ));
    InMux I__16723 (
            .O(N__74770),
            .I(N__74766));
    InMux I__16722 (
            .O(N__74769),
            .I(N__74758));
    LocalMux I__16721 (
            .O(N__74766),
            .I(N__74754));
    InMux I__16720 (
            .O(N__74765),
            .I(N__74750));
    InMux I__16719 (
            .O(N__74764),
            .I(N__74746));
    InMux I__16718 (
            .O(N__74763),
            .I(N__74742));
    InMux I__16717 (
            .O(N__74762),
            .I(N__74738));
    InMux I__16716 (
            .O(N__74761),
            .I(N__74735));
    LocalMux I__16715 (
            .O(N__74758),
            .I(N__74732));
    InMux I__16714 (
            .O(N__74757),
            .I(N__74729));
    Span4Mux_h I__16713 (
            .O(N__74754),
            .I(N__74726));
    InMux I__16712 (
            .O(N__74753),
            .I(N__74723));
    LocalMux I__16711 (
            .O(N__74750),
            .I(N__74720));
    InMux I__16710 (
            .O(N__74749),
            .I(N__74717));
    LocalMux I__16709 (
            .O(N__74746),
            .I(N__74714));
    InMux I__16708 (
            .O(N__74745),
            .I(N__74711));
    LocalMux I__16707 (
            .O(N__74742),
            .I(N__74708));
    InMux I__16706 (
            .O(N__74741),
            .I(N__74705));
    LocalMux I__16705 (
            .O(N__74738),
            .I(N__74700));
    LocalMux I__16704 (
            .O(N__74735),
            .I(N__74697));
    Span4Mux_h I__16703 (
            .O(N__74732),
            .I(N__74692));
    LocalMux I__16702 (
            .O(N__74729),
            .I(N__74692));
    Span4Mux_v I__16701 (
            .O(N__74726),
            .I(N__74689));
    LocalMux I__16700 (
            .O(N__74723),
            .I(N__74686));
    Span4Mux_h I__16699 (
            .O(N__74720),
            .I(N__74681));
    LocalMux I__16698 (
            .O(N__74717),
            .I(N__74681));
    Span4Mux_h I__16697 (
            .O(N__74714),
            .I(N__74674));
    LocalMux I__16696 (
            .O(N__74711),
            .I(N__74674));
    Span4Mux_v I__16695 (
            .O(N__74708),
            .I(N__74669));
    LocalMux I__16694 (
            .O(N__74705),
            .I(N__74669));
    InMux I__16693 (
            .O(N__74704),
            .I(N__74666));
    InMux I__16692 (
            .O(N__74703),
            .I(N__74663));
    Span12Mux_v I__16691 (
            .O(N__74700),
            .I(N__74660));
    Span4Mux_h I__16690 (
            .O(N__74697),
            .I(N__74655));
    Span4Mux_v I__16689 (
            .O(N__74692),
            .I(N__74655));
    Span4Mux_h I__16688 (
            .O(N__74689),
            .I(N__74648));
    Span4Mux_v I__16687 (
            .O(N__74686),
            .I(N__74648));
    Span4Mux_h I__16686 (
            .O(N__74681),
            .I(N__74648));
    InMux I__16685 (
            .O(N__74680),
            .I(N__74643));
    InMux I__16684 (
            .O(N__74679),
            .I(N__74643));
    Span4Mux_h I__16683 (
            .O(N__74674),
            .I(N__74634));
    Span4Mux_v I__16682 (
            .O(N__74669),
            .I(N__74634));
    LocalMux I__16681 (
            .O(N__74666),
            .I(N__74634));
    LocalMux I__16680 (
            .O(N__74663),
            .I(N__74634));
    Odrv12 I__16679 (
            .O(N__74660),
            .I(n51));
    Odrv4 I__16678 (
            .O(N__74655),
            .I(n51));
    Odrv4 I__16677 (
            .O(N__74648),
            .I(n51));
    LocalMux I__16676 (
            .O(N__74643),
            .I(n51));
    Odrv4 I__16675 (
            .O(N__74634),
            .I(n51));
    InMux I__16674 (
            .O(N__74623),
            .I(N__74617));
    InMux I__16673 (
            .O(N__74622),
            .I(N__74617));
    LocalMux I__16672 (
            .O(N__74617),
            .I(REG_mem_14_6));
    CascadeMux I__16671 (
            .O(N__74614),
            .I(N__74611));
    InMux I__16670 (
            .O(N__74611),
            .I(N__74608));
    LocalMux I__16669 (
            .O(N__74608),
            .I(N__74604));
    InMux I__16668 (
            .O(N__74607),
            .I(N__74601));
    Odrv12 I__16667 (
            .O(N__74604),
            .I(REG_mem_43_6));
    LocalMux I__16666 (
            .O(N__74601),
            .I(REG_mem_43_6));
    InMux I__16665 (
            .O(N__74596),
            .I(N__74593));
    LocalMux I__16664 (
            .O(N__74593),
            .I(N__74590));
    Span4Mux_h I__16663 (
            .O(N__74590),
            .I(N__74587));
    Span4Mux_v I__16662 (
            .O(N__74587),
            .I(N__74583));
    InMux I__16661 (
            .O(N__74586),
            .I(N__74580));
    Odrv4 I__16660 (
            .O(N__74583),
            .I(REG_mem_42_6));
    LocalMux I__16659 (
            .O(N__74580),
            .I(REG_mem_42_6));
    InMux I__16658 (
            .O(N__74575),
            .I(N__74572));
    LocalMux I__16657 (
            .O(N__74572),
            .I(N__74568));
    InMux I__16656 (
            .O(N__74571),
            .I(N__74565));
    Odrv4 I__16655 (
            .O(N__74568),
            .I(REG_mem_41_6));
    LocalMux I__16654 (
            .O(N__74565),
            .I(REG_mem_41_6));
    CascadeMux I__16653 (
            .O(N__74560),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13520_cascade_ ));
    InMux I__16652 (
            .O(N__74557),
            .I(N__74551));
    InMux I__16651 (
            .O(N__74556),
            .I(N__74551));
    LocalMux I__16650 (
            .O(N__74551),
            .I(N__74525));
    InMux I__16649 (
            .O(N__74550),
            .I(N__74510));
    InMux I__16648 (
            .O(N__74549),
            .I(N__74510));
    InMux I__16647 (
            .O(N__74548),
            .I(N__74510));
    InMux I__16646 (
            .O(N__74547),
            .I(N__74510));
    InMux I__16645 (
            .O(N__74546),
            .I(N__74510));
    InMux I__16644 (
            .O(N__74545),
            .I(N__74510));
    InMux I__16643 (
            .O(N__74544),
            .I(N__74510));
    InMux I__16642 (
            .O(N__74543),
            .I(N__74507));
    InMux I__16641 (
            .O(N__74542),
            .I(N__74498));
    InMux I__16640 (
            .O(N__74541),
            .I(N__74498));
    InMux I__16639 (
            .O(N__74540),
            .I(N__74481));
    InMux I__16638 (
            .O(N__74539),
            .I(N__74481));
    InMux I__16637 (
            .O(N__74538),
            .I(N__74481));
    InMux I__16636 (
            .O(N__74537),
            .I(N__74481));
    InMux I__16635 (
            .O(N__74536),
            .I(N__74481));
    InMux I__16634 (
            .O(N__74535),
            .I(N__74481));
    InMux I__16633 (
            .O(N__74534),
            .I(N__74481));
    InMux I__16632 (
            .O(N__74533),
            .I(N__74481));
    InMux I__16631 (
            .O(N__74532),
            .I(N__74472));
    InMux I__16630 (
            .O(N__74531),
            .I(N__74472));
    InMux I__16629 (
            .O(N__74530),
            .I(N__74472));
    InMux I__16628 (
            .O(N__74529),
            .I(N__74472));
    CascadeMux I__16627 (
            .O(N__74528),
            .I(N__74468));
    Span4Mux_v I__16626 (
            .O(N__74525),
            .I(N__74461));
    LocalMux I__16625 (
            .O(N__74510),
            .I(N__74461));
    LocalMux I__16624 (
            .O(N__74507),
            .I(N__74458));
    InMux I__16623 (
            .O(N__74506),
            .I(N__74449));
    InMux I__16622 (
            .O(N__74505),
            .I(N__74449));
    InMux I__16621 (
            .O(N__74504),
            .I(N__74449));
    InMux I__16620 (
            .O(N__74503),
            .I(N__74449));
    LocalMux I__16619 (
            .O(N__74498),
            .I(N__74442));
    LocalMux I__16618 (
            .O(N__74481),
            .I(N__74442));
    LocalMux I__16617 (
            .O(N__74472),
            .I(N__74442));
    InMux I__16616 (
            .O(N__74471),
            .I(N__74433));
    InMux I__16615 (
            .O(N__74468),
            .I(N__74433));
    InMux I__16614 (
            .O(N__74467),
            .I(N__74433));
    InMux I__16613 (
            .O(N__74466),
            .I(N__74433));
    Span4Mux_v I__16612 (
            .O(N__74461),
            .I(N__74421));
    Span4Mux_v I__16611 (
            .O(N__74458),
            .I(N__74421));
    LocalMux I__16610 (
            .O(N__74449),
            .I(N__74418));
    Span4Mux_h I__16609 (
            .O(N__74442),
            .I(N__74413));
    LocalMux I__16608 (
            .O(N__74433),
            .I(N__74413));
    InMux I__16607 (
            .O(N__74432),
            .I(N__74408));
    InMux I__16606 (
            .O(N__74431),
            .I(N__74408));
    InMux I__16605 (
            .O(N__74430),
            .I(N__74401));
    InMux I__16604 (
            .O(N__74429),
            .I(N__74401));
    InMux I__16603 (
            .O(N__74428),
            .I(N__74401));
    InMux I__16602 (
            .O(N__74427),
            .I(N__74396));
    InMux I__16601 (
            .O(N__74426),
            .I(N__74396));
    Odrv4 I__16600 (
            .O(N__74421),
            .I(wr_addr_r_1));
    Odrv4 I__16599 (
            .O(N__74418),
            .I(wr_addr_r_1));
    Odrv4 I__16598 (
            .O(N__74413),
            .I(wr_addr_r_1));
    LocalMux I__16597 (
            .O(N__74408),
            .I(wr_addr_r_1));
    LocalMux I__16596 (
            .O(N__74401),
            .I(wr_addr_r_1));
    LocalMux I__16595 (
            .O(N__74396),
            .I(wr_addr_r_1));
    CascadeMux I__16594 (
            .O(N__74383),
            .I(n32_cascade_));
    InMux I__16593 (
            .O(N__74380),
            .I(N__74373));
    InMux I__16592 (
            .O(N__74379),
            .I(N__74368));
    InMux I__16591 (
            .O(N__74378),
            .I(N__74368));
    InMux I__16590 (
            .O(N__74377),
            .I(N__74363));
    InMux I__16589 (
            .O(N__74376),
            .I(N__74363));
    LocalMux I__16588 (
            .O(N__74373),
            .I(fifo_write_cmd));
    LocalMux I__16587 (
            .O(N__74368),
            .I(fifo_write_cmd));
    LocalMux I__16586 (
            .O(N__74363),
            .I(fifo_write_cmd));
    InMux I__16585 (
            .O(N__74356),
            .I(N__74353));
    LocalMux I__16584 (
            .O(N__74353),
            .I(\tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r ));
    InMux I__16583 (
            .O(N__74350),
            .I(N__74343));
    InMux I__16582 (
            .O(N__74349),
            .I(N__74343));
    InMux I__16581 (
            .O(N__74348),
            .I(N__74340));
    LocalMux I__16580 (
            .O(N__74343),
            .I(n2207));
    LocalMux I__16579 (
            .O(N__74340),
            .I(n2207));
    InMux I__16578 (
            .O(N__74335),
            .I(N__74332));
    LocalMux I__16577 (
            .O(N__74332),
            .I(empty_o_N_1116));
    InMux I__16576 (
            .O(N__74329),
            .I(N__74322));
    InMux I__16575 (
            .O(N__74328),
            .I(N__74316));
    InMux I__16574 (
            .O(N__74327),
            .I(N__74316));
    CascadeMux I__16573 (
            .O(N__74326),
            .I(N__74312));
    CascadeMux I__16572 (
            .O(N__74325),
            .I(N__74308));
    LocalMux I__16571 (
            .O(N__74322),
            .I(N__74305));
    InMux I__16570 (
            .O(N__74321),
            .I(N__74302));
    LocalMux I__16569 (
            .O(N__74316),
            .I(N__74299));
    InMux I__16568 (
            .O(N__74315),
            .I(N__74296));
    InMux I__16567 (
            .O(N__74312),
            .I(N__74293));
    InMux I__16566 (
            .O(N__74311),
            .I(N__74288));
    InMux I__16565 (
            .O(N__74308),
            .I(N__74288));
    Odrv12 I__16564 (
            .O(N__74305),
            .I(fifo_read_cmd));
    LocalMux I__16563 (
            .O(N__74302),
            .I(fifo_read_cmd));
    Odrv4 I__16562 (
            .O(N__74299),
            .I(fifo_read_cmd));
    LocalMux I__16561 (
            .O(N__74296),
            .I(fifo_read_cmd));
    LocalMux I__16560 (
            .O(N__74293),
            .I(fifo_read_cmd));
    LocalMux I__16559 (
            .O(N__74288),
            .I(fifo_read_cmd));
    InMux I__16558 (
            .O(N__74275),
            .I(N__74269));
    InMux I__16557 (
            .O(N__74274),
            .I(N__74269));
    LocalMux I__16556 (
            .O(N__74269),
            .I(N__74265));
    CascadeMux I__16555 (
            .O(N__74268),
            .I(N__74262));
    Span4Mux_v I__16554 (
            .O(N__74265),
            .I(N__74252));
    InMux I__16553 (
            .O(N__74262),
            .I(N__74249));
    InMux I__16552 (
            .O(N__74261),
            .I(N__74246));
    InMux I__16551 (
            .O(N__74260),
            .I(N__74241));
    InMux I__16550 (
            .O(N__74259),
            .I(N__74241));
    InMux I__16549 (
            .O(N__74258),
            .I(N__74238));
    InMux I__16548 (
            .O(N__74257),
            .I(N__74235));
    InMux I__16547 (
            .O(N__74256),
            .I(N__74232));
    InMux I__16546 (
            .O(N__74255),
            .I(N__74229));
    Odrv4 I__16545 (
            .O(N__74252),
            .I(wr_addr_r_0_adj_1181));
    LocalMux I__16544 (
            .O(N__74249),
            .I(wr_addr_r_0_adj_1181));
    LocalMux I__16543 (
            .O(N__74246),
            .I(wr_addr_r_0_adj_1181));
    LocalMux I__16542 (
            .O(N__74241),
            .I(wr_addr_r_0_adj_1181));
    LocalMux I__16541 (
            .O(N__74238),
            .I(wr_addr_r_0_adj_1181));
    LocalMux I__16540 (
            .O(N__74235),
            .I(wr_addr_r_0_adj_1181));
    LocalMux I__16539 (
            .O(N__74232),
            .I(wr_addr_r_0_adj_1181));
    LocalMux I__16538 (
            .O(N__74229),
            .I(wr_addr_r_0_adj_1181));
    CascadeMux I__16537 (
            .O(N__74212),
            .I(N__74209));
    InMux I__16536 (
            .O(N__74209),
            .I(N__74206));
    LocalMux I__16535 (
            .O(N__74206),
            .I(N__74202));
    CascadeMux I__16534 (
            .O(N__74205),
            .I(N__74199));
    Span4Mux_v I__16533 (
            .O(N__74202),
            .I(N__74193));
    InMux I__16532 (
            .O(N__74199),
            .I(N__74186));
    InMux I__16531 (
            .O(N__74198),
            .I(N__74186));
    InMux I__16530 (
            .O(N__74197),
            .I(N__74186));
    InMux I__16529 (
            .O(N__74196),
            .I(N__74183));
    Odrv4 I__16528 (
            .O(N__74193),
            .I(rx_buf_byte_2));
    LocalMux I__16527 (
            .O(N__74186),
            .I(rx_buf_byte_2));
    LocalMux I__16526 (
            .O(N__74183),
            .I(rx_buf_byte_2));
    InMux I__16525 (
            .O(N__74176),
            .I(N__74173));
    LocalMux I__16524 (
            .O(N__74173),
            .I(N__74169));
    InMux I__16523 (
            .O(N__74172),
            .I(N__74166));
    Odrv4 I__16522 (
            .O(N__74169),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2 ));
    LocalMux I__16521 (
            .O(N__74166),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2 ));
    InMux I__16520 (
            .O(N__74161),
            .I(N__74158));
    LocalMux I__16519 (
            .O(N__74158),
            .I(N__74155));
    Span4Mux_h I__16518 (
            .O(N__74155),
            .I(N__74152));
    Span4Mux_v I__16517 (
            .O(N__74152),
            .I(N__74148));
    InMux I__16516 (
            .O(N__74151),
            .I(N__74145));
    Odrv4 I__16515 (
            .O(N__74148),
            .I(\spi0.multi_byte_counter_7 ));
    LocalMux I__16514 (
            .O(N__74145),
            .I(\spi0.multi_byte_counter_7 ));
    InMux I__16513 (
            .O(N__74140),
            .I(N__74137));
    LocalMux I__16512 (
            .O(N__74137),
            .I(N__74134));
    Span4Mux_h I__16511 (
            .O(N__74134),
            .I(N__74130));
    CascadeMux I__16510 (
            .O(N__74133),
            .I(N__74127));
    Span4Mux_v I__16509 (
            .O(N__74130),
            .I(N__74124));
    InMux I__16508 (
            .O(N__74127),
            .I(N__74121));
    Odrv4 I__16507 (
            .O(N__74124),
            .I(\spi0.multi_byte_counter_5 ));
    LocalMux I__16506 (
            .O(N__74121),
            .I(\spi0.multi_byte_counter_5 ));
    CascadeMux I__16505 (
            .O(N__74116),
            .I(N__74113));
    InMux I__16504 (
            .O(N__74113),
            .I(N__74110));
    LocalMux I__16503 (
            .O(N__74110),
            .I(N__74106));
    CascadeMux I__16502 (
            .O(N__74109),
            .I(N__74103));
    Span12Mux_v I__16501 (
            .O(N__74106),
            .I(N__74100));
    InMux I__16500 (
            .O(N__74103),
            .I(N__74097));
    Odrv12 I__16499 (
            .O(N__74100),
            .I(\spi0.multi_byte_counter_3 ));
    LocalMux I__16498 (
            .O(N__74097),
            .I(\spi0.multi_byte_counter_3 ));
    InMux I__16497 (
            .O(N__74092),
            .I(N__74089));
    LocalMux I__16496 (
            .O(N__74089),
            .I(N__74086));
    Span4Mux_h I__16495 (
            .O(N__74086),
            .I(N__74082));
    CascadeMux I__16494 (
            .O(N__74085),
            .I(N__74079));
    Span4Mux_v I__16493 (
            .O(N__74082),
            .I(N__74076));
    InMux I__16492 (
            .O(N__74079),
            .I(N__74073));
    Odrv4 I__16491 (
            .O(N__74076),
            .I(\spi0.multi_byte_counter_1 ));
    LocalMux I__16490 (
            .O(N__74073),
            .I(\spi0.multi_byte_counter_1 ));
    InMux I__16489 (
            .O(N__74068),
            .I(N__74065));
    LocalMux I__16488 (
            .O(N__74065),
            .I(N__74062));
    Span4Mux_v I__16487 (
            .O(N__74062),
            .I(N__74059));
    Span4Mux_h I__16486 (
            .O(N__74059),
            .I(N__74056));
    Odrv4 I__16485 (
            .O(N__74056),
            .I(\spi0.n14_adj_1140 ));
    InMux I__16484 (
            .O(N__74053),
            .I(N__74050));
    LocalMux I__16483 (
            .O(N__74050),
            .I(N__74047));
    Odrv4 I__16482 (
            .O(N__74047),
            .I(\timing_controller_inst.n62 ));
    CascadeMux I__16481 (
            .O(N__74044),
            .I(N__74041));
    InMux I__16480 (
            .O(N__74041),
            .I(N__74038));
    LocalMux I__16479 (
            .O(N__74038),
            .I(\timing_controller_inst.n49 ));
    CascadeMux I__16478 (
            .O(N__74035),
            .I(N__74032));
    InMux I__16477 (
            .O(N__74032),
            .I(N__74028));
    CascadeMux I__16476 (
            .O(N__74031),
            .I(N__74025));
    LocalMux I__16475 (
            .O(N__74028),
            .I(N__74021));
    InMux I__16474 (
            .O(N__74025),
            .I(N__74016));
    InMux I__16473 (
            .O(N__74024),
            .I(N__74016));
    Span4Mux_v I__16472 (
            .O(N__74021),
            .I(N__74011));
    LocalMux I__16471 (
            .O(N__74016),
            .I(N__74008));
    InMux I__16470 (
            .O(N__74015),
            .I(N__74005));
    InMux I__16469 (
            .O(N__74014),
            .I(N__74002));
    Odrv4 I__16468 (
            .O(N__74011),
            .I(rx_buf_byte_3));
    Odrv4 I__16467 (
            .O(N__74008),
            .I(rx_buf_byte_3));
    LocalMux I__16466 (
            .O(N__74005),
            .I(rx_buf_byte_3));
    LocalMux I__16465 (
            .O(N__74002),
            .I(rx_buf_byte_3));
    CascadeMux I__16464 (
            .O(N__73993),
            .I(N__73988));
    CascadeMux I__16463 (
            .O(N__73992),
            .I(N__73983));
    InMux I__16462 (
            .O(N__73991),
            .I(N__73977));
    InMux I__16461 (
            .O(N__73988),
            .I(N__73977));
    CascadeMux I__16460 (
            .O(N__73987),
            .I(N__73972));
    InMux I__16459 (
            .O(N__73986),
            .I(N__73965));
    InMux I__16458 (
            .O(N__73983),
            .I(N__73965));
    CascadeMux I__16457 (
            .O(N__73982),
            .I(N__73962));
    LocalMux I__16456 (
            .O(N__73977),
            .I(N__73959));
    InMux I__16455 (
            .O(N__73976),
            .I(N__73954));
    InMux I__16454 (
            .O(N__73975),
            .I(N__73954));
    InMux I__16453 (
            .O(N__73972),
            .I(N__73951));
    CascadeMux I__16452 (
            .O(N__73971),
            .I(N__73947));
    CascadeMux I__16451 (
            .O(N__73970),
            .I(N__73940));
    LocalMux I__16450 (
            .O(N__73965),
            .I(N__73937));
    InMux I__16449 (
            .O(N__73962),
            .I(N__73934));
    Span4Mux_h I__16448 (
            .O(N__73959),
            .I(N__73927));
    LocalMux I__16447 (
            .O(N__73954),
            .I(N__73927));
    LocalMux I__16446 (
            .O(N__73951),
            .I(N__73927));
    InMux I__16445 (
            .O(N__73950),
            .I(N__73924));
    InMux I__16444 (
            .O(N__73947),
            .I(N__73911));
    InMux I__16443 (
            .O(N__73946),
            .I(N__73911));
    InMux I__16442 (
            .O(N__73945),
            .I(N__73911));
    InMux I__16441 (
            .O(N__73944),
            .I(N__73911));
    InMux I__16440 (
            .O(N__73943),
            .I(N__73911));
    InMux I__16439 (
            .O(N__73940),
            .I(N__73911));
    Odrv4 I__16438 (
            .O(N__73937),
            .I(\tx_fifo.lscc_fifo_inst.n4 ));
    LocalMux I__16437 (
            .O(N__73934),
            .I(\tx_fifo.lscc_fifo_inst.n4 ));
    Odrv4 I__16436 (
            .O(N__73927),
            .I(\tx_fifo.lscc_fifo_inst.n4 ));
    LocalMux I__16435 (
            .O(N__73924),
            .I(\tx_fifo.lscc_fifo_inst.n4 ));
    LocalMux I__16434 (
            .O(N__73911),
            .I(\tx_fifo.lscc_fifo_inst.n4 ));
    CascadeMux I__16433 (
            .O(N__73900),
            .I(N__73897));
    InMux I__16432 (
            .O(N__73897),
            .I(N__73892));
    InMux I__16431 (
            .O(N__73896),
            .I(N__73889));
    CascadeMux I__16430 (
            .O(N__73895),
            .I(N__73886));
    LocalMux I__16429 (
            .O(N__73892),
            .I(N__73882));
    LocalMux I__16428 (
            .O(N__73889),
            .I(N__73879));
    InMux I__16427 (
            .O(N__73886),
            .I(N__73874));
    InMux I__16426 (
            .O(N__73885),
            .I(N__73874));
    Span4Mux_v I__16425 (
            .O(N__73882),
            .I(N__73870));
    Span4Mux_h I__16424 (
            .O(N__73879),
            .I(N__73865));
    LocalMux I__16423 (
            .O(N__73874),
            .I(N__73865));
    InMux I__16422 (
            .O(N__73873),
            .I(N__73862));
    Odrv4 I__16421 (
            .O(N__73870),
            .I(rx_buf_byte_1));
    Odrv4 I__16420 (
            .O(N__73865),
            .I(rx_buf_byte_1));
    LocalMux I__16419 (
            .O(N__73862),
            .I(rx_buf_byte_1));
    InMux I__16418 (
            .O(N__73855),
            .I(N__73851));
    InMux I__16417 (
            .O(N__73854),
            .I(N__73848));
    LocalMux I__16416 (
            .O(N__73851),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_3 ));
    LocalMux I__16415 (
            .O(N__73848),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_3 ));
    CascadeMux I__16414 (
            .O(N__73843),
            .I(N__73840));
    InMux I__16413 (
            .O(N__73840),
            .I(N__73836));
    InMux I__16412 (
            .O(N__73839),
            .I(N__73833));
    LocalMux I__16411 (
            .O(N__73836),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3 ));
    LocalMux I__16410 (
            .O(N__73833),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3 ));
    InMux I__16409 (
            .O(N__73828),
            .I(N__73825));
    LocalMux I__16408 (
            .O(N__73825),
            .I(mem_LUT_data_raw_r_4));
    InMux I__16407 (
            .O(N__73822),
            .I(N__73816));
    InMux I__16406 (
            .O(N__73821),
            .I(N__73816));
    LocalMux I__16405 (
            .O(N__73816),
            .I(fifo_temp_output_4));
    InMux I__16404 (
            .O(N__73813),
            .I(N__73810));
    LocalMux I__16403 (
            .O(N__73810),
            .I(mem_LUT_data_raw_r_5));
    InMux I__16402 (
            .O(N__73807),
            .I(N__73801));
    InMux I__16401 (
            .O(N__73806),
            .I(N__73801));
    LocalMux I__16400 (
            .O(N__73801),
            .I(fifo_temp_output_5));
    InMux I__16399 (
            .O(N__73798),
            .I(N__73795));
    LocalMux I__16398 (
            .O(N__73795),
            .I(N__73792));
    Span4Mux_v I__16397 (
            .O(N__73792),
            .I(N__73789));
    Odrv4 I__16396 (
            .O(N__73789),
            .I(mem_LUT_data_raw_r_6));
    InMux I__16395 (
            .O(N__73786),
            .I(N__73780));
    InMux I__16394 (
            .O(N__73785),
            .I(N__73780));
    LocalMux I__16393 (
            .O(N__73780),
            .I(fifo_temp_output_6));
    InMux I__16392 (
            .O(N__73777),
            .I(N__73774));
    LocalMux I__16391 (
            .O(N__73774),
            .I(N__73771));
    Odrv12 I__16390 (
            .O(N__73771),
            .I(mem_LUT_data_raw_r_7));
    InMux I__16389 (
            .O(N__73768),
            .I(N__73764));
    InMux I__16388 (
            .O(N__73767),
            .I(N__73761));
    LocalMux I__16387 (
            .O(N__73764),
            .I(fifo_temp_output_7));
    LocalMux I__16386 (
            .O(N__73761),
            .I(fifo_temp_output_7));
    SRMux I__16385 (
            .O(N__73756),
            .I(N__73751));
    SRMux I__16384 (
            .O(N__73755),
            .I(N__73748));
    SRMux I__16383 (
            .O(N__73754),
            .I(N__73743));
    LocalMux I__16382 (
            .O(N__73751),
            .I(N__73740));
    LocalMux I__16381 (
            .O(N__73748),
            .I(N__73737));
    SRMux I__16380 (
            .O(N__73747),
            .I(N__73734));
    SRMux I__16379 (
            .O(N__73746),
            .I(N__73731));
    LocalMux I__16378 (
            .O(N__73743),
            .I(N__73728));
    Span4Mux_h I__16377 (
            .O(N__73740),
            .I(N__73719));
    Span4Mux_v I__16376 (
            .O(N__73737),
            .I(N__73719));
    LocalMux I__16375 (
            .O(N__73734),
            .I(N__73719));
    LocalMux I__16374 (
            .O(N__73731),
            .I(N__73719));
    Span4Mux_h I__16373 (
            .O(N__73728),
            .I(N__73713));
    Span4Mux_h I__16372 (
            .O(N__73719),
            .I(N__73713));
    InMux I__16371 (
            .O(N__73718),
            .I(N__73705));
    Span4Mux_h I__16370 (
            .O(N__73713),
            .I(N__73701));
    SRMux I__16369 (
            .O(N__73712),
            .I(N__73698));
    SRMux I__16368 (
            .O(N__73711),
            .I(N__73695));
    SRMux I__16367 (
            .O(N__73710),
            .I(N__73692));
    SRMux I__16366 (
            .O(N__73709),
            .I(N__73686));
    InMux I__16365 (
            .O(N__73708),
            .I(N__73682));
    LocalMux I__16364 (
            .O(N__73705),
            .I(N__73678));
    SRMux I__16363 (
            .O(N__73704),
            .I(N__73675));
    Span4Mux_h I__16362 (
            .O(N__73701),
            .I(N__73670));
    LocalMux I__16361 (
            .O(N__73698),
            .I(N__73670));
    LocalMux I__16360 (
            .O(N__73695),
            .I(N__73665));
    LocalMux I__16359 (
            .O(N__73692),
            .I(N__73665));
    InMux I__16358 (
            .O(N__73691),
            .I(N__73662));
    InMux I__16357 (
            .O(N__73690),
            .I(N__73657));
    SRMux I__16356 (
            .O(N__73689),
            .I(N__73657));
    LocalMux I__16355 (
            .O(N__73686),
            .I(N__73653));
    SRMux I__16354 (
            .O(N__73685),
            .I(N__73650));
    LocalMux I__16353 (
            .O(N__73682),
            .I(N__73647));
    InMux I__16352 (
            .O(N__73681),
            .I(N__73644));
    Span4Mux_v I__16351 (
            .O(N__73678),
            .I(N__73639));
    LocalMux I__16350 (
            .O(N__73675),
            .I(N__73639));
    Span4Mux_h I__16349 (
            .O(N__73670),
            .I(N__73636));
    Span4Mux_h I__16348 (
            .O(N__73665),
            .I(N__73633));
    LocalMux I__16347 (
            .O(N__73662),
            .I(N__73630));
    LocalMux I__16346 (
            .O(N__73657),
            .I(N__73627));
    SRMux I__16345 (
            .O(N__73656),
            .I(N__73624));
    Span4Mux_h I__16344 (
            .O(N__73653),
            .I(N__73621));
    LocalMux I__16343 (
            .O(N__73650),
            .I(N__73618));
    Span12Mux_s10_h I__16342 (
            .O(N__73647),
            .I(N__73613));
    LocalMux I__16341 (
            .O(N__73644),
            .I(N__73613));
    Span4Mux_v I__16340 (
            .O(N__73639),
            .I(N__73610));
    Span4Mux_v I__16339 (
            .O(N__73636),
            .I(N__73605));
    Span4Mux_v I__16338 (
            .O(N__73633),
            .I(N__73605));
    Span4Mux_v I__16337 (
            .O(N__73630),
            .I(N__73600));
    Span4Mux_v I__16336 (
            .O(N__73627),
            .I(N__73600));
    LocalMux I__16335 (
            .O(N__73624),
            .I(N__73597));
    Span4Mux_h I__16334 (
            .O(N__73621),
            .I(N__73592));
    Span4Mux_v I__16333 (
            .O(N__73618),
            .I(N__73592));
    Span12Mux_h I__16332 (
            .O(N__73613),
            .I(N__73589));
    Span4Mux_h I__16331 (
            .O(N__73610),
            .I(N__73586));
    Span4Mux_v I__16330 (
            .O(N__73605),
            .I(N__73581));
    Span4Mux_h I__16329 (
            .O(N__73600),
            .I(N__73581));
    Span4Mux_h I__16328 (
            .O(N__73597),
            .I(N__73576));
    Span4Mux_v I__16327 (
            .O(N__73592),
            .I(N__73576));
    Odrv12 I__16326 (
            .O(N__73589),
            .I(\usb3_if_inst.reset_per_frame_latched ));
    Odrv4 I__16325 (
            .O(N__73586),
            .I(\usb3_if_inst.reset_per_frame_latched ));
    Odrv4 I__16324 (
            .O(N__73581),
            .I(\usb3_if_inst.reset_per_frame_latched ));
    Odrv4 I__16323 (
            .O(N__73576),
            .I(\usb3_if_inst.reset_per_frame_latched ));
    InMux I__16322 (
            .O(N__73567),
            .I(N__73564));
    LocalMux I__16321 (
            .O(N__73564),
            .I(reset_per_frame));
    SRMux I__16320 (
            .O(N__73561),
            .I(N__73553));
    InMux I__16319 (
            .O(N__73560),
            .I(N__73548));
    SRMux I__16318 (
            .O(N__73559),
            .I(N__73548));
    InMux I__16317 (
            .O(N__73558),
            .I(N__73545));
    SRMux I__16316 (
            .O(N__73557),
            .I(N__73542));
    SRMux I__16315 (
            .O(N__73556),
            .I(N__73539));
    LocalMux I__16314 (
            .O(N__73553),
            .I(N__73533));
    LocalMux I__16313 (
            .O(N__73548),
            .I(N__73530));
    LocalMux I__16312 (
            .O(N__73545),
            .I(N__73527));
    LocalMux I__16311 (
            .O(N__73542),
            .I(N__73524));
    LocalMux I__16310 (
            .O(N__73539),
            .I(N__73521));
    InMux I__16309 (
            .O(N__73538),
            .I(N__73518));
    InMux I__16308 (
            .O(N__73537),
            .I(N__73513));
    SRMux I__16307 (
            .O(N__73536),
            .I(N__73513));
    Span4Mux_v I__16306 (
            .O(N__73533),
            .I(N__73510));
    Span4Mux_h I__16305 (
            .O(N__73530),
            .I(N__73507));
    Span4Mux_h I__16304 (
            .O(N__73527),
            .I(N__73502));
    Span4Mux_h I__16303 (
            .O(N__73524),
            .I(N__73502));
    Span4Mux_h I__16302 (
            .O(N__73521),
            .I(N__73499));
    LocalMux I__16301 (
            .O(N__73518),
            .I(N__73494));
    LocalMux I__16300 (
            .O(N__73513),
            .I(N__73494));
    Odrv4 I__16299 (
            .O(N__73510),
            .I(buffer_switch_done));
    Odrv4 I__16298 (
            .O(N__73507),
            .I(buffer_switch_done));
    Odrv4 I__16297 (
            .O(N__73502),
            .I(buffer_switch_done));
    Odrv4 I__16296 (
            .O(N__73499),
            .I(buffer_switch_done));
    Odrv12 I__16295 (
            .O(N__73494),
            .I(buffer_switch_done));
    SRMux I__16294 (
            .O(N__73483),
            .I(N__73478));
    InMux I__16293 (
            .O(N__73482),
            .I(N__73470));
    CascadeMux I__16292 (
            .O(N__73481),
            .I(N__73453));
    LocalMux I__16291 (
            .O(N__73478),
            .I(N__73450));
    SRMux I__16290 (
            .O(N__73477),
            .I(N__73447));
    CascadeMux I__16289 (
            .O(N__73476),
            .I(N__73444));
    CascadeMux I__16288 (
            .O(N__73475),
            .I(N__73441));
    CascadeMux I__16287 (
            .O(N__73474),
            .I(N__73437));
    CascadeMux I__16286 (
            .O(N__73473),
            .I(N__73433));
    LocalMux I__16285 (
            .O(N__73470),
            .I(N__73430));
    InMux I__16284 (
            .O(N__73469),
            .I(N__73402));
    InMux I__16283 (
            .O(N__73468),
            .I(N__73402));
    InMux I__16282 (
            .O(N__73467),
            .I(N__73402));
    InMux I__16281 (
            .O(N__73466),
            .I(N__73402));
    InMux I__16280 (
            .O(N__73465),
            .I(N__73402));
    SRMux I__16279 (
            .O(N__73464),
            .I(N__73399));
    InMux I__16278 (
            .O(N__73463),
            .I(N__73396));
    InMux I__16277 (
            .O(N__73462),
            .I(N__73385));
    InMux I__16276 (
            .O(N__73461),
            .I(N__73385));
    InMux I__16275 (
            .O(N__73460),
            .I(N__73385));
    InMux I__16274 (
            .O(N__73459),
            .I(N__73385));
    InMux I__16273 (
            .O(N__73458),
            .I(N__73385));
    SRMux I__16272 (
            .O(N__73457),
            .I(N__73382));
    InMux I__16271 (
            .O(N__73456),
            .I(N__73374));
    InMux I__16270 (
            .O(N__73453),
            .I(N__73374));
    Span4Mux_h I__16269 (
            .O(N__73450),
            .I(N__73369));
    LocalMux I__16268 (
            .O(N__73447),
            .I(N__73366));
    InMux I__16267 (
            .O(N__73444),
            .I(N__73363));
    InMux I__16266 (
            .O(N__73441),
            .I(N__73352));
    InMux I__16265 (
            .O(N__73440),
            .I(N__73352));
    InMux I__16264 (
            .O(N__73437),
            .I(N__73352));
    InMux I__16263 (
            .O(N__73436),
            .I(N__73352));
    InMux I__16262 (
            .O(N__73433),
            .I(N__73352));
    Span4Mux_v I__16261 (
            .O(N__73430),
            .I(N__73349));
    InMux I__16260 (
            .O(N__73429),
            .I(N__73344));
    InMux I__16259 (
            .O(N__73428),
            .I(N__73344));
    InMux I__16258 (
            .O(N__73427),
            .I(N__73339));
    InMux I__16257 (
            .O(N__73426),
            .I(N__73339));
    InMux I__16256 (
            .O(N__73425),
            .I(N__73322));
    InMux I__16255 (
            .O(N__73424),
            .I(N__73322));
    InMux I__16254 (
            .O(N__73423),
            .I(N__73322));
    InMux I__16253 (
            .O(N__73422),
            .I(N__73322));
    InMux I__16252 (
            .O(N__73421),
            .I(N__73322));
    InMux I__16251 (
            .O(N__73420),
            .I(N__73322));
    InMux I__16250 (
            .O(N__73419),
            .I(N__73322));
    InMux I__16249 (
            .O(N__73418),
            .I(N__73322));
    InMux I__16248 (
            .O(N__73417),
            .I(N__73313));
    InMux I__16247 (
            .O(N__73416),
            .I(N__73313));
    InMux I__16246 (
            .O(N__73415),
            .I(N__73313));
    InMux I__16245 (
            .O(N__73414),
            .I(N__73313));
    SRMux I__16244 (
            .O(N__73413),
            .I(N__73310));
    LocalMux I__16243 (
            .O(N__73402),
            .I(N__73307));
    LocalMux I__16242 (
            .O(N__73399),
            .I(N__73304));
    LocalMux I__16241 (
            .O(N__73396),
            .I(N__73286));
    LocalMux I__16240 (
            .O(N__73385),
            .I(N__73286));
    LocalMux I__16239 (
            .O(N__73382),
            .I(N__73286));
    InMux I__16238 (
            .O(N__73381),
            .I(N__73279));
    InMux I__16237 (
            .O(N__73380),
            .I(N__73279));
    InMux I__16236 (
            .O(N__73379),
            .I(N__73279));
    LocalMux I__16235 (
            .O(N__73374),
            .I(N__73276));
    SRMux I__16234 (
            .O(N__73373),
            .I(N__73273));
    InMux I__16233 (
            .O(N__73372),
            .I(N__73270));
    Span4Mux_h I__16232 (
            .O(N__73369),
            .I(N__73267));
    Span4Mux_h I__16231 (
            .O(N__73366),
            .I(N__73264));
    LocalMux I__16230 (
            .O(N__73363),
            .I(N__73261));
    LocalMux I__16229 (
            .O(N__73352),
            .I(N__73258));
    Span4Mux_h I__16228 (
            .O(N__73349),
            .I(N__73245));
    LocalMux I__16227 (
            .O(N__73344),
            .I(N__73245));
    LocalMux I__16226 (
            .O(N__73339),
            .I(N__73245));
    LocalMux I__16225 (
            .O(N__73322),
            .I(N__73245));
    LocalMux I__16224 (
            .O(N__73313),
            .I(N__73245));
    LocalMux I__16223 (
            .O(N__73310),
            .I(N__73245));
    Span4Mux_v I__16222 (
            .O(N__73307),
            .I(N__73240));
    Span4Mux_v I__16221 (
            .O(N__73304),
            .I(N__73240));
    InMux I__16220 (
            .O(N__73303),
            .I(N__73237));
    InMux I__16219 (
            .O(N__73302),
            .I(N__73226));
    InMux I__16218 (
            .O(N__73301),
            .I(N__73226));
    InMux I__16217 (
            .O(N__73300),
            .I(N__73226));
    InMux I__16216 (
            .O(N__73299),
            .I(N__73226));
    InMux I__16215 (
            .O(N__73298),
            .I(N__73226));
    InMux I__16214 (
            .O(N__73297),
            .I(N__73223));
    InMux I__16213 (
            .O(N__73296),
            .I(N__73220));
    InMux I__16212 (
            .O(N__73295),
            .I(N__73213));
    InMux I__16211 (
            .O(N__73294),
            .I(N__73213));
    InMux I__16210 (
            .O(N__73293),
            .I(N__73213));
    Span4Mux_v I__16209 (
            .O(N__73286),
            .I(N__73204));
    LocalMux I__16208 (
            .O(N__73279),
            .I(N__73204));
    Span4Mux_v I__16207 (
            .O(N__73276),
            .I(N__73204));
    LocalMux I__16206 (
            .O(N__73273),
            .I(N__73204));
    LocalMux I__16205 (
            .O(N__73270),
            .I(N__73193));
    Span4Mux_h I__16204 (
            .O(N__73267),
            .I(N__73190));
    Span4Mux_h I__16203 (
            .O(N__73264),
            .I(N__73187));
    Span4Mux_v I__16202 (
            .O(N__73261),
            .I(N__73184));
    Span4Mux_v I__16201 (
            .O(N__73258),
            .I(N__73179));
    Span4Mux_v I__16200 (
            .O(N__73245),
            .I(N__73179));
    Span4Mux_h I__16199 (
            .O(N__73240),
            .I(N__73172));
    LocalMux I__16198 (
            .O(N__73237),
            .I(N__73172));
    LocalMux I__16197 (
            .O(N__73226),
            .I(N__73172));
    LocalMux I__16196 (
            .O(N__73223),
            .I(N__73165));
    LocalMux I__16195 (
            .O(N__73220),
            .I(N__73165));
    LocalMux I__16194 (
            .O(N__73213),
            .I(N__73165));
    Span4Mux_v I__16193 (
            .O(N__73204),
            .I(N__73162));
    InMux I__16192 (
            .O(N__73203),
            .I(N__73145));
    InMux I__16191 (
            .O(N__73202),
            .I(N__73145));
    InMux I__16190 (
            .O(N__73201),
            .I(N__73145));
    InMux I__16189 (
            .O(N__73200),
            .I(N__73145));
    InMux I__16188 (
            .O(N__73199),
            .I(N__73145));
    InMux I__16187 (
            .O(N__73198),
            .I(N__73145));
    InMux I__16186 (
            .O(N__73197),
            .I(N__73145));
    InMux I__16185 (
            .O(N__73196),
            .I(N__73145));
    Span12Mux_h I__16184 (
            .O(N__73193),
            .I(N__73142));
    Span4Mux_v I__16183 (
            .O(N__73190),
            .I(N__73139));
    Span4Mux_h I__16182 (
            .O(N__73187),
            .I(N__73136));
    Span4Mux_v I__16181 (
            .O(N__73184),
            .I(N__73131));
    Span4Mux_h I__16180 (
            .O(N__73179),
            .I(N__73131));
    Span4Mux_v I__16179 (
            .O(N__73172),
            .I(N__73128));
    Span12Mux_v I__16178 (
            .O(N__73165),
            .I(N__73121));
    Sp12to4 I__16177 (
            .O(N__73162),
            .I(N__73121));
    LocalMux I__16176 (
            .O(N__73145),
            .I(N__73121));
    Odrv12 I__16175 (
            .O(N__73142),
            .I(reset_all));
    Odrv4 I__16174 (
            .O(N__73139),
            .I(reset_all));
    Odrv4 I__16173 (
            .O(N__73136),
            .I(reset_all));
    Odrv4 I__16172 (
            .O(N__73131),
            .I(reset_all));
    Odrv4 I__16171 (
            .O(N__73128),
            .I(reset_all));
    Odrv12 I__16170 (
            .O(N__73121),
            .I(reset_all));
    InMux I__16169 (
            .O(N__73108),
            .I(N__73105));
    LocalMux I__16168 (
            .O(N__73105),
            .I(N__73102));
    Span4Mux_v I__16167 (
            .O(N__73102),
            .I(N__73099));
    Span4Mux_h I__16166 (
            .O(N__73099),
            .I(N__73096));
    Odrv4 I__16165 (
            .O(N__73096),
            .I(REG_out_raw_4));
    CascadeMux I__16164 (
            .O(N__73093),
            .I(\timing_controller_inst.n11375_cascade_ ));
    CEMux I__16163 (
            .O(N__73090),
            .I(N__73087));
    LocalMux I__16162 (
            .O(N__73087),
            .I(N__73084));
    Odrv4 I__16161 (
            .O(N__73084),
            .I(\timing_controller_inst.n4200 ));
    InMux I__16160 (
            .O(N__73081),
            .I(N__73078));
    LocalMux I__16159 (
            .O(N__73078),
            .I(n11376));
    CascadeMux I__16158 (
            .O(N__73075),
            .I(n11376_cascade_));
    IoInMux I__16157 (
            .O(N__73072),
            .I(N__73069));
    LocalMux I__16156 (
            .O(N__73069),
            .I(N__73066));
    IoSpan4Mux I__16155 (
            .O(N__73066),
            .I(N__73063));
    Span4Mux_s2_h I__16154 (
            .O(N__73063),
            .I(N__73060));
    Span4Mux_h I__16153 (
            .O(N__73060),
            .I(N__73057));
    Odrv4 I__16152 (
            .O(N__73057),
            .I(\timing_controller_inst.invert_N_309 ));
    InMux I__16151 (
            .O(N__73054),
            .I(N__73047));
    InMux I__16150 (
            .O(N__73053),
            .I(N__73043));
    InMux I__16149 (
            .O(N__73052),
            .I(N__73040));
    InMux I__16148 (
            .O(N__73051),
            .I(N__73037));
    InMux I__16147 (
            .O(N__73050),
            .I(N__73034));
    LocalMux I__16146 (
            .O(N__73047),
            .I(N__73029));
    InMux I__16145 (
            .O(N__73046),
            .I(N__73026));
    LocalMux I__16144 (
            .O(N__73043),
            .I(N__73022));
    LocalMux I__16143 (
            .O(N__73040),
            .I(N__73019));
    LocalMux I__16142 (
            .O(N__73037),
            .I(N__73014));
    LocalMux I__16141 (
            .O(N__73034),
            .I(N__73010));
    InMux I__16140 (
            .O(N__73033),
            .I(N__73007));
    InMux I__16139 (
            .O(N__73032),
            .I(N__73004));
    Span4Mux_h I__16138 (
            .O(N__73029),
            .I(N__73001));
    LocalMux I__16137 (
            .O(N__73026),
            .I(N__72998));
    InMux I__16136 (
            .O(N__73025),
            .I(N__72995));
    Span4Mux_h I__16135 (
            .O(N__73022),
            .I(N__72988));
    Span4Mux_h I__16134 (
            .O(N__73019),
            .I(N__72988));
    InMux I__16133 (
            .O(N__73018),
            .I(N__72985));
    InMux I__16132 (
            .O(N__73017),
            .I(N__72982));
    Span4Mux_v I__16131 (
            .O(N__73014),
            .I(N__72978));
    InMux I__16130 (
            .O(N__73013),
            .I(N__72975));
    Span4Mux_h I__16129 (
            .O(N__73010),
            .I(N__72970));
    LocalMux I__16128 (
            .O(N__73007),
            .I(N__72970));
    LocalMux I__16127 (
            .O(N__73004),
            .I(N__72967));
    Span4Mux_h I__16126 (
            .O(N__73001),
            .I(N__72960));
    Span4Mux_v I__16125 (
            .O(N__72998),
            .I(N__72960));
    LocalMux I__16124 (
            .O(N__72995),
            .I(N__72960));
    InMux I__16123 (
            .O(N__72994),
            .I(N__72957));
    InMux I__16122 (
            .O(N__72993),
            .I(N__72954));
    Span4Mux_v I__16121 (
            .O(N__72988),
            .I(N__72951));
    LocalMux I__16120 (
            .O(N__72985),
            .I(N__72948));
    LocalMux I__16119 (
            .O(N__72982),
            .I(N__72945));
    InMux I__16118 (
            .O(N__72981),
            .I(N__72942));
    Sp12to4 I__16117 (
            .O(N__72978),
            .I(N__72936));
    LocalMux I__16116 (
            .O(N__72975),
            .I(N__72936));
    Span4Mux_h I__16115 (
            .O(N__72970),
            .I(N__72931));
    Span4Mux_v I__16114 (
            .O(N__72967),
            .I(N__72931));
    Span4Mux_v I__16113 (
            .O(N__72960),
            .I(N__72928));
    LocalMux I__16112 (
            .O(N__72957),
            .I(N__72923));
    LocalMux I__16111 (
            .O(N__72954),
            .I(N__72923));
    Span4Mux_v I__16110 (
            .O(N__72951),
            .I(N__72914));
    Span4Mux_v I__16109 (
            .O(N__72948),
            .I(N__72914));
    Span4Mux_h I__16108 (
            .O(N__72945),
            .I(N__72914));
    LocalMux I__16107 (
            .O(N__72942),
            .I(N__72914));
    InMux I__16106 (
            .O(N__72941),
            .I(N__72911));
    Odrv12 I__16105 (
            .O(N__72936),
            .I(n15_adj_1184));
    Odrv4 I__16104 (
            .O(N__72931),
            .I(n15_adj_1184));
    Odrv4 I__16103 (
            .O(N__72928),
            .I(n15_adj_1184));
    Odrv12 I__16102 (
            .O(N__72923),
            .I(n15_adj_1184));
    Odrv4 I__16101 (
            .O(N__72914),
            .I(n15_adj_1184));
    LocalMux I__16100 (
            .O(N__72911),
            .I(n15_adj_1184));
    CascadeMux I__16099 (
            .O(N__72898),
            .I(N__72895));
    InMux I__16098 (
            .O(N__72895),
            .I(N__72892));
    LocalMux I__16097 (
            .O(N__72892),
            .I(N__72889));
    Span4Mux_h I__16096 (
            .O(N__72889),
            .I(N__72885));
    InMux I__16095 (
            .O(N__72888),
            .I(N__72882));
    Odrv4 I__16094 (
            .O(N__72885),
            .I(REG_mem_50_8));
    LocalMux I__16093 (
            .O(N__72882),
            .I(REG_mem_50_8));
    InMux I__16092 (
            .O(N__72877),
            .I(N__72874));
    LocalMux I__16091 (
            .O(N__72874),
            .I(N__72871));
    Span4Mux_v I__16090 (
            .O(N__72871),
            .I(N__72868));
    Span4Mux_v I__16089 (
            .O(N__72868),
            .I(N__72865));
    Odrv4 I__16088 (
            .O(N__72865),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13871 ));
    InMux I__16087 (
            .O(N__72862),
            .I(N__72859));
    LocalMux I__16086 (
            .O(N__72859),
            .I(N__72856));
    Span4Mux_v I__16085 (
            .O(N__72856),
            .I(N__72853));
    Odrv4 I__16084 (
            .O(N__72853),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13739 ));
    CascadeMux I__16083 (
            .O(N__72850),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12182_cascade_ ));
    InMux I__16082 (
            .O(N__72847),
            .I(N__72844));
    LocalMux I__16081 (
            .O(N__72844),
            .I(N__72841));
    Odrv12 I__16080 (
            .O(N__72841),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13799 ));
    InMux I__16079 (
            .O(N__72838),
            .I(N__72835));
    LocalMux I__16078 (
            .O(N__72835),
            .I(N__72832));
    Odrv4 I__16077 (
            .O(N__72832),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13787 ));
    InMux I__16076 (
            .O(N__72829),
            .I(N__72826));
    LocalMux I__16075 (
            .O(N__72826),
            .I(N__72823));
    Span4Mux_h I__16074 (
            .O(N__72823),
            .I(N__72820));
    Odrv4 I__16073 (
            .O(N__72820),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13937 ));
    InMux I__16072 (
            .O(N__72817),
            .I(N__72814));
    LocalMux I__16071 (
            .O(N__72814),
            .I(N__72811));
    Span4Mux_v I__16070 (
            .O(N__72811),
            .I(N__72808));
    Span4Mux_v I__16069 (
            .O(N__72808),
            .I(N__72805));
    Odrv4 I__16068 (
            .O(N__72805),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12066 ));
    InMux I__16067 (
            .O(N__72802),
            .I(N__72799));
    LocalMux I__16066 (
            .O(N__72799),
            .I(N__72796));
    Span4Mux_h I__16065 (
            .O(N__72796),
            .I(N__72793));
    Odrv4 I__16064 (
            .O(N__72793),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12093 ));
    InMux I__16063 (
            .O(N__72790),
            .I(N__72787));
    LocalMux I__16062 (
            .O(N__72787),
            .I(N__72784));
    Span4Mux_v I__16061 (
            .O(N__72784),
            .I(N__72781));
    Sp12to4 I__16060 (
            .O(N__72781),
            .I(N__72778));
    Span12Mux_s11_h I__16059 (
            .O(N__72778),
            .I(N__72775));
    Odrv12 I__16058 (
            .O(N__72775),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12006 ));
    CascadeMux I__16057 (
            .O(N__72772),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13610_cascade_ ));
    InMux I__16056 (
            .O(N__72769),
            .I(N__72766));
    LocalMux I__16055 (
            .O(N__72766),
            .I(N__72763));
    Span4Mux_v I__16054 (
            .O(N__72763),
            .I(N__72760));
    Odrv4 I__16053 (
            .O(N__72760),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12240 ));
    CascadeMux I__16052 (
            .O(N__72757),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12246_cascade_ ));
    InMux I__16051 (
            .O(N__72754),
            .I(N__72751));
    LocalMux I__16050 (
            .O(N__72751),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12183 ));
    CascadeMux I__16049 (
            .O(N__72748),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13442_cascade_ ));
    InMux I__16048 (
            .O(N__72745),
            .I(N__72742));
    LocalMux I__16047 (
            .O(N__72742),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12162 ));
    InMux I__16046 (
            .O(N__72739),
            .I(N__72733));
    InMux I__16045 (
            .O(N__72738),
            .I(N__72733));
    LocalMux I__16044 (
            .O(N__72733),
            .I(REG_mem_46_6));
    InMux I__16043 (
            .O(N__72730),
            .I(N__72725));
    InMux I__16042 (
            .O(N__72729),
            .I(N__72721));
    InMux I__16041 (
            .O(N__72728),
            .I(N__72717));
    LocalMux I__16040 (
            .O(N__72725),
            .I(N__72713));
    InMux I__16039 (
            .O(N__72724),
            .I(N__72706));
    LocalMux I__16038 (
            .O(N__72721),
            .I(N__72703));
    InMux I__16037 (
            .O(N__72720),
            .I(N__72697));
    LocalMux I__16036 (
            .O(N__72717),
            .I(N__72694));
    InMux I__16035 (
            .O(N__72716),
            .I(N__72691));
    Span4Mux_h I__16034 (
            .O(N__72713),
            .I(N__72688));
    InMux I__16033 (
            .O(N__72712),
            .I(N__72684));
    InMux I__16032 (
            .O(N__72711),
            .I(N__72681));
    InMux I__16031 (
            .O(N__72710),
            .I(N__72678));
    InMux I__16030 (
            .O(N__72709),
            .I(N__72675));
    LocalMux I__16029 (
            .O(N__72706),
            .I(N__72672));
    Span4Mux_h I__16028 (
            .O(N__72703),
            .I(N__72669));
    InMux I__16027 (
            .O(N__72702),
            .I(N__72664));
    InMux I__16026 (
            .O(N__72701),
            .I(N__72661));
    InMux I__16025 (
            .O(N__72700),
            .I(N__72658));
    LocalMux I__16024 (
            .O(N__72697),
            .I(N__72653));
    Span4Mux_v I__16023 (
            .O(N__72694),
            .I(N__72653));
    LocalMux I__16022 (
            .O(N__72691),
            .I(N__72648));
    Span4Mux_v I__16021 (
            .O(N__72688),
            .I(N__72648));
    InMux I__16020 (
            .O(N__72687),
            .I(N__72645));
    LocalMux I__16019 (
            .O(N__72684),
            .I(N__72640));
    LocalMux I__16018 (
            .O(N__72681),
            .I(N__72640));
    LocalMux I__16017 (
            .O(N__72678),
            .I(N__72637));
    LocalMux I__16016 (
            .O(N__72675),
            .I(N__72632));
    Span4Mux_h I__16015 (
            .O(N__72672),
            .I(N__72632));
    Span4Mux_h I__16014 (
            .O(N__72669),
            .I(N__72629));
    InMux I__16013 (
            .O(N__72668),
            .I(N__72624));
    InMux I__16012 (
            .O(N__72667),
            .I(N__72624));
    LocalMux I__16011 (
            .O(N__72664),
            .I(N__72621));
    LocalMux I__16010 (
            .O(N__72661),
            .I(N__72618));
    LocalMux I__16009 (
            .O(N__72658),
            .I(N__72615));
    Span4Mux_h I__16008 (
            .O(N__72653),
            .I(N__72610));
    Span4Mux_v I__16007 (
            .O(N__72648),
            .I(N__72610));
    LocalMux I__16006 (
            .O(N__72645),
            .I(N__72605));
    Span12Mux_h I__16005 (
            .O(N__72640),
            .I(N__72605));
    Span4Mux_h I__16004 (
            .O(N__72637),
            .I(N__72598));
    Span4Mux_v I__16003 (
            .O(N__72632),
            .I(N__72598));
    Span4Mux_h I__16002 (
            .O(N__72629),
            .I(N__72598));
    LocalMux I__16001 (
            .O(N__72624),
            .I(n61));
    Odrv4 I__16000 (
            .O(N__72621),
            .I(n61));
    Odrv12 I__15999 (
            .O(N__72618),
            .I(n61));
    Odrv12 I__15998 (
            .O(N__72615),
            .I(n61));
    Odrv4 I__15997 (
            .O(N__72610),
            .I(n61));
    Odrv12 I__15996 (
            .O(N__72605),
            .I(n61));
    Odrv4 I__15995 (
            .O(N__72598),
            .I(n61));
    InMux I__15994 (
            .O(N__72583),
            .I(N__72580));
    LocalMux I__15993 (
            .O(N__72580),
            .I(N__72576));
    InMux I__15992 (
            .O(N__72579),
            .I(N__72573));
    Odrv4 I__15991 (
            .O(N__72576),
            .I(REG_mem_4_6));
    LocalMux I__15990 (
            .O(N__72573),
            .I(REG_mem_4_6));
    InMux I__15989 (
            .O(N__72568),
            .I(N__72561));
    InMux I__15988 (
            .O(N__72567),
            .I(N__72555));
    InMux I__15987 (
            .O(N__72566),
            .I(N__72555));
    InMux I__15986 (
            .O(N__72565),
            .I(N__72552));
    InMux I__15985 (
            .O(N__72564),
            .I(N__72547));
    LocalMux I__15984 (
            .O(N__72561),
            .I(N__72544));
    InMux I__15983 (
            .O(N__72560),
            .I(N__72541));
    LocalMux I__15982 (
            .O(N__72555),
            .I(N__72536));
    LocalMux I__15981 (
            .O(N__72552),
            .I(N__72532));
    InMux I__15980 (
            .O(N__72551),
            .I(N__72529));
    InMux I__15979 (
            .O(N__72550),
            .I(N__72526));
    LocalMux I__15978 (
            .O(N__72547),
            .I(N__72523));
    Span4Mux_v I__15977 (
            .O(N__72544),
            .I(N__72520));
    LocalMux I__15976 (
            .O(N__72541),
            .I(N__72517));
    InMux I__15975 (
            .O(N__72540),
            .I(N__72511));
    InMux I__15974 (
            .O(N__72539),
            .I(N__72508));
    Span4Mux_v I__15973 (
            .O(N__72536),
            .I(N__72505));
    InMux I__15972 (
            .O(N__72535),
            .I(N__72502));
    Span4Mux_h I__15971 (
            .O(N__72532),
            .I(N__72498));
    LocalMux I__15970 (
            .O(N__72529),
            .I(N__72495));
    LocalMux I__15969 (
            .O(N__72526),
            .I(N__72492));
    Span4Mux_v I__15968 (
            .O(N__72523),
            .I(N__72488));
    Span4Mux_v I__15967 (
            .O(N__72520),
            .I(N__72485));
    Span4Mux_v I__15966 (
            .O(N__72517),
            .I(N__72482));
    InMux I__15965 (
            .O(N__72516),
            .I(N__72479));
    InMux I__15964 (
            .O(N__72515),
            .I(N__72476));
    InMux I__15963 (
            .O(N__72514),
            .I(N__72473));
    LocalMux I__15962 (
            .O(N__72511),
            .I(N__72470));
    LocalMux I__15961 (
            .O(N__72508),
            .I(N__72467));
    Span4Mux_v I__15960 (
            .O(N__72505),
            .I(N__72464));
    LocalMux I__15959 (
            .O(N__72502),
            .I(N__72461));
    InMux I__15958 (
            .O(N__72501),
            .I(N__72458));
    Span4Mux_h I__15957 (
            .O(N__72498),
            .I(N__72455));
    Span4Mux_v I__15956 (
            .O(N__72495),
            .I(N__72452));
    Span4Mux_h I__15955 (
            .O(N__72492),
            .I(N__72449));
    InMux I__15954 (
            .O(N__72491),
            .I(N__72446));
    Span4Mux_h I__15953 (
            .O(N__72488),
            .I(N__72443));
    Sp12to4 I__15952 (
            .O(N__72485),
            .I(N__72436));
    Sp12to4 I__15951 (
            .O(N__72482),
            .I(N__72436));
    LocalMux I__15950 (
            .O(N__72479),
            .I(N__72436));
    LocalMux I__15949 (
            .O(N__72476),
            .I(N__72431));
    LocalMux I__15948 (
            .O(N__72473),
            .I(N__72431));
    Span4Mux_h I__15947 (
            .O(N__72470),
            .I(N__72426));
    Span4Mux_v I__15946 (
            .O(N__72467),
            .I(N__72426));
    Span4Mux_h I__15945 (
            .O(N__72464),
            .I(N__72419));
    Span4Mux_v I__15944 (
            .O(N__72461),
            .I(N__72419));
    LocalMux I__15943 (
            .O(N__72458),
            .I(N__72419));
    Span4Mux_v I__15942 (
            .O(N__72455),
            .I(N__72410));
    Span4Mux_h I__15941 (
            .O(N__72452),
            .I(N__72410));
    Span4Mux_v I__15940 (
            .O(N__72449),
            .I(N__72410));
    LocalMux I__15939 (
            .O(N__72446),
            .I(N__72410));
    Odrv4 I__15938 (
            .O(N__72443),
            .I(n34));
    Odrv12 I__15937 (
            .O(N__72436),
            .I(n34));
    Odrv12 I__15936 (
            .O(N__72431),
            .I(n34));
    Odrv4 I__15935 (
            .O(N__72426),
            .I(n34));
    Odrv4 I__15934 (
            .O(N__72419),
            .I(n34));
    Odrv4 I__15933 (
            .O(N__72410),
            .I(n34));
    CascadeMux I__15932 (
            .O(N__72397),
            .I(N__72394));
    InMux I__15931 (
            .O(N__72394),
            .I(N__72390));
    InMux I__15930 (
            .O(N__72393),
            .I(N__72387));
    LocalMux I__15929 (
            .O(N__72390),
            .I(REG_mem_31_8));
    LocalMux I__15928 (
            .O(N__72387),
            .I(REG_mem_31_8));
    InMux I__15927 (
            .O(N__72382),
            .I(N__72376));
    InMux I__15926 (
            .O(N__72381),
            .I(N__72376));
    LocalMux I__15925 (
            .O(N__72376),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_8 ));
    CascadeMux I__15924 (
            .O(N__72373),
            .I(N__72370));
    InMux I__15923 (
            .O(N__72370),
            .I(N__72367));
    LocalMux I__15922 (
            .O(N__72367),
            .I(N__72363));
    InMux I__15921 (
            .O(N__72366),
            .I(N__72360));
    Span12Mux_h I__15920 (
            .O(N__72363),
            .I(N__72355));
    LocalMux I__15919 (
            .O(N__72360),
            .I(N__72355));
    Odrv12 I__15918 (
            .O(N__72355),
            .I(REG_mem_23_8));
    InMux I__15917 (
            .O(N__72352),
            .I(N__72348));
    CascadeMux I__15916 (
            .O(N__72351),
            .I(N__72345));
    LocalMux I__15915 (
            .O(N__72348),
            .I(N__72342));
    InMux I__15914 (
            .O(N__72345),
            .I(N__72339));
    Odrv4 I__15913 (
            .O(N__72342),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_8 ));
    LocalMux I__15912 (
            .O(N__72339),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_8 ));
    CascadeMux I__15911 (
            .O(N__72334),
            .I(N__72330));
    InMux I__15910 (
            .O(N__72333),
            .I(N__72327));
    InMux I__15909 (
            .O(N__72330),
            .I(N__72324));
    LocalMux I__15908 (
            .O(N__72327),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_8 ));
    LocalMux I__15907 (
            .O(N__72324),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_8 ));
    CascadeMux I__15906 (
            .O(N__72319),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14060_cascade_ ));
    InMux I__15905 (
            .O(N__72316),
            .I(N__72310));
    InMux I__15904 (
            .O(N__72315),
            .I(N__72310));
    LocalMux I__15903 (
            .O(N__72310),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_8 ));
    InMux I__15902 (
            .O(N__72307),
            .I(N__72304));
    LocalMux I__15901 (
            .O(N__72304),
            .I(N__72301));
    Span4Mux_v I__15900 (
            .O(N__72301),
            .I(N__72297));
    InMux I__15899 (
            .O(N__72300),
            .I(N__72294));
    Odrv4 I__15898 (
            .O(N__72297),
            .I(REG_mem_15_2));
    LocalMux I__15897 (
            .O(N__72294),
            .I(REG_mem_15_2));
    InMux I__15896 (
            .O(N__72289),
            .I(N__72286));
    LocalMux I__15895 (
            .O(N__72286),
            .I(N__72282));
    InMux I__15894 (
            .O(N__72285),
            .I(N__72279));
    Odrv12 I__15893 (
            .O(N__72282),
            .I(REG_mem_14_2));
    LocalMux I__15892 (
            .O(N__72279),
            .I(REG_mem_14_2));
    InMux I__15891 (
            .O(N__72274),
            .I(N__72271));
    LocalMux I__15890 (
            .O(N__72271),
            .I(N__72268));
    Odrv4 I__15889 (
            .O(N__72268),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11858 ));
    InMux I__15888 (
            .O(N__72265),
            .I(N__72258));
    InMux I__15887 (
            .O(N__72264),
            .I(N__72254));
    InMux I__15886 (
            .O(N__72263),
            .I(N__72251));
    InMux I__15885 (
            .O(N__72262),
            .I(N__72248));
    InMux I__15884 (
            .O(N__72261),
            .I(N__72240));
    LocalMux I__15883 (
            .O(N__72258),
            .I(N__72237));
    InMux I__15882 (
            .O(N__72257),
            .I(N__72234));
    LocalMux I__15881 (
            .O(N__72254),
            .I(N__72230));
    LocalMux I__15880 (
            .O(N__72251),
            .I(N__72225));
    LocalMux I__15879 (
            .O(N__72248),
            .I(N__72222));
    InMux I__15878 (
            .O(N__72247),
            .I(N__72219));
    InMux I__15877 (
            .O(N__72246),
            .I(N__72214));
    InMux I__15876 (
            .O(N__72245),
            .I(N__72214));
    InMux I__15875 (
            .O(N__72244),
            .I(N__72211));
    InMux I__15874 (
            .O(N__72243),
            .I(N__72208));
    LocalMux I__15873 (
            .O(N__72240),
            .I(N__72204));
    Span4Mux_h I__15872 (
            .O(N__72237),
            .I(N__72200));
    LocalMux I__15871 (
            .O(N__72234),
            .I(N__72197));
    InMux I__15870 (
            .O(N__72233),
            .I(N__72194));
    Span4Mux_v I__15869 (
            .O(N__72230),
            .I(N__72191));
    InMux I__15868 (
            .O(N__72229),
            .I(N__72188));
    InMux I__15867 (
            .O(N__72228),
            .I(N__72185));
    Span4Mux_v I__15866 (
            .O(N__72225),
            .I(N__72182));
    Span4Mux_v I__15865 (
            .O(N__72222),
            .I(N__72177));
    LocalMux I__15864 (
            .O(N__72219),
            .I(N__72177));
    LocalMux I__15863 (
            .O(N__72214),
            .I(N__72172));
    LocalMux I__15862 (
            .O(N__72211),
            .I(N__72172));
    LocalMux I__15861 (
            .O(N__72208),
            .I(N__72169));
    InMux I__15860 (
            .O(N__72207),
            .I(N__72166));
    Span4Mux_v I__15859 (
            .O(N__72204),
            .I(N__72163));
    InMux I__15858 (
            .O(N__72203),
            .I(N__72160));
    Span4Mux_h I__15857 (
            .O(N__72200),
            .I(N__72155));
    Span4Mux_v I__15856 (
            .O(N__72197),
            .I(N__72155));
    LocalMux I__15855 (
            .O(N__72194),
            .I(N__72148));
    Sp12to4 I__15854 (
            .O(N__72191),
            .I(N__72148));
    LocalMux I__15853 (
            .O(N__72188),
            .I(N__72148));
    LocalMux I__15852 (
            .O(N__72185),
            .I(N__72145));
    Span4Mux_h I__15851 (
            .O(N__72182),
            .I(N__72136));
    Span4Mux_v I__15850 (
            .O(N__72177),
            .I(N__72136));
    Span4Mux_h I__15849 (
            .O(N__72172),
            .I(N__72136));
    Span4Mux_h I__15848 (
            .O(N__72169),
            .I(N__72136));
    LocalMux I__15847 (
            .O(N__72166),
            .I(N__72133));
    Span4Mux_h I__15846 (
            .O(N__72163),
            .I(N__72128));
    LocalMux I__15845 (
            .O(N__72160),
            .I(N__72128));
    Odrv4 I__15844 (
            .O(N__72155),
            .I(n14));
    Odrv12 I__15843 (
            .O(N__72148),
            .I(n14));
    Odrv12 I__15842 (
            .O(N__72145),
            .I(n14));
    Odrv4 I__15841 (
            .O(N__72136),
            .I(n14));
    Odrv4 I__15840 (
            .O(N__72133),
            .I(n14));
    Odrv4 I__15839 (
            .O(N__72128),
            .I(n14));
    InMux I__15838 (
            .O(N__72115),
            .I(N__72106));
    InMux I__15837 (
            .O(N__72114),
            .I(N__72102));
    InMux I__15836 (
            .O(N__72113),
            .I(N__72097));
    InMux I__15835 (
            .O(N__72112),
            .I(N__72094));
    InMux I__15834 (
            .O(N__72111),
            .I(N__72089));
    InMux I__15833 (
            .O(N__72110),
            .I(N__72086));
    InMux I__15832 (
            .O(N__72109),
            .I(N__72082));
    LocalMux I__15831 (
            .O(N__72106),
            .I(N__72079));
    InMux I__15830 (
            .O(N__72105),
            .I(N__72076));
    LocalMux I__15829 (
            .O(N__72102),
            .I(N__72072));
    InMux I__15828 (
            .O(N__72101),
            .I(N__72069));
    InMux I__15827 (
            .O(N__72100),
            .I(N__72066));
    LocalMux I__15826 (
            .O(N__72097),
            .I(N__72062));
    LocalMux I__15825 (
            .O(N__72094),
            .I(N__72059));
    InMux I__15824 (
            .O(N__72093),
            .I(N__72056));
    InMux I__15823 (
            .O(N__72092),
            .I(N__72053));
    LocalMux I__15822 (
            .O(N__72089),
            .I(N__72050));
    LocalMux I__15821 (
            .O(N__72086),
            .I(N__72047));
    InMux I__15820 (
            .O(N__72085),
            .I(N__72044));
    LocalMux I__15819 (
            .O(N__72082),
            .I(N__72041));
    Span4Mux_h I__15818 (
            .O(N__72079),
            .I(N__72038));
    LocalMux I__15817 (
            .O(N__72076),
            .I(N__72035));
    InMux I__15816 (
            .O(N__72075),
            .I(N__72032));
    Span4Mux_v I__15815 (
            .O(N__72072),
            .I(N__72029));
    LocalMux I__15814 (
            .O(N__72069),
            .I(N__72026));
    LocalMux I__15813 (
            .O(N__72066),
            .I(N__72023));
    InMux I__15812 (
            .O(N__72065),
            .I(N__72020));
    Span4Mux_v I__15811 (
            .O(N__72062),
            .I(N__72016));
    Span4Mux_v I__15810 (
            .O(N__72059),
            .I(N__72013));
    LocalMux I__15809 (
            .O(N__72056),
            .I(N__72010));
    LocalMux I__15808 (
            .O(N__72053),
            .I(N__72007));
    Span4Mux_h I__15807 (
            .O(N__72050),
            .I(N__72004));
    Span4Mux_h I__15806 (
            .O(N__72047),
            .I(N__71999));
    LocalMux I__15805 (
            .O(N__72044),
            .I(N__71999));
    Span4Mux_v I__15804 (
            .O(N__72041),
            .I(N__71996));
    Span4Mux_h I__15803 (
            .O(N__72038),
            .I(N__71989));
    Span4Mux_v I__15802 (
            .O(N__72035),
            .I(N__71989));
    LocalMux I__15801 (
            .O(N__72032),
            .I(N__71989));
    Span4Mux_h I__15800 (
            .O(N__72029),
            .I(N__71980));
    Span4Mux_h I__15799 (
            .O(N__72026),
            .I(N__71980));
    Span4Mux_v I__15798 (
            .O(N__72023),
            .I(N__71980));
    LocalMux I__15797 (
            .O(N__72020),
            .I(N__71980));
    InMux I__15796 (
            .O(N__72019),
            .I(N__71977));
    Span4Mux_h I__15795 (
            .O(N__72016),
            .I(N__71974));
    Span4Mux_h I__15794 (
            .O(N__72013),
            .I(N__71969));
    Span4Mux_v I__15793 (
            .O(N__72010),
            .I(N__71969));
    Span4Mux_v I__15792 (
            .O(N__72007),
            .I(N__71966));
    Span4Mux_h I__15791 (
            .O(N__72004),
            .I(N__71961));
    Span4Mux_v I__15790 (
            .O(N__71999),
            .I(N__71961));
    Span4Mux_v I__15789 (
            .O(N__71996),
            .I(N__71952));
    Span4Mux_v I__15788 (
            .O(N__71989),
            .I(N__71952));
    Span4Mux_h I__15787 (
            .O(N__71980),
            .I(N__71952));
    LocalMux I__15786 (
            .O(N__71977),
            .I(N__71952));
    Odrv4 I__15785 (
            .O(N__71974),
            .I(n46));
    Odrv4 I__15784 (
            .O(N__71969),
            .I(n46));
    Odrv4 I__15783 (
            .O(N__71966),
            .I(n46));
    Odrv4 I__15782 (
            .O(N__71961),
            .I(n46));
    Odrv4 I__15781 (
            .O(N__71952),
            .I(n46));
    CascadeMux I__15780 (
            .O(N__71941),
            .I(N__71938));
    InMux I__15779 (
            .O(N__71938),
            .I(N__71934));
    InMux I__15778 (
            .O(N__71937),
            .I(N__71931));
    LocalMux I__15777 (
            .O(N__71934),
            .I(REG_mem_19_8));
    LocalMux I__15776 (
            .O(N__71931),
            .I(REG_mem_19_8));
    InMux I__15775 (
            .O(N__71926),
            .I(N__71923));
    LocalMux I__15774 (
            .O(N__71923),
            .I(N__71920));
    Span4Mux_v I__15773 (
            .O(N__71920),
            .I(N__71916));
    InMux I__15772 (
            .O(N__71919),
            .I(N__71913));
    Odrv4 I__15771 (
            .O(N__71916),
            .I(REG_mem_47_6));
    LocalMux I__15770 (
            .O(N__71913),
            .I(REG_mem_47_6));
    InMux I__15769 (
            .O(N__71908),
            .I(N__71905));
    LocalMux I__15768 (
            .O(N__71905),
            .I(N__71899));
    InMux I__15767 (
            .O(N__71904),
            .I(N__71896));
    InMux I__15766 (
            .O(N__71903),
            .I(N__71893));
    InMux I__15765 (
            .O(N__71902),
            .I(N__71889));
    Span4Mux_v I__15764 (
            .O(N__71899),
            .I(N__71879));
    LocalMux I__15763 (
            .O(N__71896),
            .I(N__71879));
    LocalMux I__15762 (
            .O(N__71893),
            .I(N__71875));
    InMux I__15761 (
            .O(N__71892),
            .I(N__71872));
    LocalMux I__15760 (
            .O(N__71889),
            .I(N__71869));
    InMux I__15759 (
            .O(N__71888),
            .I(N__71866));
    InMux I__15758 (
            .O(N__71887),
            .I(N__71860));
    InMux I__15757 (
            .O(N__71886),
            .I(N__71857));
    InMux I__15756 (
            .O(N__71885),
            .I(N__71854));
    InMux I__15755 (
            .O(N__71884),
            .I(N__71851));
    Span4Mux_v I__15754 (
            .O(N__71879),
            .I(N__71847));
    InMux I__15753 (
            .O(N__71878),
            .I(N__71844));
    Span4Mux_v I__15752 (
            .O(N__71875),
            .I(N__71839));
    LocalMux I__15751 (
            .O(N__71872),
            .I(N__71839));
    Span4Mux_h I__15750 (
            .O(N__71869),
            .I(N__71836));
    LocalMux I__15749 (
            .O(N__71866),
            .I(N__71833));
    InMux I__15748 (
            .O(N__71865),
            .I(N__71830));
    InMux I__15747 (
            .O(N__71864),
            .I(N__71827));
    InMux I__15746 (
            .O(N__71863),
            .I(N__71824));
    LocalMux I__15745 (
            .O(N__71860),
            .I(N__71821));
    LocalMux I__15744 (
            .O(N__71857),
            .I(N__71818));
    LocalMux I__15743 (
            .O(N__71854),
            .I(N__71813));
    LocalMux I__15742 (
            .O(N__71851),
            .I(N__71813));
    InMux I__15741 (
            .O(N__71850),
            .I(N__71810));
    Span4Mux_h I__15740 (
            .O(N__71847),
            .I(N__71806));
    LocalMux I__15739 (
            .O(N__71844),
            .I(N__71803));
    Span4Mux_v I__15738 (
            .O(N__71839),
            .I(N__71796));
    Span4Mux_h I__15737 (
            .O(N__71836),
            .I(N__71796));
    Span4Mux_v I__15736 (
            .O(N__71833),
            .I(N__71796));
    LocalMux I__15735 (
            .O(N__71830),
            .I(N__71789));
    LocalMux I__15734 (
            .O(N__71827),
            .I(N__71789));
    LocalMux I__15733 (
            .O(N__71824),
            .I(N__71789));
    Span4Mux_h I__15732 (
            .O(N__71821),
            .I(N__71780));
    Span4Mux_h I__15731 (
            .O(N__71818),
            .I(N__71780));
    Span4Mux_v I__15730 (
            .O(N__71813),
            .I(N__71780));
    LocalMux I__15729 (
            .O(N__71810),
            .I(N__71780));
    InMux I__15728 (
            .O(N__71809),
            .I(N__71777));
    Odrv4 I__15727 (
            .O(N__71806),
            .I(n20));
    Odrv12 I__15726 (
            .O(N__71803),
            .I(n20));
    Odrv4 I__15725 (
            .O(N__71796),
            .I(n20));
    Odrv12 I__15724 (
            .O(N__71789),
            .I(n20));
    Odrv4 I__15723 (
            .O(N__71780),
            .I(n20));
    LocalMux I__15722 (
            .O(N__71777),
            .I(n20));
    InMux I__15721 (
            .O(N__71764),
            .I(N__71759));
    InMux I__15720 (
            .O(N__71763),
            .I(N__71756));
    InMux I__15719 (
            .O(N__71762),
            .I(N__71752));
    LocalMux I__15718 (
            .O(N__71759),
            .I(N__71749));
    LocalMux I__15717 (
            .O(N__71756),
            .I(N__71746));
    InMux I__15716 (
            .O(N__71755),
            .I(N__71743));
    LocalMux I__15715 (
            .O(N__71752),
            .I(N__71733));
    Span4Mux_h I__15714 (
            .O(N__71749),
            .I(N__71730));
    Span4Mux_v I__15713 (
            .O(N__71746),
            .I(N__71727));
    LocalMux I__15712 (
            .O(N__71743),
            .I(N__71724));
    InMux I__15711 (
            .O(N__71742),
            .I(N__71721));
    InMux I__15710 (
            .O(N__71741),
            .I(N__71718));
    InMux I__15709 (
            .O(N__71740),
            .I(N__71715));
    InMux I__15708 (
            .O(N__71739),
            .I(N__71712));
    InMux I__15707 (
            .O(N__71738),
            .I(N__71707));
    InMux I__15706 (
            .O(N__71737),
            .I(N__71704));
    InMux I__15705 (
            .O(N__71736),
            .I(N__71700));
    Span4Mux_v I__15704 (
            .O(N__71733),
            .I(N__71696));
    Span4Mux_v I__15703 (
            .O(N__71730),
            .I(N__71689));
    Span4Mux_h I__15702 (
            .O(N__71727),
            .I(N__71689));
    Span4Mux_h I__15701 (
            .O(N__71724),
            .I(N__71689));
    LocalMux I__15700 (
            .O(N__71721),
            .I(N__71686));
    LocalMux I__15699 (
            .O(N__71718),
            .I(N__71679));
    LocalMux I__15698 (
            .O(N__71715),
            .I(N__71679));
    LocalMux I__15697 (
            .O(N__71712),
            .I(N__71679));
    InMux I__15696 (
            .O(N__71711),
            .I(N__71676));
    InMux I__15695 (
            .O(N__71710),
            .I(N__71673));
    LocalMux I__15694 (
            .O(N__71707),
            .I(N__71670));
    LocalMux I__15693 (
            .O(N__71704),
            .I(N__71667));
    InMux I__15692 (
            .O(N__71703),
            .I(N__71664));
    LocalMux I__15691 (
            .O(N__71700),
            .I(N__71661));
    InMux I__15690 (
            .O(N__71699),
            .I(N__71658));
    Span4Mux_h I__15689 (
            .O(N__71696),
            .I(N__71654));
    Sp12to4 I__15688 (
            .O(N__71689),
            .I(N__71643));
    Sp12to4 I__15687 (
            .O(N__71686),
            .I(N__71643));
    Span12Mux_h I__15686 (
            .O(N__71679),
            .I(N__71643));
    LocalMux I__15685 (
            .O(N__71676),
            .I(N__71643));
    LocalMux I__15684 (
            .O(N__71673),
            .I(N__71643));
    Span4Mux_v I__15683 (
            .O(N__71670),
            .I(N__71636));
    Span4Mux_h I__15682 (
            .O(N__71667),
            .I(N__71636));
    LocalMux I__15681 (
            .O(N__71664),
            .I(N__71636));
    Span12Mux_h I__15680 (
            .O(N__71661),
            .I(N__71631));
    LocalMux I__15679 (
            .O(N__71658),
            .I(N__71631));
    InMux I__15678 (
            .O(N__71657),
            .I(N__71628));
    Odrv4 I__15677 (
            .O(N__71654),
            .I(n21));
    Odrv12 I__15676 (
            .O(N__71643),
            .I(n21));
    Odrv4 I__15675 (
            .O(N__71636),
            .I(n21));
    Odrv12 I__15674 (
            .O(N__71631),
            .I(n21));
    LocalMux I__15673 (
            .O(N__71628),
            .I(n21));
    InMux I__15672 (
            .O(N__71617),
            .I(N__71614));
    LocalMux I__15671 (
            .O(N__71614),
            .I(N__71610));
    InMux I__15670 (
            .O(N__71613),
            .I(N__71607));
    Odrv4 I__15669 (
            .O(N__71610),
            .I(REG_mem_23_1));
    LocalMux I__15668 (
            .O(N__71607),
            .I(REG_mem_23_1));
    InMux I__15667 (
            .O(N__71602),
            .I(N__71591));
    InMux I__15666 (
            .O(N__71601),
            .I(N__71591));
    InMux I__15665 (
            .O(N__71600),
            .I(N__71588));
    InMux I__15664 (
            .O(N__71599),
            .I(N__71581));
    InMux I__15663 (
            .O(N__71598),
            .I(N__71581));
    InMux I__15662 (
            .O(N__71597),
            .I(N__71578));
    InMux I__15661 (
            .O(N__71596),
            .I(N__71575));
    LocalMux I__15660 (
            .O(N__71591),
            .I(N__71570));
    LocalMux I__15659 (
            .O(N__71588),
            .I(N__71570));
    CascadeMux I__15658 (
            .O(N__71587),
            .I(N__71565));
    CascadeMux I__15657 (
            .O(N__71586),
            .I(N__71562));
    LocalMux I__15656 (
            .O(N__71581),
            .I(N__71546));
    LocalMux I__15655 (
            .O(N__71578),
            .I(N__71546));
    LocalMux I__15654 (
            .O(N__71575),
            .I(N__71535));
    Span4Mux_v I__15653 (
            .O(N__71570),
            .I(N__71535));
    InMux I__15652 (
            .O(N__71569),
            .I(N__71532));
    CascadeMux I__15651 (
            .O(N__71568),
            .I(N__71529));
    InMux I__15650 (
            .O(N__71565),
            .I(N__71512));
    InMux I__15649 (
            .O(N__71562),
            .I(N__71512));
    InMux I__15648 (
            .O(N__71561),
            .I(N__71507));
    InMux I__15647 (
            .O(N__71560),
            .I(N__71507));
    InMux I__15646 (
            .O(N__71559),
            .I(N__71504));
    InMux I__15645 (
            .O(N__71558),
            .I(N__71499));
    InMux I__15644 (
            .O(N__71557),
            .I(N__71499));
    InMux I__15643 (
            .O(N__71556),
            .I(N__71495));
    InMux I__15642 (
            .O(N__71555),
            .I(N__71487));
    InMux I__15641 (
            .O(N__71554),
            .I(N__71487));
    InMux I__15640 (
            .O(N__71553),
            .I(N__71480));
    InMux I__15639 (
            .O(N__71552),
            .I(N__71480));
    InMux I__15638 (
            .O(N__71551),
            .I(N__71480));
    Span4Mux_v I__15637 (
            .O(N__71546),
            .I(N__71477));
    InMux I__15636 (
            .O(N__71545),
            .I(N__71472));
    InMux I__15635 (
            .O(N__71544),
            .I(N__71472));
    InMux I__15634 (
            .O(N__71543),
            .I(N__71463));
    InMux I__15633 (
            .O(N__71542),
            .I(N__71463));
    InMux I__15632 (
            .O(N__71541),
            .I(N__71463));
    InMux I__15631 (
            .O(N__71540),
            .I(N__71458));
    Span4Mux_h I__15630 (
            .O(N__71535),
            .I(N__71450));
    LocalMux I__15629 (
            .O(N__71532),
            .I(N__71450));
    InMux I__15628 (
            .O(N__71529),
            .I(N__71447));
    InMux I__15627 (
            .O(N__71528),
            .I(N__71444));
    InMux I__15626 (
            .O(N__71527),
            .I(N__71437));
    InMux I__15625 (
            .O(N__71526),
            .I(N__71437));
    InMux I__15624 (
            .O(N__71525),
            .I(N__71437));
    InMux I__15623 (
            .O(N__71524),
            .I(N__71432));
    InMux I__15622 (
            .O(N__71523),
            .I(N__71432));
    InMux I__15621 (
            .O(N__71522),
            .I(N__71425));
    InMux I__15620 (
            .O(N__71521),
            .I(N__71425));
    InMux I__15619 (
            .O(N__71520),
            .I(N__71425));
    InMux I__15618 (
            .O(N__71519),
            .I(N__71418));
    InMux I__15617 (
            .O(N__71518),
            .I(N__71418));
    InMux I__15616 (
            .O(N__71517),
            .I(N__71418));
    LocalMux I__15615 (
            .O(N__71512),
            .I(N__71409));
    LocalMux I__15614 (
            .O(N__71507),
            .I(N__71409));
    LocalMux I__15613 (
            .O(N__71504),
            .I(N__71409));
    LocalMux I__15612 (
            .O(N__71499),
            .I(N__71409));
    InMux I__15611 (
            .O(N__71498),
            .I(N__71406));
    LocalMux I__15610 (
            .O(N__71495),
            .I(N__71401));
    InMux I__15609 (
            .O(N__71494),
            .I(N__71395));
    InMux I__15608 (
            .O(N__71493),
            .I(N__71390));
    InMux I__15607 (
            .O(N__71492),
            .I(N__71390));
    LocalMux I__15606 (
            .O(N__71487),
            .I(N__71387));
    LocalMux I__15605 (
            .O(N__71480),
            .I(N__71384));
    Span4Mux_h I__15604 (
            .O(N__71477),
            .I(N__71379));
    LocalMux I__15603 (
            .O(N__71472),
            .I(N__71379));
    InMux I__15602 (
            .O(N__71471),
            .I(N__71376));
    InMux I__15601 (
            .O(N__71470),
            .I(N__71373));
    LocalMux I__15600 (
            .O(N__71463),
            .I(N__71370));
    InMux I__15599 (
            .O(N__71462),
            .I(N__71365));
    InMux I__15598 (
            .O(N__71461),
            .I(N__71365));
    LocalMux I__15597 (
            .O(N__71458),
            .I(N__71362));
    InMux I__15596 (
            .O(N__71457),
            .I(N__71359));
    InMux I__15595 (
            .O(N__71456),
            .I(N__71354));
    InMux I__15594 (
            .O(N__71455),
            .I(N__71350));
    Span4Mux_v I__15593 (
            .O(N__71450),
            .I(N__71347));
    LocalMux I__15592 (
            .O(N__71447),
            .I(N__71332));
    LocalMux I__15591 (
            .O(N__71444),
            .I(N__71332));
    LocalMux I__15590 (
            .O(N__71437),
            .I(N__71332));
    LocalMux I__15589 (
            .O(N__71432),
            .I(N__71332));
    LocalMux I__15588 (
            .O(N__71425),
            .I(N__71332));
    LocalMux I__15587 (
            .O(N__71418),
            .I(N__71332));
    Span4Mux_v I__15586 (
            .O(N__71409),
            .I(N__71332));
    LocalMux I__15585 (
            .O(N__71406),
            .I(N__71326));
    InMux I__15584 (
            .O(N__71405),
            .I(N__71322));
    InMux I__15583 (
            .O(N__71404),
            .I(N__71319));
    Span4Mux_h I__15582 (
            .O(N__71401),
            .I(N__71316));
    InMux I__15581 (
            .O(N__71400),
            .I(N__71309));
    InMux I__15580 (
            .O(N__71399),
            .I(N__71309));
    InMux I__15579 (
            .O(N__71398),
            .I(N__71309));
    LocalMux I__15578 (
            .O(N__71395),
            .I(N__71304));
    LocalMux I__15577 (
            .O(N__71390),
            .I(N__71304));
    Span4Mux_v I__15576 (
            .O(N__71387),
            .I(N__71299));
    Span4Mux_v I__15575 (
            .O(N__71384),
            .I(N__71299));
    Span4Mux_h I__15574 (
            .O(N__71379),
            .I(N__71296));
    LocalMux I__15573 (
            .O(N__71376),
            .I(N__71290));
    LocalMux I__15572 (
            .O(N__71373),
            .I(N__71290));
    Span4Mux_v I__15571 (
            .O(N__71370),
            .I(N__71285));
    LocalMux I__15570 (
            .O(N__71365),
            .I(N__71285));
    Span4Mux_v I__15569 (
            .O(N__71362),
            .I(N__71280));
    LocalMux I__15568 (
            .O(N__71359),
            .I(N__71280));
    InMux I__15567 (
            .O(N__71358),
            .I(N__71277));
    InMux I__15566 (
            .O(N__71357),
            .I(N__71274));
    LocalMux I__15565 (
            .O(N__71354),
            .I(N__71271));
    InMux I__15564 (
            .O(N__71353),
            .I(N__71268));
    LocalMux I__15563 (
            .O(N__71350),
            .I(N__71261));
    Span4Mux_h I__15562 (
            .O(N__71347),
            .I(N__71261));
    Span4Mux_v I__15561 (
            .O(N__71332),
            .I(N__71261));
    InMux I__15560 (
            .O(N__71331),
            .I(N__71258));
    InMux I__15559 (
            .O(N__71330),
            .I(N__71255));
    InMux I__15558 (
            .O(N__71329),
            .I(N__71252));
    Sp12to4 I__15557 (
            .O(N__71326),
            .I(N__71249));
    InMux I__15556 (
            .O(N__71325),
            .I(N__71246));
    LocalMux I__15555 (
            .O(N__71322),
            .I(N__71239));
    LocalMux I__15554 (
            .O(N__71319),
            .I(N__71239));
    Span4Mux_v I__15553 (
            .O(N__71316),
            .I(N__71239));
    LocalMux I__15552 (
            .O(N__71309),
            .I(N__71230));
    Span4Mux_v I__15551 (
            .O(N__71304),
            .I(N__71230));
    Span4Mux_h I__15550 (
            .O(N__71299),
            .I(N__71230));
    Span4Mux_v I__15549 (
            .O(N__71296),
            .I(N__71230));
    InMux I__15548 (
            .O(N__71295),
            .I(N__71227));
    Span4Mux_v I__15547 (
            .O(N__71290),
            .I(N__71220));
    Span4Mux_v I__15546 (
            .O(N__71285),
            .I(N__71220));
    Span4Mux_h I__15545 (
            .O(N__71280),
            .I(N__71220));
    LocalMux I__15544 (
            .O(N__71277),
            .I(N__71215));
    LocalMux I__15543 (
            .O(N__71274),
            .I(N__71215));
    Span4Mux_v I__15542 (
            .O(N__71271),
            .I(N__71212));
    LocalMux I__15541 (
            .O(N__71268),
            .I(N__71207));
    Sp12to4 I__15540 (
            .O(N__71261),
            .I(N__71207));
    LocalMux I__15539 (
            .O(N__71258),
            .I(N__71198));
    LocalMux I__15538 (
            .O(N__71255),
            .I(N__71198));
    LocalMux I__15537 (
            .O(N__71252),
            .I(N__71198));
    Span12Mux_h I__15536 (
            .O(N__71249),
            .I(N__71198));
    LocalMux I__15535 (
            .O(N__71246),
            .I(N__71191));
    Span4Mux_v I__15534 (
            .O(N__71239),
            .I(N__71191));
    Span4Mux_h I__15533 (
            .O(N__71230),
            .I(N__71191));
    LocalMux I__15532 (
            .O(N__71227),
            .I(N__71186));
    Span4Mux_h I__15531 (
            .O(N__71220),
            .I(N__71186));
    Odrv4 I__15530 (
            .O(N__71215),
            .I(dc32_fifo_data_in_0));
    Odrv4 I__15529 (
            .O(N__71212),
            .I(dc32_fifo_data_in_0));
    Odrv12 I__15528 (
            .O(N__71207),
            .I(dc32_fifo_data_in_0));
    Odrv12 I__15527 (
            .O(N__71198),
            .I(dc32_fifo_data_in_0));
    Odrv4 I__15526 (
            .O(N__71191),
            .I(dc32_fifo_data_in_0));
    Odrv4 I__15525 (
            .O(N__71186),
            .I(dc32_fifo_data_in_0));
    InMux I__15524 (
            .O(N__71173),
            .I(N__71170));
    LocalMux I__15523 (
            .O(N__71170),
            .I(N__71166));
    InMux I__15522 (
            .O(N__71169),
            .I(N__71163));
    Odrv4 I__15521 (
            .O(N__71166),
            .I(REG_mem_58_0));
    LocalMux I__15520 (
            .O(N__71163),
            .I(REG_mem_58_0));
    InMux I__15519 (
            .O(N__71158),
            .I(N__71154));
    InMux I__15518 (
            .O(N__71157),
            .I(N__71151));
    LocalMux I__15517 (
            .O(N__71154),
            .I(REG_mem_5_6));
    LocalMux I__15516 (
            .O(N__71151),
            .I(REG_mem_5_6));
    InMux I__15515 (
            .O(N__71146),
            .I(N__71143));
    LocalMux I__15514 (
            .O(N__71143),
            .I(N__71139));
    CascadeMux I__15513 (
            .O(N__71142),
            .I(N__71136));
    Span4Mux_v I__15512 (
            .O(N__71139),
            .I(N__71133));
    InMux I__15511 (
            .O(N__71136),
            .I(N__71130));
    Odrv4 I__15510 (
            .O(N__71133),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_6 ));
    LocalMux I__15509 (
            .O(N__71130),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_6 ));
    CascadeMux I__15508 (
            .O(N__71125),
            .I(N__71122));
    InMux I__15507 (
            .O(N__71122),
            .I(N__71116));
    InMux I__15506 (
            .O(N__71121),
            .I(N__71116));
    LocalMux I__15505 (
            .O(N__71116),
            .I(REG_mem_58_6));
    InMux I__15504 (
            .O(N__71113),
            .I(N__71110));
    LocalMux I__15503 (
            .O(N__71110),
            .I(N__71106));
    CascadeMux I__15502 (
            .O(N__71109),
            .I(N__71103));
    Span4Mux_v I__15501 (
            .O(N__71106),
            .I(N__71100));
    InMux I__15500 (
            .O(N__71103),
            .I(N__71097));
    Odrv4 I__15499 (
            .O(N__71100),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_2 ));
    LocalMux I__15498 (
            .O(N__71097),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_2 ));
    CascadeMux I__15497 (
            .O(N__71092),
            .I(N__71088));
    InMux I__15496 (
            .O(N__71091),
            .I(N__71083));
    InMux I__15495 (
            .O(N__71088),
            .I(N__71083));
    LocalMux I__15494 (
            .O(N__71083),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_0 ));
    InMux I__15493 (
            .O(N__71080),
            .I(N__71077));
    LocalMux I__15492 (
            .O(N__71077),
            .I(N__71074));
    Span4Mux_v I__15491 (
            .O(N__71074),
            .I(N__71071));
    Span4Mux_h I__15490 (
            .O(N__71071),
            .I(N__71068));
    Span4Mux_h I__15489 (
            .O(N__71068),
            .I(N__71065));
    Odrv4 I__15488 (
            .O(N__71065),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12008 ));
    CascadeMux I__15487 (
            .O(N__71062),
            .I(N__71058));
    InMux I__15486 (
            .O(N__71061),
            .I(N__71055));
    InMux I__15485 (
            .O(N__71058),
            .I(N__71052));
    LocalMux I__15484 (
            .O(N__71055),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_1 ));
    LocalMux I__15483 (
            .O(N__71052),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_1 ));
    CascadeMux I__15482 (
            .O(N__71047),
            .I(N__71043));
    InMux I__15481 (
            .O(N__71046),
            .I(N__71040));
    InMux I__15480 (
            .O(N__71043),
            .I(N__71037));
    LocalMux I__15479 (
            .O(N__71040),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_1 ));
    LocalMux I__15478 (
            .O(N__71037),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_1 ));
    InMux I__15477 (
            .O(N__71032),
            .I(N__71029));
    LocalMux I__15476 (
            .O(N__71029),
            .I(N__71026));
    Odrv4 I__15475 (
            .O(N__71026),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11680 ));
    InMux I__15474 (
            .O(N__71023),
            .I(N__71019));
    InMux I__15473 (
            .O(N__71022),
            .I(N__71016));
    LocalMux I__15472 (
            .O(N__71019),
            .I(REG_mem_63_6));
    LocalMux I__15471 (
            .O(N__71016),
            .I(REG_mem_63_6));
    CascadeMux I__15470 (
            .O(N__71011),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14294_cascade_ ));
    InMux I__15469 (
            .O(N__71008),
            .I(N__71000));
    InMux I__15468 (
            .O(N__71007),
            .I(N__71000));
    InMux I__15467 (
            .O(N__71006),
            .I(N__70995));
    InMux I__15466 (
            .O(N__71005),
            .I(N__70992));
    LocalMux I__15465 (
            .O(N__71000),
            .I(N__70983));
    InMux I__15464 (
            .O(N__70999),
            .I(N__70978));
    InMux I__15463 (
            .O(N__70998),
            .I(N__70978));
    LocalMux I__15462 (
            .O(N__70995),
            .I(N__70969));
    LocalMux I__15461 (
            .O(N__70992),
            .I(N__70969));
    InMux I__15460 (
            .O(N__70991),
            .I(N__70966));
    InMux I__15459 (
            .O(N__70990),
            .I(N__70961));
    InMux I__15458 (
            .O(N__70989),
            .I(N__70956));
    InMux I__15457 (
            .O(N__70988),
            .I(N__70956));
    InMux I__15456 (
            .O(N__70987),
            .I(N__70951));
    InMux I__15455 (
            .O(N__70986),
            .I(N__70951));
    Span4Mux_v I__15454 (
            .O(N__70983),
            .I(N__70945));
    LocalMux I__15453 (
            .O(N__70978),
            .I(N__70942));
    InMux I__15452 (
            .O(N__70977),
            .I(N__70939));
    InMux I__15451 (
            .O(N__70976),
            .I(N__70932));
    InMux I__15450 (
            .O(N__70975),
            .I(N__70932));
    InMux I__15449 (
            .O(N__70974),
            .I(N__70929));
    Span4Mux_h I__15448 (
            .O(N__70969),
            .I(N__70925));
    LocalMux I__15447 (
            .O(N__70966),
            .I(N__70922));
    InMux I__15446 (
            .O(N__70965),
            .I(N__70919));
    InMux I__15445 (
            .O(N__70964),
            .I(N__70916));
    LocalMux I__15444 (
            .O(N__70961),
            .I(N__70912));
    LocalMux I__15443 (
            .O(N__70956),
            .I(N__70909));
    LocalMux I__15442 (
            .O(N__70951),
            .I(N__70906));
    InMux I__15441 (
            .O(N__70950),
            .I(N__70903));
    InMux I__15440 (
            .O(N__70949),
            .I(N__70898));
    InMux I__15439 (
            .O(N__70948),
            .I(N__70898));
    Span4Mux_v I__15438 (
            .O(N__70945),
            .I(N__70889));
    Span4Mux_v I__15437 (
            .O(N__70942),
            .I(N__70889));
    LocalMux I__15436 (
            .O(N__70939),
            .I(N__70889));
    InMux I__15435 (
            .O(N__70938),
            .I(N__70886));
    InMux I__15434 (
            .O(N__70937),
            .I(N__70883));
    LocalMux I__15433 (
            .O(N__70932),
            .I(N__70879));
    LocalMux I__15432 (
            .O(N__70929),
            .I(N__70876));
    InMux I__15431 (
            .O(N__70928),
            .I(N__70873));
    Span4Mux_v I__15430 (
            .O(N__70925),
            .I(N__70864));
    Span4Mux_h I__15429 (
            .O(N__70922),
            .I(N__70864));
    LocalMux I__15428 (
            .O(N__70919),
            .I(N__70864));
    LocalMux I__15427 (
            .O(N__70916),
            .I(N__70864));
    InMux I__15426 (
            .O(N__70915),
            .I(N__70861));
    Span4Mux_h I__15425 (
            .O(N__70912),
            .I(N__70857));
    Span4Mux_v I__15424 (
            .O(N__70909),
            .I(N__70852));
    Span4Mux_h I__15423 (
            .O(N__70906),
            .I(N__70852));
    LocalMux I__15422 (
            .O(N__70903),
            .I(N__70847));
    LocalMux I__15421 (
            .O(N__70898),
            .I(N__70847));
    InMux I__15420 (
            .O(N__70897),
            .I(N__70844));
    InMux I__15419 (
            .O(N__70896),
            .I(N__70841));
    Span4Mux_h I__15418 (
            .O(N__70889),
            .I(N__70838));
    LocalMux I__15417 (
            .O(N__70886),
            .I(N__70833));
    LocalMux I__15416 (
            .O(N__70883),
            .I(N__70833));
    InMux I__15415 (
            .O(N__70882),
            .I(N__70830));
    Span4Mux_v I__15414 (
            .O(N__70879),
            .I(N__70827));
    Span4Mux_h I__15413 (
            .O(N__70876),
            .I(N__70822));
    LocalMux I__15412 (
            .O(N__70873),
            .I(N__70822));
    Span4Mux_h I__15411 (
            .O(N__70864),
            .I(N__70817));
    LocalMux I__15410 (
            .O(N__70861),
            .I(N__70817));
    InMux I__15409 (
            .O(N__70860),
            .I(N__70814));
    Span4Mux_v I__15408 (
            .O(N__70857),
            .I(N__70807));
    Span4Mux_h I__15407 (
            .O(N__70852),
            .I(N__70807));
    Span4Mux_h I__15406 (
            .O(N__70847),
            .I(N__70804));
    LocalMux I__15405 (
            .O(N__70844),
            .I(N__70799));
    LocalMux I__15404 (
            .O(N__70841),
            .I(N__70799));
    Span4Mux_h I__15403 (
            .O(N__70838),
            .I(N__70792));
    Span4Mux_v I__15402 (
            .O(N__70833),
            .I(N__70792));
    LocalMux I__15401 (
            .O(N__70830),
            .I(N__70792));
    Span4Mux_v I__15400 (
            .O(N__70827),
            .I(N__70783));
    Span4Mux_v I__15399 (
            .O(N__70822),
            .I(N__70783));
    Span4Mux_h I__15398 (
            .O(N__70817),
            .I(N__70783));
    LocalMux I__15397 (
            .O(N__70814),
            .I(N__70783));
    InMux I__15396 (
            .O(N__70813),
            .I(N__70778));
    InMux I__15395 (
            .O(N__70812),
            .I(N__70778));
    Odrv4 I__15394 (
            .O(N__70807),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n63 ));
    Odrv4 I__15393 (
            .O(N__70804),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n63 ));
    Odrv12 I__15392 (
            .O(N__70799),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n63 ));
    Odrv4 I__15391 (
            .O(N__70792),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n63 ));
    Odrv4 I__15390 (
            .O(N__70783),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n63 ));
    LocalMux I__15389 (
            .O(N__70778),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n63 ));
    CascadeMux I__15388 (
            .O(N__70765),
            .I(N__70761));
    InMux I__15387 (
            .O(N__70764),
            .I(N__70756));
    InMux I__15386 (
            .O(N__70761),
            .I(N__70756));
    LocalMux I__15385 (
            .O(N__70756),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_6 ));
    CascadeMux I__15384 (
            .O(N__70753),
            .I(N__70749));
    InMux I__15383 (
            .O(N__70752),
            .I(N__70744));
    InMux I__15382 (
            .O(N__70749),
            .I(N__70744));
    LocalMux I__15381 (
            .O(N__70744),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_6 ));
    CascadeMux I__15380 (
            .O(N__70741),
            .I(N__70737));
    InMux I__15379 (
            .O(N__70740),
            .I(N__70732));
    InMux I__15378 (
            .O(N__70737),
            .I(N__70732));
    LocalMux I__15377 (
            .O(N__70732),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_6 ));
    CascadeMux I__15376 (
            .O(N__70729),
            .I(N__70725));
    CascadeMux I__15375 (
            .O(N__70728),
            .I(N__70722));
    InMux I__15374 (
            .O(N__70725),
            .I(N__70708));
    InMux I__15373 (
            .O(N__70722),
            .I(N__70708));
    InMux I__15372 (
            .O(N__70721),
            .I(N__70702));
    CascadeMux I__15371 (
            .O(N__70720),
            .I(N__70699));
    InMux I__15370 (
            .O(N__70719),
            .I(N__70696));
    InMux I__15369 (
            .O(N__70718),
            .I(N__70693));
    CascadeMux I__15368 (
            .O(N__70717),
            .I(N__70689));
    InMux I__15367 (
            .O(N__70716),
            .I(N__70686));
    InMux I__15366 (
            .O(N__70715),
            .I(N__70683));
    CascadeMux I__15365 (
            .O(N__70714),
            .I(N__70677));
    InMux I__15364 (
            .O(N__70713),
            .I(N__70672));
    LocalMux I__15363 (
            .O(N__70708),
            .I(N__70669));
    InMux I__15362 (
            .O(N__70707),
            .I(N__70664));
    InMux I__15361 (
            .O(N__70706),
            .I(N__70664));
    InMux I__15360 (
            .O(N__70705),
            .I(N__70658));
    LocalMux I__15359 (
            .O(N__70702),
            .I(N__70655));
    InMux I__15358 (
            .O(N__70699),
            .I(N__70652));
    LocalMux I__15357 (
            .O(N__70696),
            .I(N__70649));
    LocalMux I__15356 (
            .O(N__70693),
            .I(N__70646));
    CascadeMux I__15355 (
            .O(N__70692),
            .I(N__70643));
    InMux I__15354 (
            .O(N__70689),
            .I(N__70640));
    LocalMux I__15353 (
            .O(N__70686),
            .I(N__70637));
    LocalMux I__15352 (
            .O(N__70683),
            .I(N__70634));
    InMux I__15351 (
            .O(N__70682),
            .I(N__70626));
    InMux I__15350 (
            .O(N__70681),
            .I(N__70626));
    InMux I__15349 (
            .O(N__70680),
            .I(N__70623));
    InMux I__15348 (
            .O(N__70677),
            .I(N__70620));
    InMux I__15347 (
            .O(N__70676),
            .I(N__70615));
    InMux I__15346 (
            .O(N__70675),
            .I(N__70615));
    LocalMux I__15345 (
            .O(N__70672),
            .I(N__70608));
    Span4Mux_v I__15344 (
            .O(N__70669),
            .I(N__70608));
    LocalMux I__15343 (
            .O(N__70664),
            .I(N__70608));
    InMux I__15342 (
            .O(N__70663),
            .I(N__70605));
    InMux I__15341 (
            .O(N__70662),
            .I(N__70602));
    InMux I__15340 (
            .O(N__70661),
            .I(N__70599));
    LocalMux I__15339 (
            .O(N__70658),
            .I(N__70596));
    Span4Mux_v I__15338 (
            .O(N__70655),
            .I(N__70591));
    LocalMux I__15337 (
            .O(N__70652),
            .I(N__70591));
    Span4Mux_h I__15336 (
            .O(N__70649),
            .I(N__70586));
    Span4Mux_h I__15335 (
            .O(N__70646),
            .I(N__70586));
    InMux I__15334 (
            .O(N__70643),
            .I(N__70582));
    LocalMux I__15333 (
            .O(N__70640),
            .I(N__70579));
    Span4Mux_v I__15332 (
            .O(N__70637),
            .I(N__70576));
    Span4Mux_h I__15331 (
            .O(N__70634),
            .I(N__70573));
    CascadeMux I__15330 (
            .O(N__70633),
            .I(N__70566));
    InMux I__15329 (
            .O(N__70632),
            .I(N__70560));
    InMux I__15328 (
            .O(N__70631),
            .I(N__70560));
    LocalMux I__15327 (
            .O(N__70626),
            .I(N__70557));
    LocalMux I__15326 (
            .O(N__70623),
            .I(N__70552));
    LocalMux I__15325 (
            .O(N__70620),
            .I(N__70552));
    LocalMux I__15324 (
            .O(N__70615),
            .I(N__70549));
    Span4Mux_v I__15323 (
            .O(N__70608),
            .I(N__70546));
    LocalMux I__15322 (
            .O(N__70605),
            .I(N__70543));
    LocalMux I__15321 (
            .O(N__70602),
            .I(N__70540));
    LocalMux I__15320 (
            .O(N__70599),
            .I(N__70531));
    Span4Mux_h I__15319 (
            .O(N__70596),
            .I(N__70531));
    Span4Mux_h I__15318 (
            .O(N__70591),
            .I(N__70531));
    Span4Mux_v I__15317 (
            .O(N__70586),
            .I(N__70531));
    InMux I__15316 (
            .O(N__70585),
            .I(N__70528));
    LocalMux I__15315 (
            .O(N__70582),
            .I(N__70523));
    Span4Mux_h I__15314 (
            .O(N__70579),
            .I(N__70523));
    Span4Mux_h I__15313 (
            .O(N__70576),
            .I(N__70518));
    Span4Mux_h I__15312 (
            .O(N__70573),
            .I(N__70518));
    InMux I__15311 (
            .O(N__70572),
            .I(N__70513));
    InMux I__15310 (
            .O(N__70571),
            .I(N__70513));
    InMux I__15309 (
            .O(N__70570),
            .I(N__70508));
    InMux I__15308 (
            .O(N__70569),
            .I(N__70508));
    InMux I__15307 (
            .O(N__70566),
            .I(N__70505));
    InMux I__15306 (
            .O(N__70565),
            .I(N__70502));
    LocalMux I__15305 (
            .O(N__70560),
            .I(N__70497));
    Span12Mux_h I__15304 (
            .O(N__70557),
            .I(N__70497));
    Span4Mux_h I__15303 (
            .O(N__70552),
            .I(N__70490));
    Span4Mux_h I__15302 (
            .O(N__70549),
            .I(N__70490));
    Span4Mux_h I__15301 (
            .O(N__70546),
            .I(N__70490));
    Span4Mux_h I__15300 (
            .O(N__70543),
            .I(N__70483));
    Span4Mux_h I__15299 (
            .O(N__70540),
            .I(N__70483));
    Span4Mux_h I__15298 (
            .O(N__70531),
            .I(N__70483));
    LocalMux I__15297 (
            .O(N__70528),
            .I(N__70476));
    Span4Mux_h I__15296 (
            .O(N__70523),
            .I(N__70476));
    Span4Mux_h I__15295 (
            .O(N__70518),
            .I(N__70476));
    LocalMux I__15294 (
            .O(N__70513),
            .I(N__70473));
    LocalMux I__15293 (
            .O(N__70508),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n61_adj_1154 ));
    LocalMux I__15292 (
            .O(N__70505),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n61_adj_1154 ));
    LocalMux I__15291 (
            .O(N__70502),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n61_adj_1154 ));
    Odrv12 I__15290 (
            .O(N__70497),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n61_adj_1154 ));
    Odrv4 I__15289 (
            .O(N__70490),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n61_adj_1154 ));
    Odrv4 I__15288 (
            .O(N__70483),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n61_adj_1154 ));
    Odrv4 I__15287 (
            .O(N__70476),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n61_adj_1154 ));
    Odrv12 I__15286 (
            .O(N__70473),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n61_adj_1154 ));
    InMux I__15285 (
            .O(N__70456),
            .I(N__70452));
    CascadeMux I__15284 (
            .O(N__70455),
            .I(N__70449));
    LocalMux I__15283 (
            .O(N__70452),
            .I(N__70446));
    InMux I__15282 (
            .O(N__70449),
            .I(N__70443));
    Odrv4 I__15281 (
            .O(N__70446),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_6 ));
    LocalMux I__15280 (
            .O(N__70443),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_6 ));
    CascadeMux I__15279 (
            .O(N__70438),
            .I(N__70435));
    InMux I__15278 (
            .O(N__70435),
            .I(N__70429));
    InMux I__15277 (
            .O(N__70434),
            .I(N__70429));
    LocalMux I__15276 (
            .O(N__70429),
            .I(REG_mem_31_6));
    CascadeMux I__15275 (
            .O(N__70426),
            .I(N__70423));
    InMux I__15274 (
            .O(N__70423),
            .I(N__70417));
    InMux I__15273 (
            .O(N__70422),
            .I(N__70417));
    LocalMux I__15272 (
            .O(N__70417),
            .I(REG_mem_26_6));
    InMux I__15271 (
            .O(N__70414),
            .I(N__70411));
    LocalMux I__15270 (
            .O(N__70411),
            .I(N__70408));
    Span4Mux_h I__15269 (
            .O(N__70408),
            .I(N__70405));
    Span4Mux_v I__15268 (
            .O(N__70405),
            .I(N__70401));
    InMux I__15267 (
            .O(N__70404),
            .I(N__70398));
    Odrv4 I__15266 (
            .O(N__70401),
            .I(REG_mem_31_4));
    LocalMux I__15265 (
            .O(N__70398),
            .I(REG_mem_31_4));
    InMux I__15264 (
            .O(N__70393),
            .I(N__70388));
    InMux I__15263 (
            .O(N__70392),
            .I(N__70380));
    InMux I__15262 (
            .O(N__70391),
            .I(N__70375));
    LocalMux I__15261 (
            .O(N__70388),
            .I(N__70370));
    InMux I__15260 (
            .O(N__70387),
            .I(N__70367));
    InMux I__15259 (
            .O(N__70386),
            .I(N__70364));
    InMux I__15258 (
            .O(N__70385),
            .I(N__70361));
    InMux I__15257 (
            .O(N__70384),
            .I(N__70358));
    InMux I__15256 (
            .O(N__70383),
            .I(N__70355));
    LocalMux I__15255 (
            .O(N__70380),
            .I(N__70352));
    InMux I__15254 (
            .O(N__70379),
            .I(N__70349));
    InMux I__15253 (
            .O(N__70378),
            .I(N__70346));
    LocalMux I__15252 (
            .O(N__70375),
            .I(N__70343));
    InMux I__15251 (
            .O(N__70374),
            .I(N__70340));
    InMux I__15250 (
            .O(N__70373),
            .I(N__70337));
    Span4Mux_v I__15249 (
            .O(N__70370),
            .I(N__70333));
    LocalMux I__15248 (
            .O(N__70367),
            .I(N__70330));
    LocalMux I__15247 (
            .O(N__70364),
            .I(N__70327));
    LocalMux I__15246 (
            .O(N__70361),
            .I(N__70324));
    LocalMux I__15245 (
            .O(N__70358),
            .I(N__70321));
    LocalMux I__15244 (
            .O(N__70355),
            .I(N__70318));
    Span4Mux_v I__15243 (
            .O(N__70352),
            .I(N__70314));
    LocalMux I__15242 (
            .O(N__70349),
            .I(N__70311));
    LocalMux I__15241 (
            .O(N__70346),
            .I(N__70308));
    Span4Mux_v I__15240 (
            .O(N__70343),
            .I(N__70305));
    LocalMux I__15239 (
            .O(N__70340),
            .I(N__70302));
    LocalMux I__15238 (
            .O(N__70337),
            .I(N__70299));
    InMux I__15237 (
            .O(N__70336),
            .I(N__70296));
    Span4Mux_h I__15236 (
            .O(N__70333),
            .I(N__70289));
    Span4Mux_v I__15235 (
            .O(N__70330),
            .I(N__70289));
    Span4Mux_h I__15234 (
            .O(N__70327),
            .I(N__70286));
    Span4Mux_v I__15233 (
            .O(N__70324),
            .I(N__70283));
    Span4Mux_v I__15232 (
            .O(N__70321),
            .I(N__70280));
    Span4Mux_v I__15231 (
            .O(N__70318),
            .I(N__70277));
    InMux I__15230 (
            .O(N__70317),
            .I(N__70274));
    Span4Mux_v I__15229 (
            .O(N__70314),
            .I(N__70271));
    Span4Mux_v I__15228 (
            .O(N__70311),
            .I(N__70268));
    Span4Mux_v I__15227 (
            .O(N__70308),
            .I(N__70265));
    Span4Mux_v I__15226 (
            .O(N__70305),
            .I(N__70262));
    Span4Mux_v I__15225 (
            .O(N__70302),
            .I(N__70257));
    Span4Mux_h I__15224 (
            .O(N__70299),
            .I(N__70257));
    LocalMux I__15223 (
            .O(N__70296),
            .I(N__70254));
    InMux I__15222 (
            .O(N__70295),
            .I(N__70251));
    InMux I__15221 (
            .O(N__70294),
            .I(N__70248));
    Span4Mux_h I__15220 (
            .O(N__70289),
            .I(N__70245));
    Span4Mux_v I__15219 (
            .O(N__70286),
            .I(N__70240));
    Span4Mux_h I__15218 (
            .O(N__70283),
            .I(N__70240));
    Span4Mux_v I__15217 (
            .O(N__70280),
            .I(N__70235));
    Span4Mux_h I__15216 (
            .O(N__70277),
            .I(N__70235));
    LocalMux I__15215 (
            .O(N__70274),
            .I(N__70232));
    Span4Mux_h I__15214 (
            .O(N__70271),
            .I(N__70225));
    Span4Mux_v I__15213 (
            .O(N__70268),
            .I(N__70225));
    Span4Mux_h I__15212 (
            .O(N__70265),
            .I(N__70225));
    Span4Mux_h I__15211 (
            .O(N__70262),
            .I(N__70220));
    Span4Mux_h I__15210 (
            .O(N__70257),
            .I(N__70220));
    Span12Mux_h I__15209 (
            .O(N__70254),
            .I(N__70213));
    LocalMux I__15208 (
            .O(N__70251),
            .I(N__70213));
    LocalMux I__15207 (
            .O(N__70248),
            .I(N__70213));
    Odrv4 I__15206 (
            .O(N__70245),
            .I(n39));
    Odrv4 I__15205 (
            .O(N__70240),
            .I(n39));
    Odrv4 I__15204 (
            .O(N__70235),
            .I(n39));
    Odrv12 I__15203 (
            .O(N__70232),
            .I(n39));
    Odrv4 I__15202 (
            .O(N__70225),
            .I(n39));
    Odrv4 I__15201 (
            .O(N__70220),
            .I(n39));
    Odrv12 I__15200 (
            .O(N__70213),
            .I(n39));
    CascadeMux I__15199 (
            .O(N__70198),
            .I(N__70195));
    InMux I__15198 (
            .O(N__70195),
            .I(N__70191));
    InMux I__15197 (
            .O(N__70194),
            .I(N__70188));
    LocalMux I__15196 (
            .O(N__70191),
            .I(REG_mem_26_8));
    LocalMux I__15195 (
            .O(N__70188),
            .I(REG_mem_26_8));
    InMux I__15194 (
            .O(N__70183),
            .I(N__70180));
    LocalMux I__15193 (
            .O(N__70180),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13778 ));
    CascadeMux I__15192 (
            .O(N__70177),
            .I(N__70174));
    InMux I__15191 (
            .O(N__70174),
            .I(N__70171));
    LocalMux I__15190 (
            .O(N__70171),
            .I(N__70168));
    Span4Mux_v I__15189 (
            .O(N__70168),
            .I(N__70165));
    Span4Mux_h I__15188 (
            .O(N__70165),
            .I(N__70161));
    InMux I__15187 (
            .O(N__70164),
            .I(N__70158));
    Odrv4 I__15186 (
            .O(N__70161),
            .I(REG_mem_8_6));
    LocalMux I__15185 (
            .O(N__70158),
            .I(REG_mem_8_6));
    InMux I__15184 (
            .O(N__70153),
            .I(N__70149));
    InMux I__15183 (
            .O(N__70152),
            .I(N__70146));
    LocalMux I__15182 (
            .O(N__70149),
            .I(REG_mem_9_6));
    LocalMux I__15181 (
            .O(N__70146),
            .I(REG_mem_9_6));
    InMux I__15180 (
            .O(N__70141),
            .I(N__70134));
    InMux I__15179 (
            .O(N__70140),
            .I(N__70129));
    InMux I__15178 (
            .O(N__70139),
            .I(N__70126));
    InMux I__15177 (
            .O(N__70138),
            .I(N__70123));
    CascadeMux I__15176 (
            .O(N__70137),
            .I(N__70117));
    LocalMux I__15175 (
            .O(N__70134),
            .I(N__70114));
    InMux I__15174 (
            .O(N__70133),
            .I(N__70110));
    InMux I__15173 (
            .O(N__70132),
            .I(N__70106));
    LocalMux I__15172 (
            .O(N__70129),
            .I(N__70103));
    LocalMux I__15171 (
            .O(N__70126),
            .I(N__70097));
    LocalMux I__15170 (
            .O(N__70123),
            .I(N__70094));
    InMux I__15169 (
            .O(N__70122),
            .I(N__70091));
    InMux I__15168 (
            .O(N__70121),
            .I(N__70086));
    InMux I__15167 (
            .O(N__70120),
            .I(N__70086));
    InMux I__15166 (
            .O(N__70117),
            .I(N__70083));
    Span4Mux_v I__15165 (
            .O(N__70114),
            .I(N__70080));
    InMux I__15164 (
            .O(N__70113),
            .I(N__70076));
    LocalMux I__15163 (
            .O(N__70110),
            .I(N__70073));
    InMux I__15162 (
            .O(N__70109),
            .I(N__70070));
    LocalMux I__15161 (
            .O(N__70106),
            .I(N__70067));
    Span4Mux_h I__15160 (
            .O(N__70103),
            .I(N__70064));
    InMux I__15159 (
            .O(N__70102),
            .I(N__70061));
    InMux I__15158 (
            .O(N__70101),
            .I(N__70058));
    InMux I__15157 (
            .O(N__70100),
            .I(N__70055));
    Span4Mux_h I__15156 (
            .O(N__70097),
            .I(N__70052));
    Span4Mux_h I__15155 (
            .O(N__70094),
            .I(N__70049));
    LocalMux I__15154 (
            .O(N__70091),
            .I(N__70044));
    LocalMux I__15153 (
            .O(N__70086),
            .I(N__70044));
    LocalMux I__15152 (
            .O(N__70083),
            .I(N__70039));
    Span4Mux_h I__15151 (
            .O(N__70080),
            .I(N__70039));
    InMux I__15150 (
            .O(N__70079),
            .I(N__70036));
    LocalMux I__15149 (
            .O(N__70076),
            .I(N__70033));
    Span4Mux_h I__15148 (
            .O(N__70073),
            .I(N__70030));
    LocalMux I__15147 (
            .O(N__70070),
            .I(N__70025));
    Span4Mux_v I__15146 (
            .O(N__70067),
            .I(N__70025));
    Span4Mux_h I__15145 (
            .O(N__70064),
            .I(N__70022));
    LocalMux I__15144 (
            .O(N__70061),
            .I(N__70013));
    LocalMux I__15143 (
            .O(N__70058),
            .I(N__70013));
    LocalMux I__15142 (
            .O(N__70055),
            .I(N__70013));
    Sp12to4 I__15141 (
            .O(N__70052),
            .I(N__70013));
    Span4Mux_h I__15140 (
            .O(N__70049),
            .I(N__70006));
    Span4Mux_h I__15139 (
            .O(N__70044),
            .I(N__70006));
    Span4Mux_h I__15138 (
            .O(N__70039),
            .I(N__70006));
    LocalMux I__15137 (
            .O(N__70036),
            .I(n52));
    Odrv12 I__15136 (
            .O(N__70033),
            .I(n52));
    Odrv4 I__15135 (
            .O(N__70030),
            .I(n52));
    Odrv4 I__15134 (
            .O(N__70025),
            .I(n52));
    Odrv4 I__15133 (
            .O(N__70022),
            .I(n52));
    Odrv12 I__15132 (
            .O(N__70013),
            .I(n52));
    Odrv4 I__15131 (
            .O(N__70006),
            .I(n52));
    InMux I__15130 (
            .O(N__69991),
            .I(N__69988));
    LocalMux I__15129 (
            .O(N__69988),
            .I(N__69985));
    Sp12to4 I__15128 (
            .O(N__69985),
            .I(N__69982));
    Span12Mux_v I__15127 (
            .O(N__69982),
            .I(N__69978));
    CascadeMux I__15126 (
            .O(N__69981),
            .I(N__69975));
    Span12Mux_h I__15125 (
            .O(N__69978),
            .I(N__69972));
    InMux I__15124 (
            .O(N__69975),
            .I(N__69969));
    Odrv12 I__15123 (
            .O(N__69972),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_0 ));
    LocalMux I__15122 (
            .O(N__69969),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_0 ));
    CascadeMux I__15121 (
            .O(N__69964),
            .I(rd_addr_p1_w_2_cascade_));
    IoInMux I__15120 (
            .O(N__69961),
            .I(N__69958));
    LocalMux I__15119 (
            .O(N__69958),
            .I(N__69955));
    IoSpan4Mux I__15118 (
            .O(N__69955),
            .I(N__69952));
    Sp12to4 I__15117 (
            .O(N__69952),
            .I(N__69948));
    InMux I__15116 (
            .O(N__69951),
            .I(N__69945));
    Span12Mux_v I__15115 (
            .O(N__69948),
            .I(N__69942));
    LocalMux I__15114 (
            .O(N__69945),
            .I(N__69939));
    Span12Mux_h I__15113 (
            .O(N__69942),
            .I(N__69935));
    Span4Mux_v I__15112 (
            .O(N__69939),
            .I(N__69932));
    InMux I__15111 (
            .O(N__69938),
            .I(N__69929));
    Odrv12 I__15110 (
            .O(N__69935),
            .I(RESET_c));
    Odrv4 I__15109 (
            .O(N__69932),
            .I(RESET_c));
    LocalMux I__15108 (
            .O(N__69929),
            .I(RESET_c));
    CascadeMux I__15107 (
            .O(N__69922),
            .I(\tx_fifo.lscc_fifo_inst.wr_addr_p1_w_1_cascade_ ));
    CascadeMux I__15106 (
            .O(N__69919),
            .I(N__69915));
    InMux I__15105 (
            .O(N__69918),
            .I(N__69912));
    InMux I__15104 (
            .O(N__69915),
            .I(N__69909));
    LocalMux I__15103 (
            .O(N__69912),
            .I(N__69906));
    LocalMux I__15102 (
            .O(N__69909),
            .I(N__69903));
    Odrv4 I__15101 (
            .O(N__69906),
            .I(n1));
    Odrv4 I__15100 (
            .O(N__69903),
            .I(n1));
    InMux I__15099 (
            .O(N__69898),
            .I(N__69895));
    LocalMux I__15098 (
            .O(N__69895),
            .I(n10727));
    InMux I__15097 (
            .O(N__69892),
            .I(N__69884));
    InMux I__15096 (
            .O(N__69891),
            .I(N__69884));
    InMux I__15095 (
            .O(N__69890),
            .I(N__69879));
    InMux I__15094 (
            .O(N__69889),
            .I(N__69879));
    LocalMux I__15093 (
            .O(N__69884),
            .I(wr_addr_r_2));
    LocalMux I__15092 (
            .O(N__69879),
            .I(wr_addr_r_2));
    InMux I__15091 (
            .O(N__69874),
            .I(N__69865));
    InMux I__15090 (
            .O(N__69873),
            .I(N__69865));
    InMux I__15089 (
            .O(N__69872),
            .I(N__69865));
    LocalMux I__15088 (
            .O(N__69865),
            .I(rd_addr_r_2));
    InMux I__15087 (
            .O(N__69862),
            .I(N__69859));
    LocalMux I__15086 (
            .O(N__69859),
            .I(\tx_fifo.lscc_fifo_inst.n3 ));
    CascadeMux I__15085 (
            .O(N__69856),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13598_cascade_ ));
    InMux I__15084 (
            .O(N__69853),
            .I(N__69850));
    LocalMux I__15083 (
            .O(N__69850),
            .I(N__69847));
    Span4Mux_v I__15082 (
            .O(N__69847),
            .I(N__69843));
    CascadeMux I__15081 (
            .O(N__69846),
            .I(N__69840));
    Span4Mux_h I__15080 (
            .O(N__69843),
            .I(N__69837));
    InMux I__15079 (
            .O(N__69840),
            .I(N__69834));
    Odrv4 I__15078 (
            .O(N__69837),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_6 ));
    LocalMux I__15077 (
            .O(N__69834),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_6 ));
    InMux I__15076 (
            .O(N__69829),
            .I(N__69826));
    LocalMux I__15075 (
            .O(N__69826),
            .I(N__69823));
    Span4Mux_v I__15074 (
            .O(N__69823),
            .I(N__69819));
    InMux I__15073 (
            .O(N__69822),
            .I(N__69816));
    Odrv4 I__15072 (
            .O(N__69819),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_6 ));
    LocalMux I__15071 (
            .O(N__69816),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_6 ));
    InMux I__15070 (
            .O(N__69811),
            .I(N__69808));
    LocalMux I__15069 (
            .O(N__69808),
            .I(N__69804));
    InMux I__15068 (
            .O(N__69807),
            .I(N__69801));
    Odrv12 I__15067 (
            .O(N__69804),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_6 ));
    LocalMux I__15066 (
            .O(N__69801),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_6 ));
    CascadeMux I__15065 (
            .O(N__69796),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13634_cascade_ ));
    CascadeMux I__15064 (
            .O(N__69793),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13637_cascade_ ));
    InMux I__15063 (
            .O(N__69790),
            .I(N__69787));
    LocalMux I__15062 (
            .O(N__69787),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13601 ));
    CascadeMux I__15061 (
            .O(N__69784),
            .I(n15_cascade_));
    InMux I__15060 (
            .O(N__69781),
            .I(N__69778));
    LocalMux I__15059 (
            .O(N__69778),
            .I(full_nxt_r));
    InMux I__15058 (
            .O(N__69775),
            .I(N__69769));
    InMux I__15057 (
            .O(N__69774),
            .I(N__69766));
    InMux I__15056 (
            .O(N__69773),
            .I(N__69763));
    CascadeMux I__15055 (
            .O(N__69772),
            .I(N__69760));
    LocalMux I__15054 (
            .O(N__69769),
            .I(N__69753));
    LocalMux I__15053 (
            .O(N__69766),
            .I(N__69753));
    LocalMux I__15052 (
            .O(N__69763),
            .I(N__69753));
    InMux I__15051 (
            .O(N__69760),
            .I(N__69750));
    Span4Mux_v I__15050 (
            .O(N__69753),
            .I(N__69744));
    LocalMux I__15049 (
            .O(N__69750),
            .I(N__69744));
    InMux I__15048 (
            .O(N__69749),
            .I(N__69741));
    Odrv4 I__15047 (
            .O(N__69744),
            .I(rx_buf_byte_4));
    LocalMux I__15046 (
            .O(N__69741),
            .I(rx_buf_byte_4));
    InMux I__15045 (
            .O(N__69736),
            .I(N__69732));
    CascadeMux I__15044 (
            .O(N__69735),
            .I(N__69729));
    LocalMux I__15043 (
            .O(N__69732),
            .I(N__69726));
    InMux I__15042 (
            .O(N__69729),
            .I(N__69723));
    Odrv12 I__15041 (
            .O(N__69726),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4 ));
    LocalMux I__15040 (
            .O(N__69723),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4 ));
    InMux I__15039 (
            .O(N__69718),
            .I(N__69715));
    LocalMux I__15038 (
            .O(N__69715),
            .I(N__69712));
    Span4Mux_h I__15037 (
            .O(N__69712),
            .I(N__69709));
    Odrv4 I__15036 (
            .O(N__69709),
            .I(spi_rx_byte_ready));
    InMux I__15035 (
            .O(N__69706),
            .I(N__69696));
    InMux I__15034 (
            .O(N__69705),
            .I(N__69696));
    InMux I__15033 (
            .O(N__69704),
            .I(N__69687));
    InMux I__15032 (
            .O(N__69703),
            .I(N__69687));
    InMux I__15031 (
            .O(N__69702),
            .I(N__69687));
    InMux I__15030 (
            .O(N__69701),
            .I(N__69687));
    LocalMux I__15029 (
            .O(N__69696),
            .I(is_tx_fifo_full_flag));
    LocalMux I__15028 (
            .O(N__69687),
            .I(is_tx_fifo_full_flag));
    InMux I__15027 (
            .O(N__69682),
            .I(N__69679));
    LocalMux I__15026 (
            .O(N__69679),
            .I(rd_addr_p1_w_1));
    CascadeMux I__15025 (
            .O(N__69676),
            .I(N__69673));
    InMux I__15024 (
            .O(N__69673),
            .I(N__69670));
    LocalMux I__15023 (
            .O(N__69670),
            .I(rd_addr_p1_w_2));
    InMux I__15022 (
            .O(N__69667),
            .I(N__69664));
    LocalMux I__15021 (
            .O(N__69664),
            .I(N__69660));
    InMux I__15020 (
            .O(N__69663),
            .I(N__69657));
    Odrv4 I__15019 (
            .O(N__69660),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5 ));
    LocalMux I__15018 (
            .O(N__69657),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5 ));
    InMux I__15017 (
            .O(N__69652),
            .I(N__69649));
    LocalMux I__15016 (
            .O(N__69649),
            .I(N__69645));
    InMux I__15015 (
            .O(N__69648),
            .I(N__69642));
    Odrv4 I__15014 (
            .O(N__69645),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_4 ));
    LocalMux I__15013 (
            .O(N__69642),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_4 ));
    CascadeMux I__15012 (
            .O(N__69637),
            .I(\tx_fifo.lscc_fifo_inst.n3_adj_1136_cascade_ ));
    CascadeMux I__15011 (
            .O(N__69634),
            .I(\tx_fifo.lscc_fifo_inst.n4_cascade_ ));
    InMux I__15010 (
            .O(N__69631),
            .I(N__69625));
    InMux I__15009 (
            .O(N__69630),
            .I(N__69625));
    LocalMux I__15008 (
            .O(N__69625),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0 ));
    InMux I__15007 (
            .O(N__69622),
            .I(N__69606));
    InMux I__15006 (
            .O(N__69621),
            .I(N__69606));
    CascadeMux I__15005 (
            .O(N__69620),
            .I(N__69601));
    InMux I__15004 (
            .O(N__69619),
            .I(N__69586));
    InMux I__15003 (
            .O(N__69618),
            .I(N__69586));
    InMux I__15002 (
            .O(N__69617),
            .I(N__69586));
    InMux I__15001 (
            .O(N__69616),
            .I(N__69586));
    InMux I__15000 (
            .O(N__69615),
            .I(N__69586));
    InMux I__14999 (
            .O(N__69614),
            .I(N__69586));
    InMux I__14998 (
            .O(N__69613),
            .I(N__69586));
    CascadeMux I__14997 (
            .O(N__69612),
            .I(N__69582));
    CascadeMux I__14996 (
            .O(N__69611),
            .I(N__69579));
    LocalMux I__14995 (
            .O(N__69606),
            .I(N__69576));
    InMux I__14994 (
            .O(N__69605),
            .I(N__69569));
    InMux I__14993 (
            .O(N__69604),
            .I(N__69569));
    InMux I__14992 (
            .O(N__69601),
            .I(N__69569));
    LocalMux I__14991 (
            .O(N__69586),
            .I(N__69566));
    InMux I__14990 (
            .O(N__69585),
            .I(N__69563));
    InMux I__14989 (
            .O(N__69582),
            .I(N__69558));
    InMux I__14988 (
            .O(N__69579),
            .I(N__69558));
    Odrv4 I__14987 (
            .O(N__69576),
            .I(\tx_fifo.lscc_fifo_inst.n3_adj_1136 ));
    LocalMux I__14986 (
            .O(N__69569),
            .I(\tx_fifo.lscc_fifo_inst.n3_adj_1136 ));
    Odrv4 I__14985 (
            .O(N__69566),
            .I(\tx_fifo.lscc_fifo_inst.n3_adj_1136 ));
    LocalMux I__14984 (
            .O(N__69563),
            .I(\tx_fifo.lscc_fifo_inst.n3_adj_1136 ));
    LocalMux I__14983 (
            .O(N__69558),
            .I(\tx_fifo.lscc_fifo_inst.n3_adj_1136 ));
    InMux I__14982 (
            .O(N__69547),
            .I(N__69540));
    InMux I__14981 (
            .O(N__69546),
            .I(N__69533));
    InMux I__14980 (
            .O(N__69545),
            .I(N__69533));
    InMux I__14979 (
            .O(N__69544),
            .I(N__69533));
    InMux I__14978 (
            .O(N__69543),
            .I(N__69530));
    LocalMux I__14977 (
            .O(N__69540),
            .I(rx_buf_byte_0));
    LocalMux I__14976 (
            .O(N__69533),
            .I(rx_buf_byte_0));
    LocalMux I__14975 (
            .O(N__69530),
            .I(rx_buf_byte_0));
    InMux I__14974 (
            .O(N__69523),
            .I(N__69517));
    InMux I__14973 (
            .O(N__69522),
            .I(N__69517));
    LocalMux I__14972 (
            .O(N__69517),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_0 ));
    CascadeMux I__14971 (
            .O(N__69514),
            .I(n11424_cascade_));
    InMux I__14970 (
            .O(N__69511),
            .I(N__69507));
    InMux I__14969 (
            .O(N__69510),
            .I(N__69504));
    LocalMux I__14968 (
            .O(N__69507),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2 ));
    LocalMux I__14967 (
            .O(N__69504),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2 ));
    InMux I__14966 (
            .O(N__69499),
            .I(N__69495));
    InMux I__14965 (
            .O(N__69498),
            .I(N__69492));
    LocalMux I__14964 (
            .O(N__69495),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_4 ));
    LocalMux I__14963 (
            .O(N__69492),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_4 ));
    InMux I__14962 (
            .O(N__69487),
            .I(N__69483));
    CascadeMux I__14961 (
            .O(N__69486),
            .I(N__69480));
    LocalMux I__14960 (
            .O(N__69483),
            .I(N__69477));
    InMux I__14959 (
            .O(N__69480),
            .I(N__69474));
    Odrv4 I__14958 (
            .O(N__69477),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4 ));
    LocalMux I__14957 (
            .O(N__69474),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4 ));
    InMux I__14956 (
            .O(N__69469),
            .I(N__69462));
    InMux I__14955 (
            .O(N__69468),
            .I(N__69453));
    InMux I__14954 (
            .O(N__69467),
            .I(N__69453));
    InMux I__14953 (
            .O(N__69466),
            .I(N__69453));
    InMux I__14952 (
            .O(N__69465),
            .I(N__69453));
    LocalMux I__14951 (
            .O(N__69462),
            .I(rx_buf_byte_7));
    LocalMux I__14950 (
            .O(N__69453),
            .I(rx_buf_byte_7));
    InMux I__14949 (
            .O(N__69448),
            .I(N__69445));
    LocalMux I__14948 (
            .O(N__69445),
            .I(N__69440));
    InMux I__14947 (
            .O(N__69444),
            .I(N__69437));
    InMux I__14946 (
            .O(N__69443),
            .I(N__69434));
    Span4Mux_v I__14945 (
            .O(N__69440),
            .I(N__69430));
    LocalMux I__14944 (
            .O(N__69437),
            .I(N__69427));
    LocalMux I__14943 (
            .O(N__69434),
            .I(N__69424));
    InMux I__14942 (
            .O(N__69433),
            .I(N__69421));
    Odrv4 I__14941 (
            .O(N__69430),
            .I(tx_data_byte_4));
    Odrv4 I__14940 (
            .O(N__69427),
            .I(tx_data_byte_4));
    Odrv4 I__14939 (
            .O(N__69424),
            .I(tx_data_byte_4));
    LocalMux I__14938 (
            .O(N__69421),
            .I(tx_data_byte_4));
    InMux I__14937 (
            .O(N__69412),
            .I(N__69409));
    LocalMux I__14936 (
            .O(N__69409),
            .I(N__69397));
    InMux I__14935 (
            .O(N__69408),
            .I(N__69386));
    InMux I__14934 (
            .O(N__69407),
            .I(N__69386));
    InMux I__14933 (
            .O(N__69406),
            .I(N__69386));
    InMux I__14932 (
            .O(N__69405),
            .I(N__69386));
    InMux I__14931 (
            .O(N__69404),
            .I(N__69386));
    InMux I__14930 (
            .O(N__69403),
            .I(N__69383));
    InMux I__14929 (
            .O(N__69402),
            .I(N__69380));
    InMux I__14928 (
            .O(N__69401),
            .I(N__69370));
    InMux I__14927 (
            .O(N__69400),
            .I(N__69370));
    Span4Mux_v I__14926 (
            .O(N__69397),
            .I(N__69363));
    LocalMux I__14925 (
            .O(N__69386),
            .I(N__69356));
    LocalMux I__14924 (
            .O(N__69383),
            .I(N__69356));
    LocalMux I__14923 (
            .O(N__69380),
            .I(N__69356));
    InMux I__14922 (
            .O(N__69379),
            .I(N__69353));
    InMux I__14921 (
            .O(N__69378),
            .I(N__69344));
    InMux I__14920 (
            .O(N__69377),
            .I(N__69344));
    InMux I__14919 (
            .O(N__69376),
            .I(N__69344));
    InMux I__14918 (
            .O(N__69375),
            .I(N__69344));
    LocalMux I__14917 (
            .O(N__69370),
            .I(N__69341));
    InMux I__14916 (
            .O(N__69369),
            .I(N__69332));
    InMux I__14915 (
            .O(N__69368),
            .I(N__69332));
    InMux I__14914 (
            .O(N__69367),
            .I(N__69332));
    InMux I__14913 (
            .O(N__69366),
            .I(N__69332));
    Odrv4 I__14912 (
            .O(N__69363),
            .I(uart_rx_complete_rising_edge));
    Odrv4 I__14911 (
            .O(N__69356),
            .I(uart_rx_complete_rising_edge));
    LocalMux I__14910 (
            .O(N__69353),
            .I(uart_rx_complete_rising_edge));
    LocalMux I__14909 (
            .O(N__69344),
            .I(uart_rx_complete_rising_edge));
    Odrv4 I__14908 (
            .O(N__69341),
            .I(uart_rx_complete_rising_edge));
    LocalMux I__14907 (
            .O(N__69332),
            .I(uart_rx_complete_rising_edge));
    InMux I__14906 (
            .O(N__69319),
            .I(N__69316));
    LocalMux I__14905 (
            .O(N__69316),
            .I(N__69313));
    Span4Mux_v I__14904 (
            .O(N__69313),
            .I(N__69309));
    InMux I__14903 (
            .O(N__69312),
            .I(N__69306));
    Odrv4 I__14902 (
            .O(N__69309),
            .I(tx_addr_byte_4));
    LocalMux I__14901 (
            .O(N__69306),
            .I(tx_addr_byte_4));
    InMux I__14900 (
            .O(N__69301),
            .I(N__69298));
    LocalMux I__14899 (
            .O(N__69298),
            .I(N__69294));
    InMux I__14898 (
            .O(N__69297),
            .I(N__69291));
    Odrv4 I__14897 (
            .O(N__69294),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_5 ));
    LocalMux I__14896 (
            .O(N__69291),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_5 ));
    InMux I__14895 (
            .O(N__69286),
            .I(N__69283));
    LocalMux I__14894 (
            .O(N__69283),
            .I(N__69279));
    InMux I__14893 (
            .O(N__69282),
            .I(N__69276));
    Odrv12 I__14892 (
            .O(N__69279),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5 ));
    LocalMux I__14891 (
            .O(N__69276),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5 ));
    CascadeMux I__14890 (
            .O(N__69271),
            .I(N__69266));
    CascadeMux I__14889 (
            .O(N__69270),
            .I(N__69262));
    CascadeMux I__14888 (
            .O(N__69269),
            .I(N__69259));
    InMux I__14887 (
            .O(N__69266),
            .I(N__69256));
    InMux I__14886 (
            .O(N__69265),
            .I(N__69248));
    InMux I__14885 (
            .O(N__69262),
            .I(N__69248));
    InMux I__14884 (
            .O(N__69259),
            .I(N__69248));
    LocalMux I__14883 (
            .O(N__69256),
            .I(N__69245));
    InMux I__14882 (
            .O(N__69255),
            .I(N__69242));
    LocalMux I__14881 (
            .O(N__69248),
            .I(rx_buf_byte_5));
    Odrv4 I__14880 (
            .O(N__69245),
            .I(rx_buf_byte_5));
    LocalMux I__14879 (
            .O(N__69242),
            .I(rx_buf_byte_5));
    CascadeMux I__14878 (
            .O(N__69235),
            .I(\tx_fifo.lscc_fifo_inst.n13694_cascade_ ));
    InMux I__14877 (
            .O(N__69232),
            .I(N__69229));
    LocalMux I__14876 (
            .O(N__69229),
            .I(N__69225));
    InMux I__14875 (
            .O(N__69228),
            .I(N__69222));
    Odrv4 I__14874 (
            .O(N__69225),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_5 ));
    LocalMux I__14873 (
            .O(N__69222),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_5 ));
    CascadeMux I__14872 (
            .O(N__69217),
            .I(\tx_fifo.lscc_fifo_inst.n13766_cascade_ ));
    CascadeMux I__14871 (
            .O(N__69214),
            .I(N__69210));
    InMux I__14870 (
            .O(N__69213),
            .I(N__69207));
    InMux I__14869 (
            .O(N__69210),
            .I(N__69204));
    LocalMux I__14868 (
            .O(N__69207),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_2 ));
    LocalMux I__14867 (
            .O(N__69204),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_2 ));
    InMux I__14866 (
            .O(N__69199),
            .I(N__69195));
    InMux I__14865 (
            .O(N__69198),
            .I(N__69192));
    LocalMux I__14864 (
            .O(N__69195),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_2 ));
    LocalMux I__14863 (
            .O(N__69192),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_2 ));
    SRMux I__14862 (
            .O(N__69187),
            .I(N__69184));
    LocalMux I__14861 (
            .O(N__69184),
            .I(N__69181));
    Span4Mux_h I__14860 (
            .O(N__69181),
            .I(N__69178));
    Odrv4 I__14859 (
            .O(N__69178),
            .I(\bluejay_data_inst.n7424 ));
    CEMux I__14858 (
            .O(N__69175),
            .I(N__69172));
    LocalMux I__14857 (
            .O(N__69172),
            .I(N__69165));
    CEMux I__14856 (
            .O(N__69171),
            .I(N__69162));
    CEMux I__14855 (
            .O(N__69170),
            .I(N__69159));
    CEMux I__14854 (
            .O(N__69169),
            .I(N__69156));
    CEMux I__14853 (
            .O(N__69168),
            .I(N__69149));
    Span4Mux_v I__14852 (
            .O(N__69165),
            .I(N__69146));
    LocalMux I__14851 (
            .O(N__69162),
            .I(N__69139));
    LocalMux I__14850 (
            .O(N__69159),
            .I(N__69139));
    LocalMux I__14849 (
            .O(N__69156),
            .I(N__69139));
    InMux I__14848 (
            .O(N__69155),
            .I(N__69136));
    InMux I__14847 (
            .O(N__69154),
            .I(N__69131));
    InMux I__14846 (
            .O(N__69153),
            .I(N__69131));
    CEMux I__14845 (
            .O(N__69152),
            .I(N__69128));
    LocalMux I__14844 (
            .O(N__69149),
            .I(N__69125));
    Span4Mux_h I__14843 (
            .O(N__69146),
            .I(N__69120));
    Span4Mux_v I__14842 (
            .O(N__69139),
            .I(N__69120));
    LocalMux I__14841 (
            .O(N__69136),
            .I(N__69113));
    LocalMux I__14840 (
            .O(N__69131),
            .I(N__69113));
    LocalMux I__14839 (
            .O(N__69128),
            .I(N__69113));
    Odrv4 I__14838 (
            .O(N__69125),
            .I(\bluejay_data_inst.n4062 ));
    Odrv4 I__14837 (
            .O(N__69120),
            .I(\bluejay_data_inst.n4062 ));
    Odrv12 I__14836 (
            .O(N__69113),
            .I(\bluejay_data_inst.n4062 ));
    IoInMux I__14835 (
            .O(N__69106),
            .I(N__69103));
    LocalMux I__14834 (
            .O(N__69103),
            .I(N__69100));
    Span4Mux_s3_h I__14833 (
            .O(N__69100),
            .I(N__69097));
    Span4Mux_h I__14832 (
            .O(N__69097),
            .I(N__69093));
    CascadeMux I__14831 (
            .O(N__69096),
            .I(N__69089));
    Span4Mux_h I__14830 (
            .O(N__69093),
            .I(N__69086));
    InMux I__14829 (
            .O(N__69092),
            .I(N__69083));
    InMux I__14828 (
            .O(N__69089),
            .I(N__69080));
    Odrv4 I__14827 (
            .O(N__69086),
            .I(\bluejay_data_inst.bluejay_data_out_31__N_701 ));
    LocalMux I__14826 (
            .O(N__69083),
            .I(\bluejay_data_inst.bluejay_data_out_31__N_701 ));
    LocalMux I__14825 (
            .O(N__69080),
            .I(\bluejay_data_inst.bluejay_data_out_31__N_701 ));
    SRMux I__14824 (
            .O(N__69073),
            .I(N__69070));
    LocalMux I__14823 (
            .O(N__69070),
            .I(N__69067));
    Span4Mux_h I__14822 (
            .O(N__69067),
            .I(N__69064));
    Odrv4 I__14821 (
            .O(N__69064),
            .I(\bluejay_data_inst.n4442 ));
    InMux I__14820 (
            .O(N__69061),
            .I(N__69056));
    InMux I__14819 (
            .O(N__69060),
            .I(N__69051));
    InMux I__14818 (
            .O(N__69059),
            .I(N__69051));
    LocalMux I__14817 (
            .O(N__69056),
            .I(\bluejay_data_inst.bluejay_data_out_31__N_702 ));
    LocalMux I__14816 (
            .O(N__69051),
            .I(\bluejay_data_inst.bluejay_data_out_31__N_702 ));
    InMux I__14815 (
            .O(N__69046),
            .I(N__69043));
    LocalMux I__14814 (
            .O(N__69043),
            .I(N__69040));
    Span4Mux_v I__14813 (
            .O(N__69040),
            .I(N__69033));
    InMux I__14812 (
            .O(N__69039),
            .I(N__69024));
    InMux I__14811 (
            .O(N__69038),
            .I(N__69024));
    InMux I__14810 (
            .O(N__69037),
            .I(N__69024));
    InMux I__14809 (
            .O(N__69036),
            .I(N__69024));
    Sp12to4 I__14808 (
            .O(N__69033),
            .I(N__69019));
    LocalMux I__14807 (
            .O(N__69024),
            .I(N__69019));
    Odrv12 I__14806 (
            .O(N__69019),
            .I(get_next_word));
    InMux I__14805 (
            .O(N__69016),
            .I(N__68992));
    InMux I__14804 (
            .O(N__69015),
            .I(N__68992));
    InMux I__14803 (
            .O(N__69014),
            .I(N__68992));
    InMux I__14802 (
            .O(N__69013),
            .I(N__68992));
    InMux I__14801 (
            .O(N__69012),
            .I(N__68992));
    InMux I__14800 (
            .O(N__69011),
            .I(N__68992));
    InMux I__14799 (
            .O(N__69010),
            .I(N__68992));
    InMux I__14798 (
            .O(N__69009),
            .I(N__68992));
    LocalMux I__14797 (
            .O(N__68992),
            .I(N__68982));
    InMux I__14796 (
            .O(N__68991),
            .I(N__68966));
    InMux I__14795 (
            .O(N__68990),
            .I(N__68966));
    InMux I__14794 (
            .O(N__68989),
            .I(N__68966));
    InMux I__14793 (
            .O(N__68988),
            .I(N__68966));
    InMux I__14792 (
            .O(N__68987),
            .I(N__68966));
    InMux I__14791 (
            .O(N__68986),
            .I(N__68966));
    InMux I__14790 (
            .O(N__68985),
            .I(N__68966));
    Span12Mux_v I__14789 (
            .O(N__68982),
            .I(N__68960));
    InMux I__14788 (
            .O(N__68981),
            .I(N__68957));
    LocalMux I__14787 (
            .O(N__68966),
            .I(N__68954));
    InMux I__14786 (
            .O(N__68965),
            .I(N__68947));
    InMux I__14785 (
            .O(N__68964),
            .I(N__68947));
    InMux I__14784 (
            .O(N__68963),
            .I(N__68947));
    Odrv12 I__14783 (
            .O(N__68960),
            .I(bluejay_data_out_31__N_704));
    LocalMux I__14782 (
            .O(N__68957),
            .I(bluejay_data_out_31__N_704));
    Odrv4 I__14781 (
            .O(N__68954),
            .I(bluejay_data_out_31__N_704));
    LocalMux I__14780 (
            .O(N__68947),
            .I(bluejay_data_out_31__N_704));
    InMux I__14779 (
            .O(N__68938),
            .I(N__68935));
    LocalMux I__14778 (
            .O(N__68935),
            .I(N__68932));
    Span4Mux_v I__14777 (
            .O(N__68932),
            .I(N__68928));
    CascadeMux I__14776 (
            .O(N__68931),
            .I(N__68925));
    Span4Mux_h I__14775 (
            .O(N__68928),
            .I(N__68922));
    InMux I__14774 (
            .O(N__68925),
            .I(N__68919));
    Odrv4 I__14773 (
            .O(N__68922),
            .I(fifo_data_out_14));
    LocalMux I__14772 (
            .O(N__68919),
            .I(fifo_data_out_14));
    InMux I__14771 (
            .O(N__68914),
            .I(N__68884));
    InMux I__14770 (
            .O(N__68913),
            .I(N__68884));
    InMux I__14769 (
            .O(N__68912),
            .I(N__68884));
    InMux I__14768 (
            .O(N__68911),
            .I(N__68884));
    InMux I__14767 (
            .O(N__68910),
            .I(N__68884));
    InMux I__14766 (
            .O(N__68909),
            .I(N__68884));
    InMux I__14765 (
            .O(N__68908),
            .I(N__68884));
    InMux I__14764 (
            .O(N__68907),
            .I(N__68884));
    InMux I__14763 (
            .O(N__68906),
            .I(N__68879));
    InMux I__14762 (
            .O(N__68905),
            .I(N__68879));
    InMux I__14761 (
            .O(N__68904),
            .I(N__68870));
    InMux I__14760 (
            .O(N__68903),
            .I(N__68870));
    InMux I__14759 (
            .O(N__68902),
            .I(N__68870));
    InMux I__14758 (
            .O(N__68901),
            .I(N__68870));
    LocalMux I__14757 (
            .O(N__68884),
            .I(N__68860));
    LocalMux I__14756 (
            .O(N__68879),
            .I(N__68855));
    LocalMux I__14755 (
            .O(N__68870),
            .I(N__68855));
    InMux I__14754 (
            .O(N__68869),
            .I(N__68846));
    InMux I__14753 (
            .O(N__68868),
            .I(N__68846));
    InMux I__14752 (
            .O(N__68867),
            .I(N__68846));
    InMux I__14751 (
            .O(N__68866),
            .I(N__68846));
    InMux I__14750 (
            .O(N__68865),
            .I(N__68839));
    InMux I__14749 (
            .O(N__68864),
            .I(N__68839));
    InMux I__14748 (
            .O(N__68863),
            .I(N__68839));
    Odrv12 I__14747 (
            .O(N__68860),
            .I(bluejay_data_out_31__N_703));
    Odrv4 I__14746 (
            .O(N__68855),
            .I(bluejay_data_out_31__N_703));
    LocalMux I__14745 (
            .O(N__68846),
            .I(bluejay_data_out_31__N_703));
    LocalMux I__14744 (
            .O(N__68839),
            .I(bluejay_data_out_31__N_703));
    IoInMux I__14743 (
            .O(N__68830),
            .I(N__68826));
    IoInMux I__14742 (
            .O(N__68829),
            .I(N__68823));
    LocalMux I__14741 (
            .O(N__68826),
            .I(N__68820));
    LocalMux I__14740 (
            .O(N__68823),
            .I(N__68817));
    Span4Mux_s3_h I__14739 (
            .O(N__68820),
            .I(N__68814));
    Sp12to4 I__14738 (
            .O(N__68817),
            .I(N__68811));
    Span4Mux_h I__14737 (
            .O(N__68814),
            .I(N__68808));
    Span12Mux_v I__14736 (
            .O(N__68811),
            .I(N__68805));
    Span4Mux_v I__14735 (
            .O(N__68808),
            .I(N__68802));
    Span12Mux_h I__14734 (
            .O(N__68805),
            .I(N__68799));
    Span4Mux_v I__14733 (
            .O(N__68802),
            .I(N__68796));
    Odrv12 I__14732 (
            .O(N__68799),
            .I(DATA14_c));
    Odrv4 I__14731 (
            .O(N__68796),
            .I(DATA14_c));
    CascadeMux I__14730 (
            .O(N__68791),
            .I(\tx_fifo.lscc_fifo_inst.n13544_cascade_ ));
    CascadeMux I__14729 (
            .O(N__68788),
            .I(\bluejay_data_inst.n11418_cascade_ ));
    CascadeMux I__14728 (
            .O(N__68785),
            .I(N__68782));
    InMux I__14727 (
            .O(N__68782),
            .I(N__68779));
    LocalMux I__14726 (
            .O(N__68779),
            .I(\bluejay_data_inst.n11330 ));
    InMux I__14725 (
            .O(N__68776),
            .I(N__68772));
    CascadeMux I__14724 (
            .O(N__68775),
            .I(N__68769));
    LocalMux I__14723 (
            .O(N__68772),
            .I(N__68766));
    InMux I__14722 (
            .O(N__68769),
            .I(N__68763));
    Odrv4 I__14721 (
            .O(N__68766),
            .I(\bluejay_data_inst.v_counter_2 ));
    LocalMux I__14720 (
            .O(N__68763),
            .I(\bluejay_data_inst.v_counter_2 ));
    InMux I__14719 (
            .O(N__68758),
            .I(N__68754));
    CascadeMux I__14718 (
            .O(N__68757),
            .I(N__68751));
    LocalMux I__14717 (
            .O(N__68754),
            .I(N__68748));
    InMux I__14716 (
            .O(N__68751),
            .I(N__68745));
    Odrv4 I__14715 (
            .O(N__68748),
            .I(\bluejay_data_inst.v_counter_4 ));
    LocalMux I__14714 (
            .O(N__68745),
            .I(\bluejay_data_inst.v_counter_4 ));
    InMux I__14713 (
            .O(N__68740),
            .I(N__68736));
    InMux I__14712 (
            .O(N__68739),
            .I(N__68733));
    LocalMux I__14711 (
            .O(N__68736),
            .I(\bluejay_data_inst.v_counter_8 ));
    LocalMux I__14710 (
            .O(N__68733),
            .I(\bluejay_data_inst.v_counter_8 ));
    InMux I__14709 (
            .O(N__68728),
            .I(N__68725));
    LocalMux I__14708 (
            .O(N__68725),
            .I(N__68721));
    InMux I__14707 (
            .O(N__68724),
            .I(N__68718));
    Odrv4 I__14706 (
            .O(N__68721),
            .I(\bluejay_data_inst.v_counter_0 ));
    LocalMux I__14705 (
            .O(N__68718),
            .I(\bluejay_data_inst.v_counter_0 ));
    CascadeMux I__14704 (
            .O(N__68713),
            .I(\bluejay_data_inst.n10_adj_1180_cascade_ ));
    InMux I__14703 (
            .O(N__68710),
            .I(N__68707));
    LocalMux I__14702 (
            .O(N__68707),
            .I(\bluejay_data_inst.n14 ));
    InMux I__14701 (
            .O(N__68704),
            .I(N__68701));
    LocalMux I__14700 (
            .O(N__68701),
            .I(\bluejay_data_inst.n10 ));
    InMux I__14699 (
            .O(N__68698),
            .I(N__68692));
    InMux I__14698 (
            .O(N__68697),
            .I(N__68692));
    LocalMux I__14697 (
            .O(N__68692),
            .I(N__68688));
    InMux I__14696 (
            .O(N__68691),
            .I(N__68685));
    Odrv4 I__14695 (
            .O(N__68688),
            .I(\bluejay_data_inst.v_counter_5 ));
    LocalMux I__14694 (
            .O(N__68685),
            .I(\bluejay_data_inst.v_counter_5 ));
    InMux I__14693 (
            .O(N__68680),
            .I(N__68676));
    InMux I__14692 (
            .O(N__68679),
            .I(N__68673));
    LocalMux I__14691 (
            .O(N__68676),
            .I(N__68667));
    LocalMux I__14690 (
            .O(N__68673),
            .I(N__68667));
    InMux I__14689 (
            .O(N__68672),
            .I(N__68664));
    Odrv12 I__14688 (
            .O(N__68667),
            .I(\bluejay_data_inst.v_counter_3 ));
    LocalMux I__14687 (
            .O(N__68664),
            .I(\bluejay_data_inst.v_counter_3 ));
    CascadeMux I__14686 (
            .O(N__68659),
            .I(\bluejay_data_inst.n10_cascade_ ));
    InMux I__14685 (
            .O(N__68656),
            .I(N__68649));
    InMux I__14684 (
            .O(N__68655),
            .I(N__68649));
    CascadeMux I__14683 (
            .O(N__68654),
            .I(N__68646));
    LocalMux I__14682 (
            .O(N__68649),
            .I(N__68643));
    InMux I__14681 (
            .O(N__68646),
            .I(N__68640));
    Odrv4 I__14680 (
            .O(N__68643),
            .I(\bluejay_data_inst.v_counter_6 ));
    LocalMux I__14679 (
            .O(N__68640),
            .I(\bluejay_data_inst.v_counter_6 ));
    InMux I__14678 (
            .O(N__68635),
            .I(N__68632));
    LocalMux I__14677 (
            .O(N__68632),
            .I(N__68629));
    Odrv4 I__14676 (
            .O(N__68629),
            .I(\bluejay_data_inst.n10781 ));
    CEMux I__14675 (
            .O(N__68626),
            .I(N__68623));
    LocalMux I__14674 (
            .O(N__68623),
            .I(N__68619));
    CEMux I__14673 (
            .O(N__68622),
            .I(N__68616));
    Span4Mux_v I__14672 (
            .O(N__68619),
            .I(N__68611));
    LocalMux I__14671 (
            .O(N__68616),
            .I(N__68611));
    Span4Mux_h I__14670 (
            .O(N__68611),
            .I(N__68608));
    Odrv4 I__14669 (
            .O(N__68608),
            .I(\bluejay_data_inst.n4162 ));
    InMux I__14668 (
            .O(N__68605),
            .I(N__68595));
    InMux I__14667 (
            .O(N__68604),
            .I(N__68592));
    InMux I__14666 (
            .O(N__68603),
            .I(N__68581));
    InMux I__14665 (
            .O(N__68602),
            .I(N__68581));
    InMux I__14664 (
            .O(N__68601),
            .I(N__68581));
    InMux I__14663 (
            .O(N__68600),
            .I(N__68581));
    InMux I__14662 (
            .O(N__68599),
            .I(N__68581));
    CascadeMux I__14661 (
            .O(N__68598),
            .I(N__68576));
    LocalMux I__14660 (
            .O(N__68595),
            .I(N__68572));
    LocalMux I__14659 (
            .O(N__68592),
            .I(N__68567));
    LocalMux I__14658 (
            .O(N__68581),
            .I(N__68567));
    InMux I__14657 (
            .O(N__68580),
            .I(N__68558));
    InMux I__14656 (
            .O(N__68579),
            .I(N__68558));
    InMux I__14655 (
            .O(N__68576),
            .I(N__68558));
    InMux I__14654 (
            .O(N__68575),
            .I(N__68558));
    Span4Mux_v I__14653 (
            .O(N__68572),
            .I(N__68555));
    Span4Mux_v I__14652 (
            .O(N__68567),
            .I(N__68552));
    LocalMux I__14651 (
            .O(N__68558),
            .I(N__68549));
    Odrv4 I__14650 (
            .O(N__68555),
            .I(buffer_switch_done_latched));
    Odrv4 I__14649 (
            .O(N__68552),
            .I(buffer_switch_done_latched));
    Odrv4 I__14648 (
            .O(N__68549),
            .I(buffer_switch_done_latched));
    CascadeMux I__14647 (
            .O(N__68542),
            .I(N__68539));
    InMux I__14646 (
            .O(N__68539),
            .I(N__68535));
    CascadeMux I__14645 (
            .O(N__68538),
            .I(N__68532));
    LocalMux I__14644 (
            .O(N__68535),
            .I(N__68529));
    InMux I__14643 (
            .O(N__68532),
            .I(N__68524));
    Span4Mux_v I__14642 (
            .O(N__68529),
            .I(N__68521));
    InMux I__14641 (
            .O(N__68528),
            .I(N__68516));
    InMux I__14640 (
            .O(N__68527),
            .I(N__68516));
    LocalMux I__14639 (
            .O(N__68524),
            .I(N__68513));
    Odrv4 I__14638 (
            .O(N__68521),
            .I(\bluejay_data_inst.n21 ));
    LocalMux I__14637 (
            .O(N__68516),
            .I(\bluejay_data_inst.n21 ));
    Odrv4 I__14636 (
            .O(N__68513),
            .I(\bluejay_data_inst.n21 ));
    InMux I__14635 (
            .O(N__68506),
            .I(N__68503));
    LocalMux I__14634 (
            .O(N__68503),
            .I(N__68500));
    Span4Mux_v I__14633 (
            .O(N__68500),
            .I(N__68497));
    Sp12to4 I__14632 (
            .O(N__68497),
            .I(N__68493));
    InMux I__14631 (
            .O(N__68496),
            .I(N__68490));
    Odrv12 I__14630 (
            .O(N__68493),
            .I(fifo_data_out_13));
    LocalMux I__14629 (
            .O(N__68490),
            .I(fifo_data_out_13));
    IoInMux I__14628 (
            .O(N__68485),
            .I(N__68482));
    LocalMux I__14627 (
            .O(N__68482),
            .I(N__68478));
    IoInMux I__14626 (
            .O(N__68481),
            .I(N__68475));
    IoSpan4Mux I__14625 (
            .O(N__68478),
            .I(N__68472));
    LocalMux I__14624 (
            .O(N__68475),
            .I(N__68469));
    Span4Mux_s0_v I__14623 (
            .O(N__68472),
            .I(N__68466));
    IoSpan4Mux I__14622 (
            .O(N__68469),
            .I(N__68463));
    Sp12to4 I__14621 (
            .O(N__68466),
            .I(N__68460));
    Span4Mux_s3_h I__14620 (
            .O(N__68463),
            .I(N__68457));
    Span12Mux_v I__14619 (
            .O(N__68460),
            .I(N__68454));
    Span4Mux_h I__14618 (
            .O(N__68457),
            .I(N__68451));
    Span12Mux_h I__14617 (
            .O(N__68454),
            .I(N__68448));
    Span4Mux_v I__14616 (
            .O(N__68451),
            .I(N__68445));
    Odrv12 I__14615 (
            .O(N__68448),
            .I(DATA13_c));
    Odrv4 I__14614 (
            .O(N__68445),
            .I(DATA13_c));
    InMux I__14613 (
            .O(N__68440),
            .I(N__68437));
    LocalMux I__14612 (
            .O(N__68437),
            .I(N__68434));
    Span4Mux_v I__14611 (
            .O(N__68434),
            .I(N__68430));
    InMux I__14610 (
            .O(N__68433),
            .I(N__68427));
    Odrv4 I__14609 (
            .O(N__68430),
            .I(fifo_data_out_12));
    LocalMux I__14608 (
            .O(N__68427),
            .I(fifo_data_out_12));
    IoInMux I__14607 (
            .O(N__68422),
            .I(N__68419));
    LocalMux I__14606 (
            .O(N__68419),
            .I(N__68416));
    IoSpan4Mux I__14605 (
            .O(N__68416),
            .I(N__68413));
    Span4Mux_s0_v I__14604 (
            .O(N__68413),
            .I(N__68410));
    Sp12to4 I__14603 (
            .O(N__68410),
            .I(N__68407));
    Span12Mux_s11_v I__14602 (
            .O(N__68407),
            .I(N__68403));
    IoInMux I__14601 (
            .O(N__68406),
            .I(N__68400));
    Span12Mux_h I__14600 (
            .O(N__68403),
            .I(N__68395));
    LocalMux I__14599 (
            .O(N__68400),
            .I(N__68395));
    Span12Mux_s10_h I__14598 (
            .O(N__68395),
            .I(N__68392));
    Odrv12 I__14597 (
            .O(N__68392),
            .I(DATA12_c));
    InMux I__14596 (
            .O(N__68389),
            .I(\bluejay_data_inst.n10646 ));
    InMux I__14595 (
            .O(N__68386),
            .I(\bluejay_data_inst.n10647 ));
    InMux I__14594 (
            .O(N__68383),
            .I(\bluejay_data_inst.n10648 ));
    InMux I__14593 (
            .O(N__68380),
            .I(\bluejay_data_inst.n10649 ));
    InMux I__14592 (
            .O(N__68377),
            .I(bfn_18_12_0_));
    InMux I__14591 (
            .O(N__68374),
            .I(\bluejay_data_inst.n10651 ));
    InMux I__14590 (
            .O(N__68371),
            .I(\bluejay_data_inst.n10652 ));
    InMux I__14589 (
            .O(N__68368),
            .I(N__68364));
    InMux I__14588 (
            .O(N__68367),
            .I(N__68361));
    LocalMux I__14587 (
            .O(N__68364),
            .I(\bluejay_data_inst.v_counter_10 ));
    LocalMux I__14586 (
            .O(N__68361),
            .I(\bluejay_data_inst.v_counter_10 ));
    InMux I__14585 (
            .O(N__68356),
            .I(N__68352));
    InMux I__14584 (
            .O(N__68355),
            .I(N__68349));
    LocalMux I__14583 (
            .O(N__68352),
            .I(\bluejay_data_inst.v_counter_9 ));
    LocalMux I__14582 (
            .O(N__68349),
            .I(\bluejay_data_inst.v_counter_9 ));
    CascadeMux I__14581 (
            .O(N__68344),
            .I(N__68341));
    InMux I__14580 (
            .O(N__68341),
            .I(N__68338));
    LocalMux I__14579 (
            .O(N__68338),
            .I(N__68334));
    InMux I__14578 (
            .O(N__68337),
            .I(N__68331));
    Odrv4 I__14577 (
            .O(N__68334),
            .I(\bluejay_data_inst.v_counter_7 ));
    LocalMux I__14576 (
            .O(N__68331),
            .I(\bluejay_data_inst.v_counter_7 ));
    InMux I__14575 (
            .O(N__68326),
            .I(N__68323));
    LocalMux I__14574 (
            .O(N__68323),
            .I(N__68319));
    InMux I__14573 (
            .O(N__68322),
            .I(N__68316));
    Odrv12 I__14572 (
            .O(N__68319),
            .I(\bluejay_data_inst.v_counter_1 ));
    LocalMux I__14571 (
            .O(N__68316),
            .I(\bluejay_data_inst.v_counter_1 ));
    CascadeMux I__14570 (
            .O(N__68311),
            .I(N__68307));
    InMux I__14569 (
            .O(N__68310),
            .I(N__68302));
    InMux I__14568 (
            .O(N__68307),
            .I(N__68302));
    LocalMux I__14567 (
            .O(N__68302),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_8 ));
    InMux I__14566 (
            .O(N__68299),
            .I(N__68289));
    InMux I__14565 (
            .O(N__68298),
            .I(N__68285));
    InMux I__14564 (
            .O(N__68297),
            .I(N__68282));
    InMux I__14563 (
            .O(N__68296),
            .I(N__68279));
    InMux I__14562 (
            .O(N__68295),
            .I(N__68275));
    InMux I__14561 (
            .O(N__68294),
            .I(N__68269));
    InMux I__14560 (
            .O(N__68293),
            .I(N__68269));
    InMux I__14559 (
            .O(N__68292),
            .I(N__68266));
    LocalMux I__14558 (
            .O(N__68289),
            .I(N__68262));
    InMux I__14557 (
            .O(N__68288),
            .I(N__68259));
    LocalMux I__14556 (
            .O(N__68285),
            .I(N__68256));
    LocalMux I__14555 (
            .O(N__68282),
            .I(N__68253));
    LocalMux I__14554 (
            .O(N__68279),
            .I(N__68250));
    InMux I__14553 (
            .O(N__68278),
            .I(N__68247));
    LocalMux I__14552 (
            .O(N__68275),
            .I(N__68241));
    InMux I__14551 (
            .O(N__68274),
            .I(N__68238));
    LocalMux I__14550 (
            .O(N__68269),
            .I(N__68232));
    LocalMux I__14549 (
            .O(N__68266),
            .I(N__68232));
    InMux I__14548 (
            .O(N__68265),
            .I(N__68229));
    Span4Mux_v I__14547 (
            .O(N__68262),
            .I(N__68226));
    LocalMux I__14546 (
            .O(N__68259),
            .I(N__68223));
    Span4Mux_v I__14545 (
            .O(N__68256),
            .I(N__68220));
    Span4Mux_v I__14544 (
            .O(N__68253),
            .I(N__68217));
    Span4Mux_v I__14543 (
            .O(N__68250),
            .I(N__68212));
    LocalMux I__14542 (
            .O(N__68247),
            .I(N__68212));
    InMux I__14541 (
            .O(N__68246),
            .I(N__68207));
    InMux I__14540 (
            .O(N__68245),
            .I(N__68207));
    InMux I__14539 (
            .O(N__68244),
            .I(N__68204));
    Span4Mux_v I__14538 (
            .O(N__68241),
            .I(N__68201));
    LocalMux I__14537 (
            .O(N__68238),
            .I(N__68198));
    InMux I__14536 (
            .O(N__68237),
            .I(N__68195));
    Span4Mux_v I__14535 (
            .O(N__68232),
            .I(N__68190));
    LocalMux I__14534 (
            .O(N__68229),
            .I(N__68190));
    Span4Mux_v I__14533 (
            .O(N__68226),
            .I(N__68185));
    Span4Mux_v I__14532 (
            .O(N__68223),
            .I(N__68185));
    Span4Mux_h I__14531 (
            .O(N__68220),
            .I(N__68178));
    Span4Mux_v I__14530 (
            .O(N__68217),
            .I(N__68178));
    Span4Mux_h I__14529 (
            .O(N__68212),
            .I(N__68178));
    LocalMux I__14528 (
            .O(N__68207),
            .I(N__68173));
    LocalMux I__14527 (
            .O(N__68204),
            .I(N__68173));
    Span4Mux_v I__14526 (
            .O(N__68201),
            .I(N__68168));
    Span4Mux_v I__14525 (
            .O(N__68198),
            .I(N__68168));
    LocalMux I__14524 (
            .O(N__68195),
            .I(N__68165));
    Span4Mux_h I__14523 (
            .O(N__68190),
            .I(N__68156));
    Span4Mux_h I__14522 (
            .O(N__68185),
            .I(N__68156));
    Span4Mux_h I__14521 (
            .O(N__68178),
            .I(N__68156));
    Span4Mux_v I__14520 (
            .O(N__68173),
            .I(N__68156));
    Odrv4 I__14519 (
            .O(N__68168),
            .I(n22));
    Odrv4 I__14518 (
            .O(N__68165),
            .I(n22));
    Odrv4 I__14517 (
            .O(N__68156),
            .I(n22));
    InMux I__14516 (
            .O(N__68149),
            .I(N__68146));
    LocalMux I__14515 (
            .O(N__68146),
            .I(N__68142));
    InMux I__14514 (
            .O(N__68145),
            .I(N__68139));
    Odrv12 I__14513 (
            .O(N__68142),
            .I(REG_mem_43_4));
    LocalMux I__14512 (
            .O(N__68139),
            .I(REG_mem_43_4));
    CascadeMux I__14511 (
            .O(N__68134),
            .I(N__68130));
    InMux I__14510 (
            .O(N__68133),
            .I(N__68125));
    InMux I__14509 (
            .O(N__68130),
            .I(N__68125));
    LocalMux I__14508 (
            .O(N__68125),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_8 ));
    InMux I__14507 (
            .O(N__68122),
            .I(N__68118));
    InMux I__14506 (
            .O(N__68121),
            .I(N__68115));
    LocalMux I__14505 (
            .O(N__68118),
            .I(REG_mem_5_4));
    LocalMux I__14504 (
            .O(N__68115),
            .I(REG_mem_5_4));
    InMux I__14503 (
            .O(N__68110),
            .I(N__68106));
    InMux I__14502 (
            .O(N__68109),
            .I(N__68103));
    LocalMux I__14501 (
            .O(N__68106),
            .I(REG_mem_4_4));
    LocalMux I__14500 (
            .O(N__68103),
            .I(REG_mem_4_4));
    InMux I__14499 (
            .O(N__68098),
            .I(N__68095));
    LocalMux I__14498 (
            .O(N__68095),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12520 ));
    InMux I__14497 (
            .O(N__68092),
            .I(N__68089));
    LocalMux I__14496 (
            .O(N__68089),
            .I(N__68082));
    InMux I__14495 (
            .O(N__68088),
            .I(N__68079));
    InMux I__14494 (
            .O(N__68087),
            .I(N__68072));
    InMux I__14493 (
            .O(N__68086),
            .I(N__68068));
    InMux I__14492 (
            .O(N__68085),
            .I(N__68065));
    Span4Mux_h I__14491 (
            .O(N__68082),
            .I(N__68060));
    LocalMux I__14490 (
            .O(N__68079),
            .I(N__68060));
    InMux I__14489 (
            .O(N__68078),
            .I(N__68057));
    InMux I__14488 (
            .O(N__68077),
            .I(N__68054));
    InMux I__14487 (
            .O(N__68076),
            .I(N__68051));
    InMux I__14486 (
            .O(N__68075),
            .I(N__68046));
    LocalMux I__14485 (
            .O(N__68072),
            .I(N__68042));
    InMux I__14484 (
            .O(N__68071),
            .I(N__68039));
    LocalMux I__14483 (
            .O(N__68068),
            .I(N__68035));
    LocalMux I__14482 (
            .O(N__68065),
            .I(N__68031));
    Span4Mux_h I__14481 (
            .O(N__68060),
            .I(N__68026));
    LocalMux I__14480 (
            .O(N__68057),
            .I(N__68026));
    LocalMux I__14479 (
            .O(N__68054),
            .I(N__68023));
    LocalMux I__14478 (
            .O(N__68051),
            .I(N__68020));
    InMux I__14477 (
            .O(N__68050),
            .I(N__68015));
    InMux I__14476 (
            .O(N__68049),
            .I(N__68015));
    LocalMux I__14475 (
            .O(N__68046),
            .I(N__68012));
    InMux I__14474 (
            .O(N__68045),
            .I(N__68009));
    Span4Mux_v I__14473 (
            .O(N__68042),
            .I(N__68004));
    LocalMux I__14472 (
            .O(N__68039),
            .I(N__68004));
    InMux I__14471 (
            .O(N__68038),
            .I(N__68001));
    Span4Mux_h I__14470 (
            .O(N__68035),
            .I(N__67997));
    InMux I__14469 (
            .O(N__68034),
            .I(N__67994));
    Span4Mux_v I__14468 (
            .O(N__68031),
            .I(N__67991));
    Span4Mux_v I__14467 (
            .O(N__68026),
            .I(N__67988));
    Span4Mux_v I__14466 (
            .O(N__68023),
            .I(N__67985));
    Span4Mux_v I__14465 (
            .O(N__68020),
            .I(N__67980));
    LocalMux I__14464 (
            .O(N__68015),
            .I(N__67980));
    Span4Mux_h I__14463 (
            .O(N__68012),
            .I(N__67977));
    LocalMux I__14462 (
            .O(N__68009),
            .I(N__67974));
    Span4Mux_h I__14461 (
            .O(N__68004),
            .I(N__67969));
    LocalMux I__14460 (
            .O(N__68001),
            .I(N__67969));
    InMux I__14459 (
            .O(N__68000),
            .I(N__67966));
    Span4Mux_h I__14458 (
            .O(N__67997),
            .I(N__67961));
    LocalMux I__14457 (
            .O(N__67994),
            .I(N__67961));
    Span4Mux_h I__14456 (
            .O(N__67991),
            .I(N__67952));
    Span4Mux_h I__14455 (
            .O(N__67988),
            .I(N__67952));
    Span4Mux_v I__14454 (
            .O(N__67985),
            .I(N__67952));
    Span4Mux_h I__14453 (
            .O(N__67980),
            .I(N__67952));
    Span4Mux_v I__14452 (
            .O(N__67977),
            .I(N__67947));
    Span4Mux_h I__14451 (
            .O(N__67974),
            .I(N__67947));
    Span4Mux_v I__14450 (
            .O(N__67969),
            .I(N__67940));
    LocalMux I__14449 (
            .O(N__67966),
            .I(N__67940));
    Span4Mux_h I__14448 (
            .O(N__67961),
            .I(N__67940));
    Odrv4 I__14447 (
            .O(N__67952),
            .I(n23));
    Odrv4 I__14446 (
            .O(N__67947),
            .I(n23));
    Odrv4 I__14445 (
            .O(N__67940),
            .I(n23));
    InMux I__14444 (
            .O(N__67933),
            .I(bfn_18_11_0_));
    InMux I__14443 (
            .O(N__67930),
            .I(\bluejay_data_inst.n10643 ));
    InMux I__14442 (
            .O(N__67927),
            .I(\bluejay_data_inst.n10644 ));
    InMux I__14441 (
            .O(N__67924),
            .I(\bluejay_data_inst.n10645 ));
    CascadeMux I__14440 (
            .O(N__67921),
            .I(N__67918));
    InMux I__14439 (
            .O(N__67918),
            .I(N__67915));
    LocalMux I__14438 (
            .O(N__67915),
            .I(N__67912));
    Odrv4 I__14437 (
            .O(N__67912),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12521 ));
    InMux I__14436 (
            .O(N__67909),
            .I(N__67906));
    LocalMux I__14435 (
            .O(N__67906),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12515 ));
    CascadeMux I__14434 (
            .O(N__67903),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13784_cascade_ ));
    InMux I__14433 (
            .O(N__67900),
            .I(N__67897));
    LocalMux I__14432 (
            .O(N__67897),
            .I(N__67894));
    Span4Mux_v I__14431 (
            .O(N__67894),
            .I(N__67891));
    Odrv4 I__14430 (
            .O(N__67891),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12514 ));
    InMux I__14429 (
            .O(N__67888),
            .I(N__67884));
    InMux I__14428 (
            .O(N__67887),
            .I(N__67880));
    LocalMux I__14427 (
            .O(N__67884),
            .I(N__67876));
    InMux I__14426 (
            .O(N__67883),
            .I(N__67870));
    LocalMux I__14425 (
            .O(N__67880),
            .I(N__67865));
    InMux I__14424 (
            .O(N__67879),
            .I(N__67861));
    Span4Mux_v I__14423 (
            .O(N__67876),
            .I(N__67858));
    InMux I__14422 (
            .O(N__67875),
            .I(N__67855));
    InMux I__14421 (
            .O(N__67874),
            .I(N__67851));
    InMux I__14420 (
            .O(N__67873),
            .I(N__67848));
    LocalMux I__14419 (
            .O(N__67870),
            .I(N__67843));
    InMux I__14418 (
            .O(N__67869),
            .I(N__67840));
    InMux I__14417 (
            .O(N__67868),
            .I(N__67837));
    Span4Mux_h I__14416 (
            .O(N__67865),
            .I(N__67834));
    InMux I__14415 (
            .O(N__67864),
            .I(N__67831));
    LocalMux I__14414 (
            .O(N__67861),
            .I(N__67828));
    Span4Mux_h I__14413 (
            .O(N__67858),
            .I(N__67823));
    LocalMux I__14412 (
            .O(N__67855),
            .I(N__67823));
    InMux I__14411 (
            .O(N__67854),
            .I(N__67820));
    LocalMux I__14410 (
            .O(N__67851),
            .I(N__67815));
    LocalMux I__14409 (
            .O(N__67848),
            .I(N__67815));
    InMux I__14408 (
            .O(N__67847),
            .I(N__67812));
    InMux I__14407 (
            .O(N__67846),
            .I(N__67809));
    Span4Mux_v I__14406 (
            .O(N__67843),
            .I(N__67804));
    LocalMux I__14405 (
            .O(N__67840),
            .I(N__67804));
    LocalMux I__14404 (
            .O(N__67837),
            .I(N__67801));
    Span4Mux_v I__14403 (
            .O(N__67834),
            .I(N__67795));
    LocalMux I__14402 (
            .O(N__67831),
            .I(N__67792));
    Span4Mux_h I__14401 (
            .O(N__67828),
            .I(N__67789));
    Span4Mux_h I__14400 (
            .O(N__67823),
            .I(N__67786));
    LocalMux I__14399 (
            .O(N__67820),
            .I(N__67783));
    Span12Mux_h I__14398 (
            .O(N__67815),
            .I(N__67776));
    LocalMux I__14397 (
            .O(N__67812),
            .I(N__67776));
    LocalMux I__14396 (
            .O(N__67809),
            .I(N__67776));
    Span4Mux_v I__14395 (
            .O(N__67804),
            .I(N__67771));
    Span4Mux_h I__14394 (
            .O(N__67801),
            .I(N__67771));
    InMux I__14393 (
            .O(N__67800),
            .I(N__67768));
    InMux I__14392 (
            .O(N__67799),
            .I(N__67765));
    InMux I__14391 (
            .O(N__67798),
            .I(N__67762));
    Odrv4 I__14390 (
            .O(N__67795),
            .I(n60));
    Odrv12 I__14389 (
            .O(N__67792),
            .I(n60));
    Odrv4 I__14388 (
            .O(N__67789),
            .I(n60));
    Odrv4 I__14387 (
            .O(N__67786),
            .I(n60));
    Odrv12 I__14386 (
            .O(N__67783),
            .I(n60));
    Odrv12 I__14385 (
            .O(N__67776),
            .I(n60));
    Odrv4 I__14384 (
            .O(N__67771),
            .I(n60));
    LocalMux I__14383 (
            .O(N__67768),
            .I(n60));
    LocalMux I__14382 (
            .O(N__67765),
            .I(n60));
    LocalMux I__14381 (
            .O(N__67762),
            .I(n60));
    CascadeMux I__14380 (
            .O(N__67741),
            .I(N__67737));
    InMux I__14379 (
            .O(N__67740),
            .I(N__67732));
    InMux I__14378 (
            .O(N__67737),
            .I(N__67732));
    LocalMux I__14377 (
            .O(N__67732),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_4 ));
    CascadeMux I__14376 (
            .O(N__67729),
            .I(N__67725));
    InMux I__14375 (
            .O(N__67728),
            .I(N__67720));
    InMux I__14374 (
            .O(N__67725),
            .I(N__67720));
    LocalMux I__14373 (
            .O(N__67720),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_4 ));
    InMux I__14372 (
            .O(N__67717),
            .I(N__67711));
    InMux I__14371 (
            .O(N__67716),
            .I(N__67708));
    InMux I__14370 (
            .O(N__67715),
            .I(N__67704));
    InMux I__14369 (
            .O(N__67714),
            .I(N__67701));
    LocalMux I__14368 (
            .O(N__67711),
            .I(N__67697));
    LocalMux I__14367 (
            .O(N__67708),
            .I(N__67693));
    InMux I__14366 (
            .O(N__67707),
            .I(N__67690));
    LocalMux I__14365 (
            .O(N__67704),
            .I(N__67687));
    LocalMux I__14364 (
            .O(N__67701),
            .I(N__67684));
    InMux I__14363 (
            .O(N__67700),
            .I(N__67681));
    Span4Mux_h I__14362 (
            .O(N__67697),
            .I(N__67678));
    InMux I__14361 (
            .O(N__67696),
            .I(N__67675));
    Span4Mux_v I__14360 (
            .O(N__67693),
            .I(N__67664));
    LocalMux I__14359 (
            .O(N__67690),
            .I(N__67661));
    Span4Mux_h I__14358 (
            .O(N__67687),
            .I(N__67658));
    Span4Mux_h I__14357 (
            .O(N__67684),
            .I(N__67653));
    LocalMux I__14356 (
            .O(N__67681),
            .I(N__67653));
    Span4Mux_v I__14355 (
            .O(N__67678),
            .I(N__67650));
    LocalMux I__14354 (
            .O(N__67675),
            .I(N__67647));
    InMux I__14353 (
            .O(N__67674),
            .I(N__67644));
    InMux I__14352 (
            .O(N__67673),
            .I(N__67641));
    InMux I__14351 (
            .O(N__67672),
            .I(N__67638));
    InMux I__14350 (
            .O(N__67671),
            .I(N__67633));
    InMux I__14349 (
            .O(N__67670),
            .I(N__67633));
    InMux I__14348 (
            .O(N__67669),
            .I(N__67630));
    InMux I__14347 (
            .O(N__67668),
            .I(N__67627));
    InMux I__14346 (
            .O(N__67667),
            .I(N__67624));
    Span4Mux_h I__14345 (
            .O(N__67664),
            .I(N__67618));
    Span4Mux_v I__14344 (
            .O(N__67661),
            .I(N__67618));
    Span4Mux_v I__14343 (
            .O(N__67658),
            .I(N__67613));
    Span4Mux_h I__14342 (
            .O(N__67653),
            .I(N__67613));
    Span4Mux_v I__14341 (
            .O(N__67650),
            .I(N__67608));
    Span4Mux_v I__14340 (
            .O(N__67647),
            .I(N__67608));
    LocalMux I__14339 (
            .O(N__67644),
            .I(N__67603));
    LocalMux I__14338 (
            .O(N__67641),
            .I(N__67603));
    LocalMux I__14337 (
            .O(N__67638),
            .I(N__67594));
    LocalMux I__14336 (
            .O(N__67633),
            .I(N__67594));
    LocalMux I__14335 (
            .O(N__67630),
            .I(N__67594));
    LocalMux I__14334 (
            .O(N__67627),
            .I(N__67594));
    LocalMux I__14333 (
            .O(N__67624),
            .I(N__67591));
    InMux I__14332 (
            .O(N__67623),
            .I(N__67588));
    Odrv4 I__14331 (
            .O(N__67618),
            .I(n2));
    Odrv4 I__14330 (
            .O(N__67613),
            .I(n2));
    Odrv4 I__14329 (
            .O(N__67608),
            .I(n2));
    Odrv12 I__14328 (
            .O(N__67603),
            .I(n2));
    Odrv12 I__14327 (
            .O(N__67594),
            .I(n2));
    Odrv4 I__14326 (
            .O(N__67591),
            .I(n2));
    LocalMux I__14325 (
            .O(N__67588),
            .I(n2));
    InMux I__14324 (
            .O(N__67573),
            .I(N__67569));
    InMux I__14323 (
            .O(N__67572),
            .I(N__67566));
    LocalMux I__14322 (
            .O(N__67569),
            .I(REG_mem_63_8));
    LocalMux I__14321 (
            .O(N__67566),
            .I(REG_mem_63_8));
    InMux I__14320 (
            .O(N__67561),
            .I(N__67558));
    LocalMux I__14319 (
            .O(N__67558),
            .I(N__67554));
    InMux I__14318 (
            .O(N__67557),
            .I(N__67551));
    Odrv12 I__14317 (
            .O(N__67554),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_8 ));
    LocalMux I__14316 (
            .O(N__67551),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_8 ));
    CascadeMux I__14315 (
            .O(N__67546),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13382_cascade_ ));
    InMux I__14314 (
            .O(N__67543),
            .I(N__67537));
    InMux I__14313 (
            .O(N__67542),
            .I(N__67537));
    LocalMux I__14312 (
            .O(N__67537),
            .I(N__67534));
    Odrv4 I__14311 (
            .O(N__67534),
            .I(REG_mem_17_8));
    CascadeMux I__14310 (
            .O(N__67531),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14108_cascade_ ));
    InMux I__14309 (
            .O(N__67528),
            .I(N__67525));
    LocalMux I__14308 (
            .O(N__67525),
            .I(N__67521));
    InMux I__14307 (
            .O(N__67524),
            .I(N__67518));
    Odrv12 I__14306 (
            .O(N__67521),
            .I(REG_mem_16_8));
    LocalMux I__14305 (
            .O(N__67518),
            .I(REG_mem_16_8));
    InMux I__14304 (
            .O(N__67513),
            .I(N__67506));
    CascadeMux I__14303 (
            .O(N__67512),
            .I(N__67500));
    InMux I__14302 (
            .O(N__67511),
            .I(N__67496));
    InMux I__14301 (
            .O(N__67510),
            .I(N__67493));
    InMux I__14300 (
            .O(N__67509),
            .I(N__67487));
    LocalMux I__14299 (
            .O(N__67506),
            .I(N__67483));
    InMux I__14298 (
            .O(N__67505),
            .I(N__67480));
    InMux I__14297 (
            .O(N__67504),
            .I(N__67477));
    InMux I__14296 (
            .O(N__67503),
            .I(N__67474));
    InMux I__14295 (
            .O(N__67500),
            .I(N__67471));
    InMux I__14294 (
            .O(N__67499),
            .I(N__67468));
    LocalMux I__14293 (
            .O(N__67496),
            .I(N__67464));
    LocalMux I__14292 (
            .O(N__67493),
            .I(N__67461));
    InMux I__14291 (
            .O(N__67492),
            .I(N__67455));
    InMux I__14290 (
            .O(N__67491),
            .I(N__67455));
    InMux I__14289 (
            .O(N__67490),
            .I(N__67452));
    LocalMux I__14288 (
            .O(N__67487),
            .I(N__67449));
    InMux I__14287 (
            .O(N__67486),
            .I(N__67446));
    Span4Mux_h I__14286 (
            .O(N__67483),
            .I(N__67441));
    LocalMux I__14285 (
            .O(N__67480),
            .I(N__67441));
    LocalMux I__14284 (
            .O(N__67477),
            .I(N__67438));
    LocalMux I__14283 (
            .O(N__67474),
            .I(N__67435));
    LocalMux I__14282 (
            .O(N__67471),
            .I(N__67430));
    LocalMux I__14281 (
            .O(N__67468),
            .I(N__67430));
    InMux I__14280 (
            .O(N__67467),
            .I(N__67427));
    Span4Mux_h I__14279 (
            .O(N__67464),
            .I(N__67422));
    Span4Mux_v I__14278 (
            .O(N__67461),
            .I(N__67422));
    InMux I__14277 (
            .O(N__67460),
            .I(N__67418));
    LocalMux I__14276 (
            .O(N__67455),
            .I(N__67415));
    LocalMux I__14275 (
            .O(N__67452),
            .I(N__67412));
    Span4Mux_h I__14274 (
            .O(N__67449),
            .I(N__67409));
    LocalMux I__14273 (
            .O(N__67446),
            .I(N__67404));
    Span4Mux_v I__14272 (
            .O(N__67441),
            .I(N__67404));
    Span4Mux_v I__14271 (
            .O(N__67438),
            .I(N__67401));
    Span4Mux_h I__14270 (
            .O(N__67435),
            .I(N__67398));
    Span4Mux_h I__14269 (
            .O(N__67430),
            .I(N__67395));
    LocalMux I__14268 (
            .O(N__67427),
            .I(N__67390));
    Span4Mux_h I__14267 (
            .O(N__67422),
            .I(N__67390));
    InMux I__14266 (
            .O(N__67421),
            .I(N__67387));
    LocalMux I__14265 (
            .O(N__67418),
            .I(N__67384));
    Span4Mux_v I__14264 (
            .O(N__67415),
            .I(N__67381));
    Span4Mux_v I__14263 (
            .O(N__67412),
            .I(N__67372));
    Span4Mux_h I__14262 (
            .O(N__67409),
            .I(N__67372));
    Span4Mux_h I__14261 (
            .O(N__67404),
            .I(N__67372));
    Span4Mux_v I__14260 (
            .O(N__67401),
            .I(N__67372));
    Span4Mux_h I__14259 (
            .O(N__67398),
            .I(N__67365));
    Span4Mux_h I__14258 (
            .O(N__67395),
            .I(N__67365));
    Span4Mux_v I__14257 (
            .O(N__67390),
            .I(N__67365));
    LocalMux I__14256 (
            .O(N__67387),
            .I(n47));
    Odrv12 I__14255 (
            .O(N__67384),
            .I(n47));
    Odrv4 I__14254 (
            .O(N__67381),
            .I(n47));
    Odrv4 I__14253 (
            .O(N__67372),
            .I(n47));
    Odrv4 I__14252 (
            .O(N__67365),
            .I(n47));
    InMux I__14251 (
            .O(N__67354),
            .I(N__67348));
    InMux I__14250 (
            .O(N__67353),
            .I(N__67348));
    LocalMux I__14249 (
            .O(N__67348),
            .I(REG_mem_18_8));
    InMux I__14248 (
            .O(N__67345),
            .I(N__67341));
    InMux I__14247 (
            .O(N__67344),
            .I(N__67333));
    LocalMux I__14246 (
            .O(N__67341),
            .I(N__67330));
    InMux I__14245 (
            .O(N__67340),
            .I(N__67327));
    InMux I__14244 (
            .O(N__67339),
            .I(N__67323));
    InMux I__14243 (
            .O(N__67338),
            .I(N__67319));
    InMux I__14242 (
            .O(N__67337),
            .I(N__67316));
    InMux I__14241 (
            .O(N__67336),
            .I(N__67313));
    LocalMux I__14240 (
            .O(N__67333),
            .I(N__67308));
    Span4Mux_h I__14239 (
            .O(N__67330),
            .I(N__67305));
    LocalMux I__14238 (
            .O(N__67327),
            .I(N__67302));
    InMux I__14237 (
            .O(N__67326),
            .I(N__67298));
    LocalMux I__14236 (
            .O(N__67323),
            .I(N__67295));
    InMux I__14235 (
            .O(N__67322),
            .I(N__67292));
    LocalMux I__14234 (
            .O(N__67319),
            .I(N__67285));
    LocalMux I__14233 (
            .O(N__67316),
            .I(N__67285));
    LocalMux I__14232 (
            .O(N__67313),
            .I(N__67285));
    InMux I__14231 (
            .O(N__67312),
            .I(N__67282));
    InMux I__14230 (
            .O(N__67311),
            .I(N__67279));
    Span4Mux_h I__14229 (
            .O(N__67308),
            .I(N__67275));
    Span4Mux_h I__14228 (
            .O(N__67305),
            .I(N__67270));
    Span4Mux_v I__14227 (
            .O(N__67302),
            .I(N__67270));
    InMux I__14226 (
            .O(N__67301),
            .I(N__67267));
    LocalMux I__14225 (
            .O(N__67298),
            .I(N__67263));
    Span4Mux_h I__14224 (
            .O(N__67295),
            .I(N__67260));
    LocalMux I__14223 (
            .O(N__67292),
            .I(N__67257));
    Span4Mux_h I__14222 (
            .O(N__67285),
            .I(N__67250));
    LocalMux I__14221 (
            .O(N__67282),
            .I(N__67250));
    LocalMux I__14220 (
            .O(N__67279),
            .I(N__67250));
    InMux I__14219 (
            .O(N__67278),
            .I(N__67247));
    Span4Mux_v I__14218 (
            .O(N__67275),
            .I(N__67240));
    Span4Mux_h I__14217 (
            .O(N__67270),
            .I(N__67240));
    LocalMux I__14216 (
            .O(N__67267),
            .I(N__67240));
    InMux I__14215 (
            .O(N__67266),
            .I(N__67237));
    Span4Mux_v I__14214 (
            .O(N__67263),
            .I(N__67232));
    Span4Mux_h I__14213 (
            .O(N__67260),
            .I(N__67227));
    Span4Mux_h I__14212 (
            .O(N__67257),
            .I(N__67227));
    Span4Mux_h I__14211 (
            .O(N__67250),
            .I(N__67224));
    LocalMux I__14210 (
            .O(N__67247),
            .I(N__67217));
    Sp12to4 I__14209 (
            .O(N__67240),
            .I(N__67217));
    LocalMux I__14208 (
            .O(N__67237),
            .I(N__67217));
    InMux I__14207 (
            .O(N__67236),
            .I(N__67214));
    InMux I__14206 (
            .O(N__67235),
            .I(N__67211));
    Odrv4 I__14205 (
            .O(N__67232),
            .I(n57));
    Odrv4 I__14204 (
            .O(N__67227),
            .I(n57));
    Odrv4 I__14203 (
            .O(N__67224),
            .I(n57));
    Odrv12 I__14202 (
            .O(N__67217),
            .I(n57));
    LocalMux I__14201 (
            .O(N__67214),
            .I(n57));
    LocalMux I__14200 (
            .O(N__67211),
            .I(n57));
    InMux I__14199 (
            .O(N__67198),
            .I(N__67189));
    InMux I__14198 (
            .O(N__67197),
            .I(N__67184));
    InMux I__14197 (
            .O(N__67196),
            .I(N__67179));
    InMux I__14196 (
            .O(N__67195),
            .I(N__67179));
    InMux I__14195 (
            .O(N__67194),
            .I(N__67176));
    InMux I__14194 (
            .O(N__67193),
            .I(N__67173));
    InMux I__14193 (
            .O(N__67192),
            .I(N__67170));
    LocalMux I__14192 (
            .O(N__67189),
            .I(N__67167));
    InMux I__14191 (
            .O(N__67188),
            .I(N__67164));
    InMux I__14190 (
            .O(N__67187),
            .I(N__67160));
    LocalMux I__14189 (
            .O(N__67184),
            .I(N__67157));
    LocalMux I__14188 (
            .O(N__67179),
            .I(N__67150));
    LocalMux I__14187 (
            .O(N__67176),
            .I(N__67147));
    LocalMux I__14186 (
            .O(N__67173),
            .I(N__67142));
    LocalMux I__14185 (
            .O(N__67170),
            .I(N__67142));
    Span4Mux_h I__14184 (
            .O(N__67167),
            .I(N__67137));
    LocalMux I__14183 (
            .O(N__67164),
            .I(N__67137));
    InMux I__14182 (
            .O(N__67163),
            .I(N__67134));
    LocalMux I__14181 (
            .O(N__67160),
            .I(N__67130));
    Span4Mux_h I__14180 (
            .O(N__67157),
            .I(N__67127));
    InMux I__14179 (
            .O(N__67156),
            .I(N__67124));
    InMux I__14178 (
            .O(N__67155),
            .I(N__67121));
    InMux I__14177 (
            .O(N__67154),
            .I(N__67118));
    InMux I__14176 (
            .O(N__67153),
            .I(N__67115));
    Span4Mux_v I__14175 (
            .O(N__67150),
            .I(N__67110));
    Span4Mux_h I__14174 (
            .O(N__67147),
            .I(N__67110));
    Span4Mux_h I__14173 (
            .O(N__67142),
            .I(N__67107));
    Span4Mux_h I__14172 (
            .O(N__67137),
            .I(N__67102));
    LocalMux I__14171 (
            .O(N__67134),
            .I(N__67102));
    InMux I__14170 (
            .O(N__67133),
            .I(N__67099));
    Span12Mux_v I__14169 (
            .O(N__67130),
            .I(N__67095));
    Sp12to4 I__14168 (
            .O(N__67127),
            .I(N__67090));
    LocalMux I__14167 (
            .O(N__67124),
            .I(N__67090));
    LocalMux I__14166 (
            .O(N__67121),
            .I(N__67087));
    LocalMux I__14165 (
            .O(N__67118),
            .I(N__67082));
    LocalMux I__14164 (
            .O(N__67115),
            .I(N__67082));
    Span4Mux_v I__14163 (
            .O(N__67110),
            .I(N__67073));
    Span4Mux_h I__14162 (
            .O(N__67107),
            .I(N__67073));
    Span4Mux_v I__14161 (
            .O(N__67102),
            .I(N__67073));
    LocalMux I__14160 (
            .O(N__67099),
            .I(N__67073));
    InMux I__14159 (
            .O(N__67098),
            .I(N__67070));
    Odrv12 I__14158 (
            .O(N__67095),
            .I(n56));
    Odrv12 I__14157 (
            .O(N__67090),
            .I(n56));
    Odrv4 I__14156 (
            .O(N__67087),
            .I(n56));
    Odrv4 I__14155 (
            .O(N__67082),
            .I(n56));
    Odrv4 I__14154 (
            .O(N__67073),
            .I(n56));
    LocalMux I__14153 (
            .O(N__67070),
            .I(n56));
    InMux I__14152 (
            .O(N__67057),
            .I(N__67053));
    InMux I__14151 (
            .O(N__67056),
            .I(N__67050));
    LocalMux I__14150 (
            .O(N__67053),
            .I(REG_mem_37_8));
    LocalMux I__14149 (
            .O(N__67050),
            .I(REG_mem_37_8));
    CascadeMux I__14148 (
            .O(N__67045),
            .I(N__67042));
    InMux I__14147 (
            .O(N__67042),
            .I(N__67039));
    LocalMux I__14146 (
            .O(N__67039),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13808 ));
    InMux I__14145 (
            .O(N__67036),
            .I(N__67033));
    LocalMux I__14144 (
            .O(N__67033),
            .I(N__67029));
    InMux I__14143 (
            .O(N__67032),
            .I(N__67026));
    Odrv12 I__14142 (
            .O(N__67029),
            .I(REG_mem_36_8));
    LocalMux I__14141 (
            .O(N__67026),
            .I(REG_mem_36_8));
    InMux I__14140 (
            .O(N__67021),
            .I(N__67018));
    LocalMux I__14139 (
            .O(N__67018),
            .I(N__67015));
    Odrv12 I__14138 (
            .O(N__67015),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11857 ));
    CascadeMux I__14137 (
            .O(N__67012),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13238_cascade_ ));
    InMux I__14136 (
            .O(N__67009),
            .I(N__67006));
    LocalMux I__14135 (
            .O(N__67006),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11807 ));
    InMux I__14134 (
            .O(N__67003),
            .I(N__67000));
    LocalMux I__14133 (
            .O(N__67000),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12347 ));
    InMux I__14132 (
            .O(N__66997),
            .I(N__66992));
    InMux I__14131 (
            .O(N__66996),
            .I(N__66989));
    InMux I__14130 (
            .O(N__66995),
            .I(N__66986));
    LocalMux I__14129 (
            .O(N__66992),
            .I(N__66981));
    LocalMux I__14128 (
            .O(N__66989),
            .I(N__66975));
    LocalMux I__14127 (
            .O(N__66986),
            .I(N__66968));
    InMux I__14126 (
            .O(N__66985),
            .I(N__66965));
    InMux I__14125 (
            .O(N__66984),
            .I(N__66962));
    Span4Mux_h I__14124 (
            .O(N__66981),
            .I(N__66956));
    InMux I__14123 (
            .O(N__66980),
            .I(N__66953));
    InMux I__14122 (
            .O(N__66979),
            .I(N__66948));
    InMux I__14121 (
            .O(N__66978),
            .I(N__66948));
    Span4Mux_v I__14120 (
            .O(N__66975),
            .I(N__66945));
    InMux I__14119 (
            .O(N__66974),
            .I(N__66942));
    InMux I__14118 (
            .O(N__66973),
            .I(N__66939));
    InMux I__14117 (
            .O(N__66972),
            .I(N__66934));
    InMux I__14116 (
            .O(N__66971),
            .I(N__66934));
    Span4Mux_v I__14115 (
            .O(N__66968),
            .I(N__66931));
    LocalMux I__14114 (
            .O(N__66965),
            .I(N__66928));
    LocalMux I__14113 (
            .O(N__66962),
            .I(N__66925));
    InMux I__14112 (
            .O(N__66961),
            .I(N__66922));
    InMux I__14111 (
            .O(N__66960),
            .I(N__66919));
    InMux I__14110 (
            .O(N__66959),
            .I(N__66916));
    Span4Mux_v I__14109 (
            .O(N__66956),
            .I(N__66910));
    LocalMux I__14108 (
            .O(N__66953),
            .I(N__66910));
    LocalMux I__14107 (
            .O(N__66948),
            .I(N__66907));
    Span4Mux_v I__14106 (
            .O(N__66945),
            .I(N__66904));
    LocalMux I__14105 (
            .O(N__66942),
            .I(N__66901));
    LocalMux I__14104 (
            .O(N__66939),
            .I(N__66898));
    LocalMux I__14103 (
            .O(N__66934),
            .I(N__66895));
    Span4Mux_h I__14102 (
            .O(N__66931),
            .I(N__66890));
    Span4Mux_v I__14101 (
            .O(N__66928),
            .I(N__66890));
    Span4Mux_v I__14100 (
            .O(N__66925),
            .I(N__66887));
    LocalMux I__14099 (
            .O(N__66922),
            .I(N__66882));
    LocalMux I__14098 (
            .O(N__66919),
            .I(N__66882));
    LocalMux I__14097 (
            .O(N__66916),
            .I(N__66879));
    InMux I__14096 (
            .O(N__66915),
            .I(N__66876));
    Span4Mux_h I__14095 (
            .O(N__66910),
            .I(N__66871));
    Span4Mux_v I__14094 (
            .O(N__66907),
            .I(N__66871));
    Span4Mux_h I__14093 (
            .O(N__66904),
            .I(N__66864));
    Span4Mux_v I__14092 (
            .O(N__66901),
            .I(N__66864));
    Span4Mux_h I__14091 (
            .O(N__66898),
            .I(N__66864));
    Span4Mux_h I__14090 (
            .O(N__66895),
            .I(N__66861));
    Span4Mux_h I__14089 (
            .O(N__66890),
            .I(N__66854));
    Span4Mux_v I__14088 (
            .O(N__66887),
            .I(N__66854));
    Span4Mux_v I__14087 (
            .O(N__66882),
            .I(N__66854));
    Span12Mux_v I__14086 (
            .O(N__66879),
            .I(N__66849));
    LocalMux I__14085 (
            .O(N__66876),
            .I(N__66849));
    Odrv4 I__14084 (
            .O(N__66871),
            .I(n55));
    Odrv4 I__14083 (
            .O(N__66864),
            .I(n55));
    Odrv4 I__14082 (
            .O(N__66861),
            .I(n55));
    Odrv4 I__14081 (
            .O(N__66854),
            .I(n55));
    Odrv12 I__14080 (
            .O(N__66849),
            .I(n55));
    InMux I__14079 (
            .O(N__66838),
            .I(N__66832));
    InMux I__14078 (
            .O(N__66837),
            .I(N__66832));
    LocalMux I__14077 (
            .O(N__66832),
            .I(REG_mem_10_2));
    InMux I__14076 (
            .O(N__66829),
            .I(N__66822));
    InMux I__14075 (
            .O(N__66828),
            .I(N__66819));
    InMux I__14074 (
            .O(N__66827),
            .I(N__66813));
    InMux I__14073 (
            .O(N__66826),
            .I(N__66809));
    InMux I__14072 (
            .O(N__66825),
            .I(N__66805));
    LocalMux I__14071 (
            .O(N__66822),
            .I(N__66799));
    LocalMux I__14070 (
            .O(N__66819),
            .I(N__66796));
    InMux I__14069 (
            .O(N__66818),
            .I(N__66793));
    InMux I__14068 (
            .O(N__66817),
            .I(N__66790));
    InMux I__14067 (
            .O(N__66816),
            .I(N__66787));
    LocalMux I__14066 (
            .O(N__66813),
            .I(N__66784));
    InMux I__14065 (
            .O(N__66812),
            .I(N__66781));
    LocalMux I__14064 (
            .O(N__66809),
            .I(N__66778));
    InMux I__14063 (
            .O(N__66808),
            .I(N__66775));
    LocalMux I__14062 (
            .O(N__66805),
            .I(N__66772));
    InMux I__14061 (
            .O(N__66804),
            .I(N__66769));
    InMux I__14060 (
            .O(N__66803),
            .I(N__66766));
    InMux I__14059 (
            .O(N__66802),
            .I(N__66763));
    Span4Mux_v I__14058 (
            .O(N__66799),
            .I(N__66758));
    Span4Mux_h I__14057 (
            .O(N__66796),
            .I(N__66755));
    LocalMux I__14056 (
            .O(N__66793),
            .I(N__66750));
    LocalMux I__14055 (
            .O(N__66790),
            .I(N__66750));
    LocalMux I__14054 (
            .O(N__66787),
            .I(N__66747));
    Span4Mux_v I__14053 (
            .O(N__66784),
            .I(N__66742));
    LocalMux I__14052 (
            .O(N__66781),
            .I(N__66742));
    Span4Mux_h I__14051 (
            .O(N__66778),
            .I(N__66739));
    LocalMux I__14050 (
            .O(N__66775),
            .I(N__66736));
    Span4Mux_v I__14049 (
            .O(N__66772),
            .I(N__66733));
    LocalMux I__14048 (
            .O(N__66769),
            .I(N__66730));
    LocalMux I__14047 (
            .O(N__66766),
            .I(N__66727));
    LocalMux I__14046 (
            .O(N__66763),
            .I(N__66724));
    InMux I__14045 (
            .O(N__66762),
            .I(N__66721));
    InMux I__14044 (
            .O(N__66761),
            .I(N__66718));
    Span4Mux_h I__14043 (
            .O(N__66758),
            .I(N__66710));
    Span4Mux_v I__14042 (
            .O(N__66755),
            .I(N__66710));
    Span4Mux_v I__14041 (
            .O(N__66750),
            .I(N__66710));
    Span4Mux_v I__14040 (
            .O(N__66747),
            .I(N__66705));
    Span4Mux_v I__14039 (
            .O(N__66742),
            .I(N__66705));
    Span4Mux_h I__14038 (
            .O(N__66739),
            .I(N__66700));
    Span4Mux_h I__14037 (
            .O(N__66736),
            .I(N__66700));
    Span4Mux_h I__14036 (
            .O(N__66733),
            .I(N__66691));
    Span4Mux_v I__14035 (
            .O(N__66730),
            .I(N__66691));
    Span4Mux_v I__14034 (
            .O(N__66727),
            .I(N__66691));
    Span4Mux_h I__14033 (
            .O(N__66724),
            .I(N__66691));
    LocalMux I__14032 (
            .O(N__66721),
            .I(N__66688));
    LocalMux I__14031 (
            .O(N__66718),
            .I(N__66685));
    InMux I__14030 (
            .O(N__66717),
            .I(N__66682));
    Odrv4 I__14029 (
            .O(N__66710),
            .I(n54));
    Odrv4 I__14028 (
            .O(N__66705),
            .I(n54));
    Odrv4 I__14027 (
            .O(N__66700),
            .I(n54));
    Odrv4 I__14026 (
            .O(N__66691),
            .I(n54));
    Odrv4 I__14025 (
            .O(N__66688),
            .I(n54));
    Odrv12 I__14024 (
            .O(N__66685),
            .I(n54));
    LocalMux I__14023 (
            .O(N__66682),
            .I(n54));
    InMux I__14022 (
            .O(N__66667),
            .I(N__66661));
    InMux I__14021 (
            .O(N__66666),
            .I(N__66661));
    LocalMux I__14020 (
            .O(N__66661),
            .I(REG_mem_11_2));
    InMux I__14019 (
            .O(N__66658),
            .I(N__66655));
    LocalMux I__14018 (
            .O(N__66655),
            .I(N__66652));
    Span4Mux_v I__14017 (
            .O(N__66652),
            .I(N__66649));
    Span4Mux_h I__14016 (
            .O(N__66649),
            .I(N__66645));
    InMux I__14015 (
            .O(N__66648),
            .I(N__66642));
    Odrv4 I__14014 (
            .O(N__66645),
            .I(REG_mem_8_2));
    LocalMux I__14013 (
            .O(N__66642),
            .I(REG_mem_8_2));
    InMux I__14012 (
            .O(N__66637),
            .I(N__66633));
    InMux I__14011 (
            .O(N__66636),
            .I(N__66630));
    LocalMux I__14010 (
            .O(N__66633),
            .I(REG_mem_9_2));
    LocalMux I__14009 (
            .O(N__66630),
            .I(REG_mem_9_2));
    InMux I__14008 (
            .O(N__66625),
            .I(N__66622));
    LocalMux I__14007 (
            .O(N__66622),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11806 ));
    CascadeMux I__14006 (
            .O(N__66619),
            .I(N__66616));
    InMux I__14005 (
            .O(N__66616),
            .I(N__66612));
    InMux I__14004 (
            .O(N__66615),
            .I(N__66609));
    LocalMux I__14003 (
            .O(N__66612),
            .I(REG_mem_50_4));
    LocalMux I__14002 (
            .O(N__66609),
            .I(REG_mem_50_4));
    InMux I__14001 (
            .O(N__66604),
            .I(N__66598));
    InMux I__14000 (
            .O(N__66603),
            .I(N__66598));
    LocalMux I__13999 (
            .O(N__66598),
            .I(REG_mem_51_4));
    InMux I__13998 (
            .O(N__66595),
            .I(N__66592));
    LocalMux I__13997 (
            .O(N__66592),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14348 ));
    InMux I__13996 (
            .O(N__66589),
            .I(N__66583));
    InMux I__13995 (
            .O(N__66588),
            .I(N__66574));
    InMux I__13994 (
            .O(N__66587),
            .I(N__66570));
    InMux I__13993 (
            .O(N__66586),
            .I(N__66567));
    LocalMux I__13992 (
            .O(N__66583),
            .I(N__66563));
    InMux I__13991 (
            .O(N__66582),
            .I(N__66560));
    InMux I__13990 (
            .O(N__66581),
            .I(N__66557));
    InMux I__13989 (
            .O(N__66580),
            .I(N__66554));
    InMux I__13988 (
            .O(N__66579),
            .I(N__66551));
    InMux I__13987 (
            .O(N__66578),
            .I(N__66548));
    InMux I__13986 (
            .O(N__66577),
            .I(N__66545));
    LocalMux I__13985 (
            .O(N__66574),
            .I(N__66542));
    InMux I__13984 (
            .O(N__66573),
            .I(N__66539));
    LocalMux I__13983 (
            .O(N__66570),
            .I(N__66534));
    LocalMux I__13982 (
            .O(N__66567),
            .I(N__66534));
    InMux I__13981 (
            .O(N__66566),
            .I(N__66531));
    Span4Mux_h I__13980 (
            .O(N__66563),
            .I(N__66526));
    LocalMux I__13979 (
            .O(N__66560),
            .I(N__66523));
    LocalMux I__13978 (
            .O(N__66557),
            .I(N__66520));
    LocalMux I__13977 (
            .O(N__66554),
            .I(N__66517));
    LocalMux I__13976 (
            .O(N__66551),
            .I(N__66514));
    LocalMux I__13975 (
            .O(N__66548),
            .I(N__66511));
    LocalMux I__13974 (
            .O(N__66545),
            .I(N__66508));
    Span4Mux_h I__13973 (
            .O(N__66542),
            .I(N__66505));
    LocalMux I__13972 (
            .O(N__66539),
            .I(N__66502));
    Span4Mux_v I__13971 (
            .O(N__66534),
            .I(N__66497));
    LocalMux I__13970 (
            .O(N__66531),
            .I(N__66497));
    InMux I__13969 (
            .O(N__66530),
            .I(N__66494));
    InMux I__13968 (
            .O(N__66529),
            .I(N__66491));
    Span4Mux_h I__13967 (
            .O(N__66526),
            .I(N__66486));
    Span4Mux_h I__13966 (
            .O(N__66523),
            .I(N__66483));
    Span4Mux_v I__13965 (
            .O(N__66520),
            .I(N__66480));
    Span4Mux_h I__13964 (
            .O(N__66517),
            .I(N__66477));
    Span4Mux_h I__13963 (
            .O(N__66514),
            .I(N__66474));
    Span4Mux_h I__13962 (
            .O(N__66511),
            .I(N__66469));
    Span4Mux_h I__13961 (
            .O(N__66508),
            .I(N__66469));
    Span4Mux_h I__13960 (
            .O(N__66505),
            .I(N__66462));
    Span4Mux_h I__13959 (
            .O(N__66502),
            .I(N__66462));
    Span4Mux_v I__13958 (
            .O(N__66497),
            .I(N__66462));
    LocalMux I__13957 (
            .O(N__66494),
            .I(N__66457));
    LocalMux I__13956 (
            .O(N__66491),
            .I(N__66457));
    InMux I__13955 (
            .O(N__66490),
            .I(N__66454));
    InMux I__13954 (
            .O(N__66489),
            .I(N__66451));
    Odrv4 I__13953 (
            .O(N__66486),
            .I(n48));
    Odrv4 I__13952 (
            .O(N__66483),
            .I(n48));
    Odrv4 I__13951 (
            .O(N__66480),
            .I(n48));
    Odrv4 I__13950 (
            .O(N__66477),
            .I(n48));
    Odrv4 I__13949 (
            .O(N__66474),
            .I(n48));
    Odrv4 I__13948 (
            .O(N__66469),
            .I(n48));
    Odrv4 I__13947 (
            .O(N__66462),
            .I(n48));
    Odrv12 I__13946 (
            .O(N__66457),
            .I(n48));
    LocalMux I__13945 (
            .O(N__66454),
            .I(n48));
    LocalMux I__13944 (
            .O(N__66451),
            .I(n48));
    InMux I__13943 (
            .O(N__66430),
            .I(N__66426));
    InMux I__13942 (
            .O(N__66429),
            .I(N__66417));
    LocalMux I__13941 (
            .O(N__66426),
            .I(N__66409));
    InMux I__13940 (
            .O(N__66425),
            .I(N__66406));
    InMux I__13939 (
            .O(N__66424),
            .I(N__66403));
    InMux I__13938 (
            .O(N__66423),
            .I(N__66399));
    InMux I__13937 (
            .O(N__66422),
            .I(N__66396));
    InMux I__13936 (
            .O(N__66421),
            .I(N__66391));
    InMux I__13935 (
            .O(N__66420),
            .I(N__66391));
    LocalMux I__13934 (
            .O(N__66417),
            .I(N__66388));
    InMux I__13933 (
            .O(N__66416),
            .I(N__66384));
    InMux I__13932 (
            .O(N__66415),
            .I(N__66381));
    InMux I__13931 (
            .O(N__66414),
            .I(N__66376));
    InMux I__13930 (
            .O(N__66413),
            .I(N__66376));
    InMux I__13929 (
            .O(N__66412),
            .I(N__66373));
    Span4Mux_v I__13928 (
            .O(N__66409),
            .I(N__66370));
    LocalMux I__13927 (
            .O(N__66406),
            .I(N__66367));
    LocalMux I__13926 (
            .O(N__66403),
            .I(N__66364));
    InMux I__13925 (
            .O(N__66402),
            .I(N__66361));
    LocalMux I__13924 (
            .O(N__66399),
            .I(N__66358));
    LocalMux I__13923 (
            .O(N__66396),
            .I(N__66355));
    LocalMux I__13922 (
            .O(N__66391),
            .I(N__66352));
    Span4Mux_v I__13921 (
            .O(N__66388),
            .I(N__66349));
    InMux I__13920 (
            .O(N__66387),
            .I(N__66345));
    LocalMux I__13919 (
            .O(N__66384),
            .I(N__66342));
    LocalMux I__13918 (
            .O(N__66381),
            .I(N__66339));
    LocalMux I__13917 (
            .O(N__66376),
            .I(N__66336));
    LocalMux I__13916 (
            .O(N__66373),
            .I(N__66333));
    Span4Mux_h I__13915 (
            .O(N__66370),
            .I(N__66328));
    Span4Mux_v I__13914 (
            .O(N__66367),
            .I(N__66328));
    Span4Mux_v I__13913 (
            .O(N__66364),
            .I(N__66325));
    LocalMux I__13912 (
            .O(N__66361),
            .I(N__66320));
    Span4Mux_v I__13911 (
            .O(N__66358),
            .I(N__66320));
    Span4Mux_h I__13910 (
            .O(N__66355),
            .I(N__66313));
    Span4Mux_v I__13909 (
            .O(N__66352),
            .I(N__66313));
    Span4Mux_h I__13908 (
            .O(N__66349),
            .I(N__66313));
    InMux I__13907 (
            .O(N__66348),
            .I(N__66310));
    LocalMux I__13906 (
            .O(N__66345),
            .I(N__66307));
    Span4Mux_h I__13905 (
            .O(N__66342),
            .I(N__66304));
    Span4Mux_v I__13904 (
            .O(N__66339),
            .I(N__66301));
    Span4Mux_v I__13903 (
            .O(N__66336),
            .I(N__66298));
    Span4Mux_v I__13902 (
            .O(N__66333),
            .I(N__66287));
    Span4Mux_h I__13901 (
            .O(N__66328),
            .I(N__66287));
    Span4Mux_v I__13900 (
            .O(N__66325),
            .I(N__66287));
    Span4Mux_v I__13899 (
            .O(N__66320),
            .I(N__66287));
    Span4Mux_h I__13898 (
            .O(N__66313),
            .I(N__66287));
    LocalMux I__13897 (
            .O(N__66310),
            .I(n59));
    Odrv12 I__13896 (
            .O(N__66307),
            .I(n59));
    Odrv4 I__13895 (
            .O(N__66304),
            .I(n59));
    Odrv4 I__13894 (
            .O(N__66301),
            .I(n59));
    Odrv4 I__13893 (
            .O(N__66298),
            .I(n59));
    Odrv4 I__13892 (
            .O(N__66287),
            .I(n59));
    InMux I__13891 (
            .O(N__66274),
            .I(N__66271));
    LocalMux I__13890 (
            .O(N__66271),
            .I(N__66263));
    InMux I__13889 (
            .O(N__66270),
            .I(N__66260));
    InMux I__13888 (
            .O(N__66269),
            .I(N__66256));
    InMux I__13887 (
            .O(N__66268),
            .I(N__66252));
    InMux I__13886 (
            .O(N__66267),
            .I(N__66247));
    InMux I__13885 (
            .O(N__66266),
            .I(N__66244));
    Span4Mux_h I__13884 (
            .O(N__66263),
            .I(N__66239));
    LocalMux I__13883 (
            .O(N__66260),
            .I(N__66239));
    InMux I__13882 (
            .O(N__66259),
            .I(N__66236));
    LocalMux I__13881 (
            .O(N__66256),
            .I(N__66233));
    InMux I__13880 (
            .O(N__66255),
            .I(N__66230));
    LocalMux I__13879 (
            .O(N__66252),
            .I(N__66227));
    InMux I__13878 (
            .O(N__66251),
            .I(N__66224));
    InMux I__13877 (
            .O(N__66250),
            .I(N__66221));
    LocalMux I__13876 (
            .O(N__66247),
            .I(N__66215));
    LocalMux I__13875 (
            .O(N__66244),
            .I(N__66212));
    Span4Mux_h I__13874 (
            .O(N__66239),
            .I(N__66209));
    LocalMux I__13873 (
            .O(N__66236),
            .I(N__66206));
    Span4Mux_h I__13872 (
            .O(N__66233),
            .I(N__66203));
    LocalMux I__13871 (
            .O(N__66230),
            .I(N__66200));
    Span4Mux_v I__13870 (
            .O(N__66227),
            .I(N__66197));
    LocalMux I__13869 (
            .O(N__66224),
            .I(N__66194));
    LocalMux I__13868 (
            .O(N__66221),
            .I(N__66191));
    InMux I__13867 (
            .O(N__66220),
            .I(N__66184));
    InMux I__13866 (
            .O(N__66219),
            .I(N__66184));
    InMux I__13865 (
            .O(N__66218),
            .I(N__66184));
    Span4Mux_v I__13864 (
            .O(N__66215),
            .I(N__66178));
    Span4Mux_h I__13863 (
            .O(N__66212),
            .I(N__66175));
    Span4Mux_v I__13862 (
            .O(N__66209),
            .I(N__66172));
    Span4Mux_v I__13861 (
            .O(N__66206),
            .I(N__66169));
    Span4Mux_v I__13860 (
            .O(N__66203),
            .I(N__66164));
    Span4Mux_h I__13859 (
            .O(N__66200),
            .I(N__66164));
    Span4Mux_v I__13858 (
            .O(N__66197),
            .I(N__66155));
    Span4Mux_h I__13857 (
            .O(N__66194),
            .I(N__66155));
    Span4Mux_v I__13856 (
            .O(N__66191),
            .I(N__66155));
    LocalMux I__13855 (
            .O(N__66184),
            .I(N__66155));
    InMux I__13854 (
            .O(N__66183),
            .I(N__66152));
    InMux I__13853 (
            .O(N__66182),
            .I(N__66147));
    InMux I__13852 (
            .O(N__66181),
            .I(N__66147));
    Odrv4 I__13851 (
            .O(N__66178),
            .I(n18));
    Odrv4 I__13850 (
            .O(N__66175),
            .I(n18));
    Odrv4 I__13849 (
            .O(N__66172),
            .I(n18));
    Odrv4 I__13848 (
            .O(N__66169),
            .I(n18));
    Odrv4 I__13847 (
            .O(N__66164),
            .I(n18));
    Odrv4 I__13846 (
            .O(N__66155),
            .I(n18));
    LocalMux I__13845 (
            .O(N__66152),
            .I(n18));
    LocalMux I__13844 (
            .O(N__66147),
            .I(n18));
    InMux I__13843 (
            .O(N__66130),
            .I(N__66127));
    LocalMux I__13842 (
            .O(N__66127),
            .I(N__66123));
    CascadeMux I__13841 (
            .O(N__66126),
            .I(N__66120));
    Span4Mux_v I__13840 (
            .O(N__66123),
            .I(N__66117));
    InMux I__13839 (
            .O(N__66120),
            .I(N__66114));
    Odrv4 I__13838 (
            .O(N__66117),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_1 ));
    LocalMux I__13837 (
            .O(N__66114),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_1 ));
    CascadeMux I__13836 (
            .O(N__66109),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11681_cascade_ ));
    CascadeMux I__13835 (
            .O(N__66106),
            .I(N__66103));
    InMux I__13834 (
            .O(N__66103),
            .I(N__66100));
    LocalMux I__13833 (
            .O(N__66100),
            .I(N__66097));
    Span4Mux_v I__13832 (
            .O(N__66097),
            .I(N__66094));
    Odrv4 I__13831 (
            .O(N__66094),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13352 ));
    CascadeMux I__13830 (
            .O(N__66091),
            .I(N__66088));
    InMux I__13829 (
            .O(N__66088),
            .I(N__66082));
    InMux I__13828 (
            .O(N__66087),
            .I(N__66082));
    LocalMux I__13827 (
            .O(N__66082),
            .I(REG_mem_19_6));
    CascadeMux I__13826 (
            .O(N__66079),
            .I(N__66076));
    InMux I__13825 (
            .O(N__66076),
            .I(N__66073));
    LocalMux I__13824 (
            .O(N__66073),
            .I(N__66069));
    InMux I__13823 (
            .O(N__66072),
            .I(N__66066));
    Odrv4 I__13822 (
            .O(N__66069),
            .I(REG_mem_10_6));
    LocalMux I__13821 (
            .O(N__66066),
            .I(REG_mem_10_6));
    InMux I__13820 (
            .O(N__66061),
            .I(N__66058));
    LocalMux I__13819 (
            .O(N__66058),
            .I(N__66054));
    InMux I__13818 (
            .O(N__66057),
            .I(N__66051));
    Odrv12 I__13817 (
            .O(N__66054),
            .I(REG_mem_11_6));
    LocalMux I__13816 (
            .O(N__66051),
            .I(REG_mem_11_6));
    InMux I__13815 (
            .O(N__66046),
            .I(N__66042));
    CascadeMux I__13814 (
            .O(N__66045),
            .I(N__66039));
    LocalMux I__13813 (
            .O(N__66042),
            .I(N__66036));
    InMux I__13812 (
            .O(N__66039),
            .I(N__66033));
    Odrv4 I__13811 (
            .O(N__66036),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_2 ));
    LocalMux I__13810 (
            .O(N__66033),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_2 ));
    InMux I__13809 (
            .O(N__66028),
            .I(N__66023));
    InMux I__13808 (
            .O(N__66027),
            .I(N__66018));
    InMux I__13807 (
            .O(N__66026),
            .I(N__66012));
    LocalMux I__13806 (
            .O(N__66023),
            .I(N__66009));
    InMux I__13805 (
            .O(N__66022),
            .I(N__66000));
    InMux I__13804 (
            .O(N__66021),
            .I(N__65997));
    LocalMux I__13803 (
            .O(N__66018),
            .I(N__65994));
    InMux I__13802 (
            .O(N__66017),
            .I(N__65990));
    InMux I__13801 (
            .O(N__66016),
            .I(N__65985));
    InMux I__13800 (
            .O(N__66015),
            .I(N__65985));
    LocalMux I__13799 (
            .O(N__66012),
            .I(N__65980));
    Span4Mux_v I__13798 (
            .O(N__66009),
            .I(N__65980));
    InMux I__13797 (
            .O(N__66008),
            .I(N__65976));
    InMux I__13796 (
            .O(N__66007),
            .I(N__65973));
    InMux I__13795 (
            .O(N__66006),
            .I(N__65970));
    InMux I__13794 (
            .O(N__66005),
            .I(N__65967));
    InMux I__13793 (
            .O(N__66004),
            .I(N__65964));
    InMux I__13792 (
            .O(N__66003),
            .I(N__65961));
    LocalMux I__13791 (
            .O(N__66000),
            .I(N__65954));
    LocalMux I__13790 (
            .O(N__65997),
            .I(N__65954));
    Span4Mux_v I__13789 (
            .O(N__65994),
            .I(N__65954));
    InMux I__13788 (
            .O(N__65993),
            .I(N__65951));
    LocalMux I__13787 (
            .O(N__65990),
            .I(N__65948));
    LocalMux I__13786 (
            .O(N__65985),
            .I(N__65943));
    Span4Mux_h I__13785 (
            .O(N__65980),
            .I(N__65943));
    InMux I__13784 (
            .O(N__65979),
            .I(N__65940));
    LocalMux I__13783 (
            .O(N__65976),
            .I(N__65935));
    LocalMux I__13782 (
            .O(N__65973),
            .I(N__65935));
    LocalMux I__13781 (
            .O(N__65970),
            .I(N__65932));
    LocalMux I__13780 (
            .O(N__65967),
            .I(N__65927));
    LocalMux I__13779 (
            .O(N__65964),
            .I(N__65927));
    LocalMux I__13778 (
            .O(N__65961),
            .I(N__65922));
    Span4Mux_v I__13777 (
            .O(N__65954),
            .I(N__65922));
    LocalMux I__13776 (
            .O(N__65951),
            .I(N__65915));
    Span4Mux_v I__13775 (
            .O(N__65948),
            .I(N__65915));
    Span4Mux_h I__13774 (
            .O(N__65943),
            .I(N__65915));
    LocalMux I__13773 (
            .O(N__65940),
            .I(n24_adj_1185));
    Odrv4 I__13772 (
            .O(N__65935),
            .I(n24_adj_1185));
    Odrv12 I__13771 (
            .O(N__65932),
            .I(n24_adj_1185));
    Odrv12 I__13770 (
            .O(N__65927),
            .I(n24_adj_1185));
    Odrv4 I__13769 (
            .O(N__65922),
            .I(n24_adj_1185));
    Odrv4 I__13768 (
            .O(N__65915),
            .I(n24_adj_1185));
    InMux I__13767 (
            .O(N__65902),
            .I(N__65898));
    InMux I__13766 (
            .O(N__65901),
            .I(N__65893));
    LocalMux I__13765 (
            .O(N__65898),
            .I(N__65889));
    InMux I__13764 (
            .O(N__65897),
            .I(N__65884));
    InMux I__13763 (
            .O(N__65896),
            .I(N__65881));
    LocalMux I__13762 (
            .O(N__65893),
            .I(N__65873));
    InMux I__13761 (
            .O(N__65892),
            .I(N__65870));
    Span4Mux_h I__13760 (
            .O(N__65889),
            .I(N__65867));
    InMux I__13759 (
            .O(N__65888),
            .I(N__65864));
    InMux I__13758 (
            .O(N__65887),
            .I(N__65861));
    LocalMux I__13757 (
            .O(N__65884),
            .I(N__65855));
    LocalMux I__13756 (
            .O(N__65881),
            .I(N__65855));
    InMux I__13755 (
            .O(N__65880),
            .I(N__65852));
    InMux I__13754 (
            .O(N__65879),
            .I(N__65849));
    InMux I__13753 (
            .O(N__65878),
            .I(N__65846));
    InMux I__13752 (
            .O(N__65877),
            .I(N__65843));
    InMux I__13751 (
            .O(N__65876),
            .I(N__65840));
    Span4Mux_h I__13750 (
            .O(N__65873),
            .I(N__65836));
    LocalMux I__13749 (
            .O(N__65870),
            .I(N__65833));
    Span4Mux_h I__13748 (
            .O(N__65867),
            .I(N__65830));
    LocalMux I__13747 (
            .O(N__65864),
            .I(N__65825));
    LocalMux I__13746 (
            .O(N__65861),
            .I(N__65825));
    InMux I__13745 (
            .O(N__65860),
            .I(N__65822));
    Span4Mux_v I__13744 (
            .O(N__65855),
            .I(N__65815));
    LocalMux I__13743 (
            .O(N__65852),
            .I(N__65815));
    LocalMux I__13742 (
            .O(N__65849),
            .I(N__65815));
    LocalMux I__13741 (
            .O(N__65846),
            .I(N__65808));
    LocalMux I__13740 (
            .O(N__65843),
            .I(N__65808));
    LocalMux I__13739 (
            .O(N__65840),
            .I(N__65808));
    InMux I__13738 (
            .O(N__65839),
            .I(N__65805));
    Span4Mux_v I__13737 (
            .O(N__65836),
            .I(N__65798));
    Span4Mux_v I__13736 (
            .O(N__65833),
            .I(N__65798));
    Span4Mux_h I__13735 (
            .O(N__65830),
            .I(N__65793));
    Span4Mux_v I__13734 (
            .O(N__65825),
            .I(N__65793));
    LocalMux I__13733 (
            .O(N__65822),
            .I(N__65790));
    Span4Mux_v I__13732 (
            .O(N__65815),
            .I(N__65783));
    Span4Mux_h I__13731 (
            .O(N__65808),
            .I(N__65783));
    LocalMux I__13730 (
            .O(N__65805),
            .I(N__65783));
    InMux I__13729 (
            .O(N__65804),
            .I(N__65780));
    InMux I__13728 (
            .O(N__65803),
            .I(N__65777));
    Odrv4 I__13727 (
            .O(N__65798),
            .I(n25));
    Odrv4 I__13726 (
            .O(N__65793),
            .I(n25));
    Odrv4 I__13725 (
            .O(N__65790),
            .I(n25));
    Odrv4 I__13724 (
            .O(N__65783),
            .I(n25));
    LocalMux I__13723 (
            .O(N__65780),
            .I(n25));
    LocalMux I__13722 (
            .O(N__65777),
            .I(n25));
    InMux I__13721 (
            .O(N__65764),
            .I(N__65761));
    LocalMux I__13720 (
            .O(N__65761),
            .I(N__65758));
    Span12Mux_h I__13719 (
            .O(N__65758),
            .I(N__65755));
    Odrv12 I__13718 (
            .O(N__65755),
            .I(FIFO_D8_c_8));
    InMux I__13717 (
            .O(N__65752),
            .I(N__65749));
    LocalMux I__13716 (
            .O(N__65749),
            .I(N__65746));
    Span4Mux_h I__13715 (
            .O(N__65746),
            .I(N__65743));
    Span4Mux_v I__13714 (
            .O(N__65743),
            .I(N__65740));
    Odrv4 I__13713 (
            .O(N__65740),
            .I(FIFO_D2_c_2));
    InMux I__13712 (
            .O(N__65737),
            .I(N__65734));
    LocalMux I__13711 (
            .O(N__65734),
            .I(\usb3_if_inst.usb3_data_in_latched_2 ));
    InMux I__13710 (
            .O(N__65731),
            .I(N__65728));
    LocalMux I__13709 (
            .O(N__65728),
            .I(N__65725));
    Span4Mux_h I__13708 (
            .O(N__65725),
            .I(N__65722));
    Span4Mux_v I__13707 (
            .O(N__65722),
            .I(N__65719));
    Odrv4 I__13706 (
            .O(N__65719),
            .I(FIFO_D1_c_1));
    InMux I__13705 (
            .O(N__65716),
            .I(N__65713));
    LocalMux I__13704 (
            .O(N__65713),
            .I(\usb3_if_inst.usb3_data_in_latched_1 ));
    InMux I__13703 (
            .O(N__65710),
            .I(N__65707));
    LocalMux I__13702 (
            .O(N__65707),
            .I(\usb3_if_inst.usb3_data_in_latched_8 ));
    InMux I__13701 (
            .O(N__65704),
            .I(N__65698));
    InMux I__13700 (
            .O(N__65703),
            .I(N__65698));
    LocalMux I__13699 (
            .O(N__65698),
            .I(REG_mem_17_6));
    CascadeMux I__13698 (
            .O(N__65695),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13658_cascade_ ));
    InMux I__13697 (
            .O(N__65692),
            .I(N__65689));
    LocalMux I__13696 (
            .O(N__65689),
            .I(N__65682));
    InMux I__13695 (
            .O(N__65688),
            .I(N__65679));
    InMux I__13694 (
            .O(N__65687),
            .I(N__65673));
    InMux I__13693 (
            .O(N__65686),
            .I(N__65670));
    InMux I__13692 (
            .O(N__65685),
            .I(N__65666));
    Span4Mux_h I__13691 (
            .O(N__65682),
            .I(N__65659));
    LocalMux I__13690 (
            .O(N__65679),
            .I(N__65659));
    InMux I__13689 (
            .O(N__65678),
            .I(N__65654));
    InMux I__13688 (
            .O(N__65677),
            .I(N__65654));
    InMux I__13687 (
            .O(N__65676),
            .I(N__65651));
    LocalMux I__13686 (
            .O(N__65673),
            .I(N__65647));
    LocalMux I__13685 (
            .O(N__65670),
            .I(N__65644));
    InMux I__13684 (
            .O(N__65669),
            .I(N__65641));
    LocalMux I__13683 (
            .O(N__65666),
            .I(N__65637));
    InMux I__13682 (
            .O(N__65665),
            .I(N__65634));
    InMux I__13681 (
            .O(N__65664),
            .I(N__65631));
    Span4Mux_h I__13680 (
            .O(N__65659),
            .I(N__65628));
    LocalMux I__13679 (
            .O(N__65654),
            .I(N__65625));
    LocalMux I__13678 (
            .O(N__65651),
            .I(N__65622));
    InMux I__13677 (
            .O(N__65650),
            .I(N__65619));
    Span4Mux_v I__13676 (
            .O(N__65647),
            .I(N__65615));
    Span4Mux_v I__13675 (
            .O(N__65644),
            .I(N__65612));
    LocalMux I__13674 (
            .O(N__65641),
            .I(N__65609));
    InMux I__13673 (
            .O(N__65640),
            .I(N__65606));
    Span4Mux_h I__13672 (
            .O(N__65637),
            .I(N__65601));
    LocalMux I__13671 (
            .O(N__65634),
            .I(N__65596));
    LocalMux I__13670 (
            .O(N__65631),
            .I(N__65596));
    Span4Mux_v I__13669 (
            .O(N__65628),
            .I(N__65587));
    Span4Mux_v I__13668 (
            .O(N__65625),
            .I(N__65587));
    Span4Mux_h I__13667 (
            .O(N__65622),
            .I(N__65587));
    LocalMux I__13666 (
            .O(N__65619),
            .I(N__65587));
    InMux I__13665 (
            .O(N__65618),
            .I(N__65584));
    Span4Mux_h I__13664 (
            .O(N__65615),
            .I(N__65575));
    Span4Mux_h I__13663 (
            .O(N__65612),
            .I(N__65575));
    Span4Mux_v I__13662 (
            .O(N__65609),
            .I(N__65575));
    LocalMux I__13661 (
            .O(N__65606),
            .I(N__65575));
    InMux I__13660 (
            .O(N__65605),
            .I(N__65572));
    InMux I__13659 (
            .O(N__65604),
            .I(N__65569));
    Odrv4 I__13658 (
            .O(N__65601),
            .I(n49));
    Odrv12 I__13657 (
            .O(N__65596),
            .I(n49));
    Odrv4 I__13656 (
            .O(N__65587),
            .I(n49));
    LocalMux I__13655 (
            .O(N__65584),
            .I(n49));
    Odrv4 I__13654 (
            .O(N__65575),
            .I(n49));
    LocalMux I__13653 (
            .O(N__65572),
            .I(n49));
    LocalMux I__13652 (
            .O(N__65569),
            .I(n49));
    InMux I__13651 (
            .O(N__65554),
            .I(N__65548));
    InMux I__13650 (
            .O(N__65553),
            .I(N__65548));
    LocalMux I__13649 (
            .O(N__65548),
            .I(REG_mem_16_6));
    InMux I__13648 (
            .O(N__65545),
            .I(N__65539));
    InMux I__13647 (
            .O(N__65544),
            .I(N__65539));
    LocalMux I__13646 (
            .O(N__65539),
            .I(REG_mem_18_6));
    InMux I__13645 (
            .O(N__65536),
            .I(N__65533));
    LocalMux I__13644 (
            .O(N__65533),
            .I(N__65529));
    InMux I__13643 (
            .O(N__65532),
            .I(N__65526));
    Span4Mux_v I__13642 (
            .O(N__65529),
            .I(N__65523));
    LocalMux I__13641 (
            .O(N__65526),
            .I(N__65520));
    Odrv4 I__13640 (
            .O(N__65523),
            .I(fifo_data_out_3));
    Odrv12 I__13639 (
            .O(N__65520),
            .I(fifo_data_out_3));
    IoInMux I__13638 (
            .O(N__65515),
            .I(N__65512));
    LocalMux I__13637 (
            .O(N__65512),
            .I(N__65509));
    IoSpan4Mux I__13636 (
            .O(N__65509),
            .I(N__65505));
    IoInMux I__13635 (
            .O(N__65508),
            .I(N__65502));
    IoSpan4Mux I__13634 (
            .O(N__65505),
            .I(N__65499));
    LocalMux I__13633 (
            .O(N__65502),
            .I(N__65496));
    Span4Mux_s3_v I__13632 (
            .O(N__65499),
            .I(N__65493));
    Span4Mux_s3_v I__13631 (
            .O(N__65496),
            .I(N__65490));
    Span4Mux_v I__13630 (
            .O(N__65493),
            .I(N__65485));
    Span4Mux_v I__13629 (
            .O(N__65490),
            .I(N__65485));
    Odrv4 I__13628 (
            .O(N__65485),
            .I(DATA19_c));
    InMux I__13627 (
            .O(N__65482),
            .I(N__65479));
    LocalMux I__13626 (
            .O(N__65479),
            .I(N__65476));
    Span4Mux_v I__13625 (
            .O(N__65476),
            .I(N__65472));
    InMux I__13624 (
            .O(N__65475),
            .I(N__65469));
    Odrv4 I__13623 (
            .O(N__65472),
            .I(fifo_data_out_2));
    LocalMux I__13622 (
            .O(N__65469),
            .I(fifo_data_out_2));
    IoInMux I__13621 (
            .O(N__65464),
            .I(N__65461));
    LocalMux I__13620 (
            .O(N__65461),
            .I(N__65458));
    IoSpan4Mux I__13619 (
            .O(N__65458),
            .I(N__65454));
    IoInMux I__13618 (
            .O(N__65457),
            .I(N__65451));
    IoSpan4Mux I__13617 (
            .O(N__65454),
            .I(N__65448));
    LocalMux I__13616 (
            .O(N__65451),
            .I(N__65445));
    Span4Mux_s3_v I__13615 (
            .O(N__65448),
            .I(N__65442));
    Span4Mux_s3_v I__13614 (
            .O(N__65445),
            .I(N__65439));
    Span4Mux_h I__13613 (
            .O(N__65442),
            .I(N__65434));
    Span4Mux_h I__13612 (
            .O(N__65439),
            .I(N__65434));
    Span4Mux_v I__13611 (
            .O(N__65434),
            .I(N__65431));
    Odrv4 I__13610 (
            .O(N__65431),
            .I(DATA18_c));
    InMux I__13609 (
            .O(N__65428),
            .I(N__65425));
    LocalMux I__13608 (
            .O(N__65425),
            .I(N__65421));
    InMux I__13607 (
            .O(N__65424),
            .I(N__65418));
    Odrv4 I__13606 (
            .O(N__65421),
            .I(fifo_data_out_1));
    LocalMux I__13605 (
            .O(N__65418),
            .I(fifo_data_out_1));
    IoInMux I__13604 (
            .O(N__65413),
            .I(N__65409));
    IoInMux I__13603 (
            .O(N__65412),
            .I(N__65406));
    LocalMux I__13602 (
            .O(N__65409),
            .I(N__65403));
    LocalMux I__13601 (
            .O(N__65406),
            .I(N__65400));
    Span4Mux_s2_v I__13600 (
            .O(N__65403),
            .I(N__65397));
    Span12Mux_s7_v I__13599 (
            .O(N__65400),
            .I(N__65394));
    Sp12to4 I__13598 (
            .O(N__65397),
            .I(N__65391));
    Span12Mux_h I__13597 (
            .O(N__65394),
            .I(N__65388));
    Span12Mux_s11_h I__13596 (
            .O(N__65391),
            .I(N__65385));
    Odrv12 I__13595 (
            .O(N__65388),
            .I(DATA17_c));
    Odrv12 I__13594 (
            .O(N__65385),
            .I(DATA17_c));
    InMux I__13593 (
            .O(N__65380),
            .I(N__65377));
    LocalMux I__13592 (
            .O(N__65377),
            .I(N__65374));
    Span12Mux_h I__13591 (
            .O(N__65374),
            .I(N__65370));
    InMux I__13590 (
            .O(N__65373),
            .I(N__65367));
    Odrv12 I__13589 (
            .O(N__65370),
            .I(fifo_data_out_5));
    LocalMux I__13588 (
            .O(N__65367),
            .I(fifo_data_out_5));
    IoInMux I__13587 (
            .O(N__65362),
            .I(N__65359));
    LocalMux I__13586 (
            .O(N__65359),
            .I(N__65355));
    IoInMux I__13585 (
            .O(N__65358),
            .I(N__65352));
    IoSpan4Mux I__13584 (
            .O(N__65355),
            .I(N__65349));
    LocalMux I__13583 (
            .O(N__65352),
            .I(N__65346));
    IoSpan4Mux I__13582 (
            .O(N__65349),
            .I(N__65343));
    Span4Mux_s3_v I__13581 (
            .O(N__65346),
            .I(N__65340));
    Span4Mux_s3_v I__13580 (
            .O(N__65343),
            .I(N__65335));
    Span4Mux_h I__13579 (
            .O(N__65340),
            .I(N__65335));
    Span4Mux_v I__13578 (
            .O(N__65335),
            .I(N__65332));
    Odrv4 I__13577 (
            .O(N__65332),
            .I(DATA5_c));
    InMux I__13576 (
            .O(N__65329),
            .I(N__65325));
    InMux I__13575 (
            .O(N__65328),
            .I(N__65322));
    LocalMux I__13574 (
            .O(N__65325),
            .I(fifo_data_out_6));
    LocalMux I__13573 (
            .O(N__65322),
            .I(fifo_data_out_6));
    IoInMux I__13572 (
            .O(N__65317),
            .I(N__65314));
    LocalMux I__13571 (
            .O(N__65314),
            .I(N__65310));
    IoInMux I__13570 (
            .O(N__65313),
            .I(N__65307));
    Span4Mux_s3_v I__13569 (
            .O(N__65310),
            .I(N__65304));
    LocalMux I__13568 (
            .O(N__65307),
            .I(N__65301));
    Span4Mux_h I__13567 (
            .O(N__65304),
            .I(N__65298));
    Span12Mux_s7_v I__13566 (
            .O(N__65301),
            .I(N__65295));
    Span4Mux_v I__13565 (
            .O(N__65298),
            .I(N__65292));
    Odrv12 I__13564 (
            .O(N__65295),
            .I(DATA6_c));
    Odrv4 I__13563 (
            .O(N__65292),
            .I(DATA6_c));
    CascadeMux I__13562 (
            .O(N__65287),
            .I(wr_addr_p1_w_2_cascade_));
    InMux I__13561 (
            .O(N__65284),
            .I(N__65278));
    InMux I__13560 (
            .O(N__65283),
            .I(N__65278));
    LocalMux I__13559 (
            .O(N__65278),
            .I(N__65275));
    Span4Mux_v I__13558 (
            .O(N__65275),
            .I(N__65272));
    Span4Mux_h I__13557 (
            .O(N__65272),
            .I(N__65269));
    Sp12to4 I__13556 (
            .O(N__65269),
            .I(N__65266));
    Span12Mux_h I__13555 (
            .O(N__65266),
            .I(N__65263));
    Odrv12 I__13554 (
            .O(N__65263),
            .I(rx_shift_reg_0));
    InMux I__13553 (
            .O(N__65260),
            .I(N__65251));
    InMux I__13552 (
            .O(N__65259),
            .I(N__65251));
    InMux I__13551 (
            .O(N__65258),
            .I(N__65251));
    LocalMux I__13550 (
            .O(N__65251),
            .I(rx_shift_reg_1));
    InMux I__13549 (
            .O(N__65248),
            .I(N__65243));
    InMux I__13548 (
            .O(N__65247),
            .I(N__65240));
    InMux I__13547 (
            .O(N__65246),
            .I(N__65237));
    LocalMux I__13546 (
            .O(N__65243),
            .I(rx_shift_reg_2));
    LocalMux I__13545 (
            .O(N__65240),
            .I(rx_shift_reg_2));
    LocalMux I__13544 (
            .O(N__65237),
            .I(rx_shift_reg_2));
    CEMux I__13543 (
            .O(N__65230),
            .I(N__65227));
    LocalMux I__13542 (
            .O(N__65227),
            .I(N__65217));
    InMux I__13541 (
            .O(N__65226),
            .I(N__65210));
    InMux I__13540 (
            .O(N__65225),
            .I(N__65210));
    InMux I__13539 (
            .O(N__65224),
            .I(N__65210));
    InMux I__13538 (
            .O(N__65223),
            .I(N__65207));
    InMux I__13537 (
            .O(N__65222),
            .I(N__65202));
    InMux I__13536 (
            .O(N__65221),
            .I(N__65202));
    InMux I__13535 (
            .O(N__65220),
            .I(N__65199));
    Span4Mux_s0_v I__13534 (
            .O(N__65217),
            .I(N__65196));
    LocalMux I__13533 (
            .O(N__65210),
            .I(N__65191));
    LocalMux I__13532 (
            .O(N__65207),
            .I(N__65191));
    LocalMux I__13531 (
            .O(N__65202),
            .I(N__65186));
    LocalMux I__13530 (
            .O(N__65199),
            .I(N__65186));
    Sp12to4 I__13529 (
            .O(N__65196),
            .I(N__65183));
    Span4Mux_v I__13528 (
            .O(N__65191),
            .I(N__65180));
    Span4Mux_h I__13527 (
            .O(N__65186),
            .I(N__65177));
    Span12Mux_h I__13526 (
            .O(N__65183),
            .I(N__65174));
    Span4Mux_h I__13525 (
            .O(N__65180),
            .I(N__65171));
    Span4Mux_h I__13524 (
            .O(N__65177),
            .I(N__65168));
    Odrv12 I__13523 (
            .O(N__65174),
            .I(n4093));
    Odrv4 I__13522 (
            .O(N__65171),
            .I(n4093));
    Odrv4 I__13521 (
            .O(N__65168),
            .I(n4093));
    InMux I__13520 (
            .O(N__65161),
            .I(N__65151));
    InMux I__13519 (
            .O(N__65160),
            .I(N__65148));
    InMux I__13518 (
            .O(N__65159),
            .I(N__65141));
    InMux I__13517 (
            .O(N__65158),
            .I(N__65141));
    InMux I__13516 (
            .O(N__65157),
            .I(N__65141));
    InMux I__13515 (
            .O(N__65156),
            .I(N__65134));
    InMux I__13514 (
            .O(N__65155),
            .I(N__65134));
    InMux I__13513 (
            .O(N__65154),
            .I(N__65134));
    LocalMux I__13512 (
            .O(N__65151),
            .I(N__65131));
    LocalMux I__13511 (
            .O(N__65148),
            .I(N__65124));
    LocalMux I__13510 (
            .O(N__65141),
            .I(N__65124));
    LocalMux I__13509 (
            .O(N__65134),
            .I(N__65124));
    Span4Mux_v I__13508 (
            .O(N__65131),
            .I(N__65121));
    Span4Mux_v I__13507 (
            .O(N__65124),
            .I(N__65118));
    Odrv4 I__13506 (
            .O(N__65121),
            .I(n3204));
    Odrv4 I__13505 (
            .O(N__65118),
            .I(n3204));
    InMux I__13504 (
            .O(N__65113),
            .I(N__65110));
    LocalMux I__13503 (
            .O(N__65110),
            .I(N__65105));
    InMux I__13502 (
            .O(N__65109),
            .I(N__65100));
    InMux I__13501 (
            .O(N__65108),
            .I(N__65100));
    Odrv4 I__13500 (
            .O(N__65105),
            .I(rx_shift_reg_3));
    LocalMux I__13499 (
            .O(N__65100),
            .I(rx_shift_reg_3));
    InMux I__13498 (
            .O(N__65095),
            .I(N__65092));
    LocalMux I__13497 (
            .O(N__65092),
            .I(N__65089));
    Span12Mux_s11_v I__13496 (
            .O(N__65089),
            .I(N__65085));
    InMux I__13495 (
            .O(N__65088),
            .I(N__65082));
    Odrv12 I__13494 (
            .O(N__65085),
            .I(fifo_data_out_8));
    LocalMux I__13493 (
            .O(N__65082),
            .I(fifo_data_out_8));
    IoInMux I__13492 (
            .O(N__65077),
            .I(N__65074));
    LocalMux I__13491 (
            .O(N__65074),
            .I(N__65070));
    IoInMux I__13490 (
            .O(N__65073),
            .I(N__65067));
    Span4Mux_s3_h I__13489 (
            .O(N__65070),
            .I(N__65064));
    LocalMux I__13488 (
            .O(N__65067),
            .I(N__65061));
    Span4Mux_h I__13487 (
            .O(N__65064),
            .I(N__65056));
    Span4Mux_s3_v I__13486 (
            .O(N__65061),
            .I(N__65056));
    Span4Mux_v I__13485 (
            .O(N__65056),
            .I(N__65053));
    Odrv4 I__13484 (
            .O(N__65053),
            .I(DATA8_c));
    InMux I__13483 (
            .O(N__65050),
            .I(N__65047));
    LocalMux I__13482 (
            .O(N__65047),
            .I(N__65044));
    Span4Mux_v I__13481 (
            .O(N__65044),
            .I(N__65040));
    CascadeMux I__13480 (
            .O(N__65043),
            .I(N__65037));
    Span4Mux_v I__13479 (
            .O(N__65040),
            .I(N__65034));
    InMux I__13478 (
            .O(N__65037),
            .I(N__65031));
    Odrv4 I__13477 (
            .O(N__65034),
            .I(fifo_data_out_7));
    LocalMux I__13476 (
            .O(N__65031),
            .I(fifo_data_out_7));
    IoInMux I__13475 (
            .O(N__65026),
            .I(N__65023));
    LocalMux I__13474 (
            .O(N__65023),
            .I(N__65020));
    IoSpan4Mux I__13473 (
            .O(N__65020),
            .I(N__65016));
    IoInMux I__13472 (
            .O(N__65019),
            .I(N__65013));
    IoSpan4Mux I__13471 (
            .O(N__65016),
            .I(N__65008));
    LocalMux I__13470 (
            .O(N__65013),
            .I(N__65008));
    IoSpan4Mux I__13469 (
            .O(N__65008),
            .I(N__65005));
    Span4Mux_s3_v I__13468 (
            .O(N__65005),
            .I(N__65002));
    Span4Mux_v I__13467 (
            .O(N__65002),
            .I(N__64999));
    Odrv4 I__13466 (
            .O(N__64999),
            .I(DATA7_c));
    InMux I__13465 (
            .O(N__64996),
            .I(N__64993));
    LocalMux I__13464 (
            .O(N__64993),
            .I(N__64990));
    Span4Mux_v I__13463 (
            .O(N__64990),
            .I(N__64986));
    CascadeMux I__13462 (
            .O(N__64989),
            .I(N__64983));
    Span4Mux_h I__13461 (
            .O(N__64986),
            .I(N__64980));
    InMux I__13460 (
            .O(N__64983),
            .I(N__64977));
    Odrv4 I__13459 (
            .O(N__64980),
            .I(fifo_data_out_4));
    LocalMux I__13458 (
            .O(N__64977),
            .I(fifo_data_out_4));
    IoInMux I__13457 (
            .O(N__64972),
            .I(N__64969));
    LocalMux I__13456 (
            .O(N__64969),
            .I(N__64965));
    IoInMux I__13455 (
            .O(N__64968),
            .I(N__64962));
    IoSpan4Mux I__13454 (
            .O(N__64965),
            .I(N__64957));
    LocalMux I__13453 (
            .O(N__64962),
            .I(N__64957));
    IoSpan4Mux I__13452 (
            .O(N__64957),
            .I(N__64954));
    Span4Mux_s3_v I__13451 (
            .O(N__64954),
            .I(N__64951));
    Span4Mux_v I__13450 (
            .O(N__64951),
            .I(N__64948));
    Odrv4 I__13449 (
            .O(N__64948),
            .I(DATA20_c));
    InMux I__13448 (
            .O(N__64945),
            .I(N__64942));
    LocalMux I__13447 (
            .O(N__64942),
            .I(N__64937));
    InMux I__13446 (
            .O(N__64941),
            .I(N__64932));
    InMux I__13445 (
            .O(N__64940),
            .I(N__64932));
    Odrv4 I__13444 (
            .O(N__64937),
            .I(rx_shift_reg_4));
    LocalMux I__13443 (
            .O(N__64932),
            .I(rx_shift_reg_4));
    CascadeMux I__13442 (
            .O(N__64927),
            .I(N__64924));
    InMux I__13441 (
            .O(N__64924),
            .I(N__64921));
    LocalMux I__13440 (
            .O(N__64921),
            .I(N__64917));
    InMux I__13439 (
            .O(N__64920),
            .I(N__64914));
    Odrv4 I__13438 (
            .O(N__64917),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7 ));
    LocalMux I__13437 (
            .O(N__64914),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7 ));
    InMux I__13436 (
            .O(N__64909),
            .I(N__64906));
    LocalMux I__13435 (
            .O(N__64906),
            .I(N__64902));
    InMux I__13434 (
            .O(N__64905),
            .I(N__64899));
    Odrv4 I__13433 (
            .O(N__64902),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_7 ));
    LocalMux I__13432 (
            .O(N__64899),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_7 ));
    InMux I__13431 (
            .O(N__64894),
            .I(N__64888));
    InMux I__13430 (
            .O(N__64893),
            .I(N__64888));
    LocalMux I__13429 (
            .O(N__64888),
            .I(rx_shift_reg_7));
    InMux I__13428 (
            .O(N__64885),
            .I(N__64878));
    InMux I__13427 (
            .O(N__64884),
            .I(N__64878));
    InMux I__13426 (
            .O(N__64883),
            .I(N__64875));
    LocalMux I__13425 (
            .O(N__64878),
            .I(rx_shift_reg_6));
    LocalMux I__13424 (
            .O(N__64875),
            .I(rx_shift_reg_6));
    CascadeMux I__13423 (
            .O(N__64870),
            .I(N__64866));
    CascadeMux I__13422 (
            .O(N__64869),
            .I(N__64861));
    InMux I__13421 (
            .O(N__64866),
            .I(N__64851));
    InMux I__13420 (
            .O(N__64865),
            .I(N__64851));
    InMux I__13419 (
            .O(N__64864),
            .I(N__64851));
    InMux I__13418 (
            .O(N__64861),
            .I(N__64851));
    InMux I__13417 (
            .O(N__64860),
            .I(N__64848));
    LocalMux I__13416 (
            .O(N__64851),
            .I(rx_buf_byte_6));
    LocalMux I__13415 (
            .O(N__64848),
            .I(rx_buf_byte_6));
    InMux I__13414 (
            .O(N__64843),
            .I(N__64840));
    LocalMux I__13413 (
            .O(N__64840),
            .I(N__64836));
    InMux I__13412 (
            .O(N__64839),
            .I(N__64833));
    Span4Mux_h I__13411 (
            .O(N__64836),
            .I(N__64830));
    LocalMux I__13410 (
            .O(N__64833),
            .I(\usb3_if_inst.num_lines_clocked_out_5 ));
    Odrv4 I__13409 (
            .O(N__64830),
            .I(\usb3_if_inst.num_lines_clocked_out_5 ));
    InMux I__13408 (
            .O(N__64825),
            .I(N__64822));
    LocalMux I__13407 (
            .O(N__64822),
            .I(N__64818));
    InMux I__13406 (
            .O(N__64821),
            .I(N__64815));
    Span4Mux_h I__13405 (
            .O(N__64818),
            .I(N__64812));
    LocalMux I__13404 (
            .O(N__64815),
            .I(\usb3_if_inst.num_lines_clocked_out_1 ));
    Odrv4 I__13403 (
            .O(N__64812),
            .I(\usb3_if_inst.num_lines_clocked_out_1 ));
    InMux I__13402 (
            .O(N__64807),
            .I(N__64804));
    LocalMux I__13401 (
            .O(N__64804),
            .I(\usb3_if_inst.n16 ));
    CascadeMux I__13400 (
            .O(N__64801),
            .I(N__64798));
    InMux I__13399 (
            .O(N__64798),
            .I(N__64794));
    InMux I__13398 (
            .O(N__64797),
            .I(N__64791));
    LocalMux I__13397 (
            .O(N__64794),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_6 ));
    LocalMux I__13396 (
            .O(N__64791),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_6 ));
    CascadeMux I__13395 (
            .O(N__64786),
            .I(N__64783));
    InMux I__13394 (
            .O(N__64783),
            .I(N__64780));
    LocalMux I__13393 (
            .O(N__64780),
            .I(N__64776));
    InMux I__13392 (
            .O(N__64779),
            .I(N__64773));
    Odrv4 I__13391 (
            .O(N__64776),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6 ));
    LocalMux I__13390 (
            .O(N__64773),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6 ));
    InMux I__13389 (
            .O(N__64768),
            .I(N__64764));
    InMux I__13388 (
            .O(N__64767),
            .I(N__64761));
    LocalMux I__13387 (
            .O(N__64764),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6 ));
    LocalMux I__13386 (
            .O(N__64761),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6 ));
    CascadeMux I__13385 (
            .O(N__64756),
            .I(N__64752));
    InMux I__13384 (
            .O(N__64755),
            .I(N__64749));
    InMux I__13383 (
            .O(N__64752),
            .I(N__64746));
    LocalMux I__13382 (
            .O(N__64749),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_6 ));
    LocalMux I__13381 (
            .O(N__64746),
            .I(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_6 ));
    InMux I__13380 (
            .O(N__64741),
            .I(N__64732));
    InMux I__13379 (
            .O(N__64740),
            .I(N__64732));
    InMux I__13378 (
            .O(N__64739),
            .I(N__64732));
    LocalMux I__13377 (
            .O(N__64732),
            .I(rx_shift_reg_5));
    CascadeMux I__13376 (
            .O(N__64729),
            .I(N__64725));
    InMux I__13375 (
            .O(N__64728),
            .I(N__64720));
    InMux I__13374 (
            .O(N__64725),
            .I(N__64720));
    LocalMux I__13373 (
            .O(N__64720),
            .I(N__64717));
    Odrv12 I__13372 (
            .O(N__64717),
            .I(dc32_fifo_almost_empty));
    CascadeMux I__13371 (
            .O(N__64714),
            .I(N__64710));
    InMux I__13370 (
            .O(N__64713),
            .I(N__64702));
    InMux I__13369 (
            .O(N__64710),
            .I(N__64702));
    InMux I__13368 (
            .O(N__64709),
            .I(N__64702));
    LocalMux I__13367 (
            .O(N__64702),
            .I(\bluejay_data_inst.n714 ));
    InMux I__13366 (
            .O(N__64699),
            .I(N__64695));
    InMux I__13365 (
            .O(N__64698),
            .I(N__64692));
    LocalMux I__13364 (
            .O(N__64695),
            .I(\bluejay_data_inst.n717 ));
    LocalMux I__13363 (
            .O(N__64692),
            .I(\bluejay_data_inst.n717 ));
    CascadeMux I__13362 (
            .O(N__64687),
            .I(\bluejay_data_inst.n108_cascade_ ));
    CascadeMux I__13361 (
            .O(N__64684),
            .I(\bluejay_data_inst.n4062_cascade_ ));
    InMux I__13360 (
            .O(N__64681),
            .I(N__64678));
    LocalMux I__13359 (
            .O(N__64678),
            .I(N__64675));
    Span4Mux_v I__13358 (
            .O(N__64675),
            .I(N__64671));
    InMux I__13357 (
            .O(N__64674),
            .I(N__64668));
    Odrv4 I__13356 (
            .O(N__64671),
            .I(\bluejay_data_inst.n108 ));
    LocalMux I__13355 (
            .O(N__64668),
            .I(\bluejay_data_inst.n108 ));
    SRMux I__13354 (
            .O(N__64663),
            .I(N__64660));
    LocalMux I__13353 (
            .O(N__64660),
            .I(N__64657));
    Span4Mux_v I__13352 (
            .O(N__64657),
            .I(N__64653));
    SRMux I__13351 (
            .O(N__64656),
            .I(N__64650));
    Span4Mux_v I__13350 (
            .O(N__64653),
            .I(N__64647));
    LocalMux I__13349 (
            .O(N__64650),
            .I(N__64644));
    Odrv4 I__13348 (
            .O(N__64647),
            .I(\bluejay_data_inst.n4519 ));
    Odrv12 I__13347 (
            .O(N__64644),
            .I(\bluejay_data_inst.n4519 ));
    InMux I__13346 (
            .O(N__64639),
            .I(N__64636));
    LocalMux I__13345 (
            .O(N__64636),
            .I(\tx_fifo.lscc_fifo_inst.n13952 ));
    InMux I__13344 (
            .O(N__64633),
            .I(N__64630));
    LocalMux I__13343 (
            .O(N__64630),
            .I(N__64626));
    InMux I__13342 (
            .O(N__64629),
            .I(N__64623));
    Span4Mux_v I__13341 (
            .O(N__64626),
            .I(N__64620));
    LocalMux I__13340 (
            .O(N__64623),
            .I(\usb3_if_inst.num_lines_clocked_out_3 ));
    Odrv4 I__13339 (
            .O(N__64620),
            .I(\usb3_if_inst.num_lines_clocked_out_3 ));
    InMux I__13338 (
            .O(N__64615),
            .I(N__64611));
    CascadeMux I__13337 (
            .O(N__64614),
            .I(N__64608));
    LocalMux I__13336 (
            .O(N__64611),
            .I(N__64605));
    InMux I__13335 (
            .O(N__64608),
            .I(N__64602));
    Span4Mux_h I__13334 (
            .O(N__64605),
            .I(N__64599));
    LocalMux I__13333 (
            .O(N__64602),
            .I(\usb3_if_inst.num_lines_clocked_out_6 ));
    Odrv4 I__13332 (
            .O(N__64599),
            .I(\usb3_if_inst.num_lines_clocked_out_6 ));
    CascadeMux I__13331 (
            .O(N__64594),
            .I(N__64591));
    InMux I__13330 (
            .O(N__64591),
            .I(N__64588));
    LocalMux I__13329 (
            .O(N__64588),
            .I(N__64584));
    InMux I__13328 (
            .O(N__64587),
            .I(N__64581));
    Span4Mux_h I__13327 (
            .O(N__64584),
            .I(N__64578));
    LocalMux I__13326 (
            .O(N__64581),
            .I(\usb3_if_inst.num_lines_clocked_out_10 ));
    Odrv4 I__13325 (
            .O(N__64578),
            .I(\usb3_if_inst.num_lines_clocked_out_10 ));
    InMux I__13324 (
            .O(N__64573),
            .I(N__64570));
    LocalMux I__13323 (
            .O(N__64570),
            .I(N__64567));
    Span12Mux_v I__13322 (
            .O(N__64567),
            .I(N__64564));
    Odrv12 I__13321 (
            .O(N__64564),
            .I(\usb3_if_inst.n18 ));
    InMux I__13320 (
            .O(N__64561),
            .I(N__64558));
    LocalMux I__13319 (
            .O(N__64558),
            .I(N__64554));
    InMux I__13318 (
            .O(N__64557),
            .I(N__64551));
    Span4Mux_h I__13317 (
            .O(N__64554),
            .I(N__64548));
    LocalMux I__13316 (
            .O(N__64551),
            .I(\usb3_if_inst.num_lines_clocked_out_8 ));
    Odrv4 I__13315 (
            .O(N__64548),
            .I(\usb3_if_inst.num_lines_clocked_out_8 ));
    InMux I__13314 (
            .O(N__64543),
            .I(N__64539));
    CascadeMux I__13313 (
            .O(N__64542),
            .I(N__64536));
    LocalMux I__13312 (
            .O(N__64539),
            .I(N__64533));
    InMux I__13311 (
            .O(N__64536),
            .I(N__64530));
    Span4Mux_h I__13310 (
            .O(N__64533),
            .I(N__64527));
    LocalMux I__13309 (
            .O(N__64530),
            .I(\usb3_if_inst.num_lines_clocked_out_4 ));
    Odrv4 I__13308 (
            .O(N__64527),
            .I(\usb3_if_inst.num_lines_clocked_out_4 ));
    CascadeMux I__13307 (
            .O(N__64522),
            .I(\usb3_if_inst.n20_cascade_ ));
    InMux I__13306 (
            .O(N__64519),
            .I(N__64511));
    InMux I__13305 (
            .O(N__64518),
            .I(N__64511));
    InMux I__13304 (
            .O(N__64517),
            .I(N__64508));
    InMux I__13303 (
            .O(N__64516),
            .I(N__64505));
    LocalMux I__13302 (
            .O(N__64511),
            .I(N__64498));
    LocalMux I__13301 (
            .O(N__64508),
            .I(N__64498));
    LocalMux I__13300 (
            .O(N__64505),
            .I(N__64498));
    Span4Mux_h I__13299 (
            .O(N__64498),
            .I(N__64495));
    Odrv4 I__13298 (
            .O(N__64495),
            .I(\usb3_if_inst.n21 ));
    CascadeMux I__13297 (
            .O(N__64492),
            .I(\bluejay_data_inst.n8_cascade_ ));
    InMux I__13296 (
            .O(N__64489),
            .I(N__64486));
    LocalMux I__13295 (
            .O(N__64486),
            .I(\bluejay_data_inst.n12_adj_1179 ));
    InMux I__13294 (
            .O(N__64483),
            .I(N__64474));
    InMux I__13293 (
            .O(N__64482),
            .I(N__64474));
    InMux I__13292 (
            .O(N__64481),
            .I(N__64474));
    LocalMux I__13291 (
            .O(N__64474),
            .I(N__64470));
    InMux I__13290 (
            .O(N__64473),
            .I(N__64467));
    Odrv4 I__13289 (
            .O(N__64470),
            .I(\bluejay_data_inst.state_timeout_counter_0 ));
    LocalMux I__13288 (
            .O(N__64467),
            .I(\bluejay_data_inst.state_timeout_counter_0 ));
    CascadeMux I__13287 (
            .O(N__64462),
            .I(N__64457));
    InMux I__13286 (
            .O(N__64461),
            .I(N__64449));
    InMux I__13285 (
            .O(N__64460),
            .I(N__64449));
    InMux I__13284 (
            .O(N__64457),
            .I(N__64449));
    InMux I__13283 (
            .O(N__64456),
            .I(N__64446));
    LocalMux I__13282 (
            .O(N__64449),
            .I(\bluejay_data_inst.state_timeout_counter_4 ));
    LocalMux I__13281 (
            .O(N__64446),
            .I(\bluejay_data_inst.state_timeout_counter_4 ));
    InMux I__13280 (
            .O(N__64441),
            .I(N__64436));
    InMux I__13279 (
            .O(N__64440),
            .I(N__64431));
    InMux I__13278 (
            .O(N__64439),
            .I(N__64431));
    LocalMux I__13277 (
            .O(N__64436),
            .I(N__64426));
    LocalMux I__13276 (
            .O(N__64431),
            .I(N__64426));
    Odrv4 I__13275 (
            .O(N__64426),
            .I(\bluejay_data_inst.n12 ));
    CascadeMux I__13274 (
            .O(N__64423),
            .I(n7_cascade_));
    InMux I__13273 (
            .O(N__64420),
            .I(N__64404));
    InMux I__13272 (
            .O(N__64419),
            .I(N__64404));
    InMux I__13271 (
            .O(N__64418),
            .I(N__64404));
    InMux I__13270 (
            .O(N__64417),
            .I(N__64404));
    InMux I__13269 (
            .O(N__64416),
            .I(N__64404));
    InMux I__13268 (
            .O(N__64415),
            .I(N__64401));
    LocalMux I__13267 (
            .O(N__64404),
            .I(state_timeout_counter_3));
    LocalMux I__13266 (
            .O(N__64401),
            .I(state_timeout_counter_3));
    CascadeMux I__13265 (
            .O(N__64396),
            .I(N__64392));
    InMux I__13264 (
            .O(N__64395),
            .I(N__64389));
    InMux I__13263 (
            .O(N__64392),
            .I(N__64386));
    LocalMux I__13262 (
            .O(N__64389),
            .I(n7));
    LocalMux I__13261 (
            .O(N__64386),
            .I(n7));
    InMux I__13260 (
            .O(N__64381),
            .I(N__64378));
    LocalMux I__13259 (
            .O(N__64378),
            .I(\bluejay_data_inst.n10745 ));
    IoInMux I__13258 (
            .O(N__64375),
            .I(N__64372));
    LocalMux I__13257 (
            .O(N__64372),
            .I(N__64369));
    Span4Mux_s1_v I__13256 (
            .O(N__64369),
            .I(N__64364));
    CascadeMux I__13255 (
            .O(N__64368),
            .I(N__64355));
    CascadeMux I__13254 (
            .O(N__64367),
            .I(N__64350));
    Span4Mux_h I__13253 (
            .O(N__64364),
            .I(N__64346));
    InMux I__13252 (
            .O(N__64363),
            .I(N__64341));
    InMux I__13251 (
            .O(N__64362),
            .I(N__64330));
    InMux I__13250 (
            .O(N__64361),
            .I(N__64330));
    InMux I__13249 (
            .O(N__64360),
            .I(N__64330));
    InMux I__13248 (
            .O(N__64359),
            .I(N__64330));
    InMux I__13247 (
            .O(N__64358),
            .I(N__64330));
    InMux I__13246 (
            .O(N__64355),
            .I(N__64325));
    InMux I__13245 (
            .O(N__64354),
            .I(N__64325));
    InMux I__13244 (
            .O(N__64353),
            .I(N__64322));
    InMux I__13243 (
            .O(N__64350),
            .I(N__64317));
    InMux I__13242 (
            .O(N__64349),
            .I(N__64317));
    Sp12to4 I__13241 (
            .O(N__64346),
            .I(N__64314));
    InMux I__13240 (
            .O(N__64345),
            .I(N__64308));
    InMux I__13239 (
            .O(N__64344),
            .I(N__64308));
    LocalMux I__13238 (
            .O(N__64341),
            .I(N__64303));
    LocalMux I__13237 (
            .O(N__64330),
            .I(N__64303));
    LocalMux I__13236 (
            .O(N__64325),
            .I(N__64300));
    LocalMux I__13235 (
            .O(N__64322),
            .I(N__64297));
    LocalMux I__13234 (
            .O(N__64317),
            .I(N__64294));
    Span12Mux_h I__13233 (
            .O(N__64314),
            .I(N__64288));
    InMux I__13232 (
            .O(N__64313),
            .I(N__64285));
    LocalMux I__13231 (
            .O(N__64308),
            .I(N__64280));
    Span4Mux_h I__13230 (
            .O(N__64303),
            .I(N__64280));
    Span4Mux_h I__13229 (
            .O(N__64300),
            .I(N__64275));
    Span4Mux_h I__13228 (
            .O(N__64297),
            .I(N__64275));
    Sp12to4 I__13227 (
            .O(N__64294),
            .I(N__64272));
    InMux I__13226 (
            .O(N__64293),
            .I(N__64265));
    InMux I__13225 (
            .O(N__64292),
            .I(N__64265));
    InMux I__13224 (
            .O(N__64291),
            .I(N__64265));
    Span12Mux_v I__13223 (
            .O(N__64288),
            .I(N__64260));
    LocalMux I__13222 (
            .O(N__64285),
            .I(N__64260));
    Span4Mux_h I__13221 (
            .O(N__64280),
            .I(N__64257));
    Span4Mux_h I__13220 (
            .O(N__64275),
            .I(N__64254));
    Odrv12 I__13219 (
            .O(N__64272),
            .I(DEBUG_9_c));
    LocalMux I__13218 (
            .O(N__64265),
            .I(DEBUG_9_c));
    Odrv12 I__13217 (
            .O(N__64260),
            .I(DEBUG_9_c));
    Odrv4 I__13216 (
            .O(N__64257),
            .I(DEBUG_9_c));
    Odrv4 I__13215 (
            .O(N__64254),
            .I(DEBUG_9_c));
    CascadeMux I__13214 (
            .O(N__64243),
            .I(N__64239));
    InMux I__13213 (
            .O(N__64242),
            .I(N__64234));
    InMux I__13212 (
            .O(N__64239),
            .I(N__64234));
    LocalMux I__13211 (
            .O(N__64234),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_4 ));
    CascadeMux I__13210 (
            .O(N__64231),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13418_cascade_ ));
    InMux I__13209 (
            .O(N__64228),
            .I(N__64225));
    LocalMux I__13208 (
            .O(N__64225),
            .I(N__64222));
    Span4Mux_h I__13207 (
            .O(N__64222),
            .I(N__64219));
    Odrv4 I__13206 (
            .O(N__64219),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13421 ));
    CascadeMux I__13205 (
            .O(N__64216),
            .I(N__64212));
    InMux I__13204 (
            .O(N__64215),
            .I(N__64207));
    InMux I__13203 (
            .O(N__64212),
            .I(N__64207));
    LocalMux I__13202 (
            .O(N__64207),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_4 ));
    CascadeMux I__13201 (
            .O(N__64204),
            .I(N__64200));
    CascadeMux I__13200 (
            .O(N__64203),
            .I(N__64197));
    InMux I__13199 (
            .O(N__64200),
            .I(N__64194));
    InMux I__13198 (
            .O(N__64197),
            .I(N__64191));
    LocalMux I__13197 (
            .O(N__64194),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_4 ));
    LocalMux I__13196 (
            .O(N__64191),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_4 ));
    CascadeMux I__13195 (
            .O(N__64186),
            .I(N__64182));
    InMux I__13194 (
            .O(N__64185),
            .I(N__64177));
    InMux I__13193 (
            .O(N__64182),
            .I(N__64177));
    LocalMux I__13192 (
            .O(N__64177),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_4 ));
    CascadeMux I__13191 (
            .O(N__64174),
            .I(N__64170));
    InMux I__13190 (
            .O(N__64173),
            .I(N__64165));
    InMux I__13189 (
            .O(N__64170),
            .I(N__64165));
    LocalMux I__13188 (
            .O(N__64165),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_4 ));
    InMux I__13187 (
            .O(N__64162),
            .I(N__64159));
    LocalMux I__13186 (
            .O(N__64159),
            .I(N__64156));
    Span4Mux_h I__13185 (
            .O(N__64156),
            .I(N__64153));
    Odrv4 I__13184 (
            .O(N__64153),
            .I(\usb3_if_inst.n534 ));
    CascadeMux I__13183 (
            .O(N__64150),
            .I(N__64146));
    InMux I__13182 (
            .O(N__64149),
            .I(N__64138));
    InMux I__13181 (
            .O(N__64146),
            .I(N__64135));
    InMux I__13180 (
            .O(N__64145),
            .I(N__64130));
    InMux I__13179 (
            .O(N__64144),
            .I(N__64130));
    InMux I__13178 (
            .O(N__64143),
            .I(N__64126));
    InMux I__13177 (
            .O(N__64142),
            .I(N__64121));
    InMux I__13176 (
            .O(N__64141),
            .I(N__64121));
    LocalMux I__13175 (
            .O(N__64138),
            .I(N__64118));
    LocalMux I__13174 (
            .O(N__64135),
            .I(N__64113));
    LocalMux I__13173 (
            .O(N__64130),
            .I(N__64113));
    CascadeMux I__13172 (
            .O(N__64129),
            .I(N__64110));
    LocalMux I__13171 (
            .O(N__64126),
            .I(N__64105));
    LocalMux I__13170 (
            .O(N__64121),
            .I(N__64098));
    Span4Mux_v I__13169 (
            .O(N__64118),
            .I(N__64098));
    Span4Mux_h I__13168 (
            .O(N__64113),
            .I(N__64098));
    InMux I__13167 (
            .O(N__64110),
            .I(N__64091));
    InMux I__13166 (
            .O(N__64109),
            .I(N__64091));
    InMux I__13165 (
            .O(N__64108),
            .I(N__64091));
    Span4Mux_v I__13164 (
            .O(N__64105),
            .I(N__64086));
    Span4Mux_h I__13163 (
            .O(N__64098),
            .I(N__64086));
    LocalMux I__13162 (
            .O(N__64091),
            .I(\usb3_if_inst.n550 ));
    Odrv4 I__13161 (
            .O(N__64086),
            .I(\usb3_if_inst.n550 ));
    InMux I__13160 (
            .O(N__64081),
            .I(N__64077));
    CascadeMux I__13159 (
            .O(N__64080),
            .I(N__64073));
    LocalMux I__13158 (
            .O(N__64077),
            .I(N__64065));
    InMux I__13157 (
            .O(N__64076),
            .I(N__64062));
    InMux I__13156 (
            .O(N__64073),
            .I(N__64057));
    InMux I__13155 (
            .O(N__64072),
            .I(N__64057));
    InMux I__13154 (
            .O(N__64071),
            .I(N__64054));
    InMux I__13153 (
            .O(N__64070),
            .I(N__64049));
    InMux I__13152 (
            .O(N__64069),
            .I(N__64049));
    InMux I__13151 (
            .O(N__64068),
            .I(N__64046));
    Span4Mux_h I__13150 (
            .O(N__64065),
            .I(N__64043));
    LocalMux I__13149 (
            .O(N__64062),
            .I(N__64034));
    LocalMux I__13148 (
            .O(N__64057),
            .I(N__64034));
    LocalMux I__13147 (
            .O(N__64054),
            .I(N__64034));
    LocalMux I__13146 (
            .O(N__64049),
            .I(N__64034));
    LocalMux I__13145 (
            .O(N__64046),
            .I(\usb3_if_inst.n553 ));
    Odrv4 I__13144 (
            .O(N__64043),
            .I(\usb3_if_inst.n553 ));
    Odrv12 I__13143 (
            .O(N__64034),
            .I(\usb3_if_inst.n553 ));
    InMux I__13142 (
            .O(N__64027),
            .I(N__64024));
    LocalMux I__13141 (
            .O(N__64024),
            .I(N__64021));
    Span4Mux_v I__13140 (
            .O(N__64021),
            .I(N__64018));
    Span4Mux_h I__13139 (
            .O(N__64018),
            .I(N__64015));
    Odrv4 I__13138 (
            .O(N__64015),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11755 ));
    InMux I__13137 (
            .O(N__64012),
            .I(N__64002));
    InMux I__13136 (
            .O(N__64011),
            .I(N__63999));
    InMux I__13135 (
            .O(N__64010),
            .I(N__63995));
    InMux I__13134 (
            .O(N__64009),
            .I(N__63992));
    InMux I__13133 (
            .O(N__64008),
            .I(N__63989));
    InMux I__13132 (
            .O(N__64007),
            .I(N__63986));
    InMux I__13131 (
            .O(N__64006),
            .I(N__63981));
    InMux I__13130 (
            .O(N__64005),
            .I(N__63977));
    LocalMux I__13129 (
            .O(N__64002),
            .I(N__63974));
    LocalMux I__13128 (
            .O(N__63999),
            .I(N__63971));
    InMux I__13127 (
            .O(N__63998),
            .I(N__63968));
    LocalMux I__13126 (
            .O(N__63995),
            .I(N__63965));
    LocalMux I__13125 (
            .O(N__63992),
            .I(N__63962));
    LocalMux I__13124 (
            .O(N__63989),
            .I(N__63959));
    LocalMux I__13123 (
            .O(N__63986),
            .I(N__63956));
    InMux I__13122 (
            .O(N__63985),
            .I(N__63949));
    InMux I__13121 (
            .O(N__63984),
            .I(N__63946));
    LocalMux I__13120 (
            .O(N__63981),
            .I(N__63943));
    InMux I__13119 (
            .O(N__63980),
            .I(N__63940));
    LocalMux I__13118 (
            .O(N__63977),
            .I(N__63937));
    Span4Mux_v I__13117 (
            .O(N__63974),
            .I(N__63934));
    Span4Mux_h I__13116 (
            .O(N__63971),
            .I(N__63931));
    LocalMux I__13115 (
            .O(N__63968),
            .I(N__63928));
    Span4Mux_v I__13114 (
            .O(N__63965),
            .I(N__63925));
    Span4Mux_v I__13113 (
            .O(N__63962),
            .I(N__63922));
    Span4Mux_h I__13112 (
            .O(N__63959),
            .I(N__63917));
    Span4Mux_v I__13111 (
            .O(N__63956),
            .I(N__63917));
    InMux I__13110 (
            .O(N__63955),
            .I(N__63912));
    InMux I__13109 (
            .O(N__63954),
            .I(N__63912));
    InMux I__13108 (
            .O(N__63953),
            .I(N__63909));
    InMux I__13107 (
            .O(N__63952),
            .I(N__63906));
    LocalMux I__13106 (
            .O(N__63949),
            .I(N__63901));
    LocalMux I__13105 (
            .O(N__63946),
            .I(N__63901));
    Span4Mux_v I__13104 (
            .O(N__63943),
            .I(N__63898));
    LocalMux I__13103 (
            .O(N__63940),
            .I(N__63895));
    Span4Mux_h I__13102 (
            .O(N__63937),
            .I(N__63890));
    Span4Mux_h I__13101 (
            .O(N__63934),
            .I(N__63890));
    Span4Mux_h I__13100 (
            .O(N__63931),
            .I(N__63887));
    Span4Mux_h I__13099 (
            .O(N__63928),
            .I(N__63878));
    Span4Mux_h I__13098 (
            .O(N__63925),
            .I(N__63878));
    Span4Mux_h I__13097 (
            .O(N__63922),
            .I(N__63878));
    Span4Mux_h I__13096 (
            .O(N__63917),
            .I(N__63878));
    LocalMux I__13095 (
            .O(N__63912),
            .I(n50));
    LocalMux I__13094 (
            .O(N__63909),
            .I(n50));
    LocalMux I__13093 (
            .O(N__63906),
            .I(n50));
    Odrv12 I__13092 (
            .O(N__63901),
            .I(n50));
    Odrv4 I__13091 (
            .O(N__63898),
            .I(n50));
    Odrv12 I__13090 (
            .O(N__63895),
            .I(n50));
    Odrv4 I__13089 (
            .O(N__63890),
            .I(n50));
    Odrv4 I__13088 (
            .O(N__63887),
            .I(n50));
    Odrv4 I__13087 (
            .O(N__63878),
            .I(n50));
    CascadeMux I__13086 (
            .O(N__63859),
            .I(N__63856));
    InMux I__13085 (
            .O(N__63856),
            .I(N__63852));
    InMux I__13084 (
            .O(N__63855),
            .I(N__63849));
    LocalMux I__13083 (
            .O(N__63852),
            .I(N__63846));
    LocalMux I__13082 (
            .O(N__63849),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_4 ));
    Odrv4 I__13081 (
            .O(N__63846),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_4 ));
    CascadeMux I__13080 (
            .O(N__63841),
            .I(N__63837));
    InMux I__13079 (
            .O(N__63840),
            .I(N__63832));
    InMux I__13078 (
            .O(N__63837),
            .I(N__63832));
    LocalMux I__13077 (
            .O(N__63832),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_4 ));
    InMux I__13076 (
            .O(N__63829),
            .I(N__63826));
    LocalMux I__13075 (
            .O(N__63826),
            .I(N__63823));
    Span4Mux_v I__13074 (
            .O(N__63823),
            .I(N__63820));
    Odrv4 I__13073 (
            .O(N__63820),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11756 ));
    InMux I__13072 (
            .O(N__63817),
            .I(N__63811));
    InMux I__13071 (
            .O(N__63816),
            .I(N__63811));
    LocalMux I__13070 (
            .O(N__63811),
            .I(REG_mem_23_4));
    CascadeMux I__13069 (
            .O(N__63808),
            .I(N__63804));
    InMux I__13068 (
            .O(N__63807),
            .I(N__63801));
    InMux I__13067 (
            .O(N__63804),
            .I(N__63798));
    LocalMux I__13066 (
            .O(N__63801),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_4 ));
    LocalMux I__13065 (
            .O(N__63798),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_4 ));
    InMux I__13064 (
            .O(N__63793),
            .I(N__63790));
    LocalMux I__13063 (
            .O(N__63790),
            .I(N__63787));
    Span4Mux_v I__13062 (
            .O(N__63787),
            .I(N__63783));
    InMux I__13061 (
            .O(N__63786),
            .I(N__63780));
    Odrv4 I__13060 (
            .O(N__63783),
            .I(REG_mem_13_2));
    LocalMux I__13059 (
            .O(N__63780),
            .I(REG_mem_13_2));
    InMux I__13058 (
            .O(N__63775),
            .I(N__63772));
    LocalMux I__13057 (
            .O(N__63772),
            .I(N__63769));
    Span4Mux_h I__13056 (
            .O(N__63769),
            .I(N__63766));
    Sp12to4 I__13055 (
            .O(N__63766),
            .I(N__63762));
    InMux I__13054 (
            .O(N__63765),
            .I(N__63759));
    Odrv12 I__13053 (
            .O(N__63762),
            .I(REG_mem_39_8));
    LocalMux I__13052 (
            .O(N__63759),
            .I(REG_mem_39_8));
    InMux I__13051 (
            .O(N__63754),
            .I(N__63751));
    LocalMux I__13050 (
            .O(N__63751),
            .I(N__63747));
    CascadeMux I__13049 (
            .O(N__63750),
            .I(N__63744));
    Span4Mux_v I__13048 (
            .O(N__63747),
            .I(N__63741));
    InMux I__13047 (
            .O(N__63744),
            .I(N__63738));
    Odrv4 I__13046 (
            .O(N__63741),
            .I(REG_mem_38_8));
    LocalMux I__13045 (
            .O(N__63738),
            .I(REG_mem_38_8));
    InMux I__13044 (
            .O(N__63733),
            .I(N__63730));
    LocalMux I__13043 (
            .O(N__63730),
            .I(N__63724));
    InMux I__13042 (
            .O(N__63729),
            .I(N__63721));
    InMux I__13041 (
            .O(N__63728),
            .I(N__63718));
    InMux I__13040 (
            .O(N__63727),
            .I(N__63714));
    Span4Mux_v I__13039 (
            .O(N__63724),
            .I(N__63708));
    LocalMux I__13038 (
            .O(N__63721),
            .I(N__63705));
    LocalMux I__13037 (
            .O(N__63718),
            .I(N__63702));
    InMux I__13036 (
            .O(N__63717),
            .I(N__63699));
    LocalMux I__13035 (
            .O(N__63714),
            .I(N__63696));
    InMux I__13034 (
            .O(N__63713),
            .I(N__63693));
    InMux I__13033 (
            .O(N__63712),
            .I(N__63690));
    InMux I__13032 (
            .O(N__63711),
            .I(N__63686));
    Span4Mux_h I__13031 (
            .O(N__63708),
            .I(N__63681));
    Span4Mux_h I__13030 (
            .O(N__63705),
            .I(N__63678));
    Span4Mux_v I__13029 (
            .O(N__63702),
            .I(N__63673));
    LocalMux I__13028 (
            .O(N__63699),
            .I(N__63670));
    Span4Mux_h I__13027 (
            .O(N__63696),
            .I(N__63667));
    LocalMux I__13026 (
            .O(N__63693),
            .I(N__63664));
    LocalMux I__13025 (
            .O(N__63690),
            .I(N__63661));
    InMux I__13024 (
            .O(N__63689),
            .I(N__63658));
    LocalMux I__13023 (
            .O(N__63686),
            .I(N__63655));
    InMux I__13022 (
            .O(N__63685),
            .I(N__63650));
    InMux I__13021 (
            .O(N__63684),
            .I(N__63650));
    Span4Mux_h I__13020 (
            .O(N__63681),
            .I(N__63643));
    Span4Mux_h I__13019 (
            .O(N__63678),
            .I(N__63643));
    InMux I__13018 (
            .O(N__63677),
            .I(N__63640));
    InMux I__13017 (
            .O(N__63676),
            .I(N__63637));
    Span4Mux_h I__13016 (
            .O(N__63673),
            .I(N__63631));
    Span4Mux_h I__13015 (
            .O(N__63670),
            .I(N__63631));
    Span4Mux_h I__13014 (
            .O(N__63667),
            .I(N__63624));
    Span4Mux_v I__13013 (
            .O(N__63664),
            .I(N__63624));
    Span4Mux_v I__13012 (
            .O(N__63661),
            .I(N__63624));
    LocalMux I__13011 (
            .O(N__63658),
            .I(N__63621));
    Span4Mux_h I__13010 (
            .O(N__63655),
            .I(N__63616));
    LocalMux I__13009 (
            .O(N__63650),
            .I(N__63616));
    InMux I__13008 (
            .O(N__63649),
            .I(N__63613));
    InMux I__13007 (
            .O(N__63648),
            .I(N__63610));
    Sp12to4 I__13006 (
            .O(N__63643),
            .I(N__63603));
    LocalMux I__13005 (
            .O(N__63640),
            .I(N__63603));
    LocalMux I__13004 (
            .O(N__63637),
            .I(N__63603));
    InMux I__13003 (
            .O(N__63636),
            .I(N__63600));
    Odrv4 I__13002 (
            .O(N__63631),
            .I(n28));
    Odrv4 I__13001 (
            .O(N__63624),
            .I(n28));
    Odrv12 I__13000 (
            .O(N__63621),
            .I(n28));
    Odrv4 I__12999 (
            .O(N__63616),
            .I(n28));
    LocalMux I__12998 (
            .O(N__63613),
            .I(n28));
    LocalMux I__12997 (
            .O(N__63610),
            .I(n28));
    Odrv12 I__12996 (
            .O(N__63603),
            .I(n28));
    LocalMux I__12995 (
            .O(N__63600),
            .I(n28));
    InMux I__12994 (
            .O(N__63583),
            .I(N__63580));
    LocalMux I__12993 (
            .O(N__63580),
            .I(N__63576));
    InMux I__12992 (
            .O(N__63579),
            .I(N__63573));
    Odrv4 I__12991 (
            .O(N__63576),
            .I(REG_mem_13_4));
    LocalMux I__12990 (
            .O(N__63573),
            .I(REG_mem_13_4));
    InMux I__12989 (
            .O(N__63568),
            .I(N__63565));
    LocalMux I__12988 (
            .O(N__63565),
            .I(N__63562));
    Span4Mux_v I__12987 (
            .O(N__63562),
            .I(N__63558));
    CascadeMux I__12986 (
            .O(N__63561),
            .I(N__63555));
    Span4Mux_v I__12985 (
            .O(N__63558),
            .I(N__63552));
    InMux I__12984 (
            .O(N__63555),
            .I(N__63549));
    Odrv4 I__12983 (
            .O(N__63552),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_7 ));
    LocalMux I__12982 (
            .O(N__63549),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_7 ));
    InMux I__12981 (
            .O(N__63544),
            .I(N__63522));
    InMux I__12980 (
            .O(N__63543),
            .I(N__63513));
    InMux I__12979 (
            .O(N__63542),
            .I(N__63513));
    InMux I__12978 (
            .O(N__63541),
            .I(N__63513));
    InMux I__12977 (
            .O(N__63540),
            .I(N__63513));
    InMux I__12976 (
            .O(N__63539),
            .I(N__63510));
    CascadeMux I__12975 (
            .O(N__63538),
            .I(N__63506));
    InMux I__12974 (
            .O(N__63537),
            .I(N__63500));
    CascadeMux I__12973 (
            .O(N__63536),
            .I(N__63497));
    CascadeMux I__12972 (
            .O(N__63535),
            .I(N__63494));
    InMux I__12971 (
            .O(N__63534),
            .I(N__63487));
    InMux I__12970 (
            .O(N__63533),
            .I(N__63482));
    InMux I__12969 (
            .O(N__63532),
            .I(N__63477));
    InMux I__12968 (
            .O(N__63531),
            .I(N__63477));
    CascadeMux I__12967 (
            .O(N__63530),
            .I(N__63474));
    InMux I__12966 (
            .O(N__63529),
            .I(N__63466));
    InMux I__12965 (
            .O(N__63528),
            .I(N__63466));
    InMux I__12964 (
            .O(N__63527),
            .I(N__63463));
    InMux I__12963 (
            .O(N__63526),
            .I(N__63458));
    InMux I__12962 (
            .O(N__63525),
            .I(N__63458));
    LocalMux I__12961 (
            .O(N__63522),
            .I(N__63455));
    LocalMux I__12960 (
            .O(N__63513),
            .I(N__63450));
    LocalMux I__12959 (
            .O(N__63510),
            .I(N__63450));
    InMux I__12958 (
            .O(N__63509),
            .I(N__63442));
    InMux I__12957 (
            .O(N__63506),
            .I(N__63433));
    InMux I__12956 (
            .O(N__63505),
            .I(N__63430));
    InMux I__12955 (
            .O(N__63504),
            .I(N__63425));
    InMux I__12954 (
            .O(N__63503),
            .I(N__63425));
    LocalMux I__12953 (
            .O(N__63500),
            .I(N__63422));
    InMux I__12952 (
            .O(N__63497),
            .I(N__63417));
    InMux I__12951 (
            .O(N__63494),
            .I(N__63417));
    InMux I__12950 (
            .O(N__63493),
            .I(N__63410));
    InMux I__12949 (
            .O(N__63492),
            .I(N__63410));
    InMux I__12948 (
            .O(N__63491),
            .I(N__63410));
    InMux I__12947 (
            .O(N__63490),
            .I(N__63407));
    LocalMux I__12946 (
            .O(N__63487),
            .I(N__63404));
    InMux I__12945 (
            .O(N__63486),
            .I(N__63399));
    InMux I__12944 (
            .O(N__63485),
            .I(N__63399));
    LocalMux I__12943 (
            .O(N__63482),
            .I(N__63393));
    LocalMux I__12942 (
            .O(N__63477),
            .I(N__63393));
    InMux I__12941 (
            .O(N__63474),
            .I(N__63386));
    InMux I__12940 (
            .O(N__63473),
            .I(N__63386));
    InMux I__12939 (
            .O(N__63472),
            .I(N__63386));
    InMux I__12938 (
            .O(N__63471),
            .I(N__63383));
    LocalMux I__12937 (
            .O(N__63466),
            .I(N__63366));
    LocalMux I__12936 (
            .O(N__63463),
            .I(N__63366));
    LocalMux I__12935 (
            .O(N__63458),
            .I(N__63366));
    Span4Mux_h I__12934 (
            .O(N__63455),
            .I(N__63366));
    Span4Mux_v I__12933 (
            .O(N__63450),
            .I(N__63366));
    InMux I__12932 (
            .O(N__63449),
            .I(N__63363));
    InMux I__12931 (
            .O(N__63448),
            .I(N__63354));
    InMux I__12930 (
            .O(N__63447),
            .I(N__63354));
    InMux I__12929 (
            .O(N__63446),
            .I(N__63354));
    InMux I__12928 (
            .O(N__63445),
            .I(N__63354));
    LocalMux I__12927 (
            .O(N__63442),
            .I(N__63350));
    CascadeMux I__12926 (
            .O(N__63441),
            .I(N__63347));
    CascadeMux I__12925 (
            .O(N__63440),
            .I(N__63344));
    InMux I__12924 (
            .O(N__63439),
            .I(N__63333));
    InMux I__12923 (
            .O(N__63438),
            .I(N__63333));
    InMux I__12922 (
            .O(N__63437),
            .I(N__63328));
    InMux I__12921 (
            .O(N__63436),
            .I(N__63328));
    LocalMux I__12920 (
            .O(N__63433),
            .I(N__63325));
    LocalMux I__12919 (
            .O(N__63430),
            .I(N__63322));
    LocalMux I__12918 (
            .O(N__63425),
            .I(N__63313));
    Span4Mux_h I__12917 (
            .O(N__63422),
            .I(N__63313));
    LocalMux I__12916 (
            .O(N__63417),
            .I(N__63313));
    LocalMux I__12915 (
            .O(N__63410),
            .I(N__63313));
    LocalMux I__12914 (
            .O(N__63407),
            .I(N__63308));
    Span4Mux_h I__12913 (
            .O(N__63404),
            .I(N__63303));
    LocalMux I__12912 (
            .O(N__63399),
            .I(N__63303));
    InMux I__12911 (
            .O(N__63398),
            .I(N__63300));
    Span4Mux_h I__12910 (
            .O(N__63393),
            .I(N__63297));
    LocalMux I__12909 (
            .O(N__63386),
            .I(N__63294));
    LocalMux I__12908 (
            .O(N__63383),
            .I(N__63291));
    InMux I__12907 (
            .O(N__63382),
            .I(N__63288));
    InMux I__12906 (
            .O(N__63381),
            .I(N__63283));
    InMux I__12905 (
            .O(N__63380),
            .I(N__63283));
    CascadeMux I__12904 (
            .O(N__63379),
            .I(N__63280));
    CascadeMux I__12903 (
            .O(N__63378),
            .I(N__63277));
    InMux I__12902 (
            .O(N__63377),
            .I(N__63273));
    Span4Mux_v I__12901 (
            .O(N__63366),
            .I(N__63268));
    LocalMux I__12900 (
            .O(N__63363),
            .I(N__63268));
    LocalMux I__12899 (
            .O(N__63354),
            .I(N__63265));
    InMux I__12898 (
            .O(N__63353),
            .I(N__63262));
    Span4Mux_h I__12897 (
            .O(N__63350),
            .I(N__63259));
    InMux I__12896 (
            .O(N__63347),
            .I(N__63247));
    InMux I__12895 (
            .O(N__63344),
            .I(N__63247));
    InMux I__12894 (
            .O(N__63343),
            .I(N__63247));
    InMux I__12893 (
            .O(N__63342),
            .I(N__63247));
    InMux I__12892 (
            .O(N__63341),
            .I(N__63247));
    InMux I__12891 (
            .O(N__63340),
            .I(N__63242));
    InMux I__12890 (
            .O(N__63339),
            .I(N__63242));
    InMux I__12889 (
            .O(N__63338),
            .I(N__63239));
    LocalMux I__12888 (
            .O(N__63333),
            .I(N__63234));
    LocalMux I__12887 (
            .O(N__63328),
            .I(N__63234));
    Span4Mux_h I__12886 (
            .O(N__63325),
            .I(N__63231));
    Span4Mux_v I__12885 (
            .O(N__63322),
            .I(N__63227));
    Span4Mux_v I__12884 (
            .O(N__63313),
            .I(N__63224));
    InMux I__12883 (
            .O(N__63312),
            .I(N__63221));
    InMux I__12882 (
            .O(N__63311),
            .I(N__63218));
    Span4Mux_h I__12881 (
            .O(N__63308),
            .I(N__63215));
    Span4Mux_h I__12880 (
            .O(N__63303),
            .I(N__63212));
    LocalMux I__12879 (
            .O(N__63300),
            .I(N__63209));
    Span4Mux_h I__12878 (
            .O(N__63297),
            .I(N__63204));
    Span4Mux_h I__12877 (
            .O(N__63294),
            .I(N__63204));
    Span4Mux_v I__12876 (
            .O(N__63291),
            .I(N__63199));
    LocalMux I__12875 (
            .O(N__63288),
            .I(N__63199));
    LocalMux I__12874 (
            .O(N__63283),
            .I(N__63196));
    InMux I__12873 (
            .O(N__63280),
            .I(N__63189));
    InMux I__12872 (
            .O(N__63277),
            .I(N__63189));
    InMux I__12871 (
            .O(N__63276),
            .I(N__63189));
    LocalMux I__12870 (
            .O(N__63273),
            .I(N__63182));
    Span4Mux_v I__12869 (
            .O(N__63268),
            .I(N__63182));
    Span4Mux_v I__12868 (
            .O(N__63265),
            .I(N__63182));
    LocalMux I__12867 (
            .O(N__63262),
            .I(N__63177));
    Span4Mux_h I__12866 (
            .O(N__63259),
            .I(N__63177));
    InMux I__12865 (
            .O(N__63258),
            .I(N__63174));
    LocalMux I__12864 (
            .O(N__63247),
            .I(N__63169));
    LocalMux I__12863 (
            .O(N__63242),
            .I(N__63169));
    LocalMux I__12862 (
            .O(N__63239),
            .I(N__63164));
    Span4Mux_h I__12861 (
            .O(N__63234),
            .I(N__63164));
    Span4Mux_h I__12860 (
            .O(N__63231),
            .I(N__63160));
    InMux I__12859 (
            .O(N__63230),
            .I(N__63157));
    Span4Mux_h I__12858 (
            .O(N__63227),
            .I(N__63154));
    Sp12to4 I__12857 (
            .O(N__63224),
            .I(N__63151));
    LocalMux I__12856 (
            .O(N__63221),
            .I(N__63148));
    LocalMux I__12855 (
            .O(N__63218),
            .I(N__63135));
    Span4Mux_h I__12854 (
            .O(N__63215),
            .I(N__63135));
    Span4Mux_h I__12853 (
            .O(N__63212),
            .I(N__63135));
    Span4Mux_h I__12852 (
            .O(N__63209),
            .I(N__63135));
    Span4Mux_v I__12851 (
            .O(N__63204),
            .I(N__63135));
    Span4Mux_h I__12850 (
            .O(N__63199),
            .I(N__63135));
    Span4Mux_v I__12849 (
            .O(N__63196),
            .I(N__63126));
    LocalMux I__12848 (
            .O(N__63189),
            .I(N__63126));
    Span4Mux_h I__12847 (
            .O(N__63182),
            .I(N__63126));
    Span4Mux_v I__12846 (
            .O(N__63177),
            .I(N__63126));
    LocalMux I__12845 (
            .O(N__63174),
            .I(N__63119));
    Span4Mux_v I__12844 (
            .O(N__63169),
            .I(N__63119));
    Span4Mux_h I__12843 (
            .O(N__63164),
            .I(N__63119));
    InMux I__12842 (
            .O(N__63163),
            .I(N__63116));
    Sp12to4 I__12841 (
            .O(N__63160),
            .I(N__63103));
    LocalMux I__12840 (
            .O(N__63157),
            .I(N__63103));
    Sp12to4 I__12839 (
            .O(N__63154),
            .I(N__63103));
    Span12Mux_s9_h I__12838 (
            .O(N__63151),
            .I(N__63103));
    Span12Mux_v I__12837 (
            .O(N__63148),
            .I(N__63103));
    Sp12to4 I__12836 (
            .O(N__63135),
            .I(N__63103));
    Span4Mux_v I__12835 (
            .O(N__63126),
            .I(N__63100));
    Span4Mux_v I__12834 (
            .O(N__63119),
            .I(N__63097));
    LocalMux I__12833 (
            .O(N__63116),
            .I(N__63092));
    Span12Mux_v I__12832 (
            .O(N__63103),
            .I(N__63092));
    Odrv4 I__12831 (
            .O(N__63100),
            .I(dc32_fifo_data_in_7));
    Odrv4 I__12830 (
            .O(N__63097),
            .I(dc32_fifo_data_in_7));
    Odrv12 I__12829 (
            .O(N__63092),
            .I(dc32_fifo_data_in_7));
    CascadeMux I__12828 (
            .O(N__63085),
            .I(N__63082));
    InMux I__12827 (
            .O(N__63082),
            .I(N__63079));
    LocalMux I__12826 (
            .O(N__63079),
            .I(N__63076));
    Span4Mux_v I__12825 (
            .O(N__63076),
            .I(N__63072));
    InMux I__12824 (
            .O(N__63075),
            .I(N__63069));
    Odrv4 I__12823 (
            .O(N__63072),
            .I(REG_mem_18_7));
    LocalMux I__12822 (
            .O(N__63069),
            .I(REG_mem_18_7));
    CascadeMux I__12821 (
            .O(N__63064),
            .I(N__63061));
    InMux I__12820 (
            .O(N__63061),
            .I(N__63057));
    InMux I__12819 (
            .O(N__63060),
            .I(N__63054));
    LocalMux I__12818 (
            .O(N__63057),
            .I(REG_mem_63_4));
    LocalMux I__12817 (
            .O(N__63054),
            .I(REG_mem_63_4));
    InMux I__12816 (
            .O(N__63049),
            .I(N__63046));
    LocalMux I__12815 (
            .O(N__63046),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14138 ));
    InMux I__12814 (
            .O(N__63043),
            .I(N__63039));
    InMux I__12813 (
            .O(N__63042),
            .I(N__63036));
    LocalMux I__12812 (
            .O(N__63039),
            .I(N__63033));
    LocalMux I__12811 (
            .O(N__63036),
            .I(REG_mem_31_2));
    Odrv4 I__12810 (
            .O(N__63033),
            .I(REG_mem_31_2));
    InMux I__12809 (
            .O(N__63028),
            .I(N__63025));
    LocalMux I__12808 (
            .O(N__63025),
            .I(N__63022));
    Span4Mux_v I__12807 (
            .O(N__63022),
            .I(N__63019));
    Span4Mux_h I__12806 (
            .O(N__63019),
            .I(N__63015));
    InMux I__12805 (
            .O(N__63018),
            .I(N__63012));
    Odrv4 I__12804 (
            .O(N__63015),
            .I(REG_mem_48_4));
    LocalMux I__12803 (
            .O(N__63012),
            .I(REG_mem_48_4));
    InMux I__12802 (
            .O(N__63007),
            .I(N__63002));
    InMux I__12801 (
            .O(N__63006),
            .I(N__62998));
    InMux I__12800 (
            .O(N__63005),
            .I(N__62993));
    LocalMux I__12799 (
            .O(N__63002),
            .I(N__62990));
    InMux I__12798 (
            .O(N__63001),
            .I(N__62980));
    LocalMux I__12797 (
            .O(N__62998),
            .I(N__62975));
    InMux I__12796 (
            .O(N__62997),
            .I(N__62972));
    InMux I__12795 (
            .O(N__62996),
            .I(N__62969));
    LocalMux I__12794 (
            .O(N__62993),
            .I(N__62966));
    Span4Mux_v I__12793 (
            .O(N__62990),
            .I(N__62963));
    InMux I__12792 (
            .O(N__62989),
            .I(N__62959));
    InMux I__12791 (
            .O(N__62988),
            .I(N__62956));
    InMux I__12790 (
            .O(N__62987),
            .I(N__62953));
    InMux I__12789 (
            .O(N__62986),
            .I(N__62950));
    InMux I__12788 (
            .O(N__62985),
            .I(N__62947));
    InMux I__12787 (
            .O(N__62984),
            .I(N__62944));
    InMux I__12786 (
            .O(N__62983),
            .I(N__62941));
    LocalMux I__12785 (
            .O(N__62980),
            .I(N__62938));
    InMux I__12784 (
            .O(N__62979),
            .I(N__62935));
    InMux I__12783 (
            .O(N__62978),
            .I(N__62932));
    Span4Mux_h I__12782 (
            .O(N__62975),
            .I(N__62927));
    LocalMux I__12781 (
            .O(N__62972),
            .I(N__62927));
    LocalMux I__12780 (
            .O(N__62969),
            .I(N__62920));
    Span4Mux_v I__12779 (
            .O(N__62966),
            .I(N__62920));
    Span4Mux_h I__12778 (
            .O(N__62963),
            .I(N__62920));
    InMux I__12777 (
            .O(N__62962),
            .I(N__62917));
    LocalMux I__12776 (
            .O(N__62959),
            .I(N__62914));
    LocalMux I__12775 (
            .O(N__62956),
            .I(N__62905));
    LocalMux I__12774 (
            .O(N__62953),
            .I(N__62905));
    LocalMux I__12773 (
            .O(N__62950),
            .I(N__62905));
    LocalMux I__12772 (
            .O(N__62947),
            .I(N__62905));
    LocalMux I__12771 (
            .O(N__62944),
            .I(N__62900));
    LocalMux I__12770 (
            .O(N__62941),
            .I(N__62900));
    Span4Mux_h I__12769 (
            .O(N__62938),
            .I(N__62897));
    LocalMux I__12768 (
            .O(N__62935),
            .I(N__62890));
    LocalMux I__12767 (
            .O(N__62932),
            .I(N__62890));
    Span4Mux_v I__12766 (
            .O(N__62927),
            .I(N__62890));
    Span4Mux_v I__12765 (
            .O(N__62920),
            .I(N__62887));
    LocalMux I__12764 (
            .O(N__62917),
            .I(n16));
    Odrv4 I__12763 (
            .O(N__62914),
            .I(n16));
    Odrv12 I__12762 (
            .O(N__62905),
            .I(n16));
    Odrv12 I__12761 (
            .O(N__62900),
            .I(n16));
    Odrv4 I__12760 (
            .O(N__62897),
            .I(n16));
    Odrv4 I__12759 (
            .O(N__62890),
            .I(n16));
    Odrv4 I__12758 (
            .O(N__62887),
            .I(n16));
    InMux I__12757 (
            .O(N__62872),
            .I(N__62866));
    InMux I__12756 (
            .O(N__62871),
            .I(N__62866));
    LocalMux I__12755 (
            .O(N__62866),
            .I(REG_mem_49_4));
    CascadeMux I__12754 (
            .O(N__62863),
            .I(N__62849));
    CascadeMux I__12753 (
            .O(N__62862),
            .I(N__62846));
    InMux I__12752 (
            .O(N__62861),
            .I(N__62839));
    InMux I__12751 (
            .O(N__62860),
            .I(N__62836));
    InMux I__12750 (
            .O(N__62859),
            .I(N__62824));
    InMux I__12749 (
            .O(N__62858),
            .I(N__62824));
    InMux I__12748 (
            .O(N__62857),
            .I(N__62824));
    InMux I__12747 (
            .O(N__62856),
            .I(N__62824));
    InMux I__12746 (
            .O(N__62855),
            .I(N__62818));
    CascadeMux I__12745 (
            .O(N__62854),
            .I(N__62814));
    InMux I__12744 (
            .O(N__62853),
            .I(N__62804));
    InMux I__12743 (
            .O(N__62852),
            .I(N__62793));
    InMux I__12742 (
            .O(N__62849),
            .I(N__62783));
    InMux I__12741 (
            .O(N__62846),
            .I(N__62783));
    InMux I__12740 (
            .O(N__62845),
            .I(N__62783));
    InMux I__12739 (
            .O(N__62844),
            .I(N__62770));
    InMux I__12738 (
            .O(N__62843),
            .I(N__62770));
    InMux I__12737 (
            .O(N__62842),
            .I(N__62770));
    LocalMux I__12736 (
            .O(N__62839),
            .I(N__62765));
    LocalMux I__12735 (
            .O(N__62836),
            .I(N__62765));
    InMux I__12734 (
            .O(N__62835),
            .I(N__62758));
    InMux I__12733 (
            .O(N__62834),
            .I(N__62758));
    InMux I__12732 (
            .O(N__62833),
            .I(N__62758));
    LocalMux I__12731 (
            .O(N__62824),
            .I(N__62755));
    InMux I__12730 (
            .O(N__62823),
            .I(N__62750));
    InMux I__12729 (
            .O(N__62822),
            .I(N__62750));
    InMux I__12728 (
            .O(N__62821),
            .I(N__62747));
    LocalMux I__12727 (
            .O(N__62818),
            .I(N__62744));
    InMux I__12726 (
            .O(N__62817),
            .I(N__62741));
    InMux I__12725 (
            .O(N__62814),
            .I(N__62734));
    InMux I__12724 (
            .O(N__62813),
            .I(N__62734));
    InMux I__12723 (
            .O(N__62812),
            .I(N__62734));
    InMux I__12722 (
            .O(N__62811),
            .I(N__62725));
    InMux I__12721 (
            .O(N__62810),
            .I(N__62725));
    InMux I__12720 (
            .O(N__62809),
            .I(N__62725));
    InMux I__12719 (
            .O(N__62808),
            .I(N__62725));
    CascadeMux I__12718 (
            .O(N__62807),
            .I(N__62720));
    LocalMux I__12717 (
            .O(N__62804),
            .I(N__62713));
    InMux I__12716 (
            .O(N__62803),
            .I(N__62710));
    InMux I__12715 (
            .O(N__62802),
            .I(N__62707));
    InMux I__12714 (
            .O(N__62801),
            .I(N__62704));
    InMux I__12713 (
            .O(N__62800),
            .I(N__62699));
    InMux I__12712 (
            .O(N__62799),
            .I(N__62699));
    InMux I__12711 (
            .O(N__62798),
            .I(N__62694));
    InMux I__12710 (
            .O(N__62797),
            .I(N__62694));
    InMux I__12709 (
            .O(N__62796),
            .I(N__62691));
    LocalMux I__12708 (
            .O(N__62793),
            .I(N__62685));
    InMux I__12707 (
            .O(N__62792),
            .I(N__62680));
    InMux I__12706 (
            .O(N__62791),
            .I(N__62680));
    InMux I__12705 (
            .O(N__62790),
            .I(N__62673));
    LocalMux I__12704 (
            .O(N__62783),
            .I(N__62670));
    InMux I__12703 (
            .O(N__62782),
            .I(N__62665));
    InMux I__12702 (
            .O(N__62781),
            .I(N__62665));
    InMux I__12701 (
            .O(N__62780),
            .I(N__62656));
    InMux I__12700 (
            .O(N__62779),
            .I(N__62656));
    InMux I__12699 (
            .O(N__62778),
            .I(N__62656));
    InMux I__12698 (
            .O(N__62777),
            .I(N__62656));
    LocalMux I__12697 (
            .O(N__62770),
            .I(N__62641));
    Span4Mux_h I__12696 (
            .O(N__62765),
            .I(N__62641));
    LocalMux I__12695 (
            .O(N__62758),
            .I(N__62641));
    Span4Mux_h I__12694 (
            .O(N__62755),
            .I(N__62641));
    LocalMux I__12693 (
            .O(N__62750),
            .I(N__62641));
    LocalMux I__12692 (
            .O(N__62747),
            .I(N__62641));
    Span4Mux_v I__12691 (
            .O(N__62744),
            .I(N__62641));
    LocalMux I__12690 (
            .O(N__62741),
            .I(N__62636));
    LocalMux I__12689 (
            .O(N__62734),
            .I(N__62636));
    LocalMux I__12688 (
            .O(N__62725),
            .I(N__62630));
    InMux I__12687 (
            .O(N__62724),
            .I(N__62625));
    InMux I__12686 (
            .O(N__62723),
            .I(N__62625));
    InMux I__12685 (
            .O(N__62720),
            .I(N__62618));
    InMux I__12684 (
            .O(N__62719),
            .I(N__62618));
    InMux I__12683 (
            .O(N__62718),
            .I(N__62618));
    InMux I__12682 (
            .O(N__62717),
            .I(N__62613));
    InMux I__12681 (
            .O(N__62716),
            .I(N__62613));
    Span4Mux_h I__12680 (
            .O(N__62713),
            .I(N__62607));
    LocalMux I__12679 (
            .O(N__62710),
            .I(N__62607));
    LocalMux I__12678 (
            .O(N__62707),
            .I(N__62596));
    LocalMux I__12677 (
            .O(N__62704),
            .I(N__62596));
    LocalMux I__12676 (
            .O(N__62699),
            .I(N__62596));
    LocalMux I__12675 (
            .O(N__62694),
            .I(N__62596));
    LocalMux I__12674 (
            .O(N__62691),
            .I(N__62596));
    InMux I__12673 (
            .O(N__62690),
            .I(N__62593));
    InMux I__12672 (
            .O(N__62689),
            .I(N__62590));
    InMux I__12671 (
            .O(N__62688),
            .I(N__62587));
    Span4Mux_h I__12670 (
            .O(N__62685),
            .I(N__62582));
    LocalMux I__12669 (
            .O(N__62680),
            .I(N__62582));
    InMux I__12668 (
            .O(N__62679),
            .I(N__62579));
    InMux I__12667 (
            .O(N__62678),
            .I(N__62576));
    InMux I__12666 (
            .O(N__62677),
            .I(N__62573));
    InMux I__12665 (
            .O(N__62676),
            .I(N__62570));
    LocalMux I__12664 (
            .O(N__62673),
            .I(N__62557));
    Span4Mux_h I__12663 (
            .O(N__62670),
            .I(N__62557));
    LocalMux I__12662 (
            .O(N__62665),
            .I(N__62557));
    LocalMux I__12661 (
            .O(N__62656),
            .I(N__62557));
    Span4Mux_v I__12660 (
            .O(N__62641),
            .I(N__62557));
    Span4Mux_h I__12659 (
            .O(N__62636),
            .I(N__62557));
    InMux I__12658 (
            .O(N__62635),
            .I(N__62550));
    InMux I__12657 (
            .O(N__62634),
            .I(N__62550));
    InMux I__12656 (
            .O(N__62633),
            .I(N__62550));
    Span4Mux_v I__12655 (
            .O(N__62630),
            .I(N__62547));
    LocalMux I__12654 (
            .O(N__62625),
            .I(N__62542));
    LocalMux I__12653 (
            .O(N__62618),
            .I(N__62542));
    LocalMux I__12652 (
            .O(N__62613),
            .I(N__62539));
    InMux I__12651 (
            .O(N__62612),
            .I(N__62536));
    Span4Mux_v I__12650 (
            .O(N__62607),
            .I(N__62531));
    Span4Mux_v I__12649 (
            .O(N__62596),
            .I(N__62531));
    LocalMux I__12648 (
            .O(N__62593),
            .I(N__62522));
    LocalMux I__12647 (
            .O(N__62590),
            .I(N__62522));
    LocalMux I__12646 (
            .O(N__62587),
            .I(N__62522));
    Sp12to4 I__12645 (
            .O(N__62582),
            .I(N__62522));
    LocalMux I__12644 (
            .O(N__62579),
            .I(N__62517));
    LocalMux I__12643 (
            .O(N__62576),
            .I(N__62517));
    LocalMux I__12642 (
            .O(N__62573),
            .I(N__62510));
    LocalMux I__12641 (
            .O(N__62570),
            .I(N__62510));
    Span4Mux_v I__12640 (
            .O(N__62557),
            .I(N__62510));
    LocalMux I__12639 (
            .O(N__62550),
            .I(N__62507));
    Span4Mux_h I__12638 (
            .O(N__62547),
            .I(N__62504));
    Span4Mux_v I__12637 (
            .O(N__62542),
            .I(N__62501));
    Span12Mux_h I__12636 (
            .O(N__62539),
            .I(N__62498));
    LocalMux I__12635 (
            .O(N__62536),
            .I(N__62491));
    Sp12to4 I__12634 (
            .O(N__62531),
            .I(N__62491));
    Span12Mux_v I__12633 (
            .O(N__62522),
            .I(N__62491));
    Span4Mux_v I__12632 (
            .O(N__62517),
            .I(N__62486));
    Span4Mux_h I__12631 (
            .O(N__62510),
            .I(N__62486));
    Span4Mux_h I__12630 (
            .O(N__62507),
            .I(N__62481));
    Span4Mux_h I__12629 (
            .O(N__62504),
            .I(N__62481));
    Odrv4 I__12628 (
            .O(N__62501),
            .I(dc32_fifo_data_in_5));
    Odrv12 I__12627 (
            .O(N__62498),
            .I(dc32_fifo_data_in_5));
    Odrv12 I__12626 (
            .O(N__62491),
            .I(dc32_fifo_data_in_5));
    Odrv4 I__12625 (
            .O(N__62486),
            .I(dc32_fifo_data_in_5));
    Odrv4 I__12624 (
            .O(N__62481),
            .I(dc32_fifo_data_in_5));
    CascadeMux I__12623 (
            .O(N__62470),
            .I(N__62467));
    InMux I__12622 (
            .O(N__62467),
            .I(N__62464));
    LocalMux I__12621 (
            .O(N__62464),
            .I(N__62460));
    CascadeMux I__12620 (
            .O(N__62463),
            .I(N__62457));
    Span4Mux_v I__12619 (
            .O(N__62460),
            .I(N__62454));
    InMux I__12618 (
            .O(N__62457),
            .I(N__62451));
    Odrv4 I__12617 (
            .O(N__62454),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_5 ));
    LocalMux I__12616 (
            .O(N__62451),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_5 ));
    InMux I__12615 (
            .O(N__62446),
            .I(N__62439));
    InMux I__12614 (
            .O(N__62445),
            .I(N__62439));
    InMux I__12613 (
            .O(N__62444),
            .I(N__62436));
    LocalMux I__12612 (
            .O(N__62439),
            .I(N__62431));
    LocalMux I__12611 (
            .O(N__62436),
            .I(N__62431));
    Span4Mux_v I__12610 (
            .O(N__62431),
            .I(N__62426));
    CascadeMux I__12609 (
            .O(N__62430),
            .I(N__62416));
    CascadeMux I__12608 (
            .O(N__62429),
            .I(N__62408));
    Span4Mux_h I__12607 (
            .O(N__62426),
            .I(N__62404));
    InMux I__12606 (
            .O(N__62425),
            .I(N__62401));
    InMux I__12605 (
            .O(N__62424),
            .I(N__62395));
    InMux I__12604 (
            .O(N__62423),
            .I(N__62395));
    InMux I__12603 (
            .O(N__62422),
            .I(N__62388));
    InMux I__12602 (
            .O(N__62421),
            .I(N__62388));
    InMux I__12601 (
            .O(N__62420),
            .I(N__62388));
    InMux I__12600 (
            .O(N__62419),
            .I(N__62385));
    InMux I__12599 (
            .O(N__62416),
            .I(N__62380));
    InMux I__12598 (
            .O(N__62415),
            .I(N__62368));
    InMux I__12597 (
            .O(N__62414),
            .I(N__62364));
    InMux I__12596 (
            .O(N__62413),
            .I(N__62361));
    InMux I__12595 (
            .O(N__62412),
            .I(N__62346));
    InMux I__12594 (
            .O(N__62411),
            .I(N__62341));
    InMux I__12593 (
            .O(N__62408),
            .I(N__62341));
    InMux I__12592 (
            .O(N__62407),
            .I(N__62338));
    Span4Mux_h I__12591 (
            .O(N__62404),
            .I(N__62333));
    LocalMux I__12590 (
            .O(N__62401),
            .I(N__62333));
    InMux I__12589 (
            .O(N__62400),
            .I(N__62326));
    LocalMux I__12588 (
            .O(N__62395),
            .I(N__62321));
    LocalMux I__12587 (
            .O(N__62388),
            .I(N__62321));
    LocalMux I__12586 (
            .O(N__62385),
            .I(N__62318));
    InMux I__12585 (
            .O(N__62384),
            .I(N__62312));
    InMux I__12584 (
            .O(N__62383),
            .I(N__62309));
    LocalMux I__12583 (
            .O(N__62380),
            .I(N__62306));
    InMux I__12582 (
            .O(N__62379),
            .I(N__62297));
    InMux I__12581 (
            .O(N__62378),
            .I(N__62297));
    InMux I__12580 (
            .O(N__62377),
            .I(N__62297));
    InMux I__12579 (
            .O(N__62376),
            .I(N__62297));
    InMux I__12578 (
            .O(N__62375),
            .I(N__62292));
    InMux I__12577 (
            .O(N__62374),
            .I(N__62292));
    InMux I__12576 (
            .O(N__62373),
            .I(N__62285));
    InMux I__12575 (
            .O(N__62372),
            .I(N__62285));
    InMux I__12574 (
            .O(N__62371),
            .I(N__62285));
    LocalMux I__12573 (
            .O(N__62368),
            .I(N__62282));
    InMux I__12572 (
            .O(N__62367),
            .I(N__62279));
    LocalMux I__12571 (
            .O(N__62364),
            .I(N__62274));
    LocalMux I__12570 (
            .O(N__62361),
            .I(N__62274));
    CascadeMux I__12569 (
            .O(N__62360),
            .I(N__62270));
    InMux I__12568 (
            .O(N__62359),
            .I(N__62263));
    InMux I__12567 (
            .O(N__62358),
            .I(N__62263));
    InMux I__12566 (
            .O(N__62357),
            .I(N__62256));
    InMux I__12565 (
            .O(N__62356),
            .I(N__62256));
    InMux I__12564 (
            .O(N__62355),
            .I(N__62256));
    InMux I__12563 (
            .O(N__62354),
            .I(N__62248));
    InMux I__12562 (
            .O(N__62353),
            .I(N__62245));
    InMux I__12561 (
            .O(N__62352),
            .I(N__62240));
    InMux I__12560 (
            .O(N__62351),
            .I(N__62237));
    InMux I__12559 (
            .O(N__62350),
            .I(N__62232));
    InMux I__12558 (
            .O(N__62349),
            .I(N__62232));
    LocalMux I__12557 (
            .O(N__62346),
            .I(N__62229));
    LocalMux I__12556 (
            .O(N__62341),
            .I(N__62222));
    LocalMux I__12555 (
            .O(N__62338),
            .I(N__62222));
    Span4Mux_v I__12554 (
            .O(N__62333),
            .I(N__62222));
    InMux I__12553 (
            .O(N__62332),
            .I(N__62219));
    InMux I__12552 (
            .O(N__62331),
            .I(N__62213));
    InMux I__12551 (
            .O(N__62330),
            .I(N__62208));
    InMux I__12550 (
            .O(N__62329),
            .I(N__62208));
    LocalMux I__12549 (
            .O(N__62326),
            .I(N__62205));
    Span4Mux_v I__12548 (
            .O(N__62321),
            .I(N__62202));
    Sp12to4 I__12547 (
            .O(N__62318),
            .I(N__62199));
    InMux I__12546 (
            .O(N__62317),
            .I(N__62195));
    InMux I__12545 (
            .O(N__62316),
            .I(N__62192));
    InMux I__12544 (
            .O(N__62315),
            .I(N__62189));
    LocalMux I__12543 (
            .O(N__62312),
            .I(N__62186));
    LocalMux I__12542 (
            .O(N__62309),
            .I(N__62179));
    Span4Mux_v I__12541 (
            .O(N__62306),
            .I(N__62179));
    LocalMux I__12540 (
            .O(N__62297),
            .I(N__62179));
    LocalMux I__12539 (
            .O(N__62292),
            .I(N__62168));
    LocalMux I__12538 (
            .O(N__62285),
            .I(N__62168));
    Span4Mux_h I__12537 (
            .O(N__62282),
            .I(N__62168));
    LocalMux I__12536 (
            .O(N__62279),
            .I(N__62168));
    Span4Mux_v I__12535 (
            .O(N__62274),
            .I(N__62168));
    InMux I__12534 (
            .O(N__62273),
            .I(N__62159));
    InMux I__12533 (
            .O(N__62270),
            .I(N__62159));
    InMux I__12532 (
            .O(N__62269),
            .I(N__62159));
    InMux I__12531 (
            .O(N__62268),
            .I(N__62159));
    LocalMux I__12530 (
            .O(N__62263),
            .I(N__62154));
    LocalMux I__12529 (
            .O(N__62256),
            .I(N__62154));
    InMux I__12528 (
            .O(N__62255),
            .I(N__62149));
    InMux I__12527 (
            .O(N__62254),
            .I(N__62149));
    InMux I__12526 (
            .O(N__62253),
            .I(N__62142));
    InMux I__12525 (
            .O(N__62252),
            .I(N__62142));
    InMux I__12524 (
            .O(N__62251),
            .I(N__62142));
    LocalMux I__12523 (
            .O(N__62248),
            .I(N__62137));
    LocalMux I__12522 (
            .O(N__62245),
            .I(N__62137));
    InMux I__12521 (
            .O(N__62244),
            .I(N__62132));
    InMux I__12520 (
            .O(N__62243),
            .I(N__62132));
    LocalMux I__12519 (
            .O(N__62240),
            .I(N__62125));
    LocalMux I__12518 (
            .O(N__62237),
            .I(N__62125));
    LocalMux I__12517 (
            .O(N__62232),
            .I(N__62125));
    Span4Mux_v I__12516 (
            .O(N__62229),
            .I(N__62118));
    Span4Mux_v I__12515 (
            .O(N__62222),
            .I(N__62118));
    LocalMux I__12514 (
            .O(N__62219),
            .I(N__62118));
    InMux I__12513 (
            .O(N__62218),
            .I(N__62111));
    InMux I__12512 (
            .O(N__62217),
            .I(N__62111));
    InMux I__12511 (
            .O(N__62216),
            .I(N__62111));
    LocalMux I__12510 (
            .O(N__62213),
            .I(N__62108));
    LocalMux I__12509 (
            .O(N__62208),
            .I(N__62103));
    Sp12to4 I__12508 (
            .O(N__62205),
            .I(N__62103));
    Sp12to4 I__12507 (
            .O(N__62202),
            .I(N__62098));
    Span12Mux_v I__12506 (
            .O(N__62199),
            .I(N__62098));
    InMux I__12505 (
            .O(N__62198),
            .I(N__62095));
    LocalMux I__12504 (
            .O(N__62195),
            .I(N__62084));
    LocalMux I__12503 (
            .O(N__62192),
            .I(N__62084));
    LocalMux I__12502 (
            .O(N__62189),
            .I(N__62084));
    Span4Mux_v I__12501 (
            .O(N__62186),
            .I(N__62084));
    Span4Mux_h I__12500 (
            .O(N__62179),
            .I(N__62084));
    Span4Mux_v I__12499 (
            .O(N__62168),
            .I(N__62081));
    LocalMux I__12498 (
            .O(N__62159),
            .I(N__62078));
    Span4Mux_v I__12497 (
            .O(N__62154),
            .I(N__62075));
    LocalMux I__12496 (
            .O(N__62149),
            .I(N__62068));
    LocalMux I__12495 (
            .O(N__62142),
            .I(N__62068));
    Span12Mux_v I__12494 (
            .O(N__62137),
            .I(N__62068));
    LocalMux I__12493 (
            .O(N__62132),
            .I(N__62061));
    Span4Mux_h I__12492 (
            .O(N__62125),
            .I(N__62061));
    Span4Mux_h I__12491 (
            .O(N__62118),
            .I(N__62061));
    LocalMux I__12490 (
            .O(N__62111),
            .I(N__62052));
    Span12Mux_h I__12489 (
            .O(N__62108),
            .I(N__62052));
    Span12Mux_v I__12488 (
            .O(N__62103),
            .I(N__62052));
    Span12Mux_h I__12487 (
            .O(N__62098),
            .I(N__62052));
    LocalMux I__12486 (
            .O(N__62095),
            .I(N__62045));
    Span4Mux_v I__12485 (
            .O(N__62084),
            .I(N__62045));
    Span4Mux_h I__12484 (
            .O(N__62081),
            .I(N__62045));
    Odrv4 I__12483 (
            .O(N__62078),
            .I(dc32_fifo_data_in_15));
    Odrv4 I__12482 (
            .O(N__62075),
            .I(dc32_fifo_data_in_15));
    Odrv12 I__12481 (
            .O(N__62068),
            .I(dc32_fifo_data_in_15));
    Odrv4 I__12480 (
            .O(N__62061),
            .I(dc32_fifo_data_in_15));
    Odrv12 I__12479 (
            .O(N__62052),
            .I(dc32_fifo_data_in_15));
    Odrv4 I__12478 (
            .O(N__62045),
            .I(dc32_fifo_data_in_15));
    InMux I__12477 (
            .O(N__62032),
            .I(N__62029));
    LocalMux I__12476 (
            .O(N__62029),
            .I(N__62026));
    Span4Mux_v I__12475 (
            .O(N__62026),
            .I(N__62023));
    Sp12to4 I__12474 (
            .O(N__62023),
            .I(N__62020));
    Span12Mux_s11_h I__12473 (
            .O(N__62020),
            .I(N__62016));
    InMux I__12472 (
            .O(N__62019),
            .I(N__62013));
    Odrv12 I__12471 (
            .O(N__62016),
            .I(REG_mem_26_15));
    LocalMux I__12470 (
            .O(N__62013),
            .I(REG_mem_26_15));
    InMux I__12469 (
            .O(N__62008),
            .I(N__62005));
    LocalMux I__12468 (
            .O(N__62005),
            .I(N__62002));
    Span4Mux_h I__12467 (
            .O(N__62002),
            .I(N__61998));
    InMux I__12466 (
            .O(N__62001),
            .I(N__61995));
    Span4Mux_h I__12465 (
            .O(N__61998),
            .I(N__61990));
    LocalMux I__12464 (
            .O(N__61995),
            .I(N__61990));
    Odrv4 I__12463 (
            .O(N__61990),
            .I(REG_mem_7_4));
    InMux I__12462 (
            .O(N__61987),
            .I(N__61981));
    InMux I__12461 (
            .O(N__61986),
            .I(N__61981));
    LocalMux I__12460 (
            .O(N__61981),
            .I(REG_mem_6_4));
    CascadeMux I__12459 (
            .O(N__61978),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12377_cascade_ ));
    InMux I__12458 (
            .O(N__61975),
            .I(N__61972));
    LocalMux I__12457 (
            .O(N__61972),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12376 ));
    InMux I__12456 (
            .O(N__61969),
            .I(N__61966));
    LocalMux I__12455 (
            .O(N__61966),
            .I(N__61963));
    Span4Mux_v I__12454 (
            .O(N__61963),
            .I(N__61960));
    Span4Mux_h I__12453 (
            .O(N__61960),
            .I(N__61957));
    Odrv4 I__12452 (
            .O(N__61957),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12346 ));
    CascadeMux I__12451 (
            .O(N__61954),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13010_cascade_ ));
    InMux I__12450 (
            .O(N__61951),
            .I(N__61948));
    LocalMux I__12449 (
            .O(N__61948),
            .I(N__61945));
    Odrv4 I__12448 (
            .O(N__61945),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13013 ));
    InMux I__12447 (
            .O(N__61942),
            .I(N__61939));
    LocalMux I__12446 (
            .O(N__61939),
            .I(N__61936));
    Span12Mux_h I__12445 (
            .O(N__61936),
            .I(N__61932));
    InMux I__12444 (
            .O(N__61935),
            .I(N__61929));
    Odrv12 I__12443 (
            .O(N__61932),
            .I(REG_mem_38_2));
    LocalMux I__12442 (
            .O(N__61929),
            .I(REG_mem_38_2));
    CascadeMux I__12441 (
            .O(N__61924),
            .I(N__61921));
    InMux I__12440 (
            .O(N__61921),
            .I(N__61918));
    LocalMux I__12439 (
            .O(N__61918),
            .I(N__61915));
    Odrv4 I__12438 (
            .O(N__61915),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14210 ));
    InMux I__12437 (
            .O(N__61912),
            .I(N__61909));
    LocalMux I__12436 (
            .O(N__61909),
            .I(N__61906));
    Span4Mux_v I__12435 (
            .O(N__61906),
            .I(N__61902));
    InMux I__12434 (
            .O(N__61905),
            .I(N__61899));
    Odrv4 I__12433 (
            .O(N__61902),
            .I(REG_mem_41_4));
    LocalMux I__12432 (
            .O(N__61899),
            .I(REG_mem_41_4));
    InMux I__12431 (
            .O(N__61894),
            .I(N__61886));
    InMux I__12430 (
            .O(N__61893),
            .I(N__61882));
    InMux I__12429 (
            .O(N__61892),
            .I(N__61875));
    InMux I__12428 (
            .O(N__61891),
            .I(N__61872));
    InMux I__12427 (
            .O(N__61890),
            .I(N__61867));
    InMux I__12426 (
            .O(N__61889),
            .I(N__61867));
    LocalMux I__12425 (
            .O(N__61886),
            .I(N__61864));
    InMux I__12424 (
            .O(N__61885),
            .I(N__61861));
    LocalMux I__12423 (
            .O(N__61882),
            .I(N__61858));
    InMux I__12422 (
            .O(N__61881),
            .I(N__61855));
    InMux I__12421 (
            .O(N__61880),
            .I(N__61852));
    InMux I__12420 (
            .O(N__61879),
            .I(N__61849));
    InMux I__12419 (
            .O(N__61878),
            .I(N__61846));
    LocalMux I__12418 (
            .O(N__61875),
            .I(N__61839));
    LocalMux I__12417 (
            .O(N__61872),
            .I(N__61839));
    LocalMux I__12416 (
            .O(N__61867),
            .I(N__61839));
    Span4Mux_h I__12415 (
            .O(N__61864),
            .I(N__61836));
    LocalMux I__12414 (
            .O(N__61861),
            .I(N__61831));
    Span4Mux_v I__12413 (
            .O(N__61858),
            .I(N__61831));
    LocalMux I__12412 (
            .O(N__61855),
            .I(N__61824));
    LocalMux I__12411 (
            .O(N__61852),
            .I(N__61821));
    LocalMux I__12410 (
            .O(N__61849),
            .I(N__61818));
    LocalMux I__12409 (
            .O(N__61846),
            .I(N__61815));
    Span4Mux_h I__12408 (
            .O(N__61839),
            .I(N__61810));
    Span4Mux_v I__12407 (
            .O(N__61836),
            .I(N__61810));
    Span4Mux_v I__12406 (
            .O(N__61831),
            .I(N__61807));
    InMux I__12405 (
            .O(N__61830),
            .I(N__61804));
    InMux I__12404 (
            .O(N__61829),
            .I(N__61801));
    InMux I__12403 (
            .O(N__61828),
            .I(N__61798));
    InMux I__12402 (
            .O(N__61827),
            .I(N__61795));
    Span4Mux_h I__12401 (
            .O(N__61824),
            .I(N__61792));
    Span4Mux_v I__12400 (
            .O(N__61821),
            .I(N__61783));
    Span4Mux_v I__12399 (
            .O(N__61818),
            .I(N__61783));
    Span4Mux_v I__12398 (
            .O(N__61815),
            .I(N__61783));
    Span4Mux_v I__12397 (
            .O(N__61810),
            .I(N__61783));
    Span4Mux_v I__12396 (
            .O(N__61807),
            .I(N__61780));
    LocalMux I__12395 (
            .O(N__61804),
            .I(n26));
    LocalMux I__12394 (
            .O(N__61801),
            .I(n26));
    LocalMux I__12393 (
            .O(N__61798),
            .I(n26));
    LocalMux I__12392 (
            .O(N__61795),
            .I(n26));
    Odrv4 I__12391 (
            .O(N__61792),
            .I(n26));
    Odrv4 I__12390 (
            .O(N__61783),
            .I(n26));
    Odrv4 I__12389 (
            .O(N__61780),
            .I(n26));
    InMux I__12388 (
            .O(N__61765),
            .I(N__61759));
    InMux I__12387 (
            .O(N__61764),
            .I(N__61759));
    LocalMux I__12386 (
            .O(N__61759),
            .I(REG_mem_39_2));
    InMux I__12385 (
            .O(N__61756),
            .I(N__61753));
    LocalMux I__12384 (
            .O(N__61753),
            .I(N__61750));
    Span4Mux_v I__12383 (
            .O(N__61750),
            .I(N__61747));
    Span4Mux_v I__12382 (
            .O(N__61747),
            .I(N__61743));
    InMux I__12381 (
            .O(N__61746),
            .I(N__61740));
    Odrv4 I__12380 (
            .O(N__61743),
            .I(REG_mem_18_2));
    LocalMux I__12379 (
            .O(N__61740),
            .I(REG_mem_18_2));
    InMux I__12378 (
            .O(N__61735),
            .I(N__61732));
    LocalMux I__12377 (
            .O(N__61732),
            .I(N__61729));
    Span4Mux_v I__12376 (
            .O(N__61729),
            .I(N__61725));
    InMux I__12375 (
            .O(N__61728),
            .I(N__61722));
    Odrv4 I__12374 (
            .O(N__61725),
            .I(REG_mem_19_2));
    LocalMux I__12373 (
            .O(N__61722),
            .I(REG_mem_19_2));
    InMux I__12372 (
            .O(N__61717),
            .I(N__61713));
    InMux I__12371 (
            .O(N__61716),
            .I(N__61710));
    LocalMux I__12370 (
            .O(N__61713),
            .I(REG_mem_26_2));
    LocalMux I__12369 (
            .O(N__61710),
            .I(REG_mem_26_2));
    CascadeMux I__12368 (
            .O(N__61705),
            .I(N__61702));
    InMux I__12367 (
            .O(N__61702),
            .I(N__61699));
    LocalMux I__12366 (
            .O(N__61699),
            .I(N__61696));
    Span4Mux_v I__12365 (
            .O(N__61696),
            .I(N__61692));
    InMux I__12364 (
            .O(N__61695),
            .I(N__61689));
    Odrv4 I__12363 (
            .O(N__61692),
            .I(REG_mem_42_2));
    LocalMux I__12362 (
            .O(N__61689),
            .I(REG_mem_42_2));
    InMux I__12361 (
            .O(N__61684),
            .I(N__61681));
    LocalMux I__12360 (
            .O(N__61681),
            .I(N__61677));
    InMux I__12359 (
            .O(N__61680),
            .I(N__61674));
    Odrv4 I__12358 (
            .O(N__61677),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_2 ));
    LocalMux I__12357 (
            .O(N__61674),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_2 ));
    InMux I__12356 (
            .O(N__61669),
            .I(N__61666));
    LocalMux I__12355 (
            .O(N__61666),
            .I(N__61662));
    InMux I__12354 (
            .O(N__61665),
            .I(N__61659));
    Odrv4 I__12353 (
            .O(N__61662),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_2 ));
    LocalMux I__12352 (
            .O(N__61659),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_2 ));
    InMux I__12351 (
            .O(N__61654),
            .I(N__61651));
    LocalMux I__12350 (
            .O(N__61651),
            .I(N__61648));
    Span4Mux_h I__12349 (
            .O(N__61648),
            .I(N__61644));
    CascadeMux I__12348 (
            .O(N__61647),
            .I(N__61641));
    Span4Mux_h I__12347 (
            .O(N__61644),
            .I(N__61638));
    InMux I__12346 (
            .O(N__61641),
            .I(N__61635));
    Odrv4 I__12345 (
            .O(N__61638),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_2 ));
    LocalMux I__12344 (
            .O(N__61635),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_2 ));
    CascadeMux I__12343 (
            .O(N__61630),
            .I(N__61627));
    InMux I__12342 (
            .O(N__61627),
            .I(N__61624));
    LocalMux I__12341 (
            .O(N__61624),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14360 ));
    CascadeMux I__12340 (
            .O(N__61621),
            .I(N__61618));
    InMux I__12339 (
            .O(N__61618),
            .I(N__61614));
    InMux I__12338 (
            .O(N__61617),
            .I(N__61611));
    LocalMux I__12337 (
            .O(N__61614),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_2 ));
    LocalMux I__12336 (
            .O(N__61611),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_2 ));
    CascadeMux I__12335 (
            .O(N__61606),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12848_cascade_ ));
    CascadeMux I__12334 (
            .O(N__61603),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12851_cascade_ ));
    InMux I__12333 (
            .O(N__61600),
            .I(N__61597));
    LocalMux I__12332 (
            .O(N__61597),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14363 ));
    InMux I__12331 (
            .O(N__61594),
            .I(N__61591));
    LocalMux I__12330 (
            .O(N__61591),
            .I(N__61588));
    Span4Mux_v I__12329 (
            .O(N__61588),
            .I(N__61585));
    Sp12to4 I__12328 (
            .O(N__61585),
            .I(N__61582));
    Odrv12 I__12327 (
            .O(N__61582),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13607 ));
    InMux I__12326 (
            .O(N__61579),
            .I(N__61576));
    LocalMux I__12325 (
            .O(N__61576),
            .I(N__61573));
    Odrv12 I__12324 (
            .O(N__61573),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13979 ));
    CascadeMux I__12323 (
            .O(N__61570),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14408_cascade_ ));
    InMux I__12322 (
            .O(N__61567),
            .I(N__61564));
    LocalMux I__12321 (
            .O(N__61564),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13913 ));
    CascadeMux I__12320 (
            .O(N__61561),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14411_cascade_ ));
    InMux I__12319 (
            .O(N__61558),
            .I(N__61555));
    LocalMux I__12318 (
            .O(N__61555),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12947 ));
    CascadeMux I__12317 (
            .O(N__61552),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11498_cascade_ ));
    CascadeMux I__12316 (
            .O(N__61549),
            .I(N__61546));
    InMux I__12315 (
            .O(N__61546),
            .I(N__61543));
    LocalMux I__12314 (
            .O(N__61543),
            .I(N__61540));
    Span4Mux_v I__12313 (
            .O(N__61540),
            .I(N__61537));
    Span4Mux_h I__12312 (
            .O(N__61537),
            .I(N__61534));
    Span4Mux_v I__12311 (
            .O(N__61534),
            .I(N__61531));
    Span4Mux_v I__12310 (
            .O(N__61531),
            .I(N__61528));
    Odrv4 I__12309 (
            .O(N__61528),
            .I(REG_out_raw_2));
    InMux I__12308 (
            .O(N__61525),
            .I(N__61522));
    LocalMux I__12307 (
            .O(N__61522),
            .I(N__61519));
    Span4Mux_v I__12306 (
            .O(N__61519),
            .I(N__61516));
    Span4Mux_v I__12305 (
            .O(N__61516),
            .I(N__61513));
    Sp12to4 I__12304 (
            .O(N__61513),
            .I(N__61509));
    InMux I__12303 (
            .O(N__61512),
            .I(N__61506));
    Odrv12 I__12302 (
            .O(N__61509),
            .I(REG_mem_36_2));
    LocalMux I__12301 (
            .O(N__61506),
            .I(REG_mem_36_2));
    InMux I__12300 (
            .O(N__61501),
            .I(N__61498));
    LocalMux I__12299 (
            .O(N__61498),
            .I(N__61495));
    Span4Mux_v I__12298 (
            .O(N__61495),
            .I(N__61491));
    InMux I__12297 (
            .O(N__61494),
            .I(N__61488));
    Odrv4 I__12296 (
            .O(N__61491),
            .I(REG_mem_37_2));
    LocalMux I__12295 (
            .O(N__61488),
            .I(REG_mem_37_2));
    InMux I__12294 (
            .O(N__61483),
            .I(N__61480));
    LocalMux I__12293 (
            .O(N__61480),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12057 ));
    CascadeMux I__12292 (
            .O(N__61477),
            .I(N__61474));
    InMux I__12291 (
            .O(N__61474),
            .I(N__61470));
    InMux I__12290 (
            .O(N__61473),
            .I(N__61467));
    LocalMux I__12289 (
            .O(N__61470),
            .I(REG_mem_58_4));
    LocalMux I__12288 (
            .O(N__61467),
            .I(REG_mem_58_4));
    InMux I__12287 (
            .O(N__61462),
            .I(N__61456));
    InMux I__12286 (
            .O(N__61461),
            .I(N__61456));
    LocalMux I__12285 (
            .O(N__61456),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_4 ));
    InMux I__12284 (
            .O(N__61453),
            .I(N__61450));
    LocalMux I__12283 (
            .O(N__61450),
            .I(N__61446));
    CascadeMux I__12282 (
            .O(N__61449),
            .I(N__61443));
    Span4Mux_v I__12281 (
            .O(N__61446),
            .I(N__61440));
    InMux I__12280 (
            .O(N__61443),
            .I(N__61437));
    Odrv4 I__12279 (
            .O(N__61440),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_4 ));
    LocalMux I__12278 (
            .O(N__61437),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_4 ));
    CascadeMux I__12277 (
            .O(N__61432),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14198_cascade_ ));
    InMux I__12276 (
            .O(N__61429),
            .I(N__61425));
    CascadeMux I__12275 (
            .O(N__61428),
            .I(N__61422));
    LocalMux I__12274 (
            .O(N__61425),
            .I(N__61419));
    InMux I__12273 (
            .O(N__61422),
            .I(N__61416));
    Odrv4 I__12272 (
            .O(N__61419),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_4 ));
    LocalMux I__12271 (
            .O(N__61416),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_4 ));
    InMux I__12270 (
            .O(N__61411),
            .I(N__61408));
    LocalMux I__12269 (
            .O(N__61408),
            .I(\usb3_if_inst.usb3_data_in_latched_3 ));
    CascadeMux I__12268 (
            .O(N__61405),
            .I(N__61400));
    InMux I__12267 (
            .O(N__61404),
            .I(N__61390));
    InMux I__12266 (
            .O(N__61403),
            .I(N__61390));
    InMux I__12265 (
            .O(N__61400),
            .I(N__61379));
    InMux I__12264 (
            .O(N__61399),
            .I(N__61379));
    InMux I__12263 (
            .O(N__61398),
            .I(N__61374));
    InMux I__12262 (
            .O(N__61397),
            .I(N__61374));
    InMux I__12261 (
            .O(N__61396),
            .I(N__61367));
    InMux I__12260 (
            .O(N__61395),
            .I(N__61367));
    LocalMux I__12259 (
            .O(N__61390),
            .I(N__61364));
    InMux I__12258 (
            .O(N__61389),
            .I(N__61359));
    InMux I__12257 (
            .O(N__61388),
            .I(N__61359));
    InMux I__12256 (
            .O(N__61387),
            .I(N__61350));
    InMux I__12255 (
            .O(N__61386),
            .I(N__61350));
    InMux I__12254 (
            .O(N__61385),
            .I(N__61350));
    InMux I__12253 (
            .O(N__61384),
            .I(N__61350));
    LocalMux I__12252 (
            .O(N__61379),
            .I(N__61337));
    LocalMux I__12251 (
            .O(N__61374),
            .I(N__61334));
    InMux I__12250 (
            .O(N__61373),
            .I(N__61329));
    InMux I__12249 (
            .O(N__61372),
            .I(N__61326));
    LocalMux I__12248 (
            .O(N__61367),
            .I(N__61317));
    Span4Mux_v I__12247 (
            .O(N__61364),
            .I(N__61317));
    LocalMux I__12246 (
            .O(N__61359),
            .I(N__61317));
    LocalMux I__12245 (
            .O(N__61350),
            .I(N__61317));
    InMux I__12244 (
            .O(N__61349),
            .I(N__61308));
    InMux I__12243 (
            .O(N__61348),
            .I(N__61308));
    InMux I__12242 (
            .O(N__61347),
            .I(N__61308));
    InMux I__12241 (
            .O(N__61346),
            .I(N__61308));
    InMux I__12240 (
            .O(N__61345),
            .I(N__61301));
    InMux I__12239 (
            .O(N__61344),
            .I(N__61296));
    InMux I__12238 (
            .O(N__61343),
            .I(N__61296));
    InMux I__12237 (
            .O(N__61342),
            .I(N__61292));
    CascadeMux I__12236 (
            .O(N__61341),
            .I(N__61283));
    InMux I__12235 (
            .O(N__61340),
            .I(N__61277));
    Span4Mux_v I__12234 (
            .O(N__61337),
            .I(N__61272));
    Span4Mux_v I__12233 (
            .O(N__61334),
            .I(N__61272));
    InMux I__12232 (
            .O(N__61333),
            .I(N__61269));
    CascadeMux I__12231 (
            .O(N__61332),
            .I(N__61265));
    LocalMux I__12230 (
            .O(N__61329),
            .I(N__61259));
    LocalMux I__12229 (
            .O(N__61326),
            .I(N__61252));
    Span4Mux_v I__12228 (
            .O(N__61317),
            .I(N__61252));
    LocalMux I__12227 (
            .O(N__61308),
            .I(N__61252));
    InMux I__12226 (
            .O(N__61307),
            .I(N__61241));
    InMux I__12225 (
            .O(N__61306),
            .I(N__61241));
    InMux I__12224 (
            .O(N__61305),
            .I(N__61234));
    InMux I__12223 (
            .O(N__61304),
            .I(N__61234));
    LocalMux I__12222 (
            .O(N__61301),
            .I(N__61231));
    LocalMux I__12221 (
            .O(N__61296),
            .I(N__61228));
    InMux I__12220 (
            .O(N__61295),
            .I(N__61225));
    LocalMux I__12219 (
            .O(N__61292),
            .I(N__61222));
    InMux I__12218 (
            .O(N__61291),
            .I(N__61217));
    InMux I__12217 (
            .O(N__61290),
            .I(N__61214));
    InMux I__12216 (
            .O(N__61289),
            .I(N__61211));
    InMux I__12215 (
            .O(N__61288),
            .I(N__61208));
    InMux I__12214 (
            .O(N__61287),
            .I(N__61203));
    InMux I__12213 (
            .O(N__61286),
            .I(N__61203));
    InMux I__12212 (
            .O(N__61283),
            .I(N__61194));
    InMux I__12211 (
            .O(N__61282),
            .I(N__61194));
    InMux I__12210 (
            .O(N__61281),
            .I(N__61194));
    InMux I__12209 (
            .O(N__61280),
            .I(N__61194));
    LocalMux I__12208 (
            .O(N__61277),
            .I(N__61187));
    Span4Mux_h I__12207 (
            .O(N__61272),
            .I(N__61187));
    LocalMux I__12206 (
            .O(N__61269),
            .I(N__61187));
    InMux I__12205 (
            .O(N__61268),
            .I(N__61184));
    InMux I__12204 (
            .O(N__61265),
            .I(N__61179));
    InMux I__12203 (
            .O(N__61264),
            .I(N__61179));
    InMux I__12202 (
            .O(N__61263),
            .I(N__61174));
    InMux I__12201 (
            .O(N__61262),
            .I(N__61174));
    Span4Mux_v I__12200 (
            .O(N__61259),
            .I(N__61169));
    Span4Mux_v I__12199 (
            .O(N__61252),
            .I(N__61169));
    InMux I__12198 (
            .O(N__61251),
            .I(N__61166));
    InMux I__12197 (
            .O(N__61250),
            .I(N__61161));
    InMux I__12196 (
            .O(N__61249),
            .I(N__61161));
    InMux I__12195 (
            .O(N__61248),
            .I(N__61158));
    InMux I__12194 (
            .O(N__61247),
            .I(N__61155));
    InMux I__12193 (
            .O(N__61246),
            .I(N__61152));
    LocalMux I__12192 (
            .O(N__61241),
            .I(N__61149));
    InMux I__12191 (
            .O(N__61240),
            .I(N__61144));
    InMux I__12190 (
            .O(N__61239),
            .I(N__61144));
    LocalMux I__12189 (
            .O(N__61234),
            .I(N__61137));
    Span4Mux_h I__12188 (
            .O(N__61231),
            .I(N__61137));
    Span4Mux_h I__12187 (
            .O(N__61228),
            .I(N__61137));
    LocalMux I__12186 (
            .O(N__61225),
            .I(N__61134));
    Span4Mux_h I__12185 (
            .O(N__61222),
            .I(N__61131));
    InMux I__12184 (
            .O(N__61221),
            .I(N__61128));
    InMux I__12183 (
            .O(N__61220),
            .I(N__61125));
    LocalMux I__12182 (
            .O(N__61217),
            .I(N__61116));
    LocalMux I__12181 (
            .O(N__61214),
            .I(N__61116));
    LocalMux I__12180 (
            .O(N__61211),
            .I(N__61116));
    LocalMux I__12179 (
            .O(N__61208),
            .I(N__61116));
    LocalMux I__12178 (
            .O(N__61203),
            .I(N__61113));
    LocalMux I__12177 (
            .O(N__61194),
            .I(N__61100));
    Span4Mux_v I__12176 (
            .O(N__61187),
            .I(N__61100));
    LocalMux I__12175 (
            .O(N__61184),
            .I(N__61100));
    LocalMux I__12174 (
            .O(N__61179),
            .I(N__61091));
    LocalMux I__12173 (
            .O(N__61174),
            .I(N__61091));
    Span4Mux_h I__12172 (
            .O(N__61169),
            .I(N__61091));
    LocalMux I__12171 (
            .O(N__61166),
            .I(N__61091));
    LocalMux I__12170 (
            .O(N__61161),
            .I(N__61088));
    LocalMux I__12169 (
            .O(N__61158),
            .I(N__61085));
    LocalMux I__12168 (
            .O(N__61155),
            .I(N__61080));
    LocalMux I__12167 (
            .O(N__61152),
            .I(N__61080));
    Span4Mux_h I__12166 (
            .O(N__61149),
            .I(N__61077));
    LocalMux I__12165 (
            .O(N__61144),
            .I(N__61072));
    Span4Mux_h I__12164 (
            .O(N__61137),
            .I(N__61072));
    Span4Mux_h I__12163 (
            .O(N__61134),
            .I(N__61069));
    Span4Mux_h I__12162 (
            .O(N__61131),
            .I(N__61064));
    LocalMux I__12161 (
            .O(N__61128),
            .I(N__61064));
    LocalMux I__12160 (
            .O(N__61125),
            .I(N__61057));
    Span4Mux_v I__12159 (
            .O(N__61116),
            .I(N__61057));
    Span4Mux_h I__12158 (
            .O(N__61113),
            .I(N__61057));
    InMux I__12157 (
            .O(N__61112),
            .I(N__61042));
    InMux I__12156 (
            .O(N__61111),
            .I(N__61042));
    InMux I__12155 (
            .O(N__61110),
            .I(N__61042));
    InMux I__12154 (
            .O(N__61109),
            .I(N__61042));
    InMux I__12153 (
            .O(N__61108),
            .I(N__61042));
    InMux I__12152 (
            .O(N__61107),
            .I(N__61042));
    Span4Mux_v I__12151 (
            .O(N__61100),
            .I(N__61035));
    Span4Mux_v I__12150 (
            .O(N__61091),
            .I(N__61035));
    Span4Mux_v I__12149 (
            .O(N__61088),
            .I(N__61035));
    Span4Mux_v I__12148 (
            .O(N__61085),
            .I(N__61030));
    Span4Mux_v I__12147 (
            .O(N__61080),
            .I(N__61030));
    Span4Mux_h I__12146 (
            .O(N__61077),
            .I(N__61027));
    Span4Mux_h I__12145 (
            .O(N__61072),
            .I(N__61024));
    Span4Mux_h I__12144 (
            .O(N__61069),
            .I(N__61021));
    Span4Mux_v I__12143 (
            .O(N__61064),
            .I(N__61018));
    Span4Mux_h I__12142 (
            .O(N__61057),
            .I(N__61015));
    InMux I__12141 (
            .O(N__61056),
            .I(N__61010));
    InMux I__12140 (
            .O(N__61055),
            .I(N__61010));
    LocalMux I__12139 (
            .O(N__61042),
            .I(N__61005));
    Sp12to4 I__12138 (
            .O(N__61035),
            .I(N__61005));
    Span4Mux_h I__12137 (
            .O(N__61030),
            .I(N__61002));
    Span4Mux_v I__12136 (
            .O(N__61027),
            .I(N__60999));
    Span4Mux_h I__12135 (
            .O(N__61024),
            .I(N__60996));
    Span4Mux_h I__12134 (
            .O(N__61021),
            .I(N__60989));
    Span4Mux_h I__12133 (
            .O(N__61018),
            .I(N__60989));
    Span4Mux_h I__12132 (
            .O(N__61015),
            .I(N__60989));
    LocalMux I__12131 (
            .O(N__61010),
            .I(N__60984));
    Span12Mux_s8_h I__12130 (
            .O(N__61005),
            .I(N__60984));
    Span4Mux_h I__12129 (
            .O(N__61002),
            .I(N__60979));
    Span4Mux_v I__12128 (
            .O(N__60999),
            .I(N__60979));
    Sp12to4 I__12127 (
            .O(N__60996),
            .I(N__60972));
    Sp12to4 I__12126 (
            .O(N__60989),
            .I(N__60972));
    Span12Mux_h I__12125 (
            .O(N__60984),
            .I(N__60972));
    Odrv4 I__12124 (
            .O(N__60979),
            .I(dc32_fifo_data_in_3));
    Odrv12 I__12123 (
            .O(N__60972),
            .I(dc32_fifo_data_in_3));
    InMux I__12122 (
            .O(N__60967),
            .I(N__60964));
    LocalMux I__12121 (
            .O(N__60964),
            .I(\usb3_if_inst.usb3_data_in_latched_4 ));
    InMux I__12120 (
            .O(N__60961),
            .I(N__60958));
    LocalMux I__12119 (
            .O(N__60958),
            .I(\usb3_if_inst.usb3_data_in_latched_5 ));
    InMux I__12118 (
            .O(N__60955),
            .I(N__60952));
    LocalMux I__12117 (
            .O(N__60952),
            .I(\usb3_if_inst.usb3_data_in_latched_6 ));
    InMux I__12116 (
            .O(N__60949),
            .I(N__60946));
    LocalMux I__12115 (
            .O(N__60946),
            .I(\usb3_if_inst.usb3_data_in_latched_7 ));
    CascadeMux I__12114 (
            .O(N__60943),
            .I(N__60940));
    InMux I__12113 (
            .O(N__60940),
            .I(N__60937));
    LocalMux I__12112 (
            .O(N__60937),
            .I(N__60934));
    Span4Mux_v I__12111 (
            .O(N__60934),
            .I(N__60931));
    Span4Mux_h I__12110 (
            .O(N__60931),
            .I(N__60928));
    Odrv4 I__12109 (
            .O(N__60928),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12030 ));
    InMux I__12108 (
            .O(N__60925),
            .I(N__60922));
    LocalMux I__12107 (
            .O(N__60922),
            .I(N__60919));
    Span4Mux_h I__12106 (
            .O(N__60919),
            .I(N__60916));
    Odrv4 I__12105 (
            .O(N__60916),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12114 ));
    CascadeMux I__12104 (
            .O(N__60913),
            .I(N__60910));
    InMux I__12103 (
            .O(N__60910),
            .I(N__60907));
    LocalMux I__12102 (
            .O(N__60907),
            .I(N__60904));
    Span4Mux_v I__12101 (
            .O(N__60904),
            .I(N__60901));
    Odrv4 I__12100 (
            .O(N__60901),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12078 ));
    InMux I__12099 (
            .O(N__60898),
            .I(N__60895));
    LocalMux I__12098 (
            .O(N__60895),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12944 ));
    CascadeMux I__12097 (
            .O(N__60892),
            .I(n10562_cascade_));
    InMux I__12096 (
            .O(N__60889),
            .I(N__60874));
    InMux I__12095 (
            .O(N__60888),
            .I(N__60874));
    InMux I__12094 (
            .O(N__60887),
            .I(N__60874));
    InMux I__12093 (
            .O(N__60886),
            .I(N__60874));
    InMux I__12092 (
            .O(N__60885),
            .I(N__60874));
    LocalMux I__12091 (
            .O(N__60874),
            .I(reset_clk_counter_1));
    InMux I__12090 (
            .O(N__60871),
            .I(N__60862));
    InMux I__12089 (
            .O(N__60870),
            .I(N__60862));
    InMux I__12088 (
            .O(N__60869),
            .I(N__60862));
    LocalMux I__12087 (
            .O(N__60862),
            .I(reset_clk_counter_3));
    CascadeMux I__12086 (
            .O(N__60859),
            .I(N__60853));
    InMux I__12085 (
            .O(N__60858),
            .I(N__60848));
    InMux I__12084 (
            .O(N__60857),
            .I(N__60848));
    InMux I__12083 (
            .O(N__60856),
            .I(N__60843));
    InMux I__12082 (
            .O(N__60853),
            .I(N__60843));
    LocalMux I__12081 (
            .O(N__60848),
            .I(reset_clk_counter_2));
    LocalMux I__12080 (
            .O(N__60843),
            .I(reset_clk_counter_2));
    CascadeMux I__12079 (
            .O(N__60838),
            .I(N__60835));
    InMux I__12078 (
            .O(N__60835),
            .I(N__60826));
    InMux I__12077 (
            .O(N__60834),
            .I(N__60826));
    InMux I__12076 (
            .O(N__60833),
            .I(N__60826));
    LocalMux I__12075 (
            .O(N__60826),
            .I(reset_all_w_N_61));
    CascadeMux I__12074 (
            .O(N__60823),
            .I(reset_all_w_N_61_cascade_));
    CascadeMux I__12073 (
            .O(N__60820),
            .I(N__60814));
    InMux I__12072 (
            .O(N__60819),
            .I(N__60799));
    InMux I__12071 (
            .O(N__60818),
            .I(N__60799));
    InMux I__12070 (
            .O(N__60817),
            .I(N__60799));
    InMux I__12069 (
            .O(N__60814),
            .I(N__60799));
    InMux I__12068 (
            .O(N__60813),
            .I(N__60799));
    InMux I__12067 (
            .O(N__60812),
            .I(N__60799));
    LocalMux I__12066 (
            .O(N__60799),
            .I(reset_clk_counter_0));
    InMux I__12065 (
            .O(N__60796),
            .I(N__60788));
    InMux I__12064 (
            .O(N__60795),
            .I(N__60788));
    InMux I__12063 (
            .O(N__60794),
            .I(N__60782));
    InMux I__12062 (
            .O(N__60793),
            .I(N__60782));
    LocalMux I__12061 (
            .O(N__60788),
            .I(N__60777));
    InMux I__12060 (
            .O(N__60787),
            .I(N__60774));
    LocalMux I__12059 (
            .O(N__60782),
            .I(N__60771));
    CascadeMux I__12058 (
            .O(N__60781),
            .I(N__60764));
    InMux I__12057 (
            .O(N__60780),
            .I(N__60761));
    Span4Mux_h I__12056 (
            .O(N__60777),
            .I(N__60754));
    LocalMux I__12055 (
            .O(N__60774),
            .I(N__60754));
    Span4Mux_v I__12054 (
            .O(N__60771),
            .I(N__60754));
    InMux I__12053 (
            .O(N__60770),
            .I(N__60751));
    InMux I__12052 (
            .O(N__60769),
            .I(N__60742));
    InMux I__12051 (
            .O(N__60768),
            .I(N__60742));
    InMux I__12050 (
            .O(N__60767),
            .I(N__60742));
    InMux I__12049 (
            .O(N__60764),
            .I(N__60742));
    LocalMux I__12048 (
            .O(N__60761),
            .I(\pc_rx.r_SM_Main_0 ));
    Odrv4 I__12047 (
            .O(N__60754),
            .I(\pc_rx.r_SM_Main_0 ));
    LocalMux I__12046 (
            .O(N__60751),
            .I(\pc_rx.r_SM_Main_0 ));
    LocalMux I__12045 (
            .O(N__60742),
            .I(\pc_rx.r_SM_Main_0 ));
    InMux I__12044 (
            .O(N__60733),
            .I(N__60730));
    LocalMux I__12043 (
            .O(N__60730),
            .I(N__60727));
    Span4Mux_v I__12042 (
            .O(N__60727),
            .I(N__60718));
    InMux I__12041 (
            .O(N__60726),
            .I(N__60713));
    InMux I__12040 (
            .O(N__60725),
            .I(N__60713));
    InMux I__12039 (
            .O(N__60724),
            .I(N__60710));
    InMux I__12038 (
            .O(N__60723),
            .I(N__60707));
    InMux I__12037 (
            .O(N__60722),
            .I(N__60702));
    InMux I__12036 (
            .O(N__60721),
            .I(N__60702));
    Span4Mux_h I__12035 (
            .O(N__60718),
            .I(N__60694));
    LocalMux I__12034 (
            .O(N__60713),
            .I(N__60691));
    LocalMux I__12033 (
            .O(N__60710),
            .I(N__60684));
    LocalMux I__12032 (
            .O(N__60707),
            .I(N__60684));
    LocalMux I__12031 (
            .O(N__60702),
            .I(N__60684));
    InMux I__12030 (
            .O(N__60701),
            .I(N__60675));
    InMux I__12029 (
            .O(N__60700),
            .I(N__60675));
    InMux I__12028 (
            .O(N__60699),
            .I(N__60675));
    InMux I__12027 (
            .O(N__60698),
            .I(N__60675));
    InMux I__12026 (
            .O(N__60697),
            .I(N__60672));
    Odrv4 I__12025 (
            .O(N__60694),
            .I(r_Rx_Data));
    Odrv12 I__12024 (
            .O(N__60691),
            .I(r_Rx_Data));
    Odrv12 I__12023 (
            .O(N__60684),
            .I(r_Rx_Data));
    LocalMux I__12022 (
            .O(N__60675),
            .I(r_Rx_Data));
    LocalMux I__12021 (
            .O(N__60672),
            .I(r_Rx_Data));
    InMux I__12020 (
            .O(N__60661),
            .I(N__60657));
    InMux I__12019 (
            .O(N__60660),
            .I(N__60654));
    LocalMux I__12018 (
            .O(N__60657),
            .I(\pc_rx.n13 ));
    LocalMux I__12017 (
            .O(N__60654),
            .I(\pc_rx.n13 ));
    CascadeMux I__12016 (
            .O(N__60649),
            .I(N__60646));
    InMux I__12015 (
            .O(N__60646),
            .I(N__60643));
    LocalMux I__12014 (
            .O(N__60643),
            .I(N__60640));
    Odrv4 I__12013 (
            .O(N__60640),
            .I(\pc_rx.n125 ));
    InMux I__12012 (
            .O(N__60637),
            .I(N__60634));
    LocalMux I__12011 (
            .O(N__60634),
            .I(N__60631));
    Span4Mux_v I__12010 (
            .O(N__60631),
            .I(N__60628));
    Odrv4 I__12009 (
            .O(N__60628),
            .I(FIFO_D4_c_4));
    InMux I__12008 (
            .O(N__60625),
            .I(N__60622));
    LocalMux I__12007 (
            .O(N__60622),
            .I(N__60619));
    Span12Mux_h I__12006 (
            .O(N__60619),
            .I(N__60616));
    Odrv12 I__12005 (
            .O(N__60616),
            .I(FIFO_D5_c_5));
    InMux I__12004 (
            .O(N__60613),
            .I(N__60610));
    LocalMux I__12003 (
            .O(N__60610),
            .I(N__60607));
    Span4Mux_h I__12002 (
            .O(N__60607),
            .I(N__60604));
    Span4Mux_h I__12001 (
            .O(N__60604),
            .I(N__60601));
    Sp12to4 I__12000 (
            .O(N__60601),
            .I(N__60598));
    Odrv12 I__11999 (
            .O(N__60598),
            .I(FIFO_D6_c_6));
    InMux I__11998 (
            .O(N__60595),
            .I(N__60592));
    LocalMux I__11997 (
            .O(N__60592),
            .I(N__60589));
    Span4Mux_h I__11996 (
            .O(N__60589),
            .I(N__60586));
    Span4Mux_v I__11995 (
            .O(N__60586),
            .I(N__60583));
    Odrv4 I__11994 (
            .O(N__60583),
            .I(FIFO_D3_c_3));
    InMux I__11993 (
            .O(N__60580),
            .I(N__60576));
    InMux I__11992 (
            .O(N__60579),
            .I(N__60573));
    LocalMux I__11991 (
            .O(N__60576),
            .I(\pc_rx.r_Clock_Count_8 ));
    LocalMux I__11990 (
            .O(N__60573),
            .I(\pc_rx.r_Clock_Count_8 ));
    InMux I__11989 (
            .O(N__60568),
            .I(N__60564));
    InMux I__11988 (
            .O(N__60567),
            .I(N__60561));
    LocalMux I__11987 (
            .O(N__60564),
            .I(\pc_rx.r_Clock_Count_7 ));
    LocalMux I__11986 (
            .O(N__60561),
            .I(\pc_rx.r_Clock_Count_7 ));
    InMux I__11985 (
            .O(N__60556),
            .I(N__60553));
    LocalMux I__11984 (
            .O(N__60553),
            .I(\pc_rx.n6 ));
    InMux I__11983 (
            .O(N__60550),
            .I(N__60543));
    InMux I__11982 (
            .O(N__60549),
            .I(N__60543));
    InMux I__11981 (
            .O(N__60548),
            .I(N__60540));
    LocalMux I__11980 (
            .O(N__60543),
            .I(\pc_rx.r_Clock_Count_4 ));
    LocalMux I__11979 (
            .O(N__60540),
            .I(\pc_rx.r_Clock_Count_4 ));
    InMux I__11978 (
            .O(N__60535),
            .I(N__60528));
    InMux I__11977 (
            .O(N__60534),
            .I(N__60528));
    InMux I__11976 (
            .O(N__60533),
            .I(N__60525));
    LocalMux I__11975 (
            .O(N__60528),
            .I(\pc_rx.r_Clock_Count_1 ));
    LocalMux I__11974 (
            .O(N__60525),
            .I(\pc_rx.r_Clock_Count_1 ));
    CascadeMux I__11973 (
            .O(N__60520),
            .I(N__60517));
    InMux I__11972 (
            .O(N__60517),
            .I(N__60510));
    InMux I__11971 (
            .O(N__60516),
            .I(N__60510));
    InMux I__11970 (
            .O(N__60515),
            .I(N__60507));
    LocalMux I__11969 (
            .O(N__60510),
            .I(\pc_rx.r_Clock_Count_0 ));
    LocalMux I__11968 (
            .O(N__60507),
            .I(\pc_rx.r_Clock_Count_0 ));
    InMux I__11967 (
            .O(N__60502),
            .I(N__60495));
    InMux I__11966 (
            .O(N__60501),
            .I(N__60495));
    InMux I__11965 (
            .O(N__60500),
            .I(N__60492));
    LocalMux I__11964 (
            .O(N__60495),
            .I(\pc_rx.r_Clock_Count_3 ));
    LocalMux I__11963 (
            .O(N__60492),
            .I(\pc_rx.r_Clock_Count_3 ));
    InMux I__11962 (
            .O(N__60487),
            .I(N__60481));
    InMux I__11961 (
            .O(N__60486),
            .I(N__60481));
    LocalMux I__11960 (
            .O(N__60481),
            .I(\pc_rx.n140 ));
    CascadeMux I__11959 (
            .O(N__60478),
            .I(\pc_rx.n8_cascade_ ));
    InMux I__11958 (
            .O(N__60475),
            .I(N__60468));
    InMux I__11957 (
            .O(N__60474),
            .I(N__60468));
    InMux I__11956 (
            .O(N__60473),
            .I(N__60465));
    LocalMux I__11955 (
            .O(N__60468),
            .I(\pc_rx.r_Clock_Count_2 ));
    LocalMux I__11954 (
            .O(N__60465),
            .I(\pc_rx.r_Clock_Count_2 ));
    CascadeMux I__11953 (
            .O(N__60460),
            .I(\pc_rx.n13_cascade_ ));
    InMux I__11952 (
            .O(N__60457),
            .I(N__60454));
    LocalMux I__11951 (
            .O(N__60454),
            .I(\pc_rx.n6500 ));
    InMux I__11950 (
            .O(N__60451),
            .I(N__60448));
    LocalMux I__11949 (
            .O(N__60448),
            .I(\pc_rx.n145 ));
    CascadeMux I__11948 (
            .O(N__60445),
            .I(\pc_rx.n145_cascade_ ));
    CEMux I__11947 (
            .O(N__60442),
            .I(N__60439));
    LocalMux I__11946 (
            .O(N__60439),
            .I(N__60436));
    Span4Mux_v I__11945 (
            .O(N__60436),
            .I(N__60432));
    CEMux I__11944 (
            .O(N__60435),
            .I(N__60429));
    Odrv4 I__11943 (
            .O(N__60432),
            .I(\pc_rx.n6490 ));
    LocalMux I__11942 (
            .O(N__60429),
            .I(\pc_rx.n6490 ));
    CascadeMux I__11941 (
            .O(N__60424),
            .I(N__60421));
    InMux I__11940 (
            .O(N__60421),
            .I(N__60418));
    LocalMux I__11939 (
            .O(N__60418),
            .I(\pc_rx.n4081 ));
    InMux I__11938 (
            .O(N__60415),
            .I(N__60411));
    CEMux I__11937 (
            .O(N__60414),
            .I(N__60408));
    LocalMux I__11936 (
            .O(N__60411),
            .I(N__60404));
    LocalMux I__11935 (
            .O(N__60408),
            .I(N__60401));
    InMux I__11934 (
            .O(N__60407),
            .I(N__60398));
    Span4Mux_v I__11933 (
            .O(N__60404),
            .I(N__60395));
    Span4Mux_h I__11932 (
            .O(N__60401),
            .I(N__60392));
    LocalMux I__11931 (
            .O(N__60398),
            .I(\pc_rx.n4140 ));
    Odrv4 I__11930 (
            .O(N__60395),
            .I(\pc_rx.n4140 ));
    Odrv4 I__11929 (
            .O(N__60392),
            .I(\pc_rx.n4140 ));
    InMux I__11928 (
            .O(N__60385),
            .I(N__60379));
    InMux I__11927 (
            .O(N__60384),
            .I(N__60379));
    LocalMux I__11926 (
            .O(N__60379),
            .I(N__60374));
    InMux I__11925 (
            .O(N__60378),
            .I(N__60369));
    InMux I__11924 (
            .O(N__60377),
            .I(N__60369));
    Span4Mux_v I__11923 (
            .O(N__60374),
            .I(N__60366));
    LocalMux I__11922 (
            .O(N__60369),
            .I(N__60363));
    Odrv4 I__11921 (
            .O(N__60366),
            .I(\pc_rx.n151 ));
    Odrv12 I__11920 (
            .O(N__60363),
            .I(\pc_rx.n151 ));
    InMux I__11919 (
            .O(N__60358),
            .I(N__60353));
    CascadeMux I__11918 (
            .O(N__60357),
            .I(N__60346));
    InMux I__11917 (
            .O(N__60356),
            .I(N__60340));
    LocalMux I__11916 (
            .O(N__60353),
            .I(N__60337));
    InMux I__11915 (
            .O(N__60352),
            .I(N__60334));
    InMux I__11914 (
            .O(N__60351),
            .I(N__60331));
    InMux I__11913 (
            .O(N__60350),
            .I(N__60318));
    InMux I__11912 (
            .O(N__60349),
            .I(N__60318));
    InMux I__11911 (
            .O(N__60346),
            .I(N__60318));
    InMux I__11910 (
            .O(N__60345),
            .I(N__60318));
    InMux I__11909 (
            .O(N__60344),
            .I(N__60318));
    InMux I__11908 (
            .O(N__60343),
            .I(N__60318));
    LocalMux I__11907 (
            .O(N__60340),
            .I(\pc_rx.r_SM_Main_1 ));
    Odrv4 I__11906 (
            .O(N__60337),
            .I(\pc_rx.r_SM_Main_1 ));
    LocalMux I__11905 (
            .O(N__60334),
            .I(\pc_rx.r_SM_Main_1 ));
    LocalMux I__11904 (
            .O(N__60331),
            .I(\pc_rx.r_SM_Main_1 ));
    LocalMux I__11903 (
            .O(N__60318),
            .I(\pc_rx.r_SM_Main_1 ));
    InMux I__11902 (
            .O(N__60307),
            .I(N__60304));
    LocalMux I__11901 (
            .O(N__60304),
            .I(\pc_rx.n6515 ));
    InMux I__11900 (
            .O(N__60301),
            .I(N__60290));
    InMux I__11899 (
            .O(N__60300),
            .I(N__60290));
    InMux I__11898 (
            .O(N__60299),
            .I(N__60279));
    InMux I__11897 (
            .O(N__60298),
            .I(N__60279));
    InMux I__11896 (
            .O(N__60297),
            .I(N__60279));
    InMux I__11895 (
            .O(N__60296),
            .I(N__60279));
    SRMux I__11894 (
            .O(N__60295),
            .I(N__60279));
    LocalMux I__11893 (
            .O(N__60290),
            .I(N__60274));
    LocalMux I__11892 (
            .O(N__60279),
            .I(N__60274));
    Odrv4 I__11891 (
            .O(N__60274),
            .I(\pc_rx.r_SM_Main_2 ));
    InMux I__11890 (
            .O(N__60271),
            .I(N__60267));
    InMux I__11889 (
            .O(N__60270),
            .I(N__60264));
    LocalMux I__11888 (
            .O(N__60267),
            .I(\pc_rx.r_Clock_Count_9 ));
    LocalMux I__11887 (
            .O(N__60264),
            .I(\pc_rx.r_Clock_Count_9 ));
    CascadeMux I__11886 (
            .O(N__60259),
            .I(N__60256));
    InMux I__11885 (
            .O(N__60256),
            .I(N__60252));
    InMux I__11884 (
            .O(N__60255),
            .I(N__60249));
    LocalMux I__11883 (
            .O(N__60252),
            .I(\pc_rx.r_Clock_Count_6 ));
    LocalMux I__11882 (
            .O(N__60249),
            .I(\pc_rx.r_Clock_Count_6 ));
    InMux I__11881 (
            .O(N__60244),
            .I(N__60240));
    InMux I__11880 (
            .O(N__60243),
            .I(N__60237));
    LocalMux I__11879 (
            .O(N__60240),
            .I(\pc_rx.r_Clock_Count_5 ));
    LocalMux I__11878 (
            .O(N__60237),
            .I(\pc_rx.r_Clock_Count_5 ));
    CascadeMux I__11877 (
            .O(N__60232),
            .I(\pc_rx.n4_adj_1145_cascade_ ));
    InMux I__11876 (
            .O(N__60229),
            .I(N__60226));
    LocalMux I__11875 (
            .O(N__60226),
            .I(N__60218));
    InMux I__11874 (
            .O(N__60225),
            .I(N__60215));
    InMux I__11873 (
            .O(N__60224),
            .I(N__60206));
    InMux I__11872 (
            .O(N__60223),
            .I(N__60206));
    InMux I__11871 (
            .O(N__60222),
            .I(N__60206));
    InMux I__11870 (
            .O(N__60221),
            .I(N__60206));
    Odrv4 I__11869 (
            .O(N__60218),
            .I(\pc_rx.r_SM_Main_2_N_732_2 ));
    LocalMux I__11868 (
            .O(N__60215),
            .I(\pc_rx.r_SM_Main_2_N_732_2 ));
    LocalMux I__11867 (
            .O(N__60206),
            .I(\pc_rx.r_SM_Main_2_N_732_2 ));
    InMux I__11866 (
            .O(N__60199),
            .I(N__60196));
    LocalMux I__11865 (
            .O(N__60196),
            .I(N__60193));
    Span4Mux_h I__11864 (
            .O(N__60193),
            .I(N__60190));
    Sp12to4 I__11863 (
            .O(N__60190),
            .I(N__60187));
    Span12Mux_v I__11862 (
            .O(N__60187),
            .I(N__60184));
    Span12Mux_v I__11861 (
            .O(N__60184),
            .I(N__60181));
    Span12Mux_h I__11860 (
            .O(N__60181),
            .I(N__60178));
    Odrv12 I__11859 (
            .O(N__60178),
            .I(\pc_rx.r_Rx_Data_R ));
    InMux I__11858 (
            .O(N__60175),
            .I(N__60169));
    InMux I__11857 (
            .O(N__60174),
            .I(N__60169));
    LocalMux I__11856 (
            .O(N__60169),
            .I(N__60165));
    CascadeMux I__11855 (
            .O(N__60168),
            .I(N__60162));
    Span4Mux_h I__11854 (
            .O(N__60165),
            .I(N__60159));
    InMux I__11853 (
            .O(N__60162),
            .I(N__60156));
    Odrv4 I__11852 (
            .O(N__60159),
            .I(n4002));
    LocalMux I__11851 (
            .O(N__60156),
            .I(n4002));
    CascadeMux I__11850 (
            .O(N__60151),
            .I(n4002_cascade_));
    InMux I__11849 (
            .O(N__60148),
            .I(N__60144));
    InMux I__11848 (
            .O(N__60147),
            .I(N__60141));
    LocalMux I__11847 (
            .O(N__60144),
            .I(n4));
    LocalMux I__11846 (
            .O(N__60141),
            .I(n4));
    InMux I__11845 (
            .O(N__60136),
            .I(N__60133));
    LocalMux I__11844 (
            .O(N__60133),
            .I(N__60129));
    InMux I__11843 (
            .O(N__60132),
            .I(N__60126));
    Odrv4 I__11842 (
            .O(N__60129),
            .I(pc_data_rx_3));
    LocalMux I__11841 (
            .O(N__60126),
            .I(pc_data_rx_3));
    CascadeMux I__11840 (
            .O(N__60121),
            .I(N__60118));
    InMux I__11839 (
            .O(N__60118),
            .I(N__60115));
    LocalMux I__11838 (
            .O(N__60115),
            .I(N__60112));
    Span4Mux_h I__11837 (
            .O(N__60112),
            .I(N__60109));
    Odrv4 I__11836 (
            .O(N__60109),
            .I(REG_out_raw_1));
    InMux I__11835 (
            .O(N__60106),
            .I(N__60090));
    InMux I__11834 (
            .O(N__60105),
            .I(N__60090));
    InMux I__11833 (
            .O(N__60104),
            .I(N__60090));
    InMux I__11832 (
            .O(N__60103),
            .I(N__60090));
    InMux I__11831 (
            .O(N__60102),
            .I(N__60090));
    InMux I__11830 (
            .O(N__60101),
            .I(N__60087));
    LocalMux I__11829 (
            .O(N__60090),
            .I(\pc_rx.r_Bit_Index_2 ));
    LocalMux I__11828 (
            .O(N__60087),
            .I(\pc_rx.r_Bit_Index_2 ));
    InMux I__11827 (
            .O(N__60082),
            .I(N__60076));
    InMux I__11826 (
            .O(N__60081),
            .I(N__60076));
    LocalMux I__11825 (
            .O(N__60076),
            .I(N__60073));
    Span4Mux_v I__11824 (
            .O(N__60073),
            .I(N__60065));
    InMux I__11823 (
            .O(N__60072),
            .I(N__60062));
    InMux I__11822 (
            .O(N__60071),
            .I(N__60057));
    InMux I__11821 (
            .O(N__60070),
            .I(N__60057));
    InMux I__11820 (
            .O(N__60069),
            .I(N__60052));
    InMux I__11819 (
            .O(N__60068),
            .I(N__60052));
    Odrv4 I__11818 (
            .O(N__60065),
            .I(\pc_rx.r_Bit_Index_0 ));
    LocalMux I__11817 (
            .O(N__60062),
            .I(\pc_rx.r_Bit_Index_0 ));
    LocalMux I__11816 (
            .O(N__60057),
            .I(\pc_rx.r_Bit_Index_0 ));
    LocalMux I__11815 (
            .O(N__60052),
            .I(\pc_rx.r_Bit_Index_0 ));
    InMux I__11814 (
            .O(N__60043),
            .I(N__60026));
    InMux I__11813 (
            .O(N__60042),
            .I(N__60026));
    InMux I__11812 (
            .O(N__60041),
            .I(N__60026));
    InMux I__11811 (
            .O(N__60040),
            .I(N__60026));
    InMux I__11810 (
            .O(N__60039),
            .I(N__60026));
    InMux I__11809 (
            .O(N__60038),
            .I(N__60021));
    InMux I__11808 (
            .O(N__60037),
            .I(N__60021));
    LocalMux I__11807 (
            .O(N__60026),
            .I(\pc_rx.r_Bit_Index_1 ));
    LocalMux I__11806 (
            .O(N__60021),
            .I(\pc_rx.r_Bit_Index_1 ));
    SRMux I__11805 (
            .O(N__60016),
            .I(N__60013));
    LocalMux I__11804 (
            .O(N__60013),
            .I(N__60010));
    Sp12to4 I__11803 (
            .O(N__60010),
            .I(N__60007));
    Odrv12 I__11802 (
            .O(N__60007),
            .I(\pc_rx.n4470 ));
    CascadeMux I__11801 (
            .O(N__60004),
            .I(\pc_rx.n55_adj_1144_cascade_ ));
    InMux I__11800 (
            .O(N__60001),
            .I(N__59998));
    LocalMux I__11799 (
            .O(N__59998),
            .I(N__59994));
    InMux I__11798 (
            .O(N__59997),
            .I(N__59991));
    Odrv4 I__11797 (
            .O(N__59994),
            .I(\bluejay_data_inst.state_timeout_counter_6 ));
    LocalMux I__11796 (
            .O(N__59991),
            .I(\bluejay_data_inst.state_timeout_counter_6 ));
    InMux I__11795 (
            .O(N__59986),
            .I(bfn_16_15_0_));
    InMux I__11794 (
            .O(N__59983),
            .I(\bluejay_data_inst.n10587 ));
    InMux I__11793 (
            .O(N__59980),
            .I(N__59977));
    LocalMux I__11792 (
            .O(N__59977),
            .I(N__59973));
    InMux I__11791 (
            .O(N__59976),
            .I(N__59970));
    Odrv4 I__11790 (
            .O(N__59973),
            .I(\bluejay_data_inst.state_timeout_counter_7 ));
    LocalMux I__11789 (
            .O(N__59970),
            .I(\bluejay_data_inst.state_timeout_counter_7 ));
    SRMux I__11788 (
            .O(N__59965),
            .I(N__59962));
    LocalMux I__11787 (
            .O(N__59962),
            .I(N__59959));
    Span4Mux_h I__11786 (
            .O(N__59959),
            .I(N__59956));
    Odrv4 I__11785 (
            .O(N__59956),
            .I(\bluejay_data_inst.n11177 ));
    InMux I__11784 (
            .O(N__59953),
            .I(N__59949));
    InMux I__11783 (
            .O(N__59952),
            .I(N__59946));
    LocalMux I__11782 (
            .O(N__59949),
            .I(\bluejay_data_inst.state_timeout_counter_5 ));
    LocalMux I__11781 (
            .O(N__59946),
            .I(\bluejay_data_inst.state_timeout_counter_5 ));
    InMux I__11780 (
            .O(N__59941),
            .I(bfn_16_14_0_));
    InMux I__11779 (
            .O(N__59938),
            .I(bfn_16_12_0_));
    InMux I__11778 (
            .O(N__59935),
            .I(bfn_16_13_0_));
    CascadeMux I__11777 (
            .O(N__59932),
            .I(N__59929));
    InMux I__11776 (
            .O(N__59929),
            .I(N__59926));
    LocalMux I__11775 (
            .O(N__59926),
            .I(N__59922));
    InMux I__11774 (
            .O(N__59925),
            .I(N__59919));
    Odrv12 I__11773 (
            .O(N__59922),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_4 ));
    LocalMux I__11772 (
            .O(N__59919),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_4 ));
    InMux I__11771 (
            .O(N__59914),
            .I(N__59911));
    LocalMux I__11770 (
            .O(N__59911),
            .I(N__59908));
    Span12Mux_v I__11769 (
            .O(N__59908),
            .I(N__59904));
    InMux I__11768 (
            .O(N__59907),
            .I(N__59901));
    Odrv12 I__11767 (
            .O(N__59904),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_4 ));
    LocalMux I__11766 (
            .O(N__59901),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_4 ));
    InMux I__11765 (
            .O(N__59896),
            .I(bfn_16_11_0_));
    InMux I__11764 (
            .O(N__59893),
            .I(N__59890));
    LocalMux I__11763 (
            .O(N__59890),
            .I(N__59887));
    Span4Mux_v I__11762 (
            .O(N__59887),
            .I(N__59883));
    InMux I__11761 (
            .O(N__59886),
            .I(N__59880));
    Odrv4 I__11760 (
            .O(N__59883),
            .I(\bluejay_data_inst.state_timeout_counter_1 ));
    LocalMux I__11759 (
            .O(N__59880),
            .I(\bluejay_data_inst.state_timeout_counter_1 ));
    InMux I__11758 (
            .O(N__59875),
            .I(\bluejay_data_inst.n10581 ));
    InMux I__11757 (
            .O(N__59872),
            .I(N__59869));
    LocalMux I__11756 (
            .O(N__59869),
            .I(N__59865));
    InMux I__11755 (
            .O(N__59868),
            .I(N__59862));
    Odrv4 I__11754 (
            .O(N__59865),
            .I(\bluejay_data_inst.state_timeout_counter_2 ));
    LocalMux I__11753 (
            .O(N__59862),
            .I(\bluejay_data_inst.state_timeout_counter_2 ));
    InMux I__11752 (
            .O(N__59857),
            .I(N__59854));
    LocalMux I__11751 (
            .O(N__59854),
            .I(N__59851));
    Odrv4 I__11750 (
            .O(N__59851),
            .I(\bluejay_data_inst.n86 ));
    InMux I__11749 (
            .O(N__59848),
            .I(\bluejay_data_inst.n10582 ));
    InMux I__11748 (
            .O(N__59845),
            .I(N__59842));
    LocalMux I__11747 (
            .O(N__59842),
            .I(N__59839));
    Span4Mux_h I__11746 (
            .O(N__59839),
            .I(N__59836));
    Span4Mux_v I__11745 (
            .O(N__59836),
            .I(N__59832));
    InMux I__11744 (
            .O(N__59835),
            .I(N__59829));
    Odrv4 I__11743 (
            .O(N__59832),
            .I(REG_mem_55_7));
    LocalMux I__11742 (
            .O(N__59829),
            .I(REG_mem_55_7));
    InMux I__11741 (
            .O(N__59824),
            .I(N__59821));
    LocalMux I__11740 (
            .O(N__59821),
            .I(N__59818));
    Span4Mux_h I__11739 (
            .O(N__59818),
            .I(N__59815));
    Span4Mux_v I__11738 (
            .O(N__59815),
            .I(N__59812));
    Odrv4 I__11737 (
            .O(N__59812),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13718 ));
    CascadeMux I__11736 (
            .O(N__59809),
            .I(N__59806));
    InMux I__11735 (
            .O(N__59806),
            .I(N__59802));
    CascadeMux I__11734 (
            .O(N__59805),
            .I(N__59799));
    LocalMux I__11733 (
            .O(N__59802),
            .I(N__59796));
    InMux I__11732 (
            .O(N__59799),
            .I(N__59793));
    Odrv4 I__11731 (
            .O(N__59796),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_7 ));
    LocalMux I__11730 (
            .O(N__59793),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_7 ));
    CascadeMux I__11729 (
            .O(N__59788),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13736_cascade_ ));
    CascadeMux I__11728 (
            .O(N__59785),
            .I(N__59781));
    InMux I__11727 (
            .O(N__59784),
            .I(N__59776));
    InMux I__11726 (
            .O(N__59781),
            .I(N__59776));
    LocalMux I__11725 (
            .O(N__59776),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_4 ));
    CascadeMux I__11724 (
            .O(N__59773),
            .I(N__59769));
    InMux I__11723 (
            .O(N__59772),
            .I(N__59764));
    InMux I__11722 (
            .O(N__59769),
            .I(N__59764));
    LocalMux I__11721 (
            .O(N__59764),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_4 ));
    CascadeMux I__11720 (
            .O(N__59761),
            .I(N__59757));
    CascadeMux I__11719 (
            .O(N__59760),
            .I(N__59754));
    InMux I__11718 (
            .O(N__59757),
            .I(N__59749));
    InMux I__11717 (
            .O(N__59754),
            .I(N__59749));
    LocalMux I__11716 (
            .O(N__59749),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_4 ));
    InMux I__11715 (
            .O(N__59746),
            .I(N__59740));
    InMux I__11714 (
            .O(N__59745),
            .I(N__59740));
    LocalMux I__11713 (
            .O(N__59740),
            .I(REG_mem_51_7));
    InMux I__11712 (
            .O(N__59737),
            .I(N__59734));
    LocalMux I__11711 (
            .O(N__59734),
            .I(N__59731));
    Span4Mux_h I__11710 (
            .O(N__59731),
            .I(N__59728));
    Sp12to4 I__11709 (
            .O(N__59728),
            .I(N__59724));
    InMux I__11708 (
            .O(N__59727),
            .I(N__59721));
    Odrv12 I__11707 (
            .O(N__59724),
            .I(REG_mem_15_8));
    LocalMux I__11706 (
            .O(N__59721),
            .I(REG_mem_15_8));
    InMux I__11705 (
            .O(N__59716),
            .I(N__59713));
    LocalMux I__11704 (
            .O(N__59713),
            .I(N__59709));
    InMux I__11703 (
            .O(N__59712),
            .I(N__59706));
    Odrv12 I__11702 (
            .O(N__59709),
            .I(REG_mem_13_5));
    LocalMux I__11701 (
            .O(N__59706),
            .I(REG_mem_13_5));
    InMux I__11700 (
            .O(N__59701),
            .I(N__59698));
    LocalMux I__11699 (
            .O(N__59698),
            .I(N__59695));
    Span4Mux_h I__11698 (
            .O(N__59695),
            .I(N__59691));
    InMux I__11697 (
            .O(N__59694),
            .I(N__59688));
    Odrv4 I__11696 (
            .O(N__59691),
            .I(REG_mem_49_8));
    LocalMux I__11695 (
            .O(N__59688),
            .I(REG_mem_49_8));
    CascadeMux I__11694 (
            .O(N__59683),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13532_cascade_ ));
    InMux I__11693 (
            .O(N__59680),
            .I(N__59674));
    InMux I__11692 (
            .O(N__59679),
            .I(N__59674));
    LocalMux I__11691 (
            .O(N__59674),
            .I(REG_mem_48_8));
    InMux I__11690 (
            .O(N__59671),
            .I(N__59665));
    InMux I__11689 (
            .O(N__59670),
            .I(N__59665));
    LocalMux I__11688 (
            .O(N__59665),
            .I(REG_mem_51_8));
    InMux I__11687 (
            .O(N__59662),
            .I(N__59659));
    LocalMux I__11686 (
            .O(N__59659),
            .I(N__59654));
    InMux I__11685 (
            .O(N__59658),
            .I(N__59648));
    InMux I__11684 (
            .O(N__59657),
            .I(N__59645));
    Span4Mux_h I__11683 (
            .O(N__59654),
            .I(N__59641));
    InMux I__11682 (
            .O(N__59653),
            .I(N__59638));
    InMux I__11681 (
            .O(N__59652),
            .I(N__59635));
    InMux I__11680 (
            .O(N__59651),
            .I(N__59629));
    LocalMux I__11679 (
            .O(N__59648),
            .I(N__59626));
    LocalMux I__11678 (
            .O(N__59645),
            .I(N__59623));
    InMux I__11677 (
            .O(N__59644),
            .I(N__59620));
    Span4Mux_h I__11676 (
            .O(N__59641),
            .I(N__59615));
    LocalMux I__11675 (
            .O(N__59638),
            .I(N__59615));
    LocalMux I__11674 (
            .O(N__59635),
            .I(N__59612));
    InMux I__11673 (
            .O(N__59634),
            .I(N__59608));
    InMux I__11672 (
            .O(N__59633),
            .I(N__59605));
    InMux I__11671 (
            .O(N__59632),
            .I(N__59602));
    LocalMux I__11670 (
            .O(N__59629),
            .I(N__59597));
    Span4Mux_v I__11669 (
            .O(N__59626),
            .I(N__59594));
    Span4Mux_v I__11668 (
            .O(N__59623),
            .I(N__59589));
    LocalMux I__11667 (
            .O(N__59620),
            .I(N__59589));
    Span4Mux_h I__11666 (
            .O(N__59615),
            .I(N__59586));
    Span4Mux_v I__11665 (
            .O(N__59612),
            .I(N__59583));
    InMux I__11664 (
            .O(N__59611),
            .I(N__59580));
    LocalMux I__11663 (
            .O(N__59608),
            .I(N__59577));
    LocalMux I__11662 (
            .O(N__59605),
            .I(N__59572));
    LocalMux I__11661 (
            .O(N__59602),
            .I(N__59572));
    InMux I__11660 (
            .O(N__59601),
            .I(N__59569));
    InMux I__11659 (
            .O(N__59600),
            .I(N__59566));
    Span12Mux_s11_v I__11658 (
            .O(N__59597),
            .I(N__59561));
    Span4Mux_h I__11657 (
            .O(N__59594),
            .I(N__59554));
    Span4Mux_v I__11656 (
            .O(N__59589),
            .I(N__59554));
    Span4Mux_v I__11655 (
            .O(N__59586),
            .I(N__59554));
    Sp12to4 I__11654 (
            .O(N__59583),
            .I(N__59549));
    LocalMux I__11653 (
            .O(N__59580),
            .I(N__59549));
    Span4Mux_h I__11652 (
            .O(N__59577),
            .I(N__59546));
    Span4Mux_v I__11651 (
            .O(N__59572),
            .I(N__59541));
    LocalMux I__11650 (
            .O(N__59569),
            .I(N__59541));
    LocalMux I__11649 (
            .O(N__59566),
            .I(N__59538));
    InMux I__11648 (
            .O(N__59565),
            .I(N__59535));
    InMux I__11647 (
            .O(N__59564),
            .I(N__59532));
    Odrv12 I__11646 (
            .O(N__59561),
            .I(n53));
    Odrv4 I__11645 (
            .O(N__59554),
            .I(n53));
    Odrv12 I__11644 (
            .O(N__59549),
            .I(n53));
    Odrv4 I__11643 (
            .O(N__59546),
            .I(n53));
    Odrv4 I__11642 (
            .O(N__59541),
            .I(n53));
    Odrv4 I__11641 (
            .O(N__59538),
            .I(n53));
    LocalMux I__11640 (
            .O(N__59535),
            .I(n53));
    LocalMux I__11639 (
            .O(N__59532),
            .I(n53));
    InMux I__11638 (
            .O(N__59515),
            .I(N__59509));
    InMux I__11637 (
            .O(N__59514),
            .I(N__59509));
    LocalMux I__11636 (
            .O(N__59509),
            .I(N__59506));
    Odrv4 I__11635 (
            .O(N__59506),
            .I(REG_mem_12_4));
    InMux I__11634 (
            .O(N__59503),
            .I(N__59500));
    LocalMux I__11633 (
            .O(N__59500),
            .I(N__59497));
    Span4Mux_v I__11632 (
            .O(N__59497),
            .I(N__59494));
    Odrv4 I__11631 (
            .O(N__59494),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11638 ));
    InMux I__11630 (
            .O(N__59491),
            .I(N__59488));
    LocalMux I__11629 (
            .O(N__59488),
            .I(N__59485));
    Span4Mux_v I__11628 (
            .O(N__59485),
            .I(N__59482));
    Span4Mux_h I__11627 (
            .O(N__59482),
            .I(N__59479));
    Span4Mux_h I__11626 (
            .O(N__59479),
            .I(N__59475));
    InMux I__11625 (
            .O(N__59478),
            .I(N__59472));
    Odrv4 I__11624 (
            .O(N__59475),
            .I(REG_mem_12_2));
    LocalMux I__11623 (
            .O(N__59472),
            .I(REG_mem_12_2));
    CascadeMux I__11622 (
            .O(N__59467),
            .I(N__59464));
    InMux I__11621 (
            .O(N__59464),
            .I(N__59461));
    LocalMux I__11620 (
            .O(N__59461),
            .I(N__59457));
    InMux I__11619 (
            .O(N__59460),
            .I(N__59454));
    Odrv4 I__11618 (
            .O(N__59457),
            .I(REG_mem_50_7));
    LocalMux I__11617 (
            .O(N__59454),
            .I(REG_mem_50_7));
    InMux I__11616 (
            .O(N__59449),
            .I(N__59443));
    InMux I__11615 (
            .O(N__59448),
            .I(N__59443));
    LocalMux I__11614 (
            .O(N__59443),
            .I(REG_mem_49_7));
    CascadeMux I__11613 (
            .O(N__59440),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13760_cascade_ ));
    InMux I__11612 (
            .O(N__59437),
            .I(N__59434));
    LocalMux I__11611 (
            .O(N__59434),
            .I(N__59431));
    Span4Mux_v I__11610 (
            .O(N__59431),
            .I(N__59428));
    Span4Mux_v I__11609 (
            .O(N__59428),
            .I(N__59425));
    Span4Mux_h I__11608 (
            .O(N__59425),
            .I(N__59422));
    Odrv4 I__11607 (
            .O(N__59422),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12210 ));
    InMux I__11606 (
            .O(N__59419),
            .I(N__59413));
    InMux I__11605 (
            .O(N__59418),
            .I(N__59413));
    LocalMux I__11604 (
            .O(N__59413),
            .I(REG_mem_48_7));
    InMux I__11603 (
            .O(N__59410),
            .I(N__59407));
    LocalMux I__11602 (
            .O(N__59407),
            .I(N__59403));
    InMux I__11601 (
            .O(N__59406),
            .I(N__59400));
    Odrv4 I__11600 (
            .O(N__59403),
            .I(REG_mem_11_8));
    LocalMux I__11599 (
            .O(N__59400),
            .I(REG_mem_11_8));
    InMux I__11598 (
            .O(N__59395),
            .I(N__59392));
    LocalMux I__11597 (
            .O(N__59392),
            .I(N__59389));
    Span4Mux_h I__11596 (
            .O(N__59389),
            .I(N__59386));
    Sp12to4 I__11595 (
            .O(N__59386),
            .I(N__59382));
    InMux I__11594 (
            .O(N__59385),
            .I(N__59379));
    Odrv12 I__11593 (
            .O(N__59382),
            .I(REG_mem_10_8));
    LocalMux I__11592 (
            .O(N__59379),
            .I(REG_mem_10_8));
    CascadeMux I__11591 (
            .O(N__59374),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13868_cascade_ ));
    CascadeMux I__11590 (
            .O(N__59371),
            .I(N__59367));
    InMux I__11589 (
            .O(N__59370),
            .I(N__59362));
    InMux I__11588 (
            .O(N__59367),
            .I(N__59362));
    LocalMux I__11587 (
            .O(N__59362),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_4 ));
    CascadeMux I__11586 (
            .O(N__59359),
            .I(N__59355));
    InMux I__11585 (
            .O(N__59358),
            .I(N__59350));
    InMux I__11584 (
            .O(N__59355),
            .I(N__59350));
    LocalMux I__11583 (
            .O(N__59350),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_4 ));
    CascadeMux I__11582 (
            .O(N__59347),
            .I(N__59343));
    InMux I__11581 (
            .O(N__59346),
            .I(N__59338));
    InMux I__11580 (
            .O(N__59343),
            .I(N__59338));
    LocalMux I__11579 (
            .O(N__59338),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_4 ));
    InMux I__11578 (
            .O(N__59335),
            .I(N__59332));
    LocalMux I__11577 (
            .O(N__59332),
            .I(N__59329));
    Span4Mux_h I__11576 (
            .O(N__59329),
            .I(N__59325));
    CascadeMux I__11575 (
            .O(N__59328),
            .I(N__59322));
    Span4Mux_h I__11574 (
            .O(N__59325),
            .I(N__59319));
    InMux I__11573 (
            .O(N__59322),
            .I(N__59316));
    Odrv4 I__11572 (
            .O(N__59319),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_0 ));
    LocalMux I__11571 (
            .O(N__59316),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_0 ));
    InMux I__11570 (
            .O(N__59311),
            .I(N__59308));
    LocalMux I__11569 (
            .O(N__59308),
            .I(N__59304));
    InMux I__11568 (
            .O(N__59307),
            .I(N__59301));
    Odrv4 I__11567 (
            .O(N__59304),
            .I(REG_mem_39_4));
    LocalMux I__11566 (
            .O(N__59301),
            .I(REG_mem_39_4));
    InMux I__11565 (
            .O(N__59296),
            .I(N__59293));
    LocalMux I__11564 (
            .O(N__59293),
            .I(N__59290));
    Sp12to4 I__11563 (
            .O(N__59290),
            .I(N__59287));
    Odrv12 I__11562 (
            .O(N__59287),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13178 ));
    InMux I__11561 (
            .O(N__59284),
            .I(N__59276));
    InMux I__11560 (
            .O(N__59283),
            .I(N__59269));
    InMux I__11559 (
            .O(N__59282),
            .I(N__59264));
    InMux I__11558 (
            .O(N__59281),
            .I(N__59264));
    InMux I__11557 (
            .O(N__59280),
            .I(N__59261));
    InMux I__11556 (
            .O(N__59279),
            .I(N__59258));
    LocalMux I__11555 (
            .O(N__59276),
            .I(N__59255));
    InMux I__11554 (
            .O(N__59275),
            .I(N__59252));
    InMux I__11553 (
            .O(N__59274),
            .I(N__59249));
    InMux I__11552 (
            .O(N__59273),
            .I(N__59244));
    InMux I__11551 (
            .O(N__59272),
            .I(N__59240));
    LocalMux I__11550 (
            .O(N__59269),
            .I(N__59236));
    LocalMux I__11549 (
            .O(N__59264),
            .I(N__59233));
    LocalMux I__11548 (
            .O(N__59261),
            .I(N__59230));
    LocalMux I__11547 (
            .O(N__59258),
            .I(N__59227));
    Span4Mux_h I__11546 (
            .O(N__59255),
            .I(N__59222));
    LocalMux I__11545 (
            .O(N__59252),
            .I(N__59222));
    LocalMux I__11544 (
            .O(N__59249),
            .I(N__59219));
    InMux I__11543 (
            .O(N__59248),
            .I(N__59216));
    InMux I__11542 (
            .O(N__59247),
            .I(N__59213));
    LocalMux I__11541 (
            .O(N__59244),
            .I(N__59210));
    InMux I__11540 (
            .O(N__59243),
            .I(N__59207));
    LocalMux I__11539 (
            .O(N__59240),
            .I(N__59203));
    InMux I__11538 (
            .O(N__59239),
            .I(N__59200));
    Span4Mux_v I__11537 (
            .O(N__59236),
            .I(N__59196));
    Span4Mux_v I__11536 (
            .O(N__59233),
            .I(N__59191));
    Span4Mux_v I__11535 (
            .O(N__59230),
            .I(N__59191));
    Span4Mux_h I__11534 (
            .O(N__59227),
            .I(N__59184));
    Span4Mux_h I__11533 (
            .O(N__59222),
            .I(N__59184));
    Span4Mux_h I__11532 (
            .O(N__59219),
            .I(N__59184));
    LocalMux I__11531 (
            .O(N__59216),
            .I(N__59179));
    LocalMux I__11530 (
            .O(N__59213),
            .I(N__59179));
    Span4Mux_v I__11529 (
            .O(N__59210),
            .I(N__59174));
    LocalMux I__11528 (
            .O(N__59207),
            .I(N__59174));
    InMux I__11527 (
            .O(N__59206),
            .I(N__59171));
    Span4Mux_h I__11526 (
            .O(N__59203),
            .I(N__59166));
    LocalMux I__11525 (
            .O(N__59200),
            .I(N__59166));
    InMux I__11524 (
            .O(N__59199),
            .I(N__59163));
    Odrv4 I__11523 (
            .O(N__59196),
            .I(n27));
    Odrv4 I__11522 (
            .O(N__59191),
            .I(n27));
    Odrv4 I__11521 (
            .O(N__59184),
            .I(n27));
    Odrv12 I__11520 (
            .O(N__59179),
            .I(n27));
    Odrv4 I__11519 (
            .O(N__59174),
            .I(n27));
    LocalMux I__11518 (
            .O(N__59171),
            .I(n27));
    Odrv4 I__11517 (
            .O(N__59166),
            .I(n27));
    LocalMux I__11516 (
            .O(N__59163),
            .I(n27));
    InMux I__11515 (
            .O(N__59146),
            .I(N__59143));
    LocalMux I__11514 (
            .O(N__59143),
            .I(N__59139));
    InMux I__11513 (
            .O(N__59142),
            .I(N__59136));
    Odrv4 I__11512 (
            .O(N__59139),
            .I(REG_mem_38_4));
    LocalMux I__11511 (
            .O(N__59136),
            .I(REG_mem_38_4));
    InMux I__11510 (
            .O(N__59131),
            .I(N__59128));
    LocalMux I__11509 (
            .O(N__59128),
            .I(N__59125));
    Span4Mux_h I__11508 (
            .O(N__59125),
            .I(N__59122));
    Span4Mux_v I__11507 (
            .O(N__59122),
            .I(N__59118));
    InMux I__11506 (
            .O(N__59121),
            .I(N__59115));
    Odrv4 I__11505 (
            .O(N__59118),
            .I(REG_mem_39_5));
    LocalMux I__11504 (
            .O(N__59115),
            .I(REG_mem_39_5));
    CascadeMux I__11503 (
            .O(N__59110),
            .I(N__59107));
    InMux I__11502 (
            .O(N__59107),
            .I(N__59104));
    LocalMux I__11501 (
            .O(N__59104),
            .I(N__59101));
    Span4Mux_v I__11500 (
            .O(N__59101),
            .I(N__59098));
    Span4Mux_h I__11499 (
            .O(N__59098),
            .I(N__59094));
    InMux I__11498 (
            .O(N__59097),
            .I(N__59091));
    Odrv4 I__11497 (
            .O(N__59094),
            .I(REG_mem_55_2));
    LocalMux I__11496 (
            .O(N__59091),
            .I(REG_mem_55_2));
    CascadeMux I__11495 (
            .O(N__59086),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13910_cascade_ ));
    CascadeMux I__11494 (
            .O(N__59083),
            .I(N__59079));
    InMux I__11493 (
            .O(N__59082),
            .I(N__59074));
    InMux I__11492 (
            .O(N__59079),
            .I(N__59074));
    LocalMux I__11491 (
            .O(N__59074),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_2 ));
    CascadeMux I__11490 (
            .O(N__59071),
            .I(N__59067));
    InMux I__11489 (
            .O(N__59070),
            .I(N__59062));
    InMux I__11488 (
            .O(N__59067),
            .I(N__59062));
    LocalMux I__11487 (
            .O(N__59062),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_2 ));
    CascadeMux I__11486 (
            .O(N__59059),
            .I(N__59055));
    InMux I__11485 (
            .O(N__59058),
            .I(N__59052));
    InMux I__11484 (
            .O(N__59055),
            .I(N__59049));
    LocalMux I__11483 (
            .O(N__59052),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_2 ));
    LocalMux I__11482 (
            .O(N__59049),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_2 ));
    InMux I__11481 (
            .O(N__59044),
            .I(N__59041));
    LocalMux I__11480 (
            .O(N__59041),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13283 ));
    InMux I__11479 (
            .O(N__59038),
            .I(N__59035));
    LocalMux I__11478 (
            .O(N__59035),
            .I(N__59032));
    Odrv12 I__11477 (
            .O(N__59032),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13067 ));
    CascadeMux I__11476 (
            .O(N__59029),
            .I(N__59026));
    InMux I__11475 (
            .O(N__59026),
            .I(N__59020));
    InMux I__11474 (
            .O(N__59025),
            .I(N__59020));
    LocalMux I__11473 (
            .O(N__59020),
            .I(REG_mem_26_4));
    InMux I__11472 (
            .O(N__59017),
            .I(N__59013));
    InMux I__11471 (
            .O(N__59016),
            .I(N__59010));
    LocalMux I__11470 (
            .O(N__59013),
            .I(REG_mem_6_1));
    LocalMux I__11469 (
            .O(N__59010),
            .I(REG_mem_6_1));
    InMux I__11468 (
            .O(N__59005),
            .I(N__59002));
    LocalMux I__11467 (
            .O(N__59002),
            .I(N__58999));
    Odrv4 I__11466 (
            .O(N__58999),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11657 ));
    InMux I__11465 (
            .O(N__58996),
            .I(N__58993));
    LocalMux I__11464 (
            .O(N__58993),
            .I(N__58989));
    CascadeMux I__11463 (
            .O(N__58992),
            .I(N__58986));
    Span4Mux_h I__11462 (
            .O(N__58989),
            .I(N__58983));
    InMux I__11461 (
            .O(N__58986),
            .I(N__58980));
    Odrv4 I__11460 (
            .O(N__58983),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_2 ));
    LocalMux I__11459 (
            .O(N__58980),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_2 ));
    CascadeMux I__11458 (
            .O(N__58975),
            .I(N__58971));
    InMux I__11457 (
            .O(N__58974),
            .I(N__58968));
    InMux I__11456 (
            .O(N__58971),
            .I(N__58965));
    LocalMux I__11455 (
            .O(N__58968),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_2 ));
    LocalMux I__11454 (
            .O(N__58965),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_2 ));
    CascadeMux I__11453 (
            .O(N__58960),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13064_cascade_ ));
    CascadeMux I__11452 (
            .O(N__58957),
            .I(N__58954));
    InMux I__11451 (
            .O(N__58954),
            .I(N__58951));
    LocalMux I__11450 (
            .O(N__58951),
            .I(N__58948));
    Odrv4 I__11449 (
            .O(N__58948),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13280 ));
    InMux I__11448 (
            .O(N__58945),
            .I(N__58939));
    InMux I__11447 (
            .O(N__58944),
            .I(N__58939));
    LocalMux I__11446 (
            .O(N__58939),
            .I(REG_mem_23_2));
    InMux I__11445 (
            .O(N__58936),
            .I(N__58933));
    LocalMux I__11444 (
            .O(N__58933),
            .I(N__58929));
    InMux I__11443 (
            .O(N__58932),
            .I(N__58926));
    Odrv4 I__11442 (
            .O(N__58929),
            .I(REG_mem_31_1));
    LocalMux I__11441 (
            .O(N__58926),
            .I(REG_mem_31_1));
    InMux I__11440 (
            .O(N__58921),
            .I(N__58918));
    LocalMux I__11439 (
            .O(N__58918),
            .I(N__58915));
    Span4Mux_h I__11438 (
            .O(N__58915),
            .I(N__58911));
    InMux I__11437 (
            .O(N__58914),
            .I(N__58908));
    Odrv4 I__11436 (
            .O(N__58911),
            .I(REG_mem_26_1));
    LocalMux I__11435 (
            .O(N__58908),
            .I(REG_mem_26_1));
    CascadeMux I__11434 (
            .O(N__58903),
            .I(N__58899));
    InMux I__11433 (
            .O(N__58902),
            .I(N__58896));
    InMux I__11432 (
            .O(N__58899),
            .I(N__58893));
    LocalMux I__11431 (
            .O(N__58896),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_1 ));
    LocalMux I__11430 (
            .O(N__58893),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_1 ));
    InMux I__11429 (
            .O(N__58888),
            .I(N__58885));
    LocalMux I__11428 (
            .O(N__58885),
            .I(N__58882));
    Odrv4 I__11427 (
            .O(N__58882),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11684 ));
    InMux I__11426 (
            .O(N__58879),
            .I(N__58876));
    LocalMux I__11425 (
            .O(N__58876),
            .I(N__58873));
    Span4Mux_v I__11424 (
            .O(N__58873),
            .I(N__58869));
    InMux I__11423 (
            .O(N__58872),
            .I(N__58866));
    Odrv4 I__11422 (
            .O(N__58869),
            .I(REG_mem_19_5));
    LocalMux I__11421 (
            .O(N__58866),
            .I(REG_mem_19_5));
    CascadeMux I__11420 (
            .O(N__58861),
            .I(N__58857));
    InMux I__11419 (
            .O(N__58860),
            .I(N__58852));
    InMux I__11418 (
            .O(N__58857),
            .I(N__58852));
    LocalMux I__11417 (
            .O(N__58852),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_1 ));
    CascadeMux I__11416 (
            .O(N__58849),
            .I(N__58846));
    InMux I__11415 (
            .O(N__58846),
            .I(N__58843));
    LocalMux I__11414 (
            .O(N__58843),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11740 ));
    InMux I__11413 (
            .O(N__58840),
            .I(N__58837));
    LocalMux I__11412 (
            .O(N__58837),
            .I(N__58834));
    Odrv4 I__11411 (
            .O(N__58834),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11741 ));
    InMux I__11410 (
            .O(N__58831),
            .I(N__58828));
    LocalMux I__11409 (
            .O(N__58828),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11726 ));
    CascadeMux I__11408 (
            .O(N__58825),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13892_cascade_ ));
    CascadeMux I__11407 (
            .O(N__58822),
            .I(N__58819));
    InMux I__11406 (
            .O(N__58819),
            .I(N__58816));
    LocalMux I__11405 (
            .O(N__58816),
            .I(N__58813));
    Span4Mux_v I__11404 (
            .O(N__58813),
            .I(N__58810));
    Odrv4 I__11403 (
            .O(N__58810),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11765 ));
    InMux I__11402 (
            .O(N__58807),
            .I(N__58801));
    InMux I__11401 (
            .O(N__58806),
            .I(N__58801));
    LocalMux I__11400 (
            .O(N__58801),
            .I(REG_mem_58_1));
    CascadeMux I__11399 (
            .O(N__58798),
            .I(N__58794));
    InMux I__11398 (
            .O(N__58797),
            .I(N__58789));
    InMux I__11397 (
            .O(N__58794),
            .I(N__58789));
    LocalMux I__11396 (
            .O(N__58789),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_1 ));
    InMux I__11395 (
            .O(N__58786),
            .I(N__58783));
    LocalMux I__11394 (
            .O(N__58783),
            .I(N__58780));
    Span12Mux_s10_v I__11393 (
            .O(N__58780),
            .I(N__58776));
    InMux I__11392 (
            .O(N__58779),
            .I(N__58773));
    Odrv12 I__11391 (
            .O(N__58776),
            .I(REG_mem_15_5));
    LocalMux I__11390 (
            .O(N__58773),
            .I(REG_mem_15_5));
    CascadeMux I__11389 (
            .O(N__58768),
            .I(N__58765));
    InMux I__11388 (
            .O(N__58765),
            .I(N__58762));
    LocalMux I__11387 (
            .O(N__58762),
            .I(N__58759));
    Span4Mux_v I__11386 (
            .O(N__58759),
            .I(N__58756));
    Span4Mux_h I__11385 (
            .O(N__58756),
            .I(N__58753));
    Span4Mux_h I__11384 (
            .O(N__58753),
            .I(N__58749));
    InMux I__11383 (
            .O(N__58752),
            .I(N__58746));
    Odrv4 I__11382 (
            .O(N__58749),
            .I(REG_mem_14_5));
    LocalMux I__11381 (
            .O(N__58746),
            .I(REG_mem_14_5));
    CascadeMux I__11380 (
            .O(N__58741),
            .I(N__58738));
    InMux I__11379 (
            .O(N__58738),
            .I(N__58735));
    LocalMux I__11378 (
            .O(N__58735),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14018 ));
    InMux I__11377 (
            .O(N__58732),
            .I(N__58729));
    LocalMux I__11376 (
            .O(N__58729),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13988 ));
    InMux I__11375 (
            .O(N__58726),
            .I(N__58723));
    LocalMux I__11374 (
            .O(N__58723),
            .I(N__58720));
    Span4Mux_v I__11373 (
            .O(N__58720),
            .I(N__58717));
    Odrv4 I__11372 (
            .O(N__58717),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11747 ));
    SRMux I__11371 (
            .O(N__58714),
            .I(N__58710));
    SRMux I__11370 (
            .O(N__58713),
            .I(N__58707));
    LocalMux I__11369 (
            .O(N__58710),
            .I(N__58704));
    LocalMux I__11368 (
            .O(N__58707),
            .I(N__58701));
    Odrv12 I__11367 (
            .O(N__58704),
            .I(\pc_rx.n6481 ));
    Odrv4 I__11366 (
            .O(N__58701),
            .I(\pc_rx.n6481 ));
    InMux I__11365 (
            .O(N__58696),
            .I(N__58693));
    LocalMux I__11364 (
            .O(N__58693),
            .I(N__58690));
    Span12Mux_h I__11363 (
            .O(N__58690),
            .I(N__58687));
    Odrv12 I__11362 (
            .O(N__58687),
            .I(FIFO_D7_c_7));
    InMux I__11361 (
            .O(N__58684),
            .I(N__58681));
    LocalMux I__11360 (
            .O(N__58681),
            .I(N__58678));
    Span4Mux_v I__11359 (
            .O(N__58678),
            .I(N__58675));
    Sp12to4 I__11358 (
            .O(N__58675),
            .I(N__58672));
    Span12Mux_h I__11357 (
            .O(N__58672),
            .I(N__58668));
    InMux I__11356 (
            .O(N__58671),
            .I(N__58665));
    Odrv12 I__11355 (
            .O(N__58668),
            .I(REG_mem_12_5));
    LocalMux I__11354 (
            .O(N__58665),
            .I(REG_mem_12_5));
    InMux I__11353 (
            .O(N__58660),
            .I(N__58657));
    LocalMux I__11352 (
            .O(N__58657),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14021 ));
    CascadeMux I__11351 (
            .O(N__58654),
            .I(N__58650));
    InMux I__11350 (
            .O(N__58653),
            .I(N__58647));
    InMux I__11349 (
            .O(N__58650),
            .I(N__58644));
    LocalMux I__11348 (
            .O(N__58647),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_1 ));
    LocalMux I__11347 (
            .O(N__58644),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_1 ));
    InMux I__11346 (
            .O(N__58639),
            .I(N__58636));
    LocalMux I__11345 (
            .O(N__58636),
            .I(N__58632));
    CascadeMux I__11344 (
            .O(N__58635),
            .I(N__58629));
    Span4Mux_h I__11343 (
            .O(N__58632),
            .I(N__58626));
    InMux I__11342 (
            .O(N__58629),
            .I(N__58623));
    Odrv4 I__11341 (
            .O(N__58626),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_1 ));
    LocalMux I__11340 (
            .O(N__58623),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_1 ));
    InMux I__11339 (
            .O(N__58618),
            .I(N__58615));
    LocalMux I__11338 (
            .O(N__58615),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11695 ));
    CascadeMux I__11337 (
            .O(N__58612),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11696_cascade_ ));
    CascadeMux I__11336 (
            .O(N__58609),
            .I(N__58605));
    InMux I__11335 (
            .O(N__58608),
            .I(N__58602));
    InMux I__11334 (
            .O(N__58605),
            .I(N__58599));
    LocalMux I__11333 (
            .O(N__58602),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_1 ));
    LocalMux I__11332 (
            .O(N__58599),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_1 ));
    InMux I__11331 (
            .O(N__58594),
            .I(N__58590));
    InMux I__11330 (
            .O(N__58593),
            .I(N__58587));
    LocalMux I__11329 (
            .O(N__58590),
            .I(REG_mem_63_1));
    LocalMux I__11328 (
            .O(N__58587),
            .I(REG_mem_63_1));
    CascadeMux I__11327 (
            .O(N__58582),
            .I(N__58578));
    InMux I__11326 (
            .O(N__58581),
            .I(N__58575));
    InMux I__11325 (
            .O(N__58578),
            .I(N__58572));
    LocalMux I__11324 (
            .O(N__58575),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_1 ));
    LocalMux I__11323 (
            .O(N__58572),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_1 ));
    CascadeMux I__11322 (
            .O(N__58567),
            .I(N__58563));
    CascadeMux I__11321 (
            .O(N__58566),
            .I(N__58560));
    InMux I__11320 (
            .O(N__58563),
            .I(N__58555));
    InMux I__11319 (
            .O(N__58560),
            .I(N__58555));
    LocalMux I__11318 (
            .O(N__58555),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_1 ));
    InMux I__11317 (
            .O(N__58552),
            .I(bfn_15_19_0_));
    InMux I__11316 (
            .O(N__58549),
            .I(\pc_rx.n10703 ));
    InMux I__11315 (
            .O(N__58546),
            .I(\pc_rx.n10704 ));
    InMux I__11314 (
            .O(N__58543),
            .I(\pc_rx.n10705 ));
    InMux I__11313 (
            .O(N__58540),
            .I(\pc_rx.n10706 ));
    InMux I__11312 (
            .O(N__58537),
            .I(\pc_rx.n10707 ));
    InMux I__11311 (
            .O(N__58534),
            .I(\pc_rx.n10708 ));
    InMux I__11310 (
            .O(N__58531),
            .I(\pc_rx.n10709 ));
    InMux I__11309 (
            .O(N__58528),
            .I(bfn_15_20_0_));
    InMux I__11308 (
            .O(N__58525),
            .I(\pc_rx.n10711 ));
    CascadeMux I__11307 (
            .O(N__58522),
            .I(\pc_rx.n149_cascade_ ));
    InMux I__11306 (
            .O(N__58519),
            .I(N__58510));
    InMux I__11305 (
            .O(N__58518),
            .I(N__58510));
    InMux I__11304 (
            .O(N__58517),
            .I(N__58510));
    LocalMux I__11303 (
            .O(N__58510),
            .I(debug_led3));
    InMux I__11302 (
            .O(N__58507),
            .I(N__58504));
    LocalMux I__11301 (
            .O(N__58504),
            .I(uart_rx_complete_prev));
    SRMux I__11300 (
            .O(N__58501),
            .I(N__58498));
    LocalMux I__11299 (
            .O(N__58498),
            .I(n4443));
    CascadeMux I__11298 (
            .O(N__58495),
            .I(N__58491));
    InMux I__11297 (
            .O(N__58494),
            .I(N__58483));
    InMux I__11296 (
            .O(N__58491),
            .I(N__58483));
    InMux I__11295 (
            .O(N__58490),
            .I(N__58483));
    LocalMux I__11294 (
            .O(N__58483),
            .I(even_byte_flag));
    InMux I__11293 (
            .O(N__58480),
            .I(N__58474));
    InMux I__11292 (
            .O(N__58479),
            .I(N__58474));
    LocalMux I__11291 (
            .O(N__58474),
            .I(N__58471));
    Span4Mux_v I__11290 (
            .O(N__58471),
            .I(N__58467));
    InMux I__11289 (
            .O(N__58470),
            .I(N__58464));
    Odrv4 I__11288 (
            .O(N__58467),
            .I(spi_start_transfer_r));
    LocalMux I__11287 (
            .O(N__58464),
            .I(spi_start_transfer_r));
    InMux I__11286 (
            .O(N__58459),
            .I(N__58455));
    InMux I__11285 (
            .O(N__58458),
            .I(N__58452));
    LocalMux I__11284 (
            .O(N__58455),
            .I(N__58445));
    LocalMux I__11283 (
            .O(N__58452),
            .I(N__58445));
    InMux I__11282 (
            .O(N__58451),
            .I(N__58442));
    InMux I__11281 (
            .O(N__58450),
            .I(N__58439));
    Odrv4 I__11280 (
            .O(N__58445),
            .I(tx_data_byte_7));
    LocalMux I__11279 (
            .O(N__58442),
            .I(tx_data_byte_7));
    LocalMux I__11278 (
            .O(N__58439),
            .I(tx_data_byte_7));
    InMux I__11277 (
            .O(N__58432),
            .I(N__58429));
    LocalMux I__11276 (
            .O(N__58429),
            .I(N__58426));
    Span4Mux_v I__11275 (
            .O(N__58426),
            .I(N__58422));
    InMux I__11274 (
            .O(N__58425),
            .I(N__58419));
    Odrv4 I__11273 (
            .O(N__58422),
            .I(tx_addr_byte_7));
    LocalMux I__11272 (
            .O(N__58419),
            .I(tx_addr_byte_7));
    InMux I__11271 (
            .O(N__58414),
            .I(N__58410));
    InMux I__11270 (
            .O(N__58413),
            .I(N__58407));
    LocalMux I__11269 (
            .O(N__58410),
            .I(pc_data_rx_1));
    LocalMux I__11268 (
            .O(N__58407),
            .I(pc_data_rx_1));
    CascadeMux I__11267 (
            .O(N__58402),
            .I(N__58398));
    CascadeMux I__11266 (
            .O(N__58401),
            .I(N__58395));
    InMux I__11265 (
            .O(N__58398),
            .I(N__58390));
    InMux I__11264 (
            .O(N__58395),
            .I(N__58390));
    LocalMux I__11263 (
            .O(N__58390),
            .I(pc_data_rx_4));
    InMux I__11262 (
            .O(N__58387),
            .I(N__58384));
    LocalMux I__11261 (
            .O(N__58384),
            .I(N__58381));
    Span4Mux_v I__11260 (
            .O(N__58381),
            .I(N__58378));
    Sp12to4 I__11259 (
            .O(N__58378),
            .I(N__58375));
    Span12Mux_h I__11258 (
            .O(N__58375),
            .I(N__58372));
    Span12Mux_v I__11257 (
            .O(N__58372),
            .I(N__58369));
    Odrv12 I__11256 (
            .O(N__58369),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14261 ));
    InMux I__11255 (
            .O(N__58366),
            .I(N__58363));
    LocalMux I__11254 (
            .O(N__58363),
            .I(N__58360));
    Span12Mux_v I__11253 (
            .O(N__58360),
            .I(N__58357));
    Odrv12 I__11252 (
            .O(N__58357),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13253 ));
    CascadeMux I__11251 (
            .O(N__58354),
            .I(N__58351));
    InMux I__11250 (
            .O(N__58351),
            .I(N__58348));
    LocalMux I__11249 (
            .O(N__58348),
            .I(N__58345));
    Span4Mux_v I__11248 (
            .O(N__58345),
            .I(N__58342));
    Span4Mux_h I__11247 (
            .O(N__58342),
            .I(N__58339));
    Odrv4 I__11246 (
            .O(N__58339),
            .I(REG_out_raw_5));
    InMux I__11245 (
            .O(N__58336),
            .I(N__58332));
    InMux I__11244 (
            .O(N__58335),
            .I(N__58329));
    LocalMux I__11243 (
            .O(N__58332),
            .I(n4_adj_1205));
    LocalMux I__11242 (
            .O(N__58329),
            .I(n4_adj_1205));
    CascadeMux I__11241 (
            .O(N__58324),
            .I(N__58321));
    InMux I__11240 (
            .O(N__58321),
            .I(N__58317));
    InMux I__11239 (
            .O(N__58320),
            .I(N__58314));
    LocalMux I__11238 (
            .O(N__58317),
            .I(N__58311));
    LocalMux I__11237 (
            .O(N__58314),
            .I(n4_adj_1206));
    Odrv4 I__11236 (
            .O(N__58311),
            .I(n4_adj_1206));
    CascadeMux I__11235 (
            .O(N__58306),
            .I(N__58302));
    InMux I__11234 (
            .O(N__58305),
            .I(N__58299));
    InMux I__11233 (
            .O(N__58302),
            .I(N__58296));
    LocalMux I__11232 (
            .O(N__58299),
            .I(n7455));
    LocalMux I__11231 (
            .O(N__58296),
            .I(n7455));
    InMux I__11230 (
            .O(N__58291),
            .I(N__58288));
    LocalMux I__11229 (
            .O(N__58288),
            .I(\pc_rx.n149 ));
    CascadeMux I__11228 (
            .O(N__58285),
            .I(N__58282));
    InMux I__11227 (
            .O(N__58282),
            .I(N__58279));
    LocalMux I__11226 (
            .O(N__58279),
            .I(N__58276));
    Span12Mux_v I__11225 (
            .O(N__58276),
            .I(N__58273));
    Span12Mux_h I__11224 (
            .O(N__58273),
            .I(N__58270));
    Odrv12 I__11223 (
            .O(N__58270),
            .I(REG_out_raw_3));
    CascadeMux I__11222 (
            .O(N__58267),
            .I(N__58264));
    InMux I__11221 (
            .O(N__58264),
            .I(N__58261));
    LocalMux I__11220 (
            .O(N__58261),
            .I(N__58258));
    Span4Mux_v I__11219 (
            .O(N__58258),
            .I(N__58255));
    Odrv4 I__11218 (
            .O(N__58255),
            .I(REG_out_raw_15));
    InMux I__11217 (
            .O(N__58252),
            .I(N__58248));
    InMux I__11216 (
            .O(N__58251),
            .I(N__58245));
    LocalMux I__11215 (
            .O(N__58248),
            .I(fifo_data_out_15));
    LocalMux I__11214 (
            .O(N__58245),
            .I(fifo_data_out_15));
    InMux I__11213 (
            .O(N__58240),
            .I(N__58236));
    InMux I__11212 (
            .O(N__58239),
            .I(N__58233));
    LocalMux I__11211 (
            .O(N__58236),
            .I(pc_data_rx_6));
    LocalMux I__11210 (
            .O(N__58233),
            .I(pc_data_rx_6));
    InMux I__11209 (
            .O(N__58228),
            .I(N__58223));
    InMux I__11208 (
            .O(N__58227),
            .I(N__58220));
    InMux I__11207 (
            .O(N__58226),
            .I(N__58216));
    LocalMux I__11206 (
            .O(N__58223),
            .I(N__58213));
    LocalMux I__11205 (
            .O(N__58220),
            .I(N__58210));
    InMux I__11204 (
            .O(N__58219),
            .I(N__58207));
    LocalMux I__11203 (
            .O(N__58216),
            .I(tx_data_byte_2));
    Odrv4 I__11202 (
            .O(N__58213),
            .I(tx_data_byte_2));
    Odrv4 I__11201 (
            .O(N__58210),
            .I(tx_data_byte_2));
    LocalMux I__11200 (
            .O(N__58207),
            .I(tx_data_byte_2));
    InMux I__11199 (
            .O(N__58198),
            .I(N__58194));
    InMux I__11198 (
            .O(N__58197),
            .I(N__58191));
    LocalMux I__11197 (
            .O(N__58194),
            .I(tx_addr_byte_2));
    LocalMux I__11196 (
            .O(N__58191),
            .I(tx_addr_byte_2));
    InMux I__11195 (
            .O(N__58186),
            .I(N__58177));
    InMux I__11194 (
            .O(N__58185),
            .I(N__58177));
    InMux I__11193 (
            .O(N__58184),
            .I(N__58177));
    LocalMux I__11192 (
            .O(N__58177),
            .I(n3997));
    CascadeMux I__11191 (
            .O(N__58174),
            .I(N__58170));
    InMux I__11190 (
            .O(N__58173),
            .I(N__58167));
    InMux I__11189 (
            .O(N__58170),
            .I(N__58164));
    LocalMux I__11188 (
            .O(N__58167),
            .I(pc_data_rx_2));
    LocalMux I__11187 (
            .O(N__58164),
            .I(pc_data_rx_2));
    SRMux I__11186 (
            .O(N__58159),
            .I(N__58156));
    LocalMux I__11185 (
            .O(N__58156),
            .I(\bluejay_data_inst.n4522 ));
    InMux I__11184 (
            .O(N__58153),
            .I(N__58150));
    LocalMux I__11183 (
            .O(N__58150),
            .I(N__58147));
    Span4Mux_v I__11182 (
            .O(N__58147),
            .I(N__58143));
    InMux I__11181 (
            .O(N__58146),
            .I(N__58140));
    Odrv4 I__11180 (
            .O(N__58143),
            .I(fifo_data_out_11));
    LocalMux I__11179 (
            .O(N__58140),
            .I(fifo_data_out_11));
    IoInMux I__11178 (
            .O(N__58135),
            .I(N__58131));
    IoInMux I__11177 (
            .O(N__58134),
            .I(N__58128));
    LocalMux I__11176 (
            .O(N__58131),
            .I(N__58125));
    LocalMux I__11175 (
            .O(N__58128),
            .I(N__58122));
    IoSpan4Mux I__11174 (
            .O(N__58125),
            .I(N__58119));
    IoSpan4Mux I__11173 (
            .O(N__58122),
            .I(N__58116));
    Sp12to4 I__11172 (
            .O(N__58119),
            .I(N__58113));
    Span4Mux_s0_h I__11171 (
            .O(N__58116),
            .I(N__58110));
    Span12Mux_v I__11170 (
            .O(N__58113),
            .I(N__58105));
    Sp12to4 I__11169 (
            .O(N__58110),
            .I(N__58105));
    Odrv12 I__11168 (
            .O(N__58105),
            .I(DATA11_c));
    InMux I__11167 (
            .O(N__58102),
            .I(N__58098));
    CascadeMux I__11166 (
            .O(N__58101),
            .I(N__58095));
    LocalMux I__11165 (
            .O(N__58098),
            .I(N__58092));
    InMux I__11164 (
            .O(N__58095),
            .I(N__58089));
    Odrv4 I__11163 (
            .O(N__58092),
            .I(fifo_data_out_10));
    LocalMux I__11162 (
            .O(N__58089),
            .I(fifo_data_out_10));
    IoInMux I__11161 (
            .O(N__58084),
            .I(N__58080));
    IoInMux I__11160 (
            .O(N__58083),
            .I(N__58077));
    LocalMux I__11159 (
            .O(N__58080),
            .I(N__58074));
    LocalMux I__11158 (
            .O(N__58077),
            .I(N__58071));
    Span12Mux_s3_h I__11157 (
            .O(N__58074),
            .I(N__58068));
    Span12Mux_s6_v I__11156 (
            .O(N__58071),
            .I(N__58065));
    Odrv12 I__11155 (
            .O(N__58068),
            .I(DATA10_c));
    Odrv12 I__11154 (
            .O(N__58065),
            .I(DATA10_c));
    IoInMux I__11153 (
            .O(N__58060),
            .I(N__58057));
    LocalMux I__11152 (
            .O(N__58057),
            .I(N__58053));
    IoInMux I__11151 (
            .O(N__58056),
            .I(N__58050));
    Span4Mux_s0_h I__11150 (
            .O(N__58053),
            .I(N__58047));
    LocalMux I__11149 (
            .O(N__58050),
            .I(N__58044));
    Span4Mux_h I__11148 (
            .O(N__58047),
            .I(N__58041));
    Span4Mux_s1_v I__11147 (
            .O(N__58044),
            .I(N__58038));
    Span4Mux_h I__11146 (
            .O(N__58041),
            .I(N__58035));
    Span4Mux_v I__11145 (
            .O(N__58038),
            .I(N__58032));
    Span4Mux_h I__11144 (
            .O(N__58035),
            .I(N__58027));
    Span4Mux_v I__11143 (
            .O(N__58032),
            .I(N__58027));
    Odrv4 I__11142 (
            .O(N__58027),
            .I(DATA9_c));
    InMux I__11141 (
            .O(N__58024),
            .I(N__58021));
    LocalMux I__11140 (
            .O(N__58021),
            .I(N__58015));
    InMux I__11139 (
            .O(N__58020),
            .I(N__58012));
    InMux I__11138 (
            .O(N__58019),
            .I(N__58007));
    InMux I__11137 (
            .O(N__58018),
            .I(N__58007));
    Odrv4 I__11136 (
            .O(N__58015),
            .I(tx_data_byte_0));
    LocalMux I__11135 (
            .O(N__58012),
            .I(tx_data_byte_0));
    LocalMux I__11134 (
            .O(N__58007),
            .I(tx_data_byte_0));
    CEMux I__11133 (
            .O(N__58000),
            .I(N__57997));
    LocalMux I__11132 (
            .O(N__57997),
            .I(N__57994));
    IoSpan4Mux I__11131 (
            .O(N__57994),
            .I(N__57991));
    IoSpan4Mux I__11130 (
            .O(N__57991),
            .I(N__57988));
    IoSpan4Mux I__11129 (
            .O(N__57988),
            .I(N__57984));
    CascadeMux I__11128 (
            .O(N__57987),
            .I(N__57981));
    IoSpan4Mux I__11127 (
            .O(N__57984),
            .I(N__57977));
    InMux I__11126 (
            .O(N__57981),
            .I(N__57974));
    CEMux I__11125 (
            .O(N__57980),
            .I(N__57971));
    Span4Mux_s3_v I__11124 (
            .O(N__57977),
            .I(N__57968));
    LocalMux I__11123 (
            .O(N__57974),
            .I(N__57963));
    LocalMux I__11122 (
            .O(N__57971),
            .I(N__57963));
    Sp12to4 I__11121 (
            .O(N__57968),
            .I(N__57957));
    Span12Mux_h I__11120 (
            .O(N__57963),
            .I(N__57957));
    CEMux I__11119 (
            .O(N__57962),
            .I(N__57954));
    Odrv12 I__11118 (
            .O(N__57957),
            .I(n4070));
    LocalMux I__11117 (
            .O(N__57954),
            .I(n4070));
    InMux I__11116 (
            .O(N__57949),
            .I(N__57946));
    LocalMux I__11115 (
            .O(N__57946),
            .I(N__57943));
    Span4Mux_h I__11114 (
            .O(N__57943),
            .I(N__57939));
    InMux I__11113 (
            .O(N__57942),
            .I(N__57936));
    Odrv4 I__11112 (
            .O(N__57939),
            .I(tx_shift_reg_0));
    LocalMux I__11111 (
            .O(N__57936),
            .I(tx_shift_reg_0));
    InMux I__11110 (
            .O(N__57931),
            .I(N__57925));
    InMux I__11109 (
            .O(N__57930),
            .I(N__57925));
    LocalMux I__11108 (
            .O(N__57925),
            .I(N__57914));
    InMux I__11107 (
            .O(N__57924),
            .I(N__57897));
    InMux I__11106 (
            .O(N__57923),
            .I(N__57897));
    InMux I__11105 (
            .O(N__57922),
            .I(N__57897));
    InMux I__11104 (
            .O(N__57921),
            .I(N__57897));
    InMux I__11103 (
            .O(N__57920),
            .I(N__57897));
    InMux I__11102 (
            .O(N__57919),
            .I(N__57897));
    InMux I__11101 (
            .O(N__57918),
            .I(N__57897));
    InMux I__11100 (
            .O(N__57917),
            .I(N__57897));
    Span4Mux_h I__11099 (
            .O(N__57914),
            .I(N__57886));
    LocalMux I__11098 (
            .O(N__57897),
            .I(N__57886));
    InMux I__11097 (
            .O(N__57896),
            .I(N__57873));
    InMux I__11096 (
            .O(N__57895),
            .I(N__57873));
    InMux I__11095 (
            .O(N__57894),
            .I(N__57873));
    InMux I__11094 (
            .O(N__57893),
            .I(N__57873));
    InMux I__11093 (
            .O(N__57892),
            .I(N__57873));
    InMux I__11092 (
            .O(N__57891),
            .I(N__57873));
    Span4Mux_v I__11091 (
            .O(N__57886),
            .I(N__57868));
    LocalMux I__11090 (
            .O(N__57873),
            .I(N__57868));
    Span4Mux_v I__11089 (
            .O(N__57868),
            .I(N__57865));
    Odrv4 I__11088 (
            .O(N__57865),
            .I(n1928));
    InMux I__11087 (
            .O(N__57862),
            .I(N__57859));
    LocalMux I__11086 (
            .O(N__57859),
            .I(\spi0.tx_shift_reg_14 ));
    IoInMux I__11085 (
            .O(N__57856),
            .I(N__57853));
    LocalMux I__11084 (
            .O(N__57853),
            .I(N__57850));
    IoSpan4Mux I__11083 (
            .O(N__57850),
            .I(N__57847));
    Span4Mux_s2_v I__11082 (
            .O(N__57847),
            .I(N__57844));
    Sp12to4 I__11081 (
            .O(N__57844),
            .I(N__57841));
    Span12Mux_h I__11080 (
            .O(N__57841),
            .I(N__57838));
    Odrv12 I__11079 (
            .O(N__57838),
            .I(\spi0.n1930 ));
    CascadeMux I__11078 (
            .O(N__57835),
            .I(N__57832));
    InMux I__11077 (
            .O(N__57832),
            .I(N__57829));
    LocalMux I__11076 (
            .O(N__57829),
            .I(N__57826));
    Span12Mux_v I__11075 (
            .O(N__57826),
            .I(N__57823));
    Odrv12 I__11074 (
            .O(N__57823),
            .I(REG_out_raw_12));
    CascadeMux I__11073 (
            .O(N__57820),
            .I(N__57816));
    InMux I__11072 (
            .O(N__57819),
            .I(N__57813));
    InMux I__11071 (
            .O(N__57816),
            .I(N__57810));
    LocalMux I__11070 (
            .O(N__57813),
            .I(pc_data_rx_7));
    LocalMux I__11069 (
            .O(N__57810),
            .I(pc_data_rx_7));
    InMux I__11068 (
            .O(N__57805),
            .I(N__57802));
    LocalMux I__11067 (
            .O(N__57802),
            .I(N__57799));
    Span4Mux_h I__11066 (
            .O(N__57799),
            .I(N__57796));
    Odrv4 I__11065 (
            .O(N__57796),
            .I(REG_out_raw_9));
    CascadeMux I__11064 (
            .O(N__57793),
            .I(N__57790));
    InMux I__11063 (
            .O(N__57790),
            .I(N__57786));
    InMux I__11062 (
            .O(N__57789),
            .I(N__57783));
    LocalMux I__11061 (
            .O(N__57786),
            .I(N__57780));
    LocalMux I__11060 (
            .O(N__57783),
            .I(fifo_data_out_9));
    Odrv4 I__11059 (
            .O(N__57780),
            .I(fifo_data_out_9));
    InMux I__11058 (
            .O(N__57775),
            .I(N__57772));
    LocalMux I__11057 (
            .O(N__57772),
            .I(N__57769));
    Odrv12 I__11056 (
            .O(N__57769),
            .I(\usb3_if_inst.n10869 ));
    IoInMux I__11055 (
            .O(N__57766),
            .I(N__57763));
    LocalMux I__11054 (
            .O(N__57763),
            .I(N__57760));
    IoSpan4Mux I__11053 (
            .O(N__57760),
            .I(N__57757));
    Span4Mux_s2_h I__11052 (
            .O(N__57757),
            .I(N__57754));
    Sp12to4 I__11051 (
            .O(N__57754),
            .I(N__57745));
    InMux I__11050 (
            .O(N__57753),
            .I(N__57740));
    InMux I__11049 (
            .O(N__57752),
            .I(N__57740));
    InMux I__11048 (
            .O(N__57751),
            .I(N__57737));
    InMux I__11047 (
            .O(N__57750),
            .I(N__57732));
    InMux I__11046 (
            .O(N__57749),
            .I(N__57732));
    CascadeMux I__11045 (
            .O(N__57748),
            .I(N__57728));
    Span12Mux_h I__11044 (
            .O(N__57745),
            .I(N__57725));
    LocalMux I__11043 (
            .O(N__57740),
            .I(N__57722));
    LocalMux I__11042 (
            .O(N__57737),
            .I(N__57717));
    LocalMux I__11041 (
            .O(N__57732),
            .I(N__57717));
    InMux I__11040 (
            .O(N__57731),
            .I(N__57712));
    InMux I__11039 (
            .O(N__57728),
            .I(N__57712));
    Span12Mux_v I__11038 (
            .O(N__57725),
            .I(N__57703));
    Span4Mux_v I__11037 (
            .O(N__57722),
            .I(N__57700));
    Span4Mux_v I__11036 (
            .O(N__57717),
            .I(N__57697));
    LocalMux I__11035 (
            .O(N__57712),
            .I(N__57694));
    InMux I__11034 (
            .O(N__57711),
            .I(N__57691));
    InMux I__11033 (
            .O(N__57710),
            .I(N__57680));
    InMux I__11032 (
            .O(N__57709),
            .I(N__57680));
    InMux I__11031 (
            .O(N__57708),
            .I(N__57680));
    InMux I__11030 (
            .O(N__57707),
            .I(N__57680));
    InMux I__11029 (
            .O(N__57706),
            .I(N__57680));
    Odrv12 I__11028 (
            .O(N__57703),
            .I(DEBUG_5_c));
    Odrv4 I__11027 (
            .O(N__57700),
            .I(DEBUG_5_c));
    Odrv4 I__11026 (
            .O(N__57697),
            .I(DEBUG_5_c));
    Odrv4 I__11025 (
            .O(N__57694),
            .I(DEBUG_5_c));
    LocalMux I__11024 (
            .O(N__57691),
            .I(DEBUG_5_c));
    LocalMux I__11023 (
            .O(N__57680),
            .I(DEBUG_5_c));
    InMux I__11022 (
            .O(N__57667),
            .I(N__57663));
    InMux I__11021 (
            .O(N__57666),
            .I(N__57660));
    LocalMux I__11020 (
            .O(N__57663),
            .I(\usb3_if_inst.n555 ));
    LocalMux I__11019 (
            .O(N__57660),
            .I(\usb3_if_inst.n555 ));
    InMux I__11018 (
            .O(N__57655),
            .I(N__57652));
    LocalMux I__11017 (
            .O(N__57652),
            .I(\usb3_if_inst.n10746 ));
    IoInMux I__11016 (
            .O(N__57649),
            .I(N__57642));
    CascadeMux I__11015 (
            .O(N__57648),
            .I(N__57639));
    CascadeMux I__11014 (
            .O(N__57647),
            .I(N__57634));
    CascadeMux I__11013 (
            .O(N__57646),
            .I(N__57631));
    CascadeMux I__11012 (
            .O(N__57645),
            .I(N__57626));
    LocalMux I__11011 (
            .O(N__57642),
            .I(N__57622));
    InMux I__11010 (
            .O(N__57639),
            .I(N__57619));
    InMux I__11009 (
            .O(N__57638),
            .I(N__57610));
    InMux I__11008 (
            .O(N__57637),
            .I(N__57610));
    InMux I__11007 (
            .O(N__57634),
            .I(N__57610));
    InMux I__11006 (
            .O(N__57631),
            .I(N__57610));
    CascadeMux I__11005 (
            .O(N__57630),
            .I(N__57607));
    InMux I__11004 (
            .O(N__57629),
            .I(N__57600));
    InMux I__11003 (
            .O(N__57626),
            .I(N__57600));
    InMux I__11002 (
            .O(N__57625),
            .I(N__57600));
    IoSpan4Mux I__11001 (
            .O(N__57622),
            .I(N__57596));
    LocalMux I__11000 (
            .O(N__57619),
            .I(N__57591));
    LocalMux I__10999 (
            .O(N__57610),
            .I(N__57591));
    InMux I__10998 (
            .O(N__57607),
            .I(N__57588));
    LocalMux I__10997 (
            .O(N__57600),
            .I(N__57585));
    CascadeMux I__10996 (
            .O(N__57599),
            .I(N__57580));
    Span4Mux_s0_h I__10995 (
            .O(N__57596),
            .I(N__57577));
    Span4Mux_v I__10994 (
            .O(N__57591),
            .I(N__57574));
    LocalMux I__10993 (
            .O(N__57588),
            .I(N__57571));
    Span4Mux_v I__10992 (
            .O(N__57585),
            .I(N__57568));
    InMux I__10991 (
            .O(N__57584),
            .I(N__57561));
    InMux I__10990 (
            .O(N__57583),
            .I(N__57561));
    InMux I__10989 (
            .O(N__57580),
            .I(N__57561));
    Span4Mux_h I__10988 (
            .O(N__57577),
            .I(N__57558));
    Span4Mux_h I__10987 (
            .O(N__57574),
            .I(N__57553));
    Span4Mux_v I__10986 (
            .O(N__57571),
            .I(N__57553));
    Span4Mux_h I__10985 (
            .O(N__57568),
            .I(N__57548));
    LocalMux I__10984 (
            .O(N__57561),
            .I(N__57548));
    Sp12to4 I__10983 (
            .O(N__57558),
            .I(N__57545));
    Span4Mux_h I__10982 (
            .O(N__57553),
            .I(N__57540));
    Span4Mux_h I__10981 (
            .O(N__57548),
            .I(N__57540));
    Span12Mux_v I__10980 (
            .O(N__57545),
            .I(N__57537));
    Span4Mux_v I__10979 (
            .O(N__57540),
            .I(N__57534));
    Span12Mux_h I__10978 (
            .O(N__57537),
            .I(N__57531));
    Span4Mux_v I__10977 (
            .O(N__57534),
            .I(N__57528));
    Span12Mux_h I__10976 (
            .O(N__57531),
            .I(N__57525));
    Sp12to4 I__10975 (
            .O(N__57528),
            .I(N__57522));
    Odrv12 I__10974 (
            .O(N__57525),
            .I(DEBUG_2_c_c));
    Odrv12 I__10973 (
            .O(N__57522),
            .I(DEBUG_2_c_c));
    InMux I__10972 (
            .O(N__57517),
            .I(N__57514));
    LocalMux I__10971 (
            .O(N__57514),
            .I(N__57510));
    InMux I__10970 (
            .O(N__57513),
            .I(N__57507));
    Odrv12 I__10969 (
            .O(N__57510),
            .I(\usb3_if_inst.n7360 ));
    LocalMux I__10968 (
            .O(N__57507),
            .I(\usb3_if_inst.n7360 ));
    InMux I__10967 (
            .O(N__57502),
            .I(N__57497));
    InMux I__10966 (
            .O(N__57501),
            .I(N__57492));
    InMux I__10965 (
            .O(N__57500),
            .I(N__57492));
    LocalMux I__10964 (
            .O(N__57497),
            .I(N__57488));
    LocalMux I__10963 (
            .O(N__57492),
            .I(N__57485));
    InMux I__10962 (
            .O(N__57491),
            .I(N__57482));
    Span4Mux_v I__10961 (
            .O(N__57488),
            .I(N__57479));
    Span4Mux_h I__10960 (
            .O(N__57485),
            .I(N__57474));
    LocalMux I__10959 (
            .O(N__57482),
            .I(N__57474));
    Span4Mux_h I__10958 (
            .O(N__57479),
            .I(N__57471));
    Span4Mux_h I__10957 (
            .O(N__57474),
            .I(N__57468));
    Odrv4 I__10956 (
            .O(N__57471),
            .I(\usb3_if_inst.state_timeout_counter_2 ));
    Odrv4 I__10955 (
            .O(N__57468),
            .I(\usb3_if_inst.state_timeout_counter_2 ));
    InMux I__10954 (
            .O(N__57463),
            .I(N__57460));
    LocalMux I__10953 (
            .O(N__57460),
            .I(\usb3_if_inst.n4 ));
    CascadeMux I__10952 (
            .O(N__57457),
            .I(\usb3_if_inst.n7360_cascade_ ));
    InMux I__10951 (
            .O(N__57454),
            .I(N__57451));
    LocalMux I__10950 (
            .O(N__57451),
            .I(\usb3_if_inst.n7505 ));
    IoInMux I__10949 (
            .O(N__57448),
            .I(N__57445));
    LocalMux I__10948 (
            .O(N__57445),
            .I(N__57441));
    IoInMux I__10947 (
            .O(N__57444),
            .I(N__57438));
    IoSpan4Mux I__10946 (
            .O(N__57441),
            .I(N__57435));
    LocalMux I__10945 (
            .O(N__57438),
            .I(N__57432));
    Span4Mux_s0_h I__10944 (
            .O(N__57435),
            .I(N__57429));
    Span12Mux_s4_v I__10943 (
            .O(N__57432),
            .I(N__57426));
    Sp12to4 I__10942 (
            .O(N__57429),
            .I(N__57423));
    Span12Mux_h I__10941 (
            .O(N__57426),
            .I(N__57418));
    Span12Mux_h I__10940 (
            .O(N__57423),
            .I(N__57418));
    Odrv12 I__10939 (
            .O(N__57418),
            .I(DATA15_c));
    IoInMux I__10938 (
            .O(N__57415),
            .I(N__57412));
    LocalMux I__10937 (
            .O(N__57412),
            .I(N__57409));
    Sp12to4 I__10936 (
            .O(N__57409),
            .I(N__57406));
    Span12Mux_h I__10935 (
            .O(N__57406),
            .I(N__57403));
    Odrv12 I__10934 (
            .O(N__57403),
            .I(\bluejay_data_inst.valid_N_707 ));
    InMux I__10933 (
            .O(N__57400),
            .I(N__57394));
    CascadeMux I__10932 (
            .O(N__57399),
            .I(N__57389));
    InMux I__10931 (
            .O(N__57398),
            .I(N__57382));
    InMux I__10930 (
            .O(N__57397),
            .I(N__57379));
    LocalMux I__10929 (
            .O(N__57394),
            .I(N__57376));
    InMux I__10928 (
            .O(N__57393),
            .I(N__57371));
    InMux I__10927 (
            .O(N__57392),
            .I(N__57371));
    InMux I__10926 (
            .O(N__57389),
            .I(N__57362));
    InMux I__10925 (
            .O(N__57388),
            .I(N__57362));
    InMux I__10924 (
            .O(N__57387),
            .I(N__57362));
    InMux I__10923 (
            .O(N__57386),
            .I(N__57362));
    InMux I__10922 (
            .O(N__57385),
            .I(N__57359));
    LocalMux I__10921 (
            .O(N__57382),
            .I(N__57356));
    LocalMux I__10920 (
            .O(N__57379),
            .I(N__57347));
    Span4Mux_v I__10919 (
            .O(N__57376),
            .I(N__57347));
    LocalMux I__10918 (
            .O(N__57371),
            .I(N__57347));
    LocalMux I__10917 (
            .O(N__57362),
            .I(N__57347));
    LocalMux I__10916 (
            .O(N__57359),
            .I(N__57344));
    Span4Mux_h I__10915 (
            .O(N__57356),
            .I(N__57341));
    Odrv4 I__10914 (
            .O(N__57347),
            .I(\usb3_if_inst.n7 ));
    Odrv4 I__10913 (
            .O(N__57344),
            .I(\usb3_if_inst.n7 ));
    Odrv4 I__10912 (
            .O(N__57341),
            .I(\usb3_if_inst.n7 ));
    CEMux I__10911 (
            .O(N__57334),
            .I(N__57330));
    CEMux I__10910 (
            .O(N__57333),
            .I(N__57327));
    LocalMux I__10909 (
            .O(N__57330),
            .I(\usb3_if_inst.n4178 ));
    LocalMux I__10908 (
            .O(N__57327),
            .I(\usb3_if_inst.n4178 ));
    InMux I__10907 (
            .O(N__57322),
            .I(N__57319));
    LocalMux I__10906 (
            .O(N__57319),
            .I(N__57316));
    Span4Mux_v I__10905 (
            .O(N__57316),
            .I(N__57312));
    InMux I__10904 (
            .O(N__57315),
            .I(N__57309));
    Odrv4 I__10903 (
            .O(N__57312),
            .I(fifo_data_out_0));
    LocalMux I__10902 (
            .O(N__57309),
            .I(fifo_data_out_0));
    IoInMux I__10901 (
            .O(N__57304),
            .I(N__57300));
    IoInMux I__10900 (
            .O(N__57303),
            .I(N__57297));
    LocalMux I__10899 (
            .O(N__57300),
            .I(N__57294));
    LocalMux I__10898 (
            .O(N__57297),
            .I(N__57291));
    Span4Mux_s0_v I__10897 (
            .O(N__57294),
            .I(N__57288));
    Span4Mux_s1_h I__10896 (
            .O(N__57291),
            .I(N__57285));
    Sp12to4 I__10895 (
            .O(N__57288),
            .I(N__57282));
    Sp12to4 I__10894 (
            .O(N__57285),
            .I(N__57279));
    Span12Mux_s11_h I__10893 (
            .O(N__57282),
            .I(N__57276));
    Span12Mux_s9_v I__10892 (
            .O(N__57279),
            .I(N__57273));
    Span12Mux_v I__10891 (
            .O(N__57276),
            .I(N__57270));
    Span12Mux_h I__10890 (
            .O(N__57273),
            .I(N__57267));
    Odrv12 I__10889 (
            .O(N__57270),
            .I(DATA16_c));
    Odrv12 I__10888 (
            .O(N__57267),
            .I(DATA16_c));
    CascadeMux I__10887 (
            .O(N__57262),
            .I(N__57258));
    InMux I__10886 (
            .O(N__57261),
            .I(N__57255));
    InMux I__10885 (
            .O(N__57258),
            .I(N__57252));
    LocalMux I__10884 (
            .O(N__57255),
            .I(N__57249));
    LocalMux I__10883 (
            .O(N__57252),
            .I(N__57246));
    Span4Mux_v I__10882 (
            .O(N__57249),
            .I(N__57243));
    Span4Mux_h I__10881 (
            .O(N__57246),
            .I(N__57240));
    Sp12to4 I__10880 (
            .O(N__57243),
            .I(N__57237));
    Span4Mux_h I__10879 (
            .O(N__57240),
            .I(N__57234));
    Span12Mux_h I__10878 (
            .O(N__57237),
            .I(N__57231));
    Odrv4 I__10877 (
            .O(N__57234),
            .I(\usb3_if_inst.n552 ));
    Odrv12 I__10876 (
            .O(N__57231),
            .I(\usb3_if_inst.n552 ));
    InMux I__10875 (
            .O(N__57226),
            .I(N__57215));
    InMux I__10874 (
            .O(N__57225),
            .I(N__57215));
    InMux I__10873 (
            .O(N__57224),
            .I(N__57215));
    InMux I__10872 (
            .O(N__57223),
            .I(N__57210));
    InMux I__10871 (
            .O(N__57222),
            .I(N__57210));
    LocalMux I__10870 (
            .O(N__57215),
            .I(\usb3_if_inst.n554 ));
    LocalMux I__10869 (
            .O(N__57210),
            .I(\usb3_if_inst.n554 ));
    InMux I__10868 (
            .O(N__57205),
            .I(N__57198));
    InMux I__10867 (
            .O(N__57204),
            .I(N__57198));
    InMux I__10866 (
            .O(N__57203),
            .I(N__57195));
    LocalMux I__10865 (
            .O(N__57198),
            .I(N__57192));
    LocalMux I__10864 (
            .O(N__57195),
            .I(\usb3_if_inst.n2798 ));
    Odrv4 I__10863 (
            .O(N__57192),
            .I(\usb3_if_inst.n2798 ));
    InMux I__10862 (
            .O(N__57187),
            .I(N__57184));
    LocalMux I__10861 (
            .O(N__57184),
            .I(\usb3_if_inst.n3973 ));
    CascadeMux I__10860 (
            .O(N__57181),
            .I(\usb3_if_inst.n3973_cascade_ ));
    SRMux I__10859 (
            .O(N__57178),
            .I(N__57175));
    LocalMux I__10858 (
            .O(N__57175),
            .I(N__57172));
    Odrv12 I__10857 (
            .O(N__57172),
            .I(\usb3_if_inst.n10751 ));
    CascadeMux I__10856 (
            .O(N__57169),
            .I(\bluejay_data_inst.n6_cascade_ ));
    CascadeMux I__10855 (
            .O(N__57166),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13934_cascade_ ));
    InMux I__10854 (
            .O(N__57163),
            .I(N__57160));
    LocalMux I__10853 (
            .O(N__57160),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11552 ));
    InMux I__10852 (
            .O(N__57157),
            .I(N__57151));
    InMux I__10851 (
            .O(N__57156),
            .I(N__57151));
    LocalMux I__10850 (
            .O(N__57151),
            .I(REG_mem_10_4));
    InMux I__10849 (
            .O(N__57148),
            .I(N__57145));
    LocalMux I__10848 (
            .O(N__57145),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13796 ));
    CascadeMux I__10847 (
            .O(N__57142),
            .I(N__57139));
    InMux I__10846 (
            .O(N__57139),
            .I(N__57136));
    LocalMux I__10845 (
            .O(N__57136),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11663 ));
    InMux I__10844 (
            .O(N__57133),
            .I(N__57130));
    LocalMux I__10843 (
            .O(N__57130),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11662 ));
    InMux I__10842 (
            .O(N__57127),
            .I(N__57124));
    LocalMux I__10841 (
            .O(N__57124),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11551 ));
    InMux I__10840 (
            .O(N__57121),
            .I(N__57115));
    InMux I__10839 (
            .O(N__57120),
            .I(N__57115));
    LocalMux I__10838 (
            .O(N__57115),
            .I(REG_mem_8_4));
    InMux I__10837 (
            .O(N__57112),
            .I(N__57108));
    InMux I__10836 (
            .O(N__57111),
            .I(N__57105));
    LocalMux I__10835 (
            .O(N__57108),
            .I(REG_mem_9_4));
    LocalMux I__10834 (
            .O(N__57105),
            .I(REG_mem_9_4));
    CascadeMux I__10833 (
            .O(N__57100),
            .I(\usb3_if_inst.n2755_cascade_ ));
    CascadeMux I__10832 (
            .O(N__57097),
            .I(\usb3_if_inst.n5_cascade_ ));
    CascadeMux I__10831 (
            .O(N__57094),
            .I(N__57091));
    InMux I__10830 (
            .O(N__57091),
            .I(N__57088));
    LocalMux I__10829 (
            .O(N__57088),
            .I(N__57085));
    Span4Mux_v I__10828 (
            .O(N__57085),
            .I(N__57082));
    Sp12to4 I__10827 (
            .O(N__57082),
            .I(N__57078));
    InMux I__10826 (
            .O(N__57081),
            .I(N__57075));
    Odrv12 I__10825 (
            .O(N__57078),
            .I(REG_mem_47_4));
    LocalMux I__10824 (
            .O(N__57075),
            .I(REG_mem_47_4));
    InMux I__10823 (
            .O(N__57070),
            .I(N__57067));
    LocalMux I__10822 (
            .O(N__57067),
            .I(N__57064));
    Span4Mux_h I__10821 (
            .O(N__57064),
            .I(N__57061));
    Span4Mux_h I__10820 (
            .O(N__57061),
            .I(N__57057));
    InMux I__10819 (
            .O(N__57060),
            .I(N__57054));
    Odrv4 I__10818 (
            .O(N__57057),
            .I(REG_mem_46_4));
    LocalMux I__10817 (
            .O(N__57054),
            .I(REG_mem_46_4));
    InMux I__10816 (
            .O(N__57049),
            .I(N__57046));
    LocalMux I__10815 (
            .O(N__57046),
            .I(N__57043));
    Span4Mux_v I__10814 (
            .O(N__57043),
            .I(N__57039));
    InMux I__10813 (
            .O(N__57042),
            .I(N__57036));
    Odrv4 I__10812 (
            .O(N__57039),
            .I(REG_mem_45_4));
    LocalMux I__10811 (
            .O(N__57036),
            .I(REG_mem_45_4));
    CascadeMux I__10810 (
            .O(N__57031),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12992_cascade_ ));
    InMux I__10809 (
            .O(N__57028),
            .I(N__57025));
    LocalMux I__10808 (
            .O(N__57025),
            .I(N__57021));
    InMux I__10807 (
            .O(N__57024),
            .I(N__57018));
    Span4Mux_v I__10806 (
            .O(N__57021),
            .I(N__57013));
    LocalMux I__10805 (
            .O(N__57018),
            .I(N__57013));
    Odrv4 I__10804 (
            .O(N__57013),
            .I(REG_mem_44_4));
    CascadeMux I__10803 (
            .O(N__57010),
            .I(N__57007));
    InMux I__10802 (
            .O(N__57007),
            .I(N__57004));
    LocalMux I__10801 (
            .O(N__57004),
            .I(N__57000));
    InMux I__10800 (
            .O(N__57003),
            .I(N__56997));
    Odrv4 I__10799 (
            .O(N__57000),
            .I(REG_mem_42_4));
    LocalMux I__10798 (
            .O(N__56997),
            .I(REG_mem_42_4));
    CascadeMux I__10797 (
            .O(N__56992),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13118_cascade_ ));
    InMux I__10796 (
            .O(N__56989),
            .I(N__56986));
    LocalMux I__10795 (
            .O(N__56986),
            .I(N__56983));
    Span4Mux_v I__10794 (
            .O(N__56983),
            .I(N__56979));
    InMux I__10793 (
            .O(N__56982),
            .I(N__56976));
    Odrv4 I__10792 (
            .O(N__56979),
            .I(REG_mem_40_4));
    LocalMux I__10791 (
            .O(N__56976),
            .I(REG_mem_40_4));
    InMux I__10790 (
            .O(N__56971),
            .I(N__56968));
    LocalMux I__10789 (
            .O(N__56968),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12995 ));
    CascadeMux I__10788 (
            .O(N__56965),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13121_cascade_ ));
    CascadeMux I__10787 (
            .O(N__56962),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13622_cascade_ ));
    CascadeMux I__10786 (
            .O(N__56959),
            .I(N__56956));
    InMux I__10785 (
            .O(N__56956),
            .I(N__56952));
    InMux I__10784 (
            .O(N__56955),
            .I(N__56949));
    LocalMux I__10783 (
            .O(N__56952),
            .I(REG_mem_36_4));
    LocalMux I__10782 (
            .O(N__56949),
            .I(REG_mem_36_4));
    InMux I__10781 (
            .O(N__56944),
            .I(N__56941));
    LocalMux I__10780 (
            .O(N__56941),
            .I(N__56937));
    InMux I__10779 (
            .O(N__56940),
            .I(N__56934));
    Odrv4 I__10778 (
            .O(N__56937),
            .I(REG_mem_37_4));
    LocalMux I__10777 (
            .O(N__56934),
            .I(REG_mem_37_4));
    InMux I__10776 (
            .O(N__56929),
            .I(N__56926));
    LocalMux I__10775 (
            .O(N__56926),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13181 ));
    InMux I__10774 (
            .O(N__56923),
            .I(N__56919));
    InMux I__10773 (
            .O(N__56922),
            .I(N__56916));
    LocalMux I__10772 (
            .O(N__56919),
            .I(REG_mem_11_4));
    LocalMux I__10771 (
            .O(N__56916),
            .I(REG_mem_11_4));
    InMux I__10770 (
            .O(N__56911),
            .I(N__56908));
    LocalMux I__10769 (
            .O(N__56908),
            .I(N__56905));
    Odrv12 I__10768 (
            .O(N__56905),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11639 ));
    InMux I__10767 (
            .O(N__56902),
            .I(N__56899));
    LocalMux I__10766 (
            .O(N__56899),
            .I(N__56895));
    InMux I__10765 (
            .O(N__56898),
            .I(N__56892));
    Odrv4 I__10764 (
            .O(N__56895),
            .I(REG_mem_63_5));
    LocalMux I__10763 (
            .O(N__56892),
            .I(REG_mem_63_5));
    CascadeMux I__10762 (
            .O(N__56887),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12986_cascade_ ));
    InMux I__10761 (
            .O(N__56884),
            .I(N__56881));
    LocalMux I__10760 (
            .O(N__56881),
            .I(N__56878));
    Sp12to4 I__10759 (
            .O(N__56878),
            .I(N__56875));
    Odrv12 I__10758 (
            .O(N__56875),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12989 ));
    CascadeMux I__10757 (
            .O(N__56872),
            .I(N__56868));
    InMux I__10756 (
            .O(N__56871),
            .I(N__56863));
    InMux I__10755 (
            .O(N__56868),
            .I(N__56863));
    LocalMux I__10754 (
            .O(N__56863),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_5 ));
    CascadeMux I__10753 (
            .O(N__56860),
            .I(N__56856));
    InMux I__10752 (
            .O(N__56859),
            .I(N__56851));
    InMux I__10751 (
            .O(N__56856),
            .I(N__56851));
    LocalMux I__10750 (
            .O(N__56851),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_5 ));
    CascadeMux I__10749 (
            .O(N__56848),
            .I(N__56844));
    InMux I__10748 (
            .O(N__56847),
            .I(N__56839));
    InMux I__10747 (
            .O(N__56844),
            .I(N__56839));
    LocalMux I__10746 (
            .O(N__56839),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_5 ));
    InMux I__10745 (
            .O(N__56836),
            .I(N__56833));
    LocalMux I__10744 (
            .O(N__56833),
            .I(N__56829));
    CascadeMux I__10743 (
            .O(N__56832),
            .I(N__56826));
    Span4Mux_v I__10742 (
            .O(N__56829),
            .I(N__56823));
    InMux I__10741 (
            .O(N__56826),
            .I(N__56820));
    Odrv4 I__10740 (
            .O(N__56823),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_5 ));
    LocalMux I__10739 (
            .O(N__56820),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_5 ));
    InMux I__10738 (
            .O(N__56815),
            .I(N__56812));
    LocalMux I__10737 (
            .O(N__56812),
            .I(N__56808));
    InMux I__10736 (
            .O(N__56811),
            .I(N__56805));
    Odrv12 I__10735 (
            .O(N__56808),
            .I(REG_mem_45_2));
    LocalMux I__10734 (
            .O(N__56805),
            .I(REG_mem_45_2));
    InMux I__10733 (
            .O(N__56800),
            .I(N__56797));
    LocalMux I__10732 (
            .O(N__56797),
            .I(N__56794));
    Span4Mux_v I__10731 (
            .O(N__56794),
            .I(N__56790));
    InMux I__10730 (
            .O(N__56793),
            .I(N__56787));
    Odrv4 I__10729 (
            .O(N__56790),
            .I(REG_mem_19_7));
    LocalMux I__10728 (
            .O(N__56787),
            .I(REG_mem_19_7));
    InMux I__10727 (
            .O(N__56782),
            .I(N__56779));
    LocalMux I__10726 (
            .O(N__56779),
            .I(N__56776));
    Span4Mux_v I__10725 (
            .O(N__56776),
            .I(N__56773));
    Odrv4 I__10724 (
            .O(N__56773),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13982 ));
    InMux I__10723 (
            .O(N__56770),
            .I(N__56767));
    LocalMux I__10722 (
            .O(N__56767),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14168 ));
    InMux I__10721 (
            .O(N__56764),
            .I(N__56760));
    InMux I__10720 (
            .O(N__56763),
            .I(N__56757));
    LocalMux I__10719 (
            .O(N__56760),
            .I(REG_mem_41_2));
    LocalMux I__10718 (
            .O(N__56757),
            .I(REG_mem_41_2));
    CascadeMux I__10717 (
            .O(N__56752),
            .I(N__56749));
    InMux I__10716 (
            .O(N__56749),
            .I(N__56745));
    InMux I__10715 (
            .O(N__56748),
            .I(N__56742));
    LocalMux I__10714 (
            .O(N__56745),
            .I(REG_mem_40_2));
    LocalMux I__10713 (
            .O(N__56742),
            .I(REG_mem_40_2));
    CascadeMux I__10712 (
            .O(N__56737),
            .I(N__56733));
    InMux I__10711 (
            .O(N__56736),
            .I(N__56728));
    InMux I__10710 (
            .O(N__56733),
            .I(N__56728));
    LocalMux I__10709 (
            .O(N__56728),
            .I(REG_mem_43_2));
    CascadeMux I__10708 (
            .O(N__56725),
            .I(N__56721));
    InMux I__10707 (
            .O(N__56724),
            .I(N__56718));
    InMux I__10706 (
            .O(N__56721),
            .I(N__56715));
    LocalMux I__10705 (
            .O(N__56718),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_5 ));
    LocalMux I__10704 (
            .O(N__56715),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_5 ));
    InMux I__10703 (
            .O(N__56710),
            .I(N__56704));
    InMux I__10702 (
            .O(N__56709),
            .I(N__56704));
    LocalMux I__10701 (
            .O(N__56704),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_2 ));
    InMux I__10700 (
            .O(N__56701),
            .I(N__56698));
    LocalMux I__10699 (
            .O(N__56698),
            .I(N__56694));
    InMux I__10698 (
            .O(N__56697),
            .I(N__56691));
    Odrv4 I__10697 (
            .O(N__56694),
            .I(REG_mem_31_5));
    LocalMux I__10696 (
            .O(N__56691),
            .I(REG_mem_31_5));
    InMux I__10695 (
            .O(N__56686),
            .I(N__56683));
    LocalMux I__10694 (
            .O(N__56683),
            .I(N__56680));
    Span4Mux_h I__10693 (
            .O(N__56680),
            .I(N__56676));
    InMux I__10692 (
            .O(N__56679),
            .I(N__56673));
    Odrv4 I__10691 (
            .O(N__56676),
            .I(REG_mem_47_2));
    LocalMux I__10690 (
            .O(N__56673),
            .I(REG_mem_47_2));
    InMux I__10689 (
            .O(N__56668),
            .I(N__56662));
    InMux I__10688 (
            .O(N__56667),
            .I(N__56662));
    LocalMux I__10687 (
            .O(N__56662),
            .I(REG_mem_44_2));
    CascadeMux I__10686 (
            .O(N__56659),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14084_cascade_ ));
    CascadeMux I__10685 (
            .O(N__56656),
            .I(N__56653));
    InMux I__10684 (
            .O(N__56653),
            .I(N__56647));
    InMux I__10683 (
            .O(N__56652),
            .I(N__56647));
    LocalMux I__10682 (
            .O(N__56647),
            .I(REG_mem_46_2));
    InMux I__10681 (
            .O(N__56644),
            .I(N__56640));
    InMux I__10680 (
            .O(N__56643),
            .I(N__56637));
    LocalMux I__10679 (
            .O(N__56640),
            .I(REG_mem_26_5));
    LocalMux I__10678 (
            .O(N__56637),
            .I(REG_mem_26_5));
    InMux I__10677 (
            .O(N__56632),
            .I(N__56629));
    LocalMux I__10676 (
            .O(N__56629),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11981 ));
    CascadeMux I__10675 (
            .O(N__56626),
            .I(N__56621));
    InMux I__10674 (
            .O(N__56625),
            .I(N__56616));
    InMux I__10673 (
            .O(N__56624),
            .I(N__56610));
    InMux I__10672 (
            .O(N__56621),
            .I(N__56607));
    CascadeMux I__10671 (
            .O(N__56620),
            .I(N__56600));
    InMux I__10670 (
            .O(N__56619),
            .I(N__56596));
    LocalMux I__10669 (
            .O(N__56616),
            .I(N__56589));
    InMux I__10668 (
            .O(N__56615),
            .I(N__56586));
    InMux I__10667 (
            .O(N__56614),
            .I(N__56583));
    InMux I__10666 (
            .O(N__56613),
            .I(N__56580));
    LocalMux I__10665 (
            .O(N__56610),
            .I(N__56575));
    LocalMux I__10664 (
            .O(N__56607),
            .I(N__56575));
    CascadeMux I__10663 (
            .O(N__56606),
            .I(N__56572));
    InMux I__10662 (
            .O(N__56605),
            .I(N__56558));
    InMux I__10661 (
            .O(N__56604),
            .I(N__56558));
    InMux I__10660 (
            .O(N__56603),
            .I(N__56558));
    InMux I__10659 (
            .O(N__56600),
            .I(N__56550));
    InMux I__10658 (
            .O(N__56599),
            .I(N__56550));
    LocalMux I__10657 (
            .O(N__56596),
            .I(N__56543));
    InMux I__10656 (
            .O(N__56595),
            .I(N__56538));
    InMux I__10655 (
            .O(N__56594),
            .I(N__56538));
    InMux I__10654 (
            .O(N__56593),
            .I(N__56535));
    InMux I__10653 (
            .O(N__56592),
            .I(N__56532));
    Span4Mux_v I__10652 (
            .O(N__56589),
            .I(N__56527));
    LocalMux I__10651 (
            .O(N__56586),
            .I(N__56527));
    LocalMux I__10650 (
            .O(N__56583),
            .I(N__56524));
    LocalMux I__10649 (
            .O(N__56580),
            .I(N__56521));
    Span4Mux_h I__10648 (
            .O(N__56575),
            .I(N__56504));
    InMux I__10647 (
            .O(N__56572),
            .I(N__56499));
    InMux I__10646 (
            .O(N__56571),
            .I(N__56499));
    InMux I__10645 (
            .O(N__56570),
            .I(N__56494));
    InMux I__10644 (
            .O(N__56569),
            .I(N__56494));
    CascadeMux I__10643 (
            .O(N__56568),
            .I(N__56491));
    InMux I__10642 (
            .O(N__56567),
            .I(N__56483));
    InMux I__10641 (
            .O(N__56566),
            .I(N__56483));
    InMux I__10640 (
            .O(N__56565),
            .I(N__56480));
    LocalMux I__10639 (
            .O(N__56558),
            .I(N__56477));
    InMux I__10638 (
            .O(N__56557),
            .I(N__56466));
    InMux I__10637 (
            .O(N__56556),
            .I(N__56466));
    InMux I__10636 (
            .O(N__56555),
            .I(N__56466));
    LocalMux I__10635 (
            .O(N__56550),
            .I(N__56463));
    CascadeMux I__10634 (
            .O(N__56549),
            .I(N__56460));
    InMux I__10633 (
            .O(N__56548),
            .I(N__56450));
    InMux I__10632 (
            .O(N__56547),
            .I(N__56450));
    InMux I__10631 (
            .O(N__56546),
            .I(N__56450));
    Span4Mux_h I__10630 (
            .O(N__56543),
            .I(N__56443));
    LocalMux I__10629 (
            .O(N__56538),
            .I(N__56443));
    LocalMux I__10628 (
            .O(N__56535),
            .I(N__56443));
    LocalMux I__10627 (
            .O(N__56532),
            .I(N__56438));
    Span4Mux_v I__10626 (
            .O(N__56527),
            .I(N__56438));
    Span4Mux_h I__10625 (
            .O(N__56524),
            .I(N__56433));
    Span4Mux_v I__10624 (
            .O(N__56521),
            .I(N__56433));
    InMux I__10623 (
            .O(N__56520),
            .I(N__56430));
    InMux I__10622 (
            .O(N__56519),
            .I(N__56421));
    InMux I__10621 (
            .O(N__56518),
            .I(N__56421));
    InMux I__10620 (
            .O(N__56517),
            .I(N__56421));
    InMux I__10619 (
            .O(N__56516),
            .I(N__56421));
    InMux I__10618 (
            .O(N__56515),
            .I(N__56416));
    InMux I__10617 (
            .O(N__56514),
            .I(N__56416));
    InMux I__10616 (
            .O(N__56513),
            .I(N__56410));
    InMux I__10615 (
            .O(N__56512),
            .I(N__56410));
    InMux I__10614 (
            .O(N__56511),
            .I(N__56403));
    InMux I__10613 (
            .O(N__56510),
            .I(N__56403));
    InMux I__10612 (
            .O(N__56509),
            .I(N__56400));
    InMux I__10611 (
            .O(N__56508),
            .I(N__56395));
    InMux I__10610 (
            .O(N__56507),
            .I(N__56395));
    Span4Mux_h I__10609 (
            .O(N__56504),
            .I(N__56388));
    LocalMux I__10608 (
            .O(N__56499),
            .I(N__56388));
    LocalMux I__10607 (
            .O(N__56494),
            .I(N__56388));
    InMux I__10606 (
            .O(N__56491),
            .I(N__56383));
    InMux I__10605 (
            .O(N__56490),
            .I(N__56383));
    InMux I__10604 (
            .O(N__56489),
            .I(N__56378));
    InMux I__10603 (
            .O(N__56488),
            .I(N__56378));
    LocalMux I__10602 (
            .O(N__56483),
            .I(N__56375));
    LocalMux I__10601 (
            .O(N__56480),
            .I(N__56370));
    Span4Mux_h I__10600 (
            .O(N__56477),
            .I(N__56370));
    InMux I__10599 (
            .O(N__56476),
            .I(N__56367));
    InMux I__10598 (
            .O(N__56475),
            .I(N__56364));
    InMux I__10597 (
            .O(N__56474),
            .I(N__56359));
    InMux I__10596 (
            .O(N__56473),
            .I(N__56359));
    LocalMux I__10595 (
            .O(N__56466),
            .I(N__56354));
    Span4Mux_v I__10594 (
            .O(N__56463),
            .I(N__56354));
    InMux I__10593 (
            .O(N__56460),
            .I(N__56343));
    InMux I__10592 (
            .O(N__56459),
            .I(N__56343));
    InMux I__10591 (
            .O(N__56458),
            .I(N__56343));
    InMux I__10590 (
            .O(N__56457),
            .I(N__56343));
    LocalMux I__10589 (
            .O(N__56450),
            .I(N__56340));
    Span4Mux_v I__10588 (
            .O(N__56443),
            .I(N__56333));
    Span4Mux_v I__10587 (
            .O(N__56438),
            .I(N__56333));
    Span4Mux_h I__10586 (
            .O(N__56433),
            .I(N__56333));
    LocalMux I__10585 (
            .O(N__56430),
            .I(N__56322));
    LocalMux I__10584 (
            .O(N__56421),
            .I(N__56322));
    LocalMux I__10583 (
            .O(N__56416),
            .I(N__56322));
    InMux I__10582 (
            .O(N__56415),
            .I(N__56319));
    LocalMux I__10581 (
            .O(N__56410),
            .I(N__56316));
    InMux I__10580 (
            .O(N__56409),
            .I(N__56313));
    InMux I__10579 (
            .O(N__56408),
            .I(N__56310));
    LocalMux I__10578 (
            .O(N__56403),
            .I(N__56301));
    LocalMux I__10577 (
            .O(N__56400),
            .I(N__56301));
    LocalMux I__10576 (
            .O(N__56395),
            .I(N__56301));
    Sp12to4 I__10575 (
            .O(N__56388),
            .I(N__56301));
    LocalMux I__10574 (
            .O(N__56383),
            .I(N__56298));
    LocalMux I__10573 (
            .O(N__56378),
            .I(N__56295));
    Span4Mux_v I__10572 (
            .O(N__56375),
            .I(N__56290));
    Span4Mux_v I__10571 (
            .O(N__56370),
            .I(N__56290));
    LocalMux I__10570 (
            .O(N__56367),
            .I(N__56281));
    LocalMux I__10569 (
            .O(N__56364),
            .I(N__56281));
    LocalMux I__10568 (
            .O(N__56359),
            .I(N__56281));
    Span4Mux_v I__10567 (
            .O(N__56354),
            .I(N__56281));
    InMux I__10566 (
            .O(N__56353),
            .I(N__56278));
    InMux I__10565 (
            .O(N__56352),
            .I(N__56275));
    LocalMux I__10564 (
            .O(N__56343),
            .I(N__56268));
    Span4Mux_v I__10563 (
            .O(N__56340),
            .I(N__56268));
    Span4Mux_h I__10562 (
            .O(N__56333),
            .I(N__56268));
    InMux I__10561 (
            .O(N__56332),
            .I(N__56263));
    InMux I__10560 (
            .O(N__56331),
            .I(N__56263));
    InMux I__10559 (
            .O(N__56330),
            .I(N__56258));
    InMux I__10558 (
            .O(N__56329),
            .I(N__56258));
    Span4Mux_v I__10557 (
            .O(N__56322),
            .I(N__56255));
    LocalMux I__10556 (
            .O(N__56319),
            .I(N__56250));
    Sp12to4 I__10555 (
            .O(N__56316),
            .I(N__56250));
    LocalMux I__10554 (
            .O(N__56313),
            .I(N__56243));
    LocalMux I__10553 (
            .O(N__56310),
            .I(N__56243));
    Span12Mux_v I__10552 (
            .O(N__56301),
            .I(N__56243));
    Span4Mux_v I__10551 (
            .O(N__56298),
            .I(N__56234));
    Span4Mux_v I__10550 (
            .O(N__56295),
            .I(N__56234));
    Span4Mux_v I__10549 (
            .O(N__56290),
            .I(N__56234));
    Span4Mux_v I__10548 (
            .O(N__56281),
            .I(N__56234));
    LocalMux I__10547 (
            .O(N__56278),
            .I(N__56227));
    LocalMux I__10546 (
            .O(N__56275),
            .I(N__56227));
    Span4Mux_h I__10545 (
            .O(N__56268),
            .I(N__56227));
    LocalMux I__10544 (
            .O(N__56263),
            .I(dc32_fifo_data_in_9));
    LocalMux I__10543 (
            .O(N__56258),
            .I(dc32_fifo_data_in_9));
    Odrv4 I__10542 (
            .O(N__56255),
            .I(dc32_fifo_data_in_9));
    Odrv12 I__10541 (
            .O(N__56250),
            .I(dc32_fifo_data_in_9));
    Odrv12 I__10540 (
            .O(N__56243),
            .I(dc32_fifo_data_in_9));
    Odrv4 I__10539 (
            .O(N__56234),
            .I(dc32_fifo_data_in_9));
    Odrv4 I__10538 (
            .O(N__56227),
            .I(dc32_fifo_data_in_9));
    InMux I__10537 (
            .O(N__56212),
            .I(N__56209));
    LocalMux I__10536 (
            .O(N__56209),
            .I(N__56206));
    Span4Mux_v I__10535 (
            .O(N__56206),
            .I(N__56203));
    Span4Mux_h I__10534 (
            .O(N__56203),
            .I(N__56199));
    InMux I__10533 (
            .O(N__56202),
            .I(N__56196));
    Odrv4 I__10532 (
            .O(N__56199),
            .I(REG_mem_6_9));
    LocalMux I__10531 (
            .O(N__56196),
            .I(REG_mem_6_9));
    InMux I__10530 (
            .O(N__56191),
            .I(N__56188));
    LocalMux I__10529 (
            .O(N__56188),
            .I(N__56184));
    CascadeMux I__10528 (
            .O(N__56187),
            .I(N__56181));
    Span4Mux_h I__10527 (
            .O(N__56184),
            .I(N__56178));
    InMux I__10526 (
            .O(N__56181),
            .I(N__56175));
    Odrv4 I__10525 (
            .O(N__56178),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_5 ));
    LocalMux I__10524 (
            .O(N__56175),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_5 ));
    InMux I__10523 (
            .O(N__56170),
            .I(N__56167));
    LocalMux I__10522 (
            .O(N__56167),
            .I(N__56164));
    Odrv4 I__10521 (
            .O(N__56164),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12025 ));
    InMux I__10520 (
            .O(N__56161),
            .I(N__56155));
    InMux I__10519 (
            .O(N__56160),
            .I(N__56155));
    LocalMux I__10518 (
            .O(N__56155),
            .I(REG_mem_63_2));
    CascadeMux I__10517 (
            .O(N__56152),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13604_cascade_ ));
    InMux I__10516 (
            .O(N__56149),
            .I(N__56146));
    LocalMux I__10515 (
            .O(N__56146),
            .I(N__56143));
    Span4Mux_v I__10514 (
            .O(N__56143),
            .I(N__56140));
    Span4Mux_h I__10513 (
            .O(N__56140),
            .I(N__56136));
    InMux I__10512 (
            .O(N__56139),
            .I(N__56133));
    Odrv4 I__10511 (
            .O(N__56136),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_2 ));
    LocalMux I__10510 (
            .O(N__56133),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_2 ));
    InMux I__10509 (
            .O(N__56128),
            .I(N__56122));
    InMux I__10508 (
            .O(N__56127),
            .I(N__56122));
    LocalMux I__10507 (
            .O(N__56122),
            .I(N__56119));
    Odrv4 I__10506 (
            .O(N__56119),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_2 ));
    InMux I__10505 (
            .O(N__56116),
            .I(N__56113));
    LocalMux I__10504 (
            .O(N__56113),
            .I(N__56110));
    Span4Mux_v I__10503 (
            .O(N__56110),
            .I(N__56106));
    InMux I__10502 (
            .O(N__56109),
            .I(N__56103));
    Odrv4 I__10501 (
            .O(N__56106),
            .I(REG_mem_11_5));
    LocalMux I__10500 (
            .O(N__56103),
            .I(REG_mem_11_5));
    InMux I__10499 (
            .O(N__56098),
            .I(N__56095));
    LocalMux I__10498 (
            .O(N__56095),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13850 ));
    InMux I__10497 (
            .O(N__56092),
            .I(N__56089));
    LocalMux I__10496 (
            .O(N__56089),
            .I(N__56086));
    Span4Mux_v I__10495 (
            .O(N__56086),
            .I(N__56082));
    InMux I__10494 (
            .O(N__56085),
            .I(N__56079));
    Odrv4 I__10493 (
            .O(N__56082),
            .I(REG_mem_17_2));
    LocalMux I__10492 (
            .O(N__56079),
            .I(REG_mem_17_2));
    InMux I__10491 (
            .O(N__56074),
            .I(N__56068));
    InMux I__10490 (
            .O(N__56073),
            .I(N__56068));
    LocalMux I__10489 (
            .O(N__56068),
            .I(REG_mem_16_2));
    InMux I__10488 (
            .O(N__56065),
            .I(N__56062));
    LocalMux I__10487 (
            .O(N__56062),
            .I(N__56058));
    InMux I__10486 (
            .O(N__56061),
            .I(N__56055));
    Odrv4 I__10485 (
            .O(N__56058),
            .I(REG_mem_9_5));
    LocalMux I__10484 (
            .O(N__56055),
            .I(REG_mem_9_5));
    CascadeMux I__10483 (
            .O(N__56050),
            .I(N__56047));
    InMux I__10482 (
            .O(N__56047),
            .I(N__56043));
    InMux I__10481 (
            .O(N__56046),
            .I(N__56040));
    LocalMux I__10480 (
            .O(N__56043),
            .I(REG_mem_8_5));
    LocalMux I__10479 (
            .O(N__56040),
            .I(REG_mem_8_5));
    InMux I__10478 (
            .O(N__56035),
            .I(N__56029));
    InMux I__10477 (
            .O(N__56034),
            .I(N__56029));
    LocalMux I__10476 (
            .O(N__56029),
            .I(REG_mem_10_5));
    CascadeMux I__10475 (
            .O(N__56026),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12026_cascade_ ));
    InMux I__10474 (
            .O(N__56023),
            .I(N__56020));
    LocalMux I__10473 (
            .O(N__56020),
            .I(N__56017));
    Odrv4 I__10472 (
            .O(N__56017),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11980 ));
    CascadeMux I__10471 (
            .O(N__56014),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14282_cascade_ ));
    InMux I__10470 (
            .O(N__56011),
            .I(N__56008));
    LocalMux I__10469 (
            .O(N__56008),
            .I(N__56005));
    Odrv4 I__10468 (
            .O(N__56005),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12512 ));
    InMux I__10467 (
            .O(N__56002),
            .I(N__55999));
    LocalMux I__10466 (
            .O(N__55999),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13853 ));
    CascadeMux I__10465 (
            .O(N__55996),
            .I(N__55993));
    InMux I__10464 (
            .O(N__55993),
            .I(N__55990));
    LocalMux I__10463 (
            .O(N__55990),
            .I(N__55987));
    Span4Mux_v I__10462 (
            .O(N__55987),
            .I(N__55984));
    Span4Mux_v I__10461 (
            .O(N__55984),
            .I(N__55981));
    Sp12to4 I__10460 (
            .O(N__55981),
            .I(N__55977));
    InMux I__10459 (
            .O(N__55980),
            .I(N__55974));
    Odrv12 I__10458 (
            .O(N__55977),
            .I(REG_mem_18_5));
    LocalMux I__10457 (
            .O(N__55974),
            .I(REG_mem_18_5));
    CascadeMux I__10456 (
            .O(N__55969),
            .I(N__55966));
    InMux I__10455 (
            .O(N__55966),
            .I(N__55963));
    LocalMux I__10454 (
            .O(N__55963),
            .I(N__55959));
    InMux I__10453 (
            .O(N__55962),
            .I(N__55956));
    Odrv4 I__10452 (
            .O(N__55959),
            .I(REG_mem_23_5));
    LocalMux I__10451 (
            .O(N__55956),
            .I(REG_mem_23_5));
    InMux I__10450 (
            .O(N__55951),
            .I(N__55948));
    LocalMux I__10449 (
            .O(N__55948),
            .I(N__55944));
    CascadeMux I__10448 (
            .O(N__55947),
            .I(N__55941));
    Span4Mux_v I__10447 (
            .O(N__55944),
            .I(N__55938));
    InMux I__10446 (
            .O(N__55941),
            .I(N__55935));
    Odrv4 I__10445 (
            .O(N__55938),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_5 ));
    LocalMux I__10444 (
            .O(N__55935),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_5 ));
    InMux I__10443 (
            .O(N__55930),
            .I(N__55927));
    LocalMux I__10442 (
            .O(N__55927),
            .I(N__55923));
    CascadeMux I__10441 (
            .O(N__55926),
            .I(N__55920));
    Span4Mux_v I__10440 (
            .O(N__55923),
            .I(N__55917));
    InMux I__10439 (
            .O(N__55920),
            .I(N__55914));
    Odrv4 I__10438 (
            .O(N__55917),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_5 ));
    LocalMux I__10437 (
            .O(N__55914),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_5 ));
    CascadeMux I__10436 (
            .O(N__55909),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12872_cascade_ ));
    InMux I__10435 (
            .O(N__55906),
            .I(N__55903));
    LocalMux I__10434 (
            .O(N__55903),
            .I(N__55900));
    Span4Mux_v I__10433 (
            .O(N__55900),
            .I(N__55896));
    CascadeMux I__10432 (
            .O(N__55899),
            .I(N__55893));
    Span4Mux_h I__10431 (
            .O(N__55896),
            .I(N__55890));
    InMux I__10430 (
            .O(N__55893),
            .I(N__55887));
    Odrv4 I__10429 (
            .O(N__55890),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_5 ));
    LocalMux I__10428 (
            .O(N__55887),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_5 ));
    CascadeMux I__10427 (
            .O(N__55882),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12875_cascade_ ));
    CascadeMux I__10426 (
            .O(N__55879),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12511_cascade_ ));
    InMux I__10425 (
            .O(N__55876),
            .I(N__55873));
    LocalMux I__10424 (
            .O(N__55873),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12500 ));
    CascadeMux I__10423 (
            .O(N__55870),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13250_cascade_ ));
    InMux I__10422 (
            .O(N__55867),
            .I(N__55864));
    LocalMux I__10421 (
            .O(N__55864),
            .I(N__55861));
    Odrv4 I__10420 (
            .O(N__55861),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12499 ));
    InMux I__10419 (
            .O(N__55858),
            .I(N__55855));
    LocalMux I__10418 (
            .O(N__55855),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13514 ));
    CascadeMux I__10417 (
            .O(N__55852),
            .I(N__55849));
    InMux I__10416 (
            .O(N__55849),
            .I(N__55846));
    LocalMux I__10415 (
            .O(N__55846),
            .I(N__55843));
    Span4Mux_v I__10414 (
            .O(N__55843),
            .I(N__55839));
    InMux I__10413 (
            .O(N__55842),
            .I(N__55836));
    Odrv4 I__10412 (
            .O(N__55839),
            .I(REG_mem_16_5));
    LocalMux I__10411 (
            .O(N__55836),
            .I(REG_mem_16_5));
    InMux I__10410 (
            .O(N__55831),
            .I(N__55828));
    LocalMux I__10409 (
            .O(N__55828),
            .I(N__55824));
    InMux I__10408 (
            .O(N__55827),
            .I(N__55821));
    Odrv12 I__10407 (
            .O(N__55824),
            .I(REG_mem_17_5));
    LocalMux I__10406 (
            .O(N__55821),
            .I(REG_mem_17_5));
    InMux I__10405 (
            .O(N__55816),
            .I(N__55813));
    LocalMux I__10404 (
            .O(N__55813),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13517 ));
    InMux I__10403 (
            .O(N__55810),
            .I(N__55807));
    LocalMux I__10402 (
            .O(N__55807),
            .I(N__55804));
    Span4Mux_v I__10401 (
            .O(N__55804),
            .I(N__55801));
    Span4Mux_h I__10400 (
            .O(N__55801),
            .I(N__55797));
    InMux I__10399 (
            .O(N__55800),
            .I(N__55794));
    Odrv4 I__10398 (
            .O(N__55797),
            .I(REG_mem_16_1));
    LocalMux I__10397 (
            .O(N__55794),
            .I(REG_mem_16_1));
    InMux I__10396 (
            .O(N__55789),
            .I(N__55786));
    LocalMux I__10395 (
            .O(N__55786),
            .I(N__55782));
    InMux I__10394 (
            .O(N__55785),
            .I(N__55779));
    Odrv4 I__10393 (
            .O(N__55782),
            .I(REG_mem_17_1));
    LocalMux I__10392 (
            .O(N__55779),
            .I(REG_mem_17_1));
    InMux I__10391 (
            .O(N__55774),
            .I(N__55771));
    LocalMux I__10390 (
            .O(N__55771),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11677 ));
    CascadeMux I__10389 (
            .O(N__55768),
            .I(N__55760));
    InMux I__10388 (
            .O(N__55767),
            .I(N__55757));
    CascadeMux I__10387 (
            .O(N__55766),
            .I(N__55753));
    CascadeMux I__10386 (
            .O(N__55765),
            .I(N__55749));
    CascadeMux I__10385 (
            .O(N__55764),
            .I(N__55745));
    CascadeMux I__10384 (
            .O(N__55763),
            .I(N__55741));
    InMux I__10383 (
            .O(N__55760),
            .I(N__55737));
    LocalMux I__10382 (
            .O(N__55757),
            .I(N__55734));
    InMux I__10381 (
            .O(N__55756),
            .I(N__55717));
    InMux I__10380 (
            .O(N__55753),
            .I(N__55717));
    InMux I__10379 (
            .O(N__55752),
            .I(N__55717));
    InMux I__10378 (
            .O(N__55749),
            .I(N__55717));
    InMux I__10377 (
            .O(N__55748),
            .I(N__55717));
    InMux I__10376 (
            .O(N__55745),
            .I(N__55717));
    InMux I__10375 (
            .O(N__55744),
            .I(N__55717));
    InMux I__10374 (
            .O(N__55741),
            .I(N__55717));
    InMux I__10373 (
            .O(N__55740),
            .I(N__55714));
    LocalMux I__10372 (
            .O(N__55737),
            .I(\spi0.n1979 ));
    Odrv4 I__10371 (
            .O(N__55734),
            .I(\spi0.n1979 ));
    LocalMux I__10370 (
            .O(N__55717),
            .I(\spi0.n1979 ));
    LocalMux I__10369 (
            .O(N__55714),
            .I(\spi0.n1979 ));
    InMux I__10368 (
            .O(N__55705),
            .I(\spi0.n10659 ));
    CEMux I__10367 (
            .O(N__55702),
            .I(N__55698));
    InMux I__10366 (
            .O(N__55701),
            .I(N__55695));
    LocalMux I__10365 (
            .O(N__55698),
            .I(N__55692));
    LocalMux I__10364 (
            .O(N__55695),
            .I(\spi0.n4281 ));
    Odrv4 I__10363 (
            .O(N__55692),
            .I(\spi0.n4281 ));
    SRMux I__10362 (
            .O(N__55687),
            .I(N__55684));
    LocalMux I__10361 (
            .O(N__55684),
            .I(N__55681));
    Odrv12 I__10360 (
            .O(N__55681),
            .I(\spi0.n4455 ));
    InMux I__10359 (
            .O(N__55678),
            .I(N__55675));
    LocalMux I__10358 (
            .O(N__55675),
            .I(N__55672));
    Odrv12 I__10357 (
            .O(N__55672),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13364 ));
    CascadeMux I__10356 (
            .O(N__55669),
            .I(N__55666));
    InMux I__10355 (
            .O(N__55666),
            .I(N__55663));
    LocalMux I__10354 (
            .O(N__55663),
            .I(N__55660));
    Span4Mux_v I__10353 (
            .O(N__55660),
            .I(N__55657));
    Odrv4 I__10352 (
            .O(N__55657),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11719 ));
    InMux I__10351 (
            .O(N__55654),
            .I(N__55651));
    LocalMux I__10350 (
            .O(N__55651),
            .I(N__55648));
    Odrv12 I__10349 (
            .O(N__55648),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13367 ));
    InMux I__10348 (
            .O(N__55645),
            .I(N__55639));
    InMux I__10347 (
            .O(N__55644),
            .I(N__55639));
    LocalMux I__10346 (
            .O(N__55639),
            .I(REG_mem_50_1));
    InMux I__10345 (
            .O(N__55636),
            .I(N__55633));
    LocalMux I__10344 (
            .O(N__55633),
            .I(N__55629));
    InMux I__10343 (
            .O(N__55632),
            .I(N__55626));
    Odrv4 I__10342 (
            .O(N__55629),
            .I(REG_mem_51_1));
    LocalMux I__10341 (
            .O(N__55626),
            .I(REG_mem_51_1));
    InMux I__10340 (
            .O(N__55621),
            .I(N__55618));
    LocalMux I__10339 (
            .O(N__55618),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11720 ));
    CascadeMux I__10338 (
            .O(N__55615),
            .I(N__55609));
    CascadeMux I__10337 (
            .O(N__55614),
            .I(N__55604));
    CascadeMux I__10336 (
            .O(N__55613),
            .I(N__55600));
    CascadeMux I__10335 (
            .O(N__55612),
            .I(N__55596));
    InMux I__10334 (
            .O(N__55609),
            .I(N__55591));
    InMux I__10333 (
            .O(N__55608),
            .I(N__55591));
    InMux I__10332 (
            .O(N__55607),
            .I(N__55574));
    InMux I__10331 (
            .O(N__55604),
            .I(N__55571));
    InMux I__10330 (
            .O(N__55603),
            .I(N__55562));
    InMux I__10329 (
            .O(N__55600),
            .I(N__55562));
    InMux I__10328 (
            .O(N__55599),
            .I(N__55562));
    InMux I__10327 (
            .O(N__55596),
            .I(N__55562));
    LocalMux I__10326 (
            .O(N__55591),
            .I(N__55559));
    InMux I__10325 (
            .O(N__55590),
            .I(N__55554));
    InMux I__10324 (
            .O(N__55589),
            .I(N__55554));
    InMux I__10323 (
            .O(N__55588),
            .I(N__55551));
    InMux I__10322 (
            .O(N__55587),
            .I(N__55544));
    InMux I__10321 (
            .O(N__55586),
            .I(N__55544));
    InMux I__10320 (
            .O(N__55585),
            .I(N__55544));
    InMux I__10319 (
            .O(N__55584),
            .I(N__55533));
    InMux I__10318 (
            .O(N__55583),
            .I(N__55533));
    InMux I__10317 (
            .O(N__55582),
            .I(N__55533));
    InMux I__10316 (
            .O(N__55581),
            .I(N__55533));
    InMux I__10315 (
            .O(N__55580),
            .I(N__55533));
    InMux I__10314 (
            .O(N__55579),
            .I(N__55526));
    InMux I__10313 (
            .O(N__55578),
            .I(N__55526));
    InMux I__10312 (
            .O(N__55577),
            .I(N__55526));
    LocalMux I__10311 (
            .O(N__55574),
            .I(\spi0.state_1 ));
    LocalMux I__10310 (
            .O(N__55571),
            .I(\spi0.state_1 ));
    LocalMux I__10309 (
            .O(N__55562),
            .I(\spi0.state_1 ));
    Odrv12 I__10308 (
            .O(N__55559),
            .I(\spi0.state_1 ));
    LocalMux I__10307 (
            .O(N__55554),
            .I(\spi0.state_1 ));
    LocalMux I__10306 (
            .O(N__55551),
            .I(\spi0.state_1 ));
    LocalMux I__10305 (
            .O(N__55544),
            .I(\spi0.state_1 ));
    LocalMux I__10304 (
            .O(N__55533),
            .I(\spi0.state_1 ));
    LocalMux I__10303 (
            .O(N__55526),
            .I(\spi0.state_1 ));
    CascadeMux I__10302 (
            .O(N__55507),
            .I(\spi0.n1979_cascade_ ));
    InMux I__10301 (
            .O(N__55504),
            .I(N__55501));
    LocalMux I__10300 (
            .O(N__55501),
            .I(\spi0.n12586 ));
    CascadeMux I__10299 (
            .O(N__55498),
            .I(N__55494));
    CascadeMux I__10298 (
            .O(N__55497),
            .I(N__55490));
    InMux I__10297 (
            .O(N__55494),
            .I(N__55484));
    InMux I__10296 (
            .O(N__55493),
            .I(N__55467));
    InMux I__10295 (
            .O(N__55490),
            .I(N__55467));
    InMux I__10294 (
            .O(N__55489),
            .I(N__55467));
    InMux I__10293 (
            .O(N__55488),
            .I(N__55467));
    InMux I__10292 (
            .O(N__55487),
            .I(N__55467));
    LocalMux I__10291 (
            .O(N__55484),
            .I(N__55456));
    InMux I__10290 (
            .O(N__55483),
            .I(N__55447));
    InMux I__10289 (
            .O(N__55482),
            .I(N__55447));
    InMux I__10288 (
            .O(N__55481),
            .I(N__55447));
    InMux I__10287 (
            .O(N__55480),
            .I(N__55447));
    InMux I__10286 (
            .O(N__55479),
            .I(N__55443));
    CascadeMux I__10285 (
            .O(N__55478),
            .I(N__55440));
    LocalMux I__10284 (
            .O(N__55467),
            .I(N__55427));
    InMux I__10283 (
            .O(N__55466),
            .I(N__55420));
    InMux I__10282 (
            .O(N__55465),
            .I(N__55420));
    InMux I__10281 (
            .O(N__55464),
            .I(N__55420));
    InMux I__10280 (
            .O(N__55463),
            .I(N__55417));
    InMux I__10279 (
            .O(N__55462),
            .I(N__55408));
    InMux I__10278 (
            .O(N__55461),
            .I(N__55408));
    InMux I__10277 (
            .O(N__55460),
            .I(N__55408));
    InMux I__10276 (
            .O(N__55459),
            .I(N__55408));
    Span4Mux_v I__10275 (
            .O(N__55456),
            .I(N__55403));
    LocalMux I__10274 (
            .O(N__55447),
            .I(N__55403));
    InMux I__10273 (
            .O(N__55446),
            .I(N__55400));
    LocalMux I__10272 (
            .O(N__55443),
            .I(N__55397));
    InMux I__10271 (
            .O(N__55440),
            .I(N__55392));
    InMux I__10270 (
            .O(N__55439),
            .I(N__55392));
    InMux I__10269 (
            .O(N__55438),
            .I(N__55383));
    InMux I__10268 (
            .O(N__55437),
            .I(N__55383));
    InMux I__10267 (
            .O(N__55436),
            .I(N__55383));
    InMux I__10266 (
            .O(N__55435),
            .I(N__55383));
    InMux I__10265 (
            .O(N__55434),
            .I(N__55372));
    InMux I__10264 (
            .O(N__55433),
            .I(N__55372));
    InMux I__10263 (
            .O(N__55432),
            .I(N__55372));
    InMux I__10262 (
            .O(N__55431),
            .I(N__55372));
    InMux I__10261 (
            .O(N__55430),
            .I(N__55372));
    Odrv4 I__10260 (
            .O(N__55427),
            .I(\spi0.state_3 ));
    LocalMux I__10259 (
            .O(N__55420),
            .I(\spi0.state_3 ));
    LocalMux I__10258 (
            .O(N__55417),
            .I(\spi0.state_3 ));
    LocalMux I__10257 (
            .O(N__55408),
            .I(\spi0.state_3 ));
    Odrv4 I__10256 (
            .O(N__55403),
            .I(\spi0.state_3 ));
    LocalMux I__10255 (
            .O(N__55400),
            .I(\spi0.state_3 ));
    Odrv4 I__10254 (
            .O(N__55397),
            .I(\spi0.state_3 ));
    LocalMux I__10253 (
            .O(N__55392),
            .I(\spi0.state_3 ));
    LocalMux I__10252 (
            .O(N__55383),
            .I(\spi0.state_3 ));
    LocalMux I__10251 (
            .O(N__55372),
            .I(\spi0.state_3 ));
    CEMux I__10250 (
            .O(N__55351),
            .I(N__55348));
    LocalMux I__10249 (
            .O(N__55348),
            .I(N__55345));
    Odrv4 I__10248 (
            .O(N__55345),
            .I(\spi0.n19_adj_1139 ));
    InMux I__10247 (
            .O(N__55342),
            .I(N__55338));
    InMux I__10246 (
            .O(N__55341),
            .I(N__55335));
    LocalMux I__10245 (
            .O(N__55338),
            .I(\spi0.multi_byte_counter_0 ));
    LocalMux I__10244 (
            .O(N__55335),
            .I(\spi0.multi_byte_counter_0 ));
    InMux I__10243 (
            .O(N__55330),
            .I(\spi0.n10653 ));
    InMux I__10242 (
            .O(N__55327),
            .I(N__55324));
    LocalMux I__10241 (
            .O(N__55324),
            .I(N__55320));
    InMux I__10240 (
            .O(N__55323),
            .I(N__55317));
    Odrv4 I__10239 (
            .O(N__55320),
            .I(\spi0.multi_byte_counter_2 ));
    LocalMux I__10238 (
            .O(N__55317),
            .I(\spi0.multi_byte_counter_2 ));
    InMux I__10237 (
            .O(N__55312),
            .I(\spi0.n10654 ));
    InMux I__10236 (
            .O(N__55309),
            .I(\spi0.n10655 ));
    InMux I__10235 (
            .O(N__55306),
            .I(N__55302));
    InMux I__10234 (
            .O(N__55305),
            .I(N__55299));
    LocalMux I__10233 (
            .O(N__55302),
            .I(\spi0.multi_byte_counter_4 ));
    LocalMux I__10232 (
            .O(N__55299),
            .I(\spi0.multi_byte_counter_4 ));
    InMux I__10231 (
            .O(N__55294),
            .I(\spi0.n10656 ));
    InMux I__10230 (
            .O(N__55291),
            .I(\spi0.n10657 ));
    InMux I__10229 (
            .O(N__55288),
            .I(N__55285));
    LocalMux I__10228 (
            .O(N__55285),
            .I(N__55281));
    InMux I__10227 (
            .O(N__55284),
            .I(N__55278));
    Odrv4 I__10226 (
            .O(N__55281),
            .I(\spi0.multi_byte_counter_6 ));
    LocalMux I__10225 (
            .O(N__55278),
            .I(\spi0.multi_byte_counter_6 ));
    InMux I__10224 (
            .O(N__55273),
            .I(\spi0.n10658 ));
    CascadeMux I__10223 (
            .O(N__55270),
            .I(N__55266));
    CascadeMux I__10222 (
            .O(N__55269),
            .I(N__55262));
    InMux I__10221 (
            .O(N__55266),
            .I(N__55244));
    InMux I__10220 (
            .O(N__55265),
            .I(N__55244));
    InMux I__10219 (
            .O(N__55262),
            .I(N__55244));
    InMux I__10218 (
            .O(N__55261),
            .I(N__55239));
    InMux I__10217 (
            .O(N__55260),
            .I(N__55239));
    CascadeMux I__10216 (
            .O(N__55259),
            .I(N__55236));
    InMux I__10215 (
            .O(N__55258),
            .I(N__55219));
    InMux I__10214 (
            .O(N__55257),
            .I(N__55219));
    InMux I__10213 (
            .O(N__55256),
            .I(N__55219));
    InMux I__10212 (
            .O(N__55255),
            .I(N__55219));
    InMux I__10211 (
            .O(N__55254),
            .I(N__55219));
    CascadeMux I__10210 (
            .O(N__55253),
            .I(N__55215));
    CascadeMux I__10209 (
            .O(N__55252),
            .I(N__55211));
    InMux I__10208 (
            .O(N__55251),
            .I(N__55207));
    LocalMux I__10207 (
            .O(N__55244),
            .I(N__55204));
    LocalMux I__10206 (
            .O(N__55239),
            .I(N__55201));
    InMux I__10205 (
            .O(N__55236),
            .I(N__55192));
    InMux I__10204 (
            .O(N__55235),
            .I(N__55192));
    InMux I__10203 (
            .O(N__55234),
            .I(N__55192));
    InMux I__10202 (
            .O(N__55233),
            .I(N__55192));
    CascadeMux I__10201 (
            .O(N__55232),
            .I(N__55189));
    CascadeMux I__10200 (
            .O(N__55231),
            .I(N__55186));
    CascadeMux I__10199 (
            .O(N__55230),
            .I(N__55180));
    LocalMux I__10198 (
            .O(N__55219),
            .I(N__55173));
    InMux I__10197 (
            .O(N__55218),
            .I(N__55170));
    InMux I__10196 (
            .O(N__55215),
            .I(N__55161));
    InMux I__10195 (
            .O(N__55214),
            .I(N__55161));
    InMux I__10194 (
            .O(N__55211),
            .I(N__55161));
    InMux I__10193 (
            .O(N__55210),
            .I(N__55161));
    LocalMux I__10192 (
            .O(N__55207),
            .I(N__55152));
    Span4Mux_h I__10191 (
            .O(N__55204),
            .I(N__55152));
    Span4Mux_h I__10190 (
            .O(N__55201),
            .I(N__55152));
    LocalMux I__10189 (
            .O(N__55192),
            .I(N__55152));
    InMux I__10188 (
            .O(N__55189),
            .I(N__55145));
    InMux I__10187 (
            .O(N__55186),
            .I(N__55145));
    InMux I__10186 (
            .O(N__55185),
            .I(N__55145));
    InMux I__10185 (
            .O(N__55184),
            .I(N__55138));
    InMux I__10184 (
            .O(N__55183),
            .I(N__55138));
    InMux I__10183 (
            .O(N__55180),
            .I(N__55138));
    InMux I__10182 (
            .O(N__55179),
            .I(N__55129));
    InMux I__10181 (
            .O(N__55178),
            .I(N__55129));
    InMux I__10180 (
            .O(N__55177),
            .I(N__55129));
    InMux I__10179 (
            .O(N__55176),
            .I(N__55129));
    Odrv4 I__10178 (
            .O(N__55173),
            .I(\spi0.state_0 ));
    LocalMux I__10177 (
            .O(N__55170),
            .I(\spi0.state_0 ));
    LocalMux I__10176 (
            .O(N__55161),
            .I(\spi0.state_0 ));
    Odrv4 I__10175 (
            .O(N__55152),
            .I(\spi0.state_0 ));
    LocalMux I__10174 (
            .O(N__55145),
            .I(\spi0.state_0 ));
    LocalMux I__10173 (
            .O(N__55138),
            .I(\spi0.state_0 ));
    LocalMux I__10172 (
            .O(N__55129),
            .I(\spi0.state_0 ));
    CascadeMux I__10171 (
            .O(N__55114),
            .I(\spi0.n12576_cascade_ ));
    InMux I__10170 (
            .O(N__55111),
            .I(N__55108));
    LocalMux I__10169 (
            .O(N__55108),
            .I(\spi0.n37 ));
    InMux I__10168 (
            .O(N__55105),
            .I(N__55102));
    LocalMux I__10167 (
            .O(N__55102),
            .I(N__55099));
    Odrv4 I__10166 (
            .O(N__55099),
            .I(\spi0.n2768 ));
    InMux I__10165 (
            .O(N__55096),
            .I(N__55093));
    LocalMux I__10164 (
            .O(N__55093),
            .I(\spi0.n6 ));
    CascadeMux I__10163 (
            .O(N__55090),
            .I(\spi0.n2768_cascade_ ));
    InMux I__10162 (
            .O(N__55087),
            .I(N__55084));
    LocalMux I__10161 (
            .O(N__55084),
            .I(\spi0.n4260 ));
    CEMux I__10160 (
            .O(N__55081),
            .I(N__55078));
    LocalMux I__10159 (
            .O(N__55078),
            .I(\spi0.n14414 ));
    InMux I__10158 (
            .O(N__55075),
            .I(N__55052));
    InMux I__10157 (
            .O(N__55074),
            .I(N__55052));
    InMux I__10156 (
            .O(N__55073),
            .I(N__55052));
    InMux I__10155 (
            .O(N__55072),
            .I(N__55038));
    InMux I__10154 (
            .O(N__55071),
            .I(N__55038));
    InMux I__10153 (
            .O(N__55070),
            .I(N__55038));
    InMux I__10152 (
            .O(N__55069),
            .I(N__55038));
    InMux I__10151 (
            .O(N__55068),
            .I(N__55029));
    InMux I__10150 (
            .O(N__55067),
            .I(N__55029));
    InMux I__10149 (
            .O(N__55066),
            .I(N__55029));
    InMux I__10148 (
            .O(N__55065),
            .I(N__55029));
    InMux I__10147 (
            .O(N__55064),
            .I(N__55016));
    InMux I__10146 (
            .O(N__55063),
            .I(N__55016));
    InMux I__10145 (
            .O(N__55062),
            .I(N__55016));
    InMux I__10144 (
            .O(N__55061),
            .I(N__55016));
    InMux I__10143 (
            .O(N__55060),
            .I(N__55016));
    InMux I__10142 (
            .O(N__55059),
            .I(N__55016));
    LocalMux I__10141 (
            .O(N__55052),
            .I(N__55005));
    InMux I__10140 (
            .O(N__55051),
            .I(N__54998));
    InMux I__10139 (
            .O(N__55050),
            .I(N__54998));
    InMux I__10138 (
            .O(N__55049),
            .I(N__54998));
    InMux I__10137 (
            .O(N__55048),
            .I(N__54993));
    InMux I__10136 (
            .O(N__55047),
            .I(N__54993));
    LocalMux I__10135 (
            .O(N__55038),
            .I(N__54986));
    LocalMux I__10134 (
            .O(N__55029),
            .I(N__54986));
    LocalMux I__10133 (
            .O(N__55016),
            .I(N__54986));
    InMux I__10132 (
            .O(N__55015),
            .I(N__54977));
    InMux I__10131 (
            .O(N__55014),
            .I(N__54977));
    InMux I__10130 (
            .O(N__55013),
            .I(N__54977));
    InMux I__10129 (
            .O(N__55012),
            .I(N__54977));
    InMux I__10128 (
            .O(N__55011),
            .I(N__54968));
    InMux I__10127 (
            .O(N__55010),
            .I(N__54968));
    InMux I__10126 (
            .O(N__55009),
            .I(N__54968));
    InMux I__10125 (
            .O(N__55008),
            .I(N__54968));
    Odrv4 I__10124 (
            .O(N__55005),
            .I(\spi0.state_2 ));
    LocalMux I__10123 (
            .O(N__54998),
            .I(\spi0.state_2 ));
    LocalMux I__10122 (
            .O(N__54993),
            .I(\spi0.state_2 ));
    Odrv4 I__10121 (
            .O(N__54986),
            .I(\spi0.state_2 ));
    LocalMux I__10120 (
            .O(N__54977),
            .I(\spi0.state_2 ));
    LocalMux I__10119 (
            .O(N__54968),
            .I(\spi0.state_2 ));
    CascadeMux I__10118 (
            .O(N__54955),
            .I(N__54952));
    InMux I__10117 (
            .O(N__54952),
            .I(N__54946));
    CascadeMux I__10116 (
            .O(N__54951),
            .I(N__54942));
    InMux I__10115 (
            .O(N__54950),
            .I(N__54937));
    InMux I__10114 (
            .O(N__54949),
            .I(N__54937));
    LocalMux I__10113 (
            .O(N__54946),
            .I(N__54934));
    InMux I__10112 (
            .O(N__54945),
            .I(N__54929));
    InMux I__10111 (
            .O(N__54942),
            .I(N__54929));
    LocalMux I__10110 (
            .O(N__54937),
            .I(N__54923));
    Span4Mux_v I__10109 (
            .O(N__54934),
            .I(N__54920));
    LocalMux I__10108 (
            .O(N__54929),
            .I(N__54917));
    InMux I__10107 (
            .O(N__54928),
            .I(N__54914));
    InMux I__10106 (
            .O(N__54927),
            .I(N__54909));
    InMux I__10105 (
            .O(N__54926),
            .I(N__54909));
    Odrv4 I__10104 (
            .O(N__54923),
            .I(\spi0.n19 ));
    Odrv4 I__10103 (
            .O(N__54920),
            .I(\spi0.n19 ));
    Odrv12 I__10102 (
            .O(N__54917),
            .I(\spi0.n19 ));
    LocalMux I__10101 (
            .O(N__54914),
            .I(\spi0.n19 ));
    LocalMux I__10100 (
            .O(N__54909),
            .I(\spi0.n19 ));
    InMux I__10099 (
            .O(N__54898),
            .I(N__54895));
    LocalMux I__10098 (
            .O(N__54895),
            .I(\spi0.n21 ));
    CascadeMux I__10097 (
            .O(N__54892),
            .I(\spi0.n10_cascade_ ));
    InMux I__10096 (
            .O(N__54889),
            .I(N__54886));
    LocalMux I__10095 (
            .O(N__54886),
            .I(N__54882));
    InMux I__10094 (
            .O(N__54885),
            .I(N__54879));
    Odrv4 I__10093 (
            .O(N__54882),
            .I(tx_addr_byte_3));
    LocalMux I__10092 (
            .O(N__54879),
            .I(tx_addr_byte_3));
    InMux I__10091 (
            .O(N__54874),
            .I(N__54871));
    LocalMux I__10090 (
            .O(N__54871),
            .I(N__54865));
    InMux I__10089 (
            .O(N__54870),
            .I(N__54862));
    InMux I__10088 (
            .O(N__54869),
            .I(N__54857));
    InMux I__10087 (
            .O(N__54868),
            .I(N__54857));
    Odrv4 I__10086 (
            .O(N__54865),
            .I(tx_data_byte_5));
    LocalMux I__10085 (
            .O(N__54862),
            .I(tx_data_byte_5));
    LocalMux I__10084 (
            .O(N__54857),
            .I(tx_data_byte_5));
    InMux I__10083 (
            .O(N__54850),
            .I(N__54847));
    LocalMux I__10082 (
            .O(N__54847),
            .I(N__54841));
    InMux I__10081 (
            .O(N__54846),
            .I(N__54838));
    InMux I__10080 (
            .O(N__54845),
            .I(N__54835));
    InMux I__10079 (
            .O(N__54844),
            .I(N__54832));
    Odrv4 I__10078 (
            .O(N__54841),
            .I(tx_data_byte_3));
    LocalMux I__10077 (
            .O(N__54838),
            .I(tx_data_byte_3));
    LocalMux I__10076 (
            .O(N__54835),
            .I(tx_data_byte_3));
    LocalMux I__10075 (
            .O(N__54832),
            .I(tx_data_byte_3));
    CascadeMux I__10074 (
            .O(N__54823),
            .I(n11412_cascade_));
    InMux I__10073 (
            .O(N__54820),
            .I(N__54817));
    LocalMux I__10072 (
            .O(N__54817),
            .I(N__54811));
    InMux I__10071 (
            .O(N__54816),
            .I(N__54808));
    InMux I__10070 (
            .O(N__54815),
            .I(N__54803));
    InMux I__10069 (
            .O(N__54814),
            .I(N__54803));
    Odrv4 I__10068 (
            .O(N__54811),
            .I(tx_data_byte_6));
    LocalMux I__10067 (
            .O(N__54808),
            .I(tx_data_byte_6));
    LocalMux I__10066 (
            .O(N__54803),
            .I(tx_data_byte_6));
    CascadeMux I__10065 (
            .O(N__54796),
            .I(n11471_cascade_));
    InMux I__10064 (
            .O(N__54793),
            .I(N__54787));
    InMux I__10063 (
            .O(N__54792),
            .I(N__54784));
    InMux I__10062 (
            .O(N__54791),
            .I(N__54781));
    InMux I__10061 (
            .O(N__54790),
            .I(N__54778));
    LocalMux I__10060 (
            .O(N__54787),
            .I(tx_data_byte_1));
    LocalMux I__10059 (
            .O(N__54784),
            .I(tx_data_byte_1));
    LocalMux I__10058 (
            .O(N__54781),
            .I(tx_data_byte_1));
    LocalMux I__10057 (
            .O(N__54778),
            .I(tx_data_byte_1));
    InMux I__10056 (
            .O(N__54769),
            .I(N__54766));
    LocalMux I__10055 (
            .O(N__54766),
            .I(\spi0.n12605 ));
    InMux I__10054 (
            .O(N__54763),
            .I(N__54760));
    LocalMux I__10053 (
            .O(N__54760),
            .I(\spi0.n10090 ));
    CascadeMux I__10052 (
            .O(N__54757),
            .I(N__54753));
    CascadeMux I__10051 (
            .O(N__54756),
            .I(N__54749));
    InMux I__10050 (
            .O(N__54753),
            .I(N__54742));
    InMux I__10049 (
            .O(N__54752),
            .I(N__54742));
    InMux I__10048 (
            .O(N__54749),
            .I(N__54742));
    LocalMux I__10047 (
            .O(N__54742),
            .I(multi_byte_spi_trans_flag_r));
    InMux I__10046 (
            .O(N__54739),
            .I(N__54736));
    LocalMux I__10045 (
            .O(N__54736),
            .I(N__54733));
    Odrv4 I__10044 (
            .O(N__54733),
            .I(\spi0.n3 ));
    InMux I__10043 (
            .O(N__54730),
            .I(N__54726));
    InMux I__10042 (
            .O(N__54729),
            .I(N__54723));
    LocalMux I__10041 (
            .O(N__54726),
            .I(tx_addr_byte_1));
    LocalMux I__10040 (
            .O(N__54723),
            .I(tx_addr_byte_1));
    CascadeMux I__10039 (
            .O(N__54718),
            .I(N__54714));
    InMux I__10038 (
            .O(N__54717),
            .I(N__54709));
    InMux I__10037 (
            .O(N__54714),
            .I(N__54709));
    LocalMux I__10036 (
            .O(N__54709),
            .I(pc_data_rx_5));
    InMux I__10035 (
            .O(N__54706),
            .I(N__54702));
    InMux I__10034 (
            .O(N__54705),
            .I(N__54699));
    LocalMux I__10033 (
            .O(N__54702),
            .I(tx_addr_byte_6));
    LocalMux I__10032 (
            .O(N__54699),
            .I(tx_addr_byte_6));
    CascadeMux I__10031 (
            .O(N__54694),
            .I(n10847_cascade_));
    InMux I__10030 (
            .O(N__54691),
            .I(N__54685));
    InMux I__10029 (
            .O(N__54690),
            .I(N__54685));
    LocalMux I__10028 (
            .O(N__54685),
            .I(pc_data_rx_0));
    InMux I__10027 (
            .O(N__54682),
            .I(N__54679));
    LocalMux I__10026 (
            .O(N__54679),
            .I(N__54675));
    InMux I__10025 (
            .O(N__54678),
            .I(N__54672));
    Odrv4 I__10024 (
            .O(N__54675),
            .I(tx_addr_byte_0));
    LocalMux I__10023 (
            .O(N__54672),
            .I(tx_addr_byte_0));
    InMux I__10022 (
            .O(N__54667),
            .I(N__54664));
    LocalMux I__10021 (
            .O(N__54664),
            .I(\spi0.tx_shift_reg_10 ));
    InMux I__10020 (
            .O(N__54661),
            .I(N__54658));
    LocalMux I__10019 (
            .O(N__54658),
            .I(\spi0.tx_shift_reg_11 ));
    InMux I__10018 (
            .O(N__54655),
            .I(N__54652));
    LocalMux I__10017 (
            .O(N__54652),
            .I(N__54649));
    Odrv4 I__10016 (
            .O(N__54649),
            .I(\spi0.tx_shift_reg_12 ));
    InMux I__10015 (
            .O(N__54646),
            .I(N__54643));
    LocalMux I__10014 (
            .O(N__54643),
            .I(\spi0.tx_shift_reg_13 ));
    InMux I__10013 (
            .O(N__54640),
            .I(N__54637));
    LocalMux I__10012 (
            .O(N__54637),
            .I(\spi0.tx_shift_reg_8 ));
    InMux I__10011 (
            .O(N__54634),
            .I(N__54631));
    LocalMux I__10010 (
            .O(N__54631),
            .I(\spi0.tx_shift_reg_6 ));
    InMux I__10009 (
            .O(N__54628),
            .I(N__54625));
    LocalMux I__10008 (
            .O(N__54625),
            .I(\spi0.tx_shift_reg_7 ));
    InMux I__10007 (
            .O(N__54622),
            .I(N__54618));
    InMux I__10006 (
            .O(N__54621),
            .I(N__54615));
    LocalMux I__10005 (
            .O(N__54618),
            .I(tx_addr_byte_5));
    LocalMux I__10004 (
            .O(N__54615),
            .I(tx_addr_byte_5));
    InMux I__10003 (
            .O(N__54610),
            .I(\usb3_if_inst.n10663 ));
    InMux I__10002 (
            .O(N__54607),
            .I(\usb3_if_inst.n10664 ));
    InMux I__10001 (
            .O(N__54604),
            .I(\usb3_if_inst.n10665 ));
    InMux I__10000 (
            .O(N__54601),
            .I(N__54598));
    LocalMux I__9999 (
            .O(N__54598),
            .I(N__54594));
    InMux I__9998 (
            .O(N__54597),
            .I(N__54591));
    Span4Mux_v I__9997 (
            .O(N__54594),
            .I(N__54588));
    LocalMux I__9996 (
            .O(N__54591),
            .I(\usb3_if_inst.num_lines_clocked_out_7 ));
    Odrv4 I__9995 (
            .O(N__54588),
            .I(\usb3_if_inst.num_lines_clocked_out_7 ));
    InMux I__9994 (
            .O(N__54583),
            .I(\usb3_if_inst.n10666 ));
    InMux I__9993 (
            .O(N__54580),
            .I(bfn_14_14_0_));
    InMux I__9992 (
            .O(N__54577),
            .I(N__54573));
    CascadeMux I__9991 (
            .O(N__54576),
            .I(N__54570));
    LocalMux I__9990 (
            .O(N__54573),
            .I(N__54567));
    InMux I__9989 (
            .O(N__54570),
            .I(N__54564));
    Span4Mux_h I__9988 (
            .O(N__54567),
            .I(N__54561));
    LocalMux I__9987 (
            .O(N__54564),
            .I(\usb3_if_inst.num_lines_clocked_out_9 ));
    Odrv4 I__9986 (
            .O(N__54561),
            .I(\usb3_if_inst.num_lines_clocked_out_9 ));
    InMux I__9985 (
            .O(N__54556),
            .I(\usb3_if_inst.n10668 ));
    InMux I__9984 (
            .O(N__54553),
            .I(\usb3_if_inst.n10669 ));
    InMux I__9983 (
            .O(N__54550),
            .I(N__54547));
    LocalMux I__9982 (
            .O(N__54547),
            .I(\spi0.tx_shift_reg_9 ));
    CascadeMux I__9981 (
            .O(N__54544),
            .I(\usb3_if_inst.n4403_cascade_ ));
    InMux I__9980 (
            .O(N__54541),
            .I(N__54538));
    LocalMux I__9979 (
            .O(N__54538),
            .I(N__54535));
    Span4Mux_h I__9978 (
            .O(N__54535),
            .I(N__54532));
    Odrv4 I__9977 (
            .O(N__54532),
            .I(\usb3_if_inst.n6904 ));
    InMux I__9976 (
            .O(N__54529),
            .I(N__54526));
    LocalMux I__9975 (
            .O(N__54526),
            .I(\usb3_if_inst.n135 ));
    CascadeMux I__9974 (
            .O(N__54523),
            .I(N__54520));
    InMux I__9973 (
            .O(N__54520),
            .I(N__54517));
    LocalMux I__9972 (
            .O(N__54517),
            .I(\usb3_if_inst.n3686 ));
    CascadeMux I__9971 (
            .O(N__54514),
            .I(N__54510));
    CascadeMux I__9970 (
            .O(N__54513),
            .I(N__54507));
    InMux I__9969 (
            .O(N__54510),
            .I(N__54504));
    InMux I__9968 (
            .O(N__54507),
            .I(N__54501));
    LocalMux I__9967 (
            .O(N__54504),
            .I(\usb3_if_inst.state_timeout_counter_3 ));
    LocalMux I__9966 (
            .O(N__54501),
            .I(\usb3_if_inst.state_timeout_counter_3 ));
    CascadeMux I__9965 (
            .O(N__54496),
            .I(\usb3_if_inst.n12582_cascade_ ));
    CEMux I__9964 (
            .O(N__54493),
            .I(N__54489));
    CEMux I__9963 (
            .O(N__54492),
            .I(N__54486));
    LocalMux I__9962 (
            .O(N__54489),
            .I(N__54483));
    LocalMux I__9961 (
            .O(N__54486),
            .I(N__54479));
    Span4Mux_h I__9960 (
            .O(N__54483),
            .I(N__54476));
    CEMux I__9959 (
            .O(N__54482),
            .I(N__54473));
    Span4Mux_h I__9958 (
            .O(N__54479),
            .I(N__54470));
    Span4Mux_h I__9957 (
            .O(N__54476),
            .I(N__54467));
    LocalMux I__9956 (
            .O(N__54473),
            .I(N__54462));
    Span4Mux_h I__9955 (
            .O(N__54470),
            .I(N__54462));
    Odrv4 I__9954 (
            .O(N__54467),
            .I(\usb3_if_inst.n4061 ));
    Odrv4 I__9953 (
            .O(N__54462),
            .I(\usb3_if_inst.n4061 ));
    CascadeMux I__9952 (
            .O(N__54457),
            .I(N__54454));
    InMux I__9951 (
            .O(N__54454),
            .I(N__54451));
    LocalMux I__9950 (
            .O(N__54451),
            .I(\usb3_if_inst.empty_o_N_599 ));
    CascadeMux I__9949 (
            .O(N__54448),
            .I(N__54445));
    InMux I__9948 (
            .O(N__54445),
            .I(N__54442));
    LocalMux I__9947 (
            .O(N__54442),
            .I(N__54438));
    InMux I__9946 (
            .O(N__54441),
            .I(N__54435));
    Span12Mux_v I__9945 (
            .O(N__54438),
            .I(N__54432));
    LocalMux I__9944 (
            .O(N__54435),
            .I(\usb3_if_inst.num_lines_clocked_out_0 ));
    Odrv12 I__9943 (
            .O(N__54432),
            .I(\usb3_if_inst.num_lines_clocked_out_0 ));
    InMux I__9942 (
            .O(N__54427),
            .I(bfn_14_13_0_));
    InMux I__9941 (
            .O(N__54424),
            .I(\usb3_if_inst.n10660 ));
    InMux I__9940 (
            .O(N__54421),
            .I(N__54417));
    CascadeMux I__9939 (
            .O(N__54420),
            .I(N__54414));
    LocalMux I__9938 (
            .O(N__54417),
            .I(N__54411));
    InMux I__9937 (
            .O(N__54414),
            .I(N__54408));
    Span4Mux_v I__9936 (
            .O(N__54411),
            .I(N__54405));
    LocalMux I__9935 (
            .O(N__54408),
            .I(\usb3_if_inst.num_lines_clocked_out_2 ));
    Odrv4 I__9934 (
            .O(N__54405),
            .I(\usb3_if_inst.num_lines_clocked_out_2 ));
    InMux I__9933 (
            .O(N__54400),
            .I(\usb3_if_inst.n10661 ));
    InMux I__9932 (
            .O(N__54397),
            .I(\usb3_if_inst.n10662 ));
    InMux I__9931 (
            .O(N__54394),
            .I(N__54388));
    InMux I__9930 (
            .O(N__54393),
            .I(N__54388));
    LocalMux I__9929 (
            .O(N__54388),
            .I(REG_mem_18_4));
    InMux I__9928 (
            .O(N__54385),
            .I(N__54379));
    InMux I__9927 (
            .O(N__54384),
            .I(N__54379));
    LocalMux I__9926 (
            .O(N__54379),
            .I(REG_mem_19_4));
    CascadeMux I__9925 (
            .O(N__54376),
            .I(N__54372));
    InMux I__9924 (
            .O(N__54375),
            .I(N__54367));
    InMux I__9923 (
            .O(N__54372),
            .I(N__54367));
    LocalMux I__9922 (
            .O(N__54367),
            .I(REG_mem_16_4));
    InMux I__9921 (
            .O(N__54364),
            .I(N__54358));
    InMux I__9920 (
            .O(N__54363),
            .I(N__54358));
    LocalMux I__9919 (
            .O(N__54358),
            .I(REG_mem_17_4));
    CascadeMux I__9918 (
            .O(N__54355),
            .I(\usb3_if_inst.n3686_cascade_ ));
    InMux I__9917 (
            .O(N__54352),
            .I(N__54345));
    InMux I__9916 (
            .O(N__54351),
            .I(N__54340));
    InMux I__9915 (
            .O(N__54350),
            .I(N__54340));
    InMux I__9914 (
            .O(N__54349),
            .I(N__54335));
    InMux I__9913 (
            .O(N__54348),
            .I(N__54335));
    LocalMux I__9912 (
            .O(N__54345),
            .I(\usb3_if_inst.state_timeout_counter_1 ));
    LocalMux I__9911 (
            .O(N__54340),
            .I(\usb3_if_inst.state_timeout_counter_1 ));
    LocalMux I__9910 (
            .O(N__54335),
            .I(\usb3_if_inst.state_timeout_counter_1 ));
    InMux I__9909 (
            .O(N__54328),
            .I(N__54319));
    InMux I__9908 (
            .O(N__54327),
            .I(N__54314));
    InMux I__9907 (
            .O(N__54326),
            .I(N__54314));
    InMux I__9906 (
            .O(N__54325),
            .I(N__54305));
    InMux I__9905 (
            .O(N__54324),
            .I(N__54305));
    InMux I__9904 (
            .O(N__54323),
            .I(N__54305));
    InMux I__9903 (
            .O(N__54322),
            .I(N__54305));
    LocalMux I__9902 (
            .O(N__54319),
            .I(\usb3_if_inst.state_timeout_counter_0 ));
    LocalMux I__9901 (
            .O(N__54314),
            .I(\usb3_if_inst.state_timeout_counter_0 ));
    LocalMux I__9900 (
            .O(N__54305),
            .I(\usb3_if_inst.state_timeout_counter_0 ));
    CascadeMux I__9899 (
            .O(N__54298),
            .I(\usb3_if_inst.n4_cascade_ ));
    InMux I__9898 (
            .O(N__54295),
            .I(N__54292));
    LocalMux I__9897 (
            .O(N__54292),
            .I(N__54288));
    CascadeMux I__9896 (
            .O(N__54291),
            .I(N__54285));
    Span4Mux_v I__9895 (
            .O(N__54288),
            .I(N__54282));
    InMux I__9894 (
            .O(N__54285),
            .I(N__54279));
    Odrv4 I__9893 (
            .O(N__54282),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_7 ));
    LocalMux I__9892 (
            .O(N__54279),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_7 ));
    InMux I__9891 (
            .O(N__54274),
            .I(N__54271));
    LocalMux I__9890 (
            .O(N__54271),
            .I(N__54267));
    InMux I__9889 (
            .O(N__54270),
            .I(N__54264));
    Odrv4 I__9888 (
            .O(N__54267),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_7 ));
    LocalMux I__9887 (
            .O(N__54264),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_7 ));
    CascadeMux I__9886 (
            .O(N__54259),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14090_cascade_ ));
    InMux I__9885 (
            .O(N__54256),
            .I(N__54253));
    LocalMux I__9884 (
            .O(N__54253),
            .I(N__54249));
    CascadeMux I__9883 (
            .O(N__54252),
            .I(N__54246));
    Span4Mux_v I__9882 (
            .O(N__54249),
            .I(N__54243));
    InMux I__9881 (
            .O(N__54246),
            .I(N__54240));
    Odrv4 I__9880 (
            .O(N__54243),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_7 ));
    LocalMux I__9879 (
            .O(N__54240),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_7 ));
    InMux I__9878 (
            .O(N__54235),
            .I(N__54232));
    LocalMux I__9877 (
            .O(N__54232),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12111 ));
    CascadeMux I__9876 (
            .O(N__54229),
            .I(N__54225));
    InMux I__9875 (
            .O(N__54228),
            .I(N__54220));
    InMux I__9874 (
            .O(N__54225),
            .I(N__54220));
    LocalMux I__9873 (
            .O(N__54220),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_7 ));
    CascadeMux I__9872 (
            .O(N__54217),
            .I(N__54214));
    InMux I__9871 (
            .O(N__54214),
            .I(N__54208));
    InMux I__9870 (
            .O(N__54213),
            .I(N__54208));
    LocalMux I__9869 (
            .O(N__54208),
            .I(REG_mem_23_7));
    CascadeMux I__9868 (
            .O(N__54205),
            .I(N__54201));
    InMux I__9867 (
            .O(N__54204),
            .I(N__54198));
    InMux I__9866 (
            .O(N__54201),
            .I(N__54195));
    LocalMux I__9865 (
            .O(N__54198),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_7 ));
    LocalMux I__9864 (
            .O(N__54195),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_7 ));
    CascadeMux I__9863 (
            .O(N__54190),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13964_cascade_ ));
    InMux I__9862 (
            .O(N__54187),
            .I(N__54183));
    InMux I__9861 (
            .O(N__54186),
            .I(N__54180));
    LocalMux I__9860 (
            .O(N__54183),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_7 ));
    LocalMux I__9859 (
            .O(N__54180),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_7 ));
    CascadeMux I__9858 (
            .O(N__54175),
            .I(N__54172));
    InMux I__9857 (
            .O(N__54172),
            .I(N__54169));
    LocalMux I__9856 (
            .O(N__54169),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12150 ));
    InMux I__9855 (
            .O(N__54166),
            .I(N__54163));
    LocalMux I__9854 (
            .O(N__54163),
            .I(N__54160));
    Sp12to4 I__9853 (
            .O(N__54160),
            .I(N__54157));
    Span12Mux_h I__9852 (
            .O(N__54157),
            .I(N__54153));
    InMux I__9851 (
            .O(N__54156),
            .I(N__54150));
    Odrv12 I__9850 (
            .O(N__54153),
            .I(REG_mem_31_15));
    LocalMux I__9849 (
            .O(N__54150),
            .I(REG_mem_31_15));
    CascadeMux I__9848 (
            .O(N__54145),
            .I(N__54142));
    InMux I__9847 (
            .O(N__54142),
            .I(N__54139));
    LocalMux I__9846 (
            .O(N__54139),
            .I(N__54136));
    Span4Mux_v I__9845 (
            .O(N__54136),
            .I(N__54133));
    Span4Mux_h I__9844 (
            .O(N__54133),
            .I(N__54130));
    Odrv4 I__9843 (
            .O(N__54130),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11996 ));
    InMux I__9842 (
            .O(N__54127),
            .I(N__54121));
    InMux I__9841 (
            .O(N__54126),
            .I(N__54121));
    LocalMux I__9840 (
            .O(N__54121),
            .I(REG_mem_38_15));
    InMux I__9839 (
            .O(N__54118),
            .I(N__54112));
    InMux I__9838 (
            .O(N__54117),
            .I(N__54112));
    LocalMux I__9837 (
            .O(N__54112),
            .I(REG_mem_39_15));
    InMux I__9836 (
            .O(N__54109),
            .I(N__54105));
    InMux I__9835 (
            .O(N__54108),
            .I(N__54102));
    LocalMux I__9834 (
            .O(N__54105),
            .I(N__54099));
    LocalMux I__9833 (
            .O(N__54102),
            .I(N__54095));
    Span4Mux_v I__9832 (
            .O(N__54099),
            .I(N__54090));
    InMux I__9831 (
            .O(N__54098),
            .I(N__54087));
    Span4Mux_v I__9830 (
            .O(N__54095),
            .I(N__54083));
    InMux I__9829 (
            .O(N__54094),
            .I(N__54077));
    InMux I__9828 (
            .O(N__54093),
            .I(N__54074));
    Span4Mux_h I__9827 (
            .O(N__54090),
            .I(N__54069));
    LocalMux I__9826 (
            .O(N__54087),
            .I(N__54066));
    InMux I__9825 (
            .O(N__54086),
            .I(N__54060));
    Span4Mux_h I__9824 (
            .O(N__54083),
            .I(N__54057));
    InMux I__9823 (
            .O(N__54082),
            .I(N__54054));
    InMux I__9822 (
            .O(N__54081),
            .I(N__54051));
    InMux I__9821 (
            .O(N__54080),
            .I(N__54048));
    LocalMux I__9820 (
            .O(N__54077),
            .I(N__54045));
    LocalMux I__9819 (
            .O(N__54074),
            .I(N__54042));
    InMux I__9818 (
            .O(N__54073),
            .I(N__54038));
    InMux I__9817 (
            .O(N__54072),
            .I(N__54035));
    Span4Mux_h I__9816 (
            .O(N__54069),
            .I(N__54030));
    Span4Mux_h I__9815 (
            .O(N__54066),
            .I(N__54030));
    InMux I__9814 (
            .O(N__54065),
            .I(N__54026));
    InMux I__9813 (
            .O(N__54064),
            .I(N__54021));
    InMux I__9812 (
            .O(N__54063),
            .I(N__54021));
    LocalMux I__9811 (
            .O(N__54060),
            .I(N__54018));
    Span4Mux_h I__9810 (
            .O(N__54057),
            .I(N__54015));
    LocalMux I__9809 (
            .O(N__54054),
            .I(N__54012));
    LocalMux I__9808 (
            .O(N__54051),
            .I(N__54007));
    LocalMux I__9807 (
            .O(N__54048),
            .I(N__54007));
    Span4Mux_h I__9806 (
            .O(N__54045),
            .I(N__54004));
    Span4Mux_h I__9805 (
            .O(N__54042),
            .I(N__54001));
    InMux I__9804 (
            .O(N__54041),
            .I(N__53998));
    LocalMux I__9803 (
            .O(N__54038),
            .I(N__53995));
    LocalMux I__9802 (
            .O(N__54035),
            .I(N__53990));
    Span4Mux_h I__9801 (
            .O(N__54030),
            .I(N__53990));
    InMux I__9800 (
            .O(N__54029),
            .I(N__53987));
    LocalMux I__9799 (
            .O(N__54026),
            .I(N__53984));
    LocalMux I__9798 (
            .O(N__54021),
            .I(N__53979));
    Span12Mux_h I__9797 (
            .O(N__54018),
            .I(N__53979));
    Span4Mux_h I__9796 (
            .O(N__54015),
            .I(N__53976));
    Span4Mux_v I__9795 (
            .O(N__54012),
            .I(N__53973));
    Span4Mux_h I__9794 (
            .O(N__54007),
            .I(N__53966));
    Span4Mux_h I__9793 (
            .O(N__54004),
            .I(N__53966));
    Span4Mux_v I__9792 (
            .O(N__54001),
            .I(N__53966));
    LocalMux I__9791 (
            .O(N__53998),
            .I(N__53959));
    Span4Mux_h I__9790 (
            .O(N__53995),
            .I(N__53959));
    Span4Mux_v I__9789 (
            .O(N__53990),
            .I(N__53959));
    LocalMux I__9788 (
            .O(N__53987),
            .I(n29));
    Odrv12 I__9787 (
            .O(N__53984),
            .I(n29));
    Odrv12 I__9786 (
            .O(N__53979),
            .I(n29));
    Odrv4 I__9785 (
            .O(N__53976),
            .I(n29));
    Odrv4 I__9784 (
            .O(N__53973),
            .I(n29));
    Odrv4 I__9783 (
            .O(N__53966),
            .I(n29));
    Odrv4 I__9782 (
            .O(N__53959),
            .I(n29));
    InMux I__9781 (
            .O(N__53944),
            .I(N__53940));
    InMux I__9780 (
            .O(N__53943),
            .I(N__53937));
    LocalMux I__9779 (
            .O(N__53940),
            .I(REG_mem_13_8));
    LocalMux I__9778 (
            .O(N__53937),
            .I(REG_mem_13_8));
    CascadeMux I__9777 (
            .O(N__53932),
            .I(N__53929));
    InMux I__9776 (
            .O(N__53929),
            .I(N__53926));
    LocalMux I__9775 (
            .O(N__53926),
            .I(N__53923));
    Span4Mux_v I__9774 (
            .O(N__53923),
            .I(N__53919));
    InMux I__9773 (
            .O(N__53922),
            .I(N__53916));
    Odrv4 I__9772 (
            .O(N__53919),
            .I(REG_mem_4_5));
    LocalMux I__9771 (
            .O(N__53916),
            .I(REG_mem_4_5));
    InMux I__9770 (
            .O(N__53911),
            .I(N__53908));
    LocalMux I__9769 (
            .O(N__53908),
            .I(N__53904));
    InMux I__9768 (
            .O(N__53907),
            .I(N__53901));
    Odrv4 I__9767 (
            .O(N__53904),
            .I(REG_mem_12_8));
    LocalMux I__9766 (
            .O(N__53901),
            .I(REG_mem_12_8));
    InMux I__9765 (
            .O(N__53896),
            .I(N__53893));
    LocalMux I__9764 (
            .O(N__53893),
            .I(N__53890));
    Span4Mux_v I__9763 (
            .O(N__53890),
            .I(N__53886));
    CascadeMux I__9762 (
            .O(N__53889),
            .I(N__53883));
    Span4Mux_v I__9761 (
            .O(N__53886),
            .I(N__53880));
    InMux I__9760 (
            .O(N__53883),
            .I(N__53877));
    Odrv4 I__9759 (
            .O(N__53880),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_1 ));
    LocalMux I__9758 (
            .O(N__53877),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_1 ));
    InMux I__9757 (
            .O(N__53872),
            .I(N__53869));
    LocalMux I__9756 (
            .O(N__53869),
            .I(N__53866));
    Span4Mux_v I__9755 (
            .O(N__53866),
            .I(N__53862));
    InMux I__9754 (
            .O(N__53865),
            .I(N__53859));
    Odrv4 I__9753 (
            .O(N__53862),
            .I(REG_mem_41_1));
    LocalMux I__9752 (
            .O(N__53859),
            .I(REG_mem_41_1));
    CascadeMux I__9751 (
            .O(N__53854),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14192_cascade_ ));
    InMux I__9750 (
            .O(N__53851),
            .I(N__53845));
    InMux I__9749 (
            .O(N__53850),
            .I(N__53845));
    LocalMux I__9748 (
            .O(N__53845),
            .I(REG_mem_14_8));
    InMux I__9747 (
            .O(N__53842),
            .I(N__53839));
    LocalMux I__9746 (
            .O(N__53839),
            .I(N__53835));
    InMux I__9745 (
            .O(N__53838),
            .I(N__53832));
    Odrv4 I__9744 (
            .O(N__53835),
            .I(REG_mem_15_9));
    LocalMux I__9743 (
            .O(N__53832),
            .I(REG_mem_15_9));
    InMux I__9742 (
            .O(N__53827),
            .I(N__53824));
    LocalMux I__9741 (
            .O(N__53824),
            .I(N__53821));
    Span4Mux_v I__9740 (
            .O(N__53821),
            .I(N__53817));
    InMux I__9739 (
            .O(N__53820),
            .I(N__53814));
    Odrv4 I__9738 (
            .O(N__53817),
            .I(REG_mem_15_1));
    LocalMux I__9737 (
            .O(N__53814),
            .I(REG_mem_15_1));
    InMux I__9736 (
            .O(N__53809),
            .I(N__53806));
    LocalMux I__9735 (
            .O(N__53806),
            .I(N__53802));
    InMux I__9734 (
            .O(N__53805),
            .I(N__53799));
    Odrv12 I__9733 (
            .O(N__53802),
            .I(REG_mem_39_0));
    LocalMux I__9732 (
            .O(N__53799),
            .I(REG_mem_39_0));
    InMux I__9731 (
            .O(N__53794),
            .I(N__53791));
    LocalMux I__9730 (
            .O(N__53791),
            .I(N__53787));
    CascadeMux I__9729 (
            .O(N__53790),
            .I(N__53784));
    Span4Mux_h I__9728 (
            .O(N__53787),
            .I(N__53781));
    InMux I__9727 (
            .O(N__53784),
            .I(N__53778));
    Odrv4 I__9726 (
            .O(N__53781),
            .I(REG_mem_37_0));
    LocalMux I__9725 (
            .O(N__53778),
            .I(REG_mem_37_0));
    CascadeMux I__9724 (
            .O(N__53773),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13016_cascade_ ));
    InMux I__9723 (
            .O(N__53770),
            .I(N__53767));
    LocalMux I__9722 (
            .O(N__53767),
            .I(N__53764));
    Span4Mux_v I__9721 (
            .O(N__53764),
            .I(N__53761));
    Span4Mux_v I__9720 (
            .O(N__53761),
            .I(N__53758));
    Span4Mux_h I__9719 (
            .O(N__53758),
            .I(N__53754));
    InMux I__9718 (
            .O(N__53757),
            .I(N__53751));
    Odrv4 I__9717 (
            .O(N__53754),
            .I(REG_mem_36_0));
    LocalMux I__9716 (
            .O(N__53751),
            .I(REG_mem_36_0));
    InMux I__9715 (
            .O(N__53746),
            .I(N__53743));
    LocalMux I__9714 (
            .O(N__53743),
            .I(N__53740));
    Span12Mux_h I__9713 (
            .O(N__53740),
            .I(N__53737));
    Odrv12 I__9712 (
            .O(N__53737),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13019 ));
    CascadeMux I__9711 (
            .O(N__53734),
            .I(N__53731));
    InMux I__9710 (
            .O(N__53731),
            .I(N__53725));
    InMux I__9709 (
            .O(N__53730),
            .I(N__53725));
    LocalMux I__9708 (
            .O(N__53725),
            .I(REG_mem_38_0));
    InMux I__9707 (
            .O(N__53722),
            .I(N__53719));
    LocalMux I__9706 (
            .O(N__53719),
            .I(N__53716));
    Span4Mux_h I__9705 (
            .O(N__53716),
            .I(N__53713));
    Span4Mux_v I__9704 (
            .O(N__53713),
            .I(N__53709));
    InMux I__9703 (
            .O(N__53712),
            .I(N__53706));
    Odrv4 I__9702 (
            .O(N__53709),
            .I(REG_mem_14_4));
    LocalMux I__9701 (
            .O(N__53706),
            .I(REG_mem_14_4));
    InMux I__9700 (
            .O(N__53701),
            .I(N__53697));
    InMux I__9699 (
            .O(N__53700),
            .I(N__53694));
    LocalMux I__9698 (
            .O(N__53697),
            .I(REG_mem_4_0));
    LocalMux I__9697 (
            .O(N__53694),
            .I(REG_mem_4_0));
    InMux I__9696 (
            .O(N__53689),
            .I(N__53686));
    LocalMux I__9695 (
            .O(N__53686),
            .I(N__53683));
    Span4Mux_v I__9694 (
            .O(N__53683),
            .I(N__53680));
    Sp12to4 I__9693 (
            .O(N__53680),
            .I(N__53676));
    InMux I__9692 (
            .O(N__53679),
            .I(N__53673));
    Odrv12 I__9691 (
            .O(N__53676),
            .I(REG_mem_46_0));
    LocalMux I__9690 (
            .O(N__53673),
            .I(REG_mem_46_0));
    InMux I__9689 (
            .O(N__53668),
            .I(N__53662));
    InMux I__9688 (
            .O(N__53667),
            .I(N__53662));
    LocalMux I__9687 (
            .O(N__53662),
            .I(REG_mem_38_6));
    CascadeMux I__9686 (
            .O(N__53659),
            .I(N__53656));
    InMux I__9685 (
            .O(N__53656),
            .I(N__53650));
    InMux I__9684 (
            .O(N__53655),
            .I(N__53650));
    LocalMux I__9683 (
            .O(N__53650),
            .I(REG_mem_39_6));
    InMux I__9682 (
            .O(N__53647),
            .I(N__53644));
    LocalMux I__9681 (
            .O(N__53644),
            .I(N__53641));
    Span4Mux_h I__9680 (
            .O(N__53641),
            .I(N__53637));
    InMux I__9679 (
            .O(N__53640),
            .I(N__53634));
    Odrv4 I__9678 (
            .O(N__53637),
            .I(REG_mem_37_5));
    LocalMux I__9677 (
            .O(N__53634),
            .I(REG_mem_37_5));
    CascadeMux I__9676 (
            .O(N__53629),
            .I(N__53626));
    InMux I__9675 (
            .O(N__53626),
            .I(N__53623));
    LocalMux I__9674 (
            .O(N__53623),
            .I(N__53620));
    Odrv4 I__9673 (
            .O(N__53620),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11671 ));
    InMux I__9672 (
            .O(N__53617),
            .I(N__53611));
    InMux I__9671 (
            .O(N__53616),
            .I(N__53611));
    LocalMux I__9670 (
            .O(N__53611),
            .I(REG_mem_12_1));
    InMux I__9669 (
            .O(N__53608),
            .I(N__53604));
    InMux I__9668 (
            .O(N__53607),
            .I(N__53601));
    LocalMux I__9667 (
            .O(N__53604),
            .I(REG_mem_13_1));
    LocalMux I__9666 (
            .O(N__53601),
            .I(REG_mem_13_1));
    InMux I__9665 (
            .O(N__53596),
            .I(N__53593));
    LocalMux I__9664 (
            .O(N__53593),
            .I(N__53590));
    Span4Mux_v I__9663 (
            .O(N__53590),
            .I(N__53586));
    InMux I__9662 (
            .O(N__53589),
            .I(N__53583));
    Odrv4 I__9661 (
            .O(N__53586),
            .I(REG_mem_42_1));
    LocalMux I__9660 (
            .O(N__53583),
            .I(REG_mem_42_1));
    InMux I__9659 (
            .O(N__53578),
            .I(N__53575));
    LocalMux I__9658 (
            .O(N__53575),
            .I(N__53572));
    Span4Mux_h I__9657 (
            .O(N__53572),
            .I(N__53568));
    InMux I__9656 (
            .O(N__53571),
            .I(N__53565));
    Odrv4 I__9655 (
            .O(N__53568),
            .I(REG_mem_38_1));
    LocalMux I__9654 (
            .O(N__53565),
            .I(REG_mem_38_1));
    InMux I__9653 (
            .O(N__53560),
            .I(N__53557));
    LocalMux I__9652 (
            .O(N__53557),
            .I(N__53553));
    InMux I__9651 (
            .O(N__53556),
            .I(N__53550));
    Odrv12 I__9650 (
            .O(N__53553),
            .I(REG_mem_39_1));
    LocalMux I__9649 (
            .O(N__53550),
            .I(REG_mem_39_1));
    InMux I__9648 (
            .O(N__53545),
            .I(N__53542));
    LocalMux I__9647 (
            .O(N__53542),
            .I(N__53539));
    Span4Mux_v I__9646 (
            .O(N__53539),
            .I(N__53536));
    Odrv4 I__9645 (
            .O(N__53536),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11702 ));
    InMux I__9644 (
            .O(N__53533),
            .I(N__53530));
    LocalMux I__9643 (
            .O(N__53530),
            .I(N__53527));
    Span4Mux_h I__9642 (
            .O(N__53527),
            .I(N__53524));
    Odrv4 I__9641 (
            .O(N__53524),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11660 ));
    InMux I__9640 (
            .O(N__53521),
            .I(N__53518));
    LocalMux I__9639 (
            .O(N__53518),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11659 ));
    CascadeMux I__9638 (
            .O(N__53515),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13994_cascade_ ));
    CascadeMux I__9637 (
            .O(N__53512),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11744_cascade_ ));
    InMux I__9636 (
            .O(N__53509),
            .I(N__53506));
    LocalMux I__9635 (
            .O(N__53506),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13349 ));
    InMux I__9634 (
            .O(N__53503),
            .I(N__53500));
    LocalMux I__9633 (
            .O(N__53500),
            .I(N__53497));
    Span4Mux_v I__9632 (
            .O(N__53497),
            .I(N__53494));
    Span4Mux_v I__9631 (
            .O(N__53494),
            .I(N__53491));
    Span4Mux_v I__9630 (
            .O(N__53491),
            .I(N__53488));
    Odrv4 I__9629 (
            .O(N__53488),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13379 ));
    InMux I__9628 (
            .O(N__53485),
            .I(N__53482));
    LocalMux I__9627 (
            .O(N__53482),
            .I(N__53479));
    Odrv12 I__9626 (
            .O(N__53479),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11678 ));
    CascadeMux I__9625 (
            .O(N__53476),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13355_cascade_ ));
    InMux I__9624 (
            .O(N__53473),
            .I(N__53470));
    LocalMux I__9623 (
            .O(N__53470),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13376 ));
    InMux I__9622 (
            .O(N__53467),
            .I(N__53463));
    InMux I__9621 (
            .O(N__53466),
            .I(N__53460));
    LocalMux I__9620 (
            .O(N__53463),
            .I(REG_mem_45_5));
    LocalMux I__9619 (
            .O(N__53460),
            .I(REG_mem_45_5));
    InMux I__9618 (
            .O(N__53455),
            .I(N__53452));
    LocalMux I__9617 (
            .O(N__53452),
            .I(N__53449));
    Span12Mux_v I__9616 (
            .O(N__53449),
            .I(N__53445));
    InMux I__9615 (
            .O(N__53448),
            .I(N__53442));
    Odrv12 I__9614 (
            .O(N__53445),
            .I(REG_mem_37_6));
    LocalMux I__9613 (
            .O(N__53442),
            .I(REG_mem_37_6));
    CascadeMux I__9612 (
            .O(N__53437),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13550_cascade_ ));
    InMux I__9611 (
            .O(N__53434),
            .I(N__53428));
    InMux I__9610 (
            .O(N__53433),
            .I(N__53428));
    LocalMux I__9609 (
            .O(N__53428),
            .I(REG_mem_36_6));
    CascadeMux I__9608 (
            .O(N__53425),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13340_cascade_ ));
    InMux I__9607 (
            .O(N__53422),
            .I(N__53419));
    LocalMux I__9606 (
            .O(N__53419),
            .I(N__53416));
    Span4Mux_v I__9605 (
            .O(N__53416),
            .I(N__53412));
    CascadeMux I__9604 (
            .O(N__53415),
            .I(N__53409));
    Span4Mux_v I__9603 (
            .O(N__53412),
            .I(N__53406));
    InMux I__9602 (
            .O(N__53409),
            .I(N__53403));
    Odrv4 I__9601 (
            .O(N__53406),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_5 ));
    LocalMux I__9600 (
            .O(N__53403),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_5 ));
    InMux I__9599 (
            .O(N__53398),
            .I(N__53395));
    LocalMux I__9598 (
            .O(N__53395),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13343 ));
    CascadeMux I__9597 (
            .O(N__53392),
            .I(N__53388));
    InMux I__9596 (
            .O(N__53391),
            .I(N__53383));
    InMux I__9595 (
            .O(N__53388),
            .I(N__53383));
    LocalMux I__9594 (
            .O(N__53383),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_5 ));
    CascadeMux I__9593 (
            .O(N__53380),
            .I(N__53376));
    CascadeMux I__9592 (
            .O(N__53379),
            .I(N__53373));
    InMux I__9591 (
            .O(N__53376),
            .I(N__53368));
    InMux I__9590 (
            .O(N__53373),
            .I(N__53368));
    LocalMux I__9589 (
            .O(N__53368),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_5 ));
    InMux I__9588 (
            .O(N__53365),
            .I(N__53362));
    LocalMux I__9587 (
            .O(N__53362),
            .I(N__53359));
    Span4Mux_v I__9586 (
            .O(N__53359),
            .I(N__53355));
    InMux I__9585 (
            .O(N__53358),
            .I(N__53352));
    Odrv4 I__9584 (
            .O(N__53355),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_15 ));
    LocalMux I__9583 (
            .O(N__53352),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_15 ));
    CascadeMux I__9582 (
            .O(N__53347),
            .I(N__53343));
    InMux I__9581 (
            .O(N__53346),
            .I(N__53340));
    InMux I__9580 (
            .O(N__53343),
            .I(N__53337));
    LocalMux I__9579 (
            .O(N__53340),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_5 ));
    LocalMux I__9578 (
            .O(N__53337),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_5 ));
    CascadeMux I__9577 (
            .O(N__53332),
            .I(N__53328));
    InMux I__9576 (
            .O(N__53331),
            .I(N__53325));
    InMux I__9575 (
            .O(N__53328),
            .I(N__53322));
    LocalMux I__9574 (
            .O(N__53325),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_5 ));
    LocalMux I__9573 (
            .O(N__53322),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_5 ));
    CascadeMux I__9572 (
            .O(N__53317),
            .I(N__53314));
    InMux I__9571 (
            .O(N__53314),
            .I(N__53311));
    LocalMux I__9570 (
            .O(N__53311),
            .I(N__53308));
    Odrv4 I__9569 (
            .O(N__53308),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11656 ));
    InMux I__9568 (
            .O(N__53305),
            .I(N__53302));
    LocalMux I__9567 (
            .O(N__53302),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11654 ));
    InMux I__9566 (
            .O(N__53299),
            .I(N__53296));
    LocalMux I__9565 (
            .O(N__53296),
            .I(N__53293));
    Span4Mux_v I__9564 (
            .O(N__53293),
            .I(N__53290));
    Span4Mux_h I__9563 (
            .O(N__53290),
            .I(N__53287));
    Odrv4 I__9562 (
            .O(N__53287),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11653 ));
    CascadeMux I__9561 (
            .O(N__53284),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13346_cascade_ ));
    InMux I__9560 (
            .O(N__53281),
            .I(N__53278));
    LocalMux I__9559 (
            .O(N__53278),
            .I(N__53275));
    Odrv4 I__9558 (
            .O(N__53275),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11672 ));
    InMux I__9557 (
            .O(N__53272),
            .I(N__53268));
    InMux I__9556 (
            .O(N__53271),
            .I(N__53265));
    LocalMux I__9555 (
            .O(N__53268),
            .I(REG_mem_14_1));
    LocalMux I__9554 (
            .O(N__53265),
            .I(REG_mem_14_1));
    InMux I__9553 (
            .O(N__53260),
            .I(N__53256));
    InMux I__9552 (
            .O(N__53259),
            .I(N__53253));
    LocalMux I__9551 (
            .O(N__53256),
            .I(REG_mem_18_1));
    LocalMux I__9550 (
            .O(N__53253),
            .I(REG_mem_18_1));
    InMux I__9549 (
            .O(N__53248),
            .I(N__53242));
    InMux I__9548 (
            .O(N__53247),
            .I(N__53242));
    LocalMux I__9547 (
            .O(N__53242),
            .I(REG_mem_19_1));
    InMux I__9546 (
            .O(N__53239),
            .I(N__53236));
    LocalMux I__9545 (
            .O(N__53236),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11555 ));
    InMux I__9544 (
            .O(N__53233),
            .I(N__53230));
    LocalMux I__9543 (
            .O(N__53230),
            .I(N__53226));
    InMux I__9542 (
            .O(N__53229),
            .I(N__53223));
    Odrv4 I__9541 (
            .O(N__53226),
            .I(REG_mem_36_1));
    LocalMux I__9540 (
            .O(N__53223),
            .I(REG_mem_36_1));
    InMux I__9539 (
            .O(N__53218),
            .I(N__53215));
    LocalMux I__9538 (
            .O(N__53215),
            .I(N__53212));
    Span4Mux_h I__9537 (
            .O(N__53212),
            .I(N__53209));
    Span4Mux_v I__9536 (
            .O(N__53209),
            .I(N__53205));
    InMux I__9535 (
            .O(N__53208),
            .I(N__53202));
    Odrv4 I__9534 (
            .O(N__53205),
            .I(REG_mem_37_1));
    LocalMux I__9533 (
            .O(N__53202),
            .I(REG_mem_37_1));
    InMux I__9532 (
            .O(N__53197),
            .I(N__53194));
    LocalMux I__9531 (
            .O(N__53194),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11701 ));
    InMux I__9530 (
            .O(N__53191),
            .I(N__53185));
    InMux I__9529 (
            .O(N__53190),
            .I(N__53185));
    LocalMux I__9528 (
            .O(N__53185),
            .I(REG_mem_58_5));
    CascadeMux I__9527 (
            .O(N__53182),
            .I(\spi0.n81_cascade_ ));
    InMux I__9526 (
            .O(N__53179),
            .I(N__53176));
    LocalMux I__9525 (
            .O(N__53176),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11699 ));
    CascadeMux I__9524 (
            .O(N__53173),
            .I(N__53169));
    InMux I__9523 (
            .O(N__53172),
            .I(N__53164));
    InMux I__9522 (
            .O(N__53169),
            .I(N__53164));
    LocalMux I__9521 (
            .O(N__53164),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_1 ));
    CascadeMux I__9520 (
            .O(N__53161),
            .I(N__53158));
    InMux I__9519 (
            .O(N__53158),
            .I(N__53155));
    LocalMux I__9518 (
            .O(N__53155),
            .I(N__53151));
    CascadeMux I__9517 (
            .O(N__53154),
            .I(N__53148));
    Span4Mux_h I__9516 (
            .O(N__53151),
            .I(N__53145));
    InMux I__9515 (
            .O(N__53148),
            .I(N__53142));
    Odrv4 I__9514 (
            .O(N__53145),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_2 ));
    LocalMux I__9513 (
            .O(N__53142),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_2 ));
    InMux I__9512 (
            .O(N__53137),
            .I(N__53134));
    LocalMux I__9511 (
            .O(N__53134),
            .I(N__53130));
    CascadeMux I__9510 (
            .O(N__53133),
            .I(N__53127));
    Span4Mux_v I__9509 (
            .O(N__53130),
            .I(N__53124));
    InMux I__9508 (
            .O(N__53127),
            .I(N__53121));
    Odrv4 I__9507 (
            .O(N__53124),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_5 ));
    LocalMux I__9506 (
            .O(N__53121),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_5 ));
    InMux I__9505 (
            .O(N__53116),
            .I(N__53110));
    InMux I__9504 (
            .O(N__53115),
            .I(N__53110));
    LocalMux I__9503 (
            .O(N__53110),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_5 ));
    InMux I__9502 (
            .O(N__53107),
            .I(N__53104));
    LocalMux I__9501 (
            .O(N__53104),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12089 ));
    InMux I__9500 (
            .O(N__53101),
            .I(N__53097));
    InMux I__9499 (
            .O(N__53100),
            .I(N__53094));
    LocalMux I__9498 (
            .O(N__53097),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_5 ));
    LocalMux I__9497 (
            .O(N__53094),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_5 ));
    InMux I__9496 (
            .O(N__53089),
            .I(N__53086));
    LocalMux I__9495 (
            .O(N__53086),
            .I(N__53083));
    Span4Mux_v I__9494 (
            .O(N__53083),
            .I(N__53079));
    CascadeMux I__9493 (
            .O(N__53082),
            .I(N__53076));
    Span4Mux_h I__9492 (
            .O(N__53079),
            .I(N__53073));
    InMux I__9491 (
            .O(N__53076),
            .I(N__53070));
    Odrv4 I__9490 (
            .O(N__53073),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_0 ));
    LocalMux I__9489 (
            .O(N__53070),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_0 ));
    InMux I__9488 (
            .O(N__53065),
            .I(N__53062));
    LocalMux I__9487 (
            .O(N__53062),
            .I(\spi0.n10106 ));
    CascadeMux I__9486 (
            .O(N__53059),
            .I(\spi0.n12598_cascade_ ));
    InMux I__9485 (
            .O(N__53056),
            .I(N__53053));
    LocalMux I__9484 (
            .O(N__53053),
            .I(N__53050));
    Odrv4 I__9483 (
            .O(N__53050),
            .I(\spi0.n14442 ));
    IoInMux I__9482 (
            .O(N__53047),
            .I(N__53044));
    LocalMux I__9481 (
            .O(N__53044),
            .I(N__53041));
    Span12Mux_s0_v I__9480 (
            .O(N__53041),
            .I(N__53038));
    Span12Mux_h I__9479 (
            .O(N__53038),
            .I(N__53035));
    Odrv12 I__9478 (
            .O(N__53035),
            .I(\spi0.CS_N_974 ));
    SRMux I__9477 (
            .O(N__53032),
            .I(N__53028));
    SRMux I__9476 (
            .O(N__53031),
            .I(N__53025));
    LocalMux I__9475 (
            .O(N__53028),
            .I(N__53022));
    LocalMux I__9474 (
            .O(N__53025),
            .I(N__53019));
    Span4Mux_h I__9473 (
            .O(N__53022),
            .I(N__53016));
    Span4Mux_v I__9472 (
            .O(N__53019),
            .I(N__53013));
    Odrv4 I__9471 (
            .O(N__53016),
            .I(\spi0.n10082 ));
    Odrv4 I__9470 (
            .O(N__53013),
            .I(\spi0.n10082 ));
    CascadeMux I__9469 (
            .O(N__53008),
            .I(\spi0.n10076_cascade_ ));
    InMux I__9468 (
            .O(N__53005),
            .I(N__53002));
    LocalMux I__9467 (
            .O(N__53002),
            .I(\spi0.n10081 ));
    InMux I__9466 (
            .O(N__52999),
            .I(N__52996));
    LocalMux I__9465 (
            .O(N__52996),
            .I(\spi0.n11398 ));
    InMux I__9464 (
            .O(N__52993),
            .I(N__52990));
    LocalMux I__9463 (
            .O(N__52990),
            .I(\spi0.n11350 ));
    CascadeMux I__9462 (
            .O(N__52987),
            .I(\spi0.n11398_cascade_ ));
    InMux I__9461 (
            .O(N__52984),
            .I(N__52981));
    LocalMux I__9460 (
            .O(N__52981),
            .I(\spi0.n81 ));
    InMux I__9459 (
            .O(N__52978),
            .I(N__52974));
    InMux I__9458 (
            .O(N__52977),
            .I(N__52971));
    LocalMux I__9457 (
            .O(N__52974),
            .I(\spi0.n11311 ));
    LocalMux I__9456 (
            .O(N__52971),
            .I(\spi0.n11311 ));
    CascadeMux I__9455 (
            .O(N__52966),
            .I(\spi0.n11311_cascade_ ));
    InMux I__9454 (
            .O(N__52963),
            .I(N__52960));
    LocalMux I__9453 (
            .O(N__52960),
            .I(\spi0.n11344 ));
    InMux I__9452 (
            .O(N__52957),
            .I(N__52951));
    InMux I__9451 (
            .O(N__52956),
            .I(N__52951));
    LocalMux I__9450 (
            .O(N__52951),
            .I(\spi0.n4105 ));
    CascadeMux I__9449 (
            .O(N__52948),
            .I(\spi0.n12607_cascade_ ));
    CEMux I__9448 (
            .O(N__52945),
            .I(N__52942));
    LocalMux I__9447 (
            .O(N__52942),
            .I(N__52939));
    Span4Mux_v I__9446 (
            .O(N__52939),
            .I(N__52935));
    CEMux I__9445 (
            .O(N__52938),
            .I(N__52932));
    Span4Mux_v I__9444 (
            .O(N__52935),
            .I(N__52927));
    LocalMux I__9443 (
            .O(N__52932),
            .I(N__52927));
    Odrv4 I__9442 (
            .O(N__52927),
            .I(\spi0.n4120 ));
    InMux I__9441 (
            .O(N__52924),
            .I(N__52921));
    LocalMux I__9440 (
            .O(N__52921),
            .I(\spi0.n12702 ));
    CascadeMux I__9439 (
            .O(N__52918),
            .I(\spi0.n4105_cascade_ ));
    CascadeMux I__9438 (
            .O(N__52915),
            .I(\spi0.n14442_cascade_ ));
    InMux I__9437 (
            .O(N__52912),
            .I(N__52909));
    LocalMux I__9436 (
            .O(N__52909),
            .I(\spi0.n10119 ));
    CEMux I__9435 (
            .O(N__52906),
            .I(N__52903));
    LocalMux I__9434 (
            .O(N__52903),
            .I(N__52900));
    Odrv4 I__9433 (
            .O(N__52900),
            .I(\spi0.n11345 ));
    CascadeMux I__9432 (
            .O(N__52897),
            .I(\spi0.n12594_cascade_ ));
    CascadeMux I__9431 (
            .O(N__52894),
            .I(\spi0.n3295_cascade_ ));
    CEMux I__9430 (
            .O(N__52891),
            .I(N__52888));
    LocalMux I__9429 (
            .O(N__52888),
            .I(\spi0.n11346 ));
    InMux I__9428 (
            .O(N__52885),
            .I(N__52882));
    LocalMux I__9427 (
            .O(N__52882),
            .I(\spi0.tx_shift_reg_3 ));
    InMux I__9426 (
            .O(N__52879),
            .I(N__52876));
    LocalMux I__9425 (
            .O(N__52876),
            .I(\spi0.tx_shift_reg_4 ));
    InMux I__9424 (
            .O(N__52873),
            .I(N__52870));
    LocalMux I__9423 (
            .O(N__52870),
            .I(\spi0.tx_shift_reg_5 ));
    InMux I__9422 (
            .O(N__52867),
            .I(N__52864));
    LocalMux I__9421 (
            .O(N__52864),
            .I(N__52860));
    InMux I__9420 (
            .O(N__52863),
            .I(N__52857));
    Span4Mux_h I__9419 (
            .O(N__52860),
            .I(N__52854));
    LocalMux I__9418 (
            .O(N__52857),
            .I(N__52847));
    Span4Mux_v I__9417 (
            .O(N__52854),
            .I(N__52847));
    InMux I__9416 (
            .O(N__52853),
            .I(N__52844));
    InMux I__9415 (
            .O(N__52852),
            .I(N__52841));
    Odrv4 I__9414 (
            .O(N__52847),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_6 ));
    LocalMux I__9413 (
            .O(N__52844),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_6 ));
    LocalMux I__9412 (
            .O(N__52841),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_6 ));
    InMux I__9411 (
            .O(N__52834),
            .I(N__52831));
    LocalMux I__9410 (
            .O(N__52831),
            .I(N__52828));
    Span4Mux_h I__9409 (
            .O(N__52828),
            .I(N__52825));
    Odrv4 I__9408 (
            .O(N__52825),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n2 ));
    CascadeMux I__9407 (
            .O(N__52822),
            .I(N__52819));
    InMux I__9406 (
            .O(N__52819),
            .I(N__52814));
    InMux I__9405 (
            .O(N__52818),
            .I(N__52809));
    InMux I__9404 (
            .O(N__52817),
            .I(N__52809));
    LocalMux I__9403 (
            .O(N__52814),
            .I(\spi0.n11317 ));
    LocalMux I__9402 (
            .O(N__52809),
            .I(\spi0.n11317 ));
    InMux I__9401 (
            .O(N__52804),
            .I(N__52801));
    LocalMux I__9400 (
            .O(N__52801),
            .I(N__52798));
    Span4Mux_h I__9399 (
            .O(N__52798),
            .I(N__52790));
    InMux I__9398 (
            .O(N__52797),
            .I(N__52783));
    InMux I__9397 (
            .O(N__52796),
            .I(N__52783));
    InMux I__9396 (
            .O(N__52795),
            .I(N__52783));
    InMux I__9395 (
            .O(N__52794),
            .I(N__52780));
    InMux I__9394 (
            .O(N__52793),
            .I(N__52777));
    Odrv4 I__9393 (
            .O(N__52790),
            .I(\spi0.counter_4 ));
    LocalMux I__9392 (
            .O(N__52783),
            .I(\spi0.counter_4 ));
    LocalMux I__9391 (
            .O(N__52780),
            .I(\spi0.counter_4 ));
    LocalMux I__9390 (
            .O(N__52777),
            .I(\spi0.counter_4 ));
    CascadeMux I__9389 (
            .O(N__52768),
            .I(\spi0.n24_cascade_ ));
    InMux I__9388 (
            .O(N__52765),
            .I(N__52762));
    LocalMux I__9387 (
            .O(N__52762),
            .I(\spi0.n16 ));
    CascadeMux I__9386 (
            .O(N__52759),
            .I(N__52756));
    InMux I__9385 (
            .O(N__52756),
            .I(N__52753));
    LocalMux I__9384 (
            .O(N__52753),
            .I(N__52750));
    Odrv4 I__9383 (
            .O(N__52750),
            .I(REG_out_raw_11));
    InMux I__9382 (
            .O(N__52747),
            .I(N__52744));
    LocalMux I__9381 (
            .O(N__52744),
            .I(N__52739));
    InMux I__9380 (
            .O(N__52743),
            .I(N__52736));
    InMux I__9379 (
            .O(N__52742),
            .I(N__52733));
    Odrv4 I__9378 (
            .O(N__52739),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_2 ));
    LocalMux I__9377 (
            .O(N__52736),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_2 ));
    LocalMux I__9376 (
            .O(N__52733),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_2 ));
    InMux I__9375 (
            .O(N__52726),
            .I(N__52723));
    LocalMux I__9374 (
            .O(N__52723),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11430 ));
    CascadeMux I__9373 (
            .O(N__52720),
            .I(N__52717));
    InMux I__9372 (
            .O(N__52717),
            .I(N__52714));
    LocalMux I__9371 (
            .O(N__52714),
            .I(N__52711));
    Span4Mux_v I__9370 (
            .O(N__52711),
            .I(N__52708));
    Odrv4 I__9369 (
            .O(N__52708),
            .I(REG_out_raw_0));
    InMux I__9368 (
            .O(N__52705),
            .I(N__52701));
    CascadeMux I__9367 (
            .O(N__52704),
            .I(N__52698));
    LocalMux I__9366 (
            .O(N__52701),
            .I(N__52693));
    InMux I__9365 (
            .O(N__52698),
            .I(N__52690));
    InMux I__9364 (
            .O(N__52697),
            .I(N__52685));
    InMux I__9363 (
            .O(N__52696),
            .I(N__52685));
    Odrv4 I__9362 (
            .O(N__52693),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_1 ));
    LocalMux I__9361 (
            .O(N__52690),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_1 ));
    LocalMux I__9360 (
            .O(N__52685),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_1 ));
    InMux I__9359 (
            .O(N__52678),
            .I(N__52675));
    LocalMux I__9358 (
            .O(N__52675),
            .I(N__52672));
    Odrv4 I__9357 (
            .O(N__52672),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_0 ));
    InMux I__9356 (
            .O(N__52669),
            .I(N__52663));
    InMux I__9355 (
            .O(N__52668),
            .I(N__52663));
    LocalMux I__9354 (
            .O(N__52663),
            .I(N__52659));
    InMux I__9353 (
            .O(N__52662),
            .I(N__52656));
    Odrv4 I__9352 (
            .O(N__52659),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_0 ));
    LocalMux I__9351 (
            .O(N__52656),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_0 ));
    InMux I__9350 (
            .O(N__52651),
            .I(N__52648));
    LocalMux I__9349 (
            .O(N__52648),
            .I(N__52645));
    Span4Mux_h I__9348 (
            .O(N__52645),
            .I(N__52641));
    InMux I__9347 (
            .O(N__52644),
            .I(N__52638));
    Odrv4 I__9346 (
            .O(N__52641),
            .I(rd_addr_nxt_c_6_N_465_1));
    LocalMux I__9345 (
            .O(N__52638),
            .I(rd_addr_nxt_c_6_N_465_1));
    InMux I__9344 (
            .O(N__52633),
            .I(N__52630));
    LocalMux I__9343 (
            .O(N__52630),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7_adj_1151 ));
    InMux I__9342 (
            .O(N__52627),
            .I(N__52624));
    LocalMux I__9341 (
            .O(N__52624),
            .I(\spi0.tx_shift_reg_1 ));
    InMux I__9340 (
            .O(N__52621),
            .I(N__52618));
    LocalMux I__9339 (
            .O(N__52618),
            .I(\spi0.tx_shift_reg_2 ));
    InMux I__9338 (
            .O(N__52615),
            .I(N__52612));
    LocalMux I__9337 (
            .O(N__52612),
            .I(N__52609));
    Odrv4 I__9336 (
            .O(N__52609),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11445 ));
    InMux I__9335 (
            .O(N__52606),
            .I(N__52603));
    LocalMux I__9334 (
            .O(N__52603),
            .I(N__52600));
    Sp12to4 I__9333 (
            .O(N__52600),
            .I(N__52597));
    Span12Mux_v I__9332 (
            .O(N__52597),
            .I(N__52594));
    Odrv12 I__9331 (
            .O(N__52594),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11408 ));
    CascadeMux I__9330 (
            .O(N__52591),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11483_cascade_ ));
    InMux I__9329 (
            .O(N__52588),
            .I(N__52585));
    LocalMux I__9328 (
            .O(N__52585),
            .I(N__52582));
    Odrv4 I__9327 (
            .O(N__52582),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10760 ));
    CascadeMux I__9326 (
            .O(N__52579),
            .I(N__52575));
    CascadeMux I__9325 (
            .O(N__52578),
            .I(N__52568));
    InMux I__9324 (
            .O(N__52575),
            .I(N__52563));
    InMux I__9323 (
            .O(N__52574),
            .I(N__52563));
    InMux I__9322 (
            .O(N__52573),
            .I(N__52553));
    InMux I__9321 (
            .O(N__52572),
            .I(N__52546));
    InMux I__9320 (
            .O(N__52571),
            .I(N__52546));
    InMux I__9319 (
            .O(N__52568),
            .I(N__52546));
    LocalMux I__9318 (
            .O(N__52563),
            .I(N__52543));
    InMux I__9317 (
            .O(N__52562),
            .I(N__52540));
    InMux I__9316 (
            .O(N__52561),
            .I(N__52527));
    InMux I__9315 (
            .O(N__52560),
            .I(N__52527));
    InMux I__9314 (
            .O(N__52559),
            .I(N__52527));
    InMux I__9313 (
            .O(N__52558),
            .I(N__52527));
    InMux I__9312 (
            .O(N__52557),
            .I(N__52527));
    InMux I__9311 (
            .O(N__52556),
            .I(N__52527));
    LocalMux I__9310 (
            .O(N__52553),
            .I(N__52522));
    LocalMux I__9309 (
            .O(N__52546),
            .I(N__52522));
    Span4Mux_h I__9308 (
            .O(N__52543),
            .I(N__52515));
    LocalMux I__9307 (
            .O(N__52540),
            .I(N__52515));
    LocalMux I__9306 (
            .O(N__52527),
            .I(N__52515));
    Span4Mux_h I__9305 (
            .O(N__52522),
            .I(N__52512));
    Span4Mux_h I__9304 (
            .O(N__52515),
            .I(N__52509));
    Span4Mux_v I__9303 (
            .O(N__52512),
            .I(N__52506));
    Span4Mux_v I__9302 (
            .O(N__52509),
            .I(N__52503));
    Odrv4 I__9301 (
            .O(N__52506),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_fifo_en_w ));
    Odrv4 I__9300 (
            .O(N__52503),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_fifo_en_w ));
    InMux I__9299 (
            .O(N__52498),
            .I(N__52495));
    LocalMux I__9298 (
            .O(N__52495),
            .I(N__52492));
    Odrv4 I__9297 (
            .O(N__52492),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7 ));
    InMux I__9296 (
            .O(N__52489),
            .I(N__52486));
    LocalMux I__9295 (
            .O(N__52486),
            .I(N__52483));
    Odrv4 I__9294 (
            .O(N__52483),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n8 ));
    InMux I__9293 (
            .O(N__52480),
            .I(N__52477));
    LocalMux I__9292 (
            .O(N__52477),
            .I(N__52474));
    Odrv4 I__9291 (
            .O(N__52474),
            .I(rd_sig_diff0_w_0));
    InMux I__9290 (
            .O(N__52471),
            .I(N__52468));
    LocalMux I__9289 (
            .O(N__52468),
            .I(N__52465));
    Odrv4 I__9288 (
            .O(N__52465),
            .I(rd_sig_diff0_w_1));
    CascadeMux I__9287 (
            .O(N__52462),
            .I(n5_cascade_));
    InMux I__9286 (
            .O(N__52459),
            .I(N__52456));
    LocalMux I__9285 (
            .O(N__52456),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.genblk16_rd_prev_r ));
    CascadeMux I__9284 (
            .O(N__52453),
            .I(\usb3_if_inst.n138_cascade_ ));
    CascadeMux I__9283 (
            .O(N__52450),
            .I(\usb3_if_inst.n2739_cascade_ ));
    InMux I__9282 (
            .O(N__52447),
            .I(N__52443));
    CascadeMux I__9281 (
            .O(N__52446),
            .I(N__52439));
    LocalMux I__9280 (
            .O(N__52443),
            .I(N__52436));
    CascadeMux I__9279 (
            .O(N__52442),
            .I(N__52431));
    InMux I__9278 (
            .O(N__52439),
            .I(N__52428));
    Span4Mux_v I__9277 (
            .O(N__52436),
            .I(N__52425));
    InMux I__9276 (
            .O(N__52435),
            .I(N__52422));
    InMux I__9275 (
            .O(N__52434),
            .I(N__52419));
    InMux I__9274 (
            .O(N__52431),
            .I(N__52416));
    LocalMux I__9273 (
            .O(N__52428),
            .I(N__52413));
    Sp12to4 I__9272 (
            .O(N__52425),
            .I(N__52406));
    LocalMux I__9271 (
            .O(N__52422),
            .I(N__52406));
    LocalMux I__9270 (
            .O(N__52419),
            .I(N__52406));
    LocalMux I__9269 (
            .O(N__52416),
            .I(wr_grey_sync_r_6));
    Odrv4 I__9268 (
            .O(N__52413),
            .I(wr_grey_sync_r_6));
    Odrv12 I__9267 (
            .O(N__52406),
            .I(wr_grey_sync_r_6));
    InMux I__9266 (
            .O(N__52399),
            .I(N__52396));
    LocalMux I__9265 (
            .O(N__52396),
            .I(wp_sync1_r_6));
    InMux I__9264 (
            .O(N__52393),
            .I(N__52390));
    LocalMux I__9263 (
            .O(N__52390),
            .I(N__52382));
    InMux I__9262 (
            .O(N__52389),
            .I(N__52379));
    InMux I__9261 (
            .O(N__52388),
            .I(N__52370));
    InMux I__9260 (
            .O(N__52387),
            .I(N__52370));
    InMux I__9259 (
            .O(N__52386),
            .I(N__52370));
    InMux I__9258 (
            .O(N__52385),
            .I(N__52370));
    Span4Mux_v I__9257 (
            .O(N__52382),
            .I(N__52363));
    LocalMux I__9256 (
            .O(N__52379),
            .I(N__52363));
    LocalMux I__9255 (
            .O(N__52370),
            .I(N__52363));
    Odrv4 I__9254 (
            .O(N__52363),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6 ));
    InMux I__9253 (
            .O(N__52360),
            .I(N__52357));
    LocalMux I__9252 (
            .O(N__52357),
            .I(N__52354));
    Span4Mux_v I__9251 (
            .O(N__52354),
            .I(N__52351));
    Span4Mux_v I__9250 (
            .O(N__52351),
            .I(N__52348));
    Span4Mux_h I__9249 (
            .O(N__52348),
            .I(N__52345));
    Odrv4 I__9248 (
            .O(N__52345),
            .I(wr_grey_sync_r_2));
    InMux I__9247 (
            .O(N__52342),
            .I(N__52339));
    LocalMux I__9246 (
            .O(N__52339),
            .I(N__52336));
    Odrv4 I__9245 (
            .O(N__52336),
            .I(wp_sync1_r_2));
    InMux I__9244 (
            .O(N__52333),
            .I(N__52330));
    LocalMux I__9243 (
            .O(N__52330),
            .I(N__52327));
    Odrv12 I__9242 (
            .O(N__52327),
            .I(REG_out_raw_7));
    InMux I__9241 (
            .O(N__52324),
            .I(N__52321));
    LocalMux I__9240 (
            .O(N__52321),
            .I(REG_out_raw_14));
    CascadeMux I__9239 (
            .O(N__52318),
            .I(N__52315));
    InMux I__9238 (
            .O(N__52315),
            .I(N__52312));
    LocalMux I__9237 (
            .O(N__52312),
            .I(N__52309));
    Span4Mux_h I__9236 (
            .O(N__52309),
            .I(N__52306));
    Span4Mux_v I__9235 (
            .O(N__52306),
            .I(N__52303));
    Odrv4 I__9234 (
            .O(N__52303),
            .I(REG_out_raw_13));
    CascadeMux I__9233 (
            .O(N__52300),
            .I(N__52296));
    InMux I__9232 (
            .O(N__52299),
            .I(N__52291));
    InMux I__9231 (
            .O(N__52296),
            .I(N__52291));
    LocalMux I__9230 (
            .O(N__52291),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_7 ));
    InMux I__9229 (
            .O(N__52288),
            .I(N__52284));
    InMux I__9228 (
            .O(N__52287),
            .I(N__52281));
    LocalMux I__9227 (
            .O(N__52284),
            .I(REG_mem_15_4));
    LocalMux I__9226 (
            .O(N__52281),
            .I(REG_mem_15_4));
    CascadeMux I__9225 (
            .O(N__52276),
            .I(\usb3_if_inst.n2912_cascade_ ));
    CascadeMux I__9224 (
            .O(N__52273),
            .I(\usb3_if_inst.n7_cascade_ ));
    InMux I__9223 (
            .O(N__52270),
            .I(N__52267));
    LocalMux I__9222 (
            .O(N__52267),
            .I(\usb3_if_inst.n137 ));
    InMux I__9221 (
            .O(N__52264),
            .I(N__52261));
    LocalMux I__9220 (
            .O(N__52261),
            .I(\usb3_if_inst.n3684 ));
    CascadeMux I__9219 (
            .O(N__52258),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12330_cascade_ ));
    CascadeMux I__9218 (
            .O(N__52255),
            .I(N__52252));
    InMux I__9217 (
            .O(N__52252),
            .I(N__52249));
    LocalMux I__9216 (
            .O(N__52249),
            .I(N__52246));
    Span4Mux_v I__9215 (
            .O(N__52246),
            .I(N__52243));
    Odrv4 I__9214 (
            .O(N__52243),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12180 ));
    InMux I__9213 (
            .O(N__52240),
            .I(N__52237));
    LocalMux I__9212 (
            .O(N__52237),
            .I(N__52234));
    Span12Mux_v I__9211 (
            .O(N__52234),
            .I(N__52231));
    Odrv12 I__9210 (
            .O(N__52231),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13466 ));
    InMux I__9209 (
            .O(N__52228),
            .I(N__52225));
    LocalMux I__9208 (
            .O(N__52225),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12288 ));
    InMux I__9207 (
            .O(N__52222),
            .I(N__52219));
    LocalMux I__9206 (
            .O(N__52219),
            .I(N__52216));
    Span12Mux_v I__9205 (
            .O(N__52216),
            .I(N__52213));
    Span12Mux_h I__9204 (
            .O(N__52213),
            .I(N__52210));
    Odrv12 I__9203 (
            .O(N__52210),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13580 ));
    CascadeMux I__9202 (
            .O(N__52207),
            .I(N__52204));
    InMux I__9201 (
            .O(N__52204),
            .I(N__52201));
    LocalMux I__9200 (
            .O(N__52201),
            .I(N__52198));
    Odrv4 I__9199 (
            .O(N__52198),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12120 ));
    InMux I__9198 (
            .O(N__52195),
            .I(N__52192));
    LocalMux I__9197 (
            .O(N__52192),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12282 ));
    CascadeMux I__9196 (
            .O(N__52189),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12258_cascade_ ));
    InMux I__9195 (
            .O(N__52186),
            .I(N__52183));
    LocalMux I__9194 (
            .O(N__52183),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13286 ));
    CascadeMux I__9193 (
            .O(N__52180),
            .I(N__52176));
    InMux I__9192 (
            .O(N__52179),
            .I(N__52171));
    InMux I__9191 (
            .O(N__52176),
            .I(N__52171));
    LocalMux I__9190 (
            .O(N__52171),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_7 ));
    CascadeMux I__9189 (
            .O(N__52168),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13880_cascade_ ));
    InMux I__9188 (
            .O(N__52165),
            .I(N__52162));
    LocalMux I__9187 (
            .O(N__52162),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12177 ));
    CascadeMux I__9186 (
            .O(N__52159),
            .I(N__52155));
    InMux I__9185 (
            .O(N__52158),
            .I(N__52150));
    InMux I__9184 (
            .O(N__52155),
            .I(N__52150));
    LocalMux I__9183 (
            .O(N__52150),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_7 ));
    InMux I__9182 (
            .O(N__52147),
            .I(N__52144));
    LocalMux I__9181 (
            .O(N__52144),
            .I(N__52140));
    InMux I__9180 (
            .O(N__52143),
            .I(N__52137));
    Odrv12 I__9179 (
            .O(N__52140),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_7 ));
    LocalMux I__9178 (
            .O(N__52137),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_7 ));
    InMux I__9177 (
            .O(N__52132),
            .I(N__52129));
    LocalMux I__9176 (
            .O(N__52129),
            .I(N__52126));
    Span4Mux_h I__9175 (
            .O(N__52126),
            .I(N__52123));
    Span4Mux_v I__9174 (
            .O(N__52123),
            .I(N__52119));
    CascadeMux I__9173 (
            .O(N__52122),
            .I(N__52116));
    Span4Mux_v I__9172 (
            .O(N__52119),
            .I(N__52113));
    InMux I__9171 (
            .O(N__52116),
            .I(N__52110));
    Odrv4 I__9170 (
            .O(N__52113),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_1 ));
    LocalMux I__9169 (
            .O(N__52110),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_1 ));
    InMux I__9168 (
            .O(N__52105),
            .I(N__52099));
    InMux I__9167 (
            .O(N__52104),
            .I(N__52099));
    LocalMux I__9166 (
            .O(N__52099),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_7 ));
    CascadeMux I__9165 (
            .O(N__52096),
            .I(N__52093));
    InMux I__9164 (
            .O(N__52093),
            .I(N__52087));
    InMux I__9163 (
            .O(N__52092),
            .I(N__52087));
    LocalMux I__9162 (
            .O(N__52087),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_7 ));
    InMux I__9161 (
            .O(N__52084),
            .I(N__52081));
    LocalMux I__9160 (
            .O(N__52081),
            .I(N__52078));
    Span4Mux_v I__9159 (
            .O(N__52078),
            .I(N__52075));
    Span4Mux_h I__9158 (
            .O(N__52075),
            .I(N__52072));
    Odrv4 I__9157 (
            .O(N__52072),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13478 ));
    InMux I__9156 (
            .O(N__52069),
            .I(N__52066));
    LocalMux I__9155 (
            .O(N__52066),
            .I(N__52063));
    Odrv4 I__9154 (
            .O(N__52063),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12144 ));
    InMux I__9153 (
            .O(N__52060),
            .I(N__52057));
    LocalMux I__9152 (
            .O(N__52057),
            .I(N__52054));
    Span4Mux_h I__9151 (
            .O(N__52054),
            .I(N__52051));
    Span4Mux_h I__9150 (
            .O(N__52051),
            .I(N__52048));
    Odrv4 I__9149 (
            .O(N__52048),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13316 ));
    CascadeMux I__9148 (
            .O(N__52045),
            .I(N__52042));
    InMux I__9147 (
            .O(N__52042),
            .I(N__52039));
    LocalMux I__9146 (
            .O(N__52039),
            .I(N__52036));
    Odrv4 I__9145 (
            .O(N__52036),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12222 ));
    CascadeMux I__9144 (
            .O(N__52033),
            .I(N__52030));
    InMux I__9143 (
            .O(N__52030),
            .I(N__52027));
    LocalMux I__9142 (
            .O(N__52027),
            .I(N__52024));
    Span4Mux_v I__9141 (
            .O(N__52024),
            .I(N__52020));
    InMux I__9140 (
            .O(N__52023),
            .I(N__52017));
    Odrv4 I__9139 (
            .O(N__52020),
            .I(REG_mem_17_7));
    LocalMux I__9138 (
            .O(N__52017),
            .I(REG_mem_17_7));
    InMux I__9137 (
            .O(N__52012),
            .I(N__52009));
    LocalMux I__9136 (
            .O(N__52009),
            .I(N__52006));
    Sp12to4 I__9135 (
            .O(N__52006),
            .I(N__52002));
    InMux I__9134 (
            .O(N__52005),
            .I(N__51999));
    Odrv12 I__9133 (
            .O(N__52002),
            .I(REG_mem_11_1));
    LocalMux I__9132 (
            .O(N__51999),
            .I(REG_mem_11_1));
    InMux I__9131 (
            .O(N__51994),
            .I(N__51988));
    InMux I__9130 (
            .O(N__51993),
            .I(N__51988));
    LocalMux I__9129 (
            .O(N__51988),
            .I(REG_mem_16_7));
    CascadeMux I__9128 (
            .O(N__51985),
            .I(N__51982));
    InMux I__9127 (
            .O(N__51982),
            .I(N__51979));
    LocalMux I__9126 (
            .O(N__51979),
            .I(N__51976));
    Span4Mux_v I__9125 (
            .O(N__51976),
            .I(N__51972));
    InMux I__9124 (
            .O(N__51975),
            .I(N__51969));
    Odrv4 I__9123 (
            .O(N__51972),
            .I(REG_mem_7_7));
    LocalMux I__9122 (
            .O(N__51969),
            .I(REG_mem_7_7));
    InMux I__9121 (
            .O(N__51964),
            .I(N__51960));
    InMux I__9120 (
            .O(N__51963),
            .I(N__51957));
    LocalMux I__9119 (
            .O(N__51960),
            .I(REG_mem_6_7));
    LocalMux I__9118 (
            .O(N__51957),
            .I(REG_mem_6_7));
    InMux I__9117 (
            .O(N__51952),
            .I(N__51948));
    InMux I__9116 (
            .O(N__51951),
            .I(N__51945));
    LocalMux I__9115 (
            .O(N__51948),
            .I(REG_mem_4_7));
    LocalMux I__9114 (
            .O(N__51945),
            .I(REG_mem_4_7));
    CascadeMux I__9113 (
            .O(N__51940),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14072_cascade_ ));
    InMux I__9112 (
            .O(N__51937),
            .I(N__51933));
    InMux I__9111 (
            .O(N__51936),
            .I(N__51930));
    LocalMux I__9110 (
            .O(N__51933),
            .I(REG_mem_5_7));
    LocalMux I__9109 (
            .O(N__51930),
            .I(REG_mem_5_7));
    CascadeMux I__9108 (
            .O(N__51925),
            .I(N__51922));
    InMux I__9107 (
            .O(N__51922),
            .I(N__51919));
    LocalMux I__9106 (
            .O(N__51919),
            .I(N__51915));
    CascadeMux I__9105 (
            .O(N__51918),
            .I(N__51912));
    Span4Mux_v I__9104 (
            .O(N__51915),
            .I(N__51909));
    InMux I__9103 (
            .O(N__51912),
            .I(N__51906));
    Odrv4 I__9102 (
            .O(N__51909),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_2 ));
    LocalMux I__9101 (
            .O(N__51906),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_2 ));
    InMux I__9100 (
            .O(N__51901),
            .I(N__51898));
    LocalMux I__9099 (
            .O(N__51898),
            .I(N__51894));
    InMux I__9098 (
            .O(N__51897),
            .I(N__51891));
    Odrv12 I__9097 (
            .O(N__51894),
            .I(REG_mem_5_5));
    LocalMux I__9096 (
            .O(N__51891),
            .I(REG_mem_5_5));
    InMux I__9095 (
            .O(N__51886),
            .I(N__51882));
    InMux I__9094 (
            .O(N__51885),
            .I(N__51879));
    LocalMux I__9093 (
            .O(N__51882),
            .I(REG_mem_5_0));
    LocalMux I__9092 (
            .O(N__51879),
            .I(REG_mem_5_0));
    CascadeMux I__9091 (
            .O(N__51874),
            .I(N__51871));
    InMux I__9090 (
            .O(N__51871),
            .I(N__51868));
    LocalMux I__9089 (
            .O(N__51868),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11761 ));
    CascadeMux I__9088 (
            .O(N__51865),
            .I(N__51862));
    InMux I__9087 (
            .O(N__51862),
            .I(N__51859));
    LocalMux I__9086 (
            .O(N__51859),
            .I(N__51855));
    InMux I__9085 (
            .O(N__51858),
            .I(N__51852));
    Odrv4 I__9084 (
            .O(N__51855),
            .I(REG_mem_9_0));
    LocalMux I__9083 (
            .O(N__51852),
            .I(REG_mem_9_0));
    InMux I__9082 (
            .O(N__51847),
            .I(N__51844));
    LocalMux I__9081 (
            .O(N__51844),
            .I(N__51841));
    Span4Mux_v I__9080 (
            .O(N__51841),
            .I(N__51838));
    Sp12to4 I__9079 (
            .O(N__51838),
            .I(N__51834));
    InMux I__9078 (
            .O(N__51837),
            .I(N__51831));
    Odrv12 I__9077 (
            .O(N__51834),
            .I(REG_mem_19_15));
    LocalMux I__9076 (
            .O(N__51831),
            .I(REG_mem_19_15));
    InMux I__9075 (
            .O(N__51826),
            .I(N__51822));
    InMux I__9074 (
            .O(N__51825),
            .I(N__51819));
    LocalMux I__9073 (
            .O(N__51822),
            .I(REG_mem_46_5));
    LocalMux I__9072 (
            .O(N__51819),
            .I(REG_mem_46_5));
    InMux I__9071 (
            .O(N__51814),
            .I(N__51811));
    LocalMux I__9070 (
            .O(N__51811),
            .I(N__51807));
    InMux I__9069 (
            .O(N__51810),
            .I(N__51804));
    Span4Mux_v I__9068 (
            .O(N__51807),
            .I(N__51799));
    LocalMux I__9067 (
            .O(N__51804),
            .I(N__51799));
    Odrv4 I__9066 (
            .O(N__51799),
            .I(REG_mem_11_0));
    CascadeMux I__9065 (
            .O(N__51796),
            .I(N__51793));
    InMux I__9064 (
            .O(N__51793),
            .I(N__51789));
    InMux I__9063 (
            .O(N__51792),
            .I(N__51786));
    LocalMux I__9062 (
            .O(N__51789),
            .I(REG_mem_10_0));
    LocalMux I__9061 (
            .O(N__51786),
            .I(REG_mem_10_0));
    InMux I__9060 (
            .O(N__51781),
            .I(N__51778));
    LocalMux I__9059 (
            .O(N__51778),
            .I(N__51775));
    Odrv4 I__9058 (
            .O(N__51775),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13856 ));
    CascadeMux I__9057 (
            .O(N__51772),
            .I(N__51769));
    InMux I__9056 (
            .O(N__51769),
            .I(N__51766));
    LocalMux I__9055 (
            .O(N__51766),
            .I(N__51763));
    Span4Mux_v I__9054 (
            .O(N__51763),
            .I(N__51760));
    Span4Mux_v I__9053 (
            .O(N__51760),
            .I(N__51756));
    InMux I__9052 (
            .O(N__51759),
            .I(N__51753));
    Odrv4 I__9051 (
            .O(N__51756),
            .I(REG_mem_43_5));
    LocalMux I__9050 (
            .O(N__51753),
            .I(REG_mem_43_5));
    CascadeMux I__9049 (
            .O(N__51748),
            .I(N__51745));
    InMux I__9048 (
            .O(N__51745),
            .I(N__51741));
    InMux I__9047 (
            .O(N__51744),
            .I(N__51738));
    LocalMux I__9046 (
            .O(N__51741),
            .I(N__51735));
    LocalMux I__9045 (
            .O(N__51738),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_2 ));
    Odrv4 I__9044 (
            .O(N__51735),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_2 ));
    InMux I__9043 (
            .O(N__51730),
            .I(N__51726));
    CascadeMux I__9042 (
            .O(N__51729),
            .I(N__51723));
    LocalMux I__9041 (
            .O(N__51726),
            .I(N__51720));
    InMux I__9040 (
            .O(N__51723),
            .I(N__51717));
    Span4Mux_v I__9039 (
            .O(N__51720),
            .I(N__51714));
    LocalMux I__9038 (
            .O(N__51717),
            .I(N__51711));
    Odrv4 I__9037 (
            .O(N__51714),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_2 ));
    Odrv4 I__9036 (
            .O(N__51711),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_2 ));
    CascadeMux I__9035 (
            .O(N__51706),
            .I(N__51702));
    InMux I__9034 (
            .O(N__51705),
            .I(N__51699));
    InMux I__9033 (
            .O(N__51702),
            .I(N__51696));
    LocalMux I__9032 (
            .O(N__51699),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_2 ));
    LocalMux I__9031 (
            .O(N__51696),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_2 ));
    InMux I__9030 (
            .O(N__51691),
            .I(N__51688));
    LocalMux I__9029 (
            .O(N__51688),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13574 ));
    InMux I__9028 (
            .O(N__51685),
            .I(N__51681));
    InMux I__9027 (
            .O(N__51684),
            .I(N__51678));
    LocalMux I__9026 (
            .O(N__51681),
            .I(REG_mem_6_0));
    LocalMux I__9025 (
            .O(N__51678),
            .I(REG_mem_6_0));
    InMux I__9024 (
            .O(N__51673),
            .I(N__51670));
    LocalMux I__9023 (
            .O(N__51670),
            .I(N__51666));
    InMux I__9022 (
            .O(N__51669),
            .I(N__51663));
    Odrv12 I__9021 (
            .O(N__51666),
            .I(REG_mem_6_5));
    LocalMux I__9020 (
            .O(N__51663),
            .I(REG_mem_6_5));
    CascadeMux I__9019 (
            .O(N__51658),
            .I(N__51655));
    InMux I__9018 (
            .O(N__51655),
            .I(N__51649));
    InMux I__9017 (
            .O(N__51654),
            .I(N__51649));
    LocalMux I__9016 (
            .O(N__51649),
            .I(REG_mem_47_5));
    InMux I__9015 (
            .O(N__51646),
            .I(N__51642));
    InMux I__9014 (
            .O(N__51645),
            .I(N__51639));
    LocalMux I__9013 (
            .O(N__51642),
            .I(REG_mem_38_7));
    LocalMux I__9012 (
            .O(N__51639),
            .I(REG_mem_38_7));
    InMux I__9011 (
            .O(N__51634),
            .I(N__51628));
    InMux I__9010 (
            .O(N__51633),
            .I(N__51628));
    LocalMux I__9009 (
            .O(N__51628),
            .I(N__51625));
    Odrv4 I__9008 (
            .O(N__51625),
            .I(REG_mem_8_1));
    InMux I__9007 (
            .O(N__51622),
            .I(N__51619));
    LocalMux I__9006 (
            .O(N__51619),
            .I(N__51616));
    Span4Mux_v I__9005 (
            .O(N__51616),
            .I(N__51613));
    Span4Mux_v I__9004 (
            .O(N__51613),
            .I(N__51610));
    Sp12to4 I__9003 (
            .O(N__51610),
            .I(N__51606));
    InMux I__9002 (
            .O(N__51609),
            .I(N__51603));
    Odrv12 I__9001 (
            .O(N__51606),
            .I(REG_mem_9_1));
    LocalMux I__9000 (
            .O(N__51603),
            .I(REG_mem_9_1));
    CascadeMux I__8999 (
            .O(N__51598),
            .I(N__51595));
    InMux I__8998 (
            .O(N__51595),
            .I(N__51592));
    LocalMux I__8997 (
            .O(N__51592),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14288 ));
    InMux I__8996 (
            .O(N__51589),
            .I(N__51586));
    LocalMux I__8995 (
            .O(N__51586),
            .I(N__51583));
    Span4Mux_v I__8994 (
            .O(N__51583),
            .I(N__51579));
    InMux I__8993 (
            .O(N__51582),
            .I(N__51576));
    Odrv4 I__8992 (
            .O(N__51579),
            .I(REG_mem_8_0));
    LocalMux I__8991 (
            .O(N__51576),
            .I(REG_mem_8_0));
    InMux I__8990 (
            .O(N__51571),
            .I(N__51568));
    LocalMux I__8989 (
            .O(N__51568),
            .I(N__51565));
    Span4Mux_v I__8988 (
            .O(N__51565),
            .I(N__51562));
    Odrv4 I__8987 (
            .O(N__51562),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13859 ));
    CascadeMux I__8986 (
            .O(N__51559),
            .I(N__51556));
    InMux I__8985 (
            .O(N__51556),
            .I(N__51553));
    LocalMux I__8984 (
            .O(N__51553),
            .I(N__51550));
    Span4Mux_v I__8983 (
            .O(N__51550),
            .I(N__51547));
    Sp12to4 I__8982 (
            .O(N__51547),
            .I(N__51543));
    InMux I__8981 (
            .O(N__51546),
            .I(N__51540));
    Odrv12 I__8980 (
            .O(N__51543),
            .I(REG_mem_44_5));
    LocalMux I__8979 (
            .O(N__51540),
            .I(REG_mem_44_5));
    InMux I__8978 (
            .O(N__51535),
            .I(N__51532));
    LocalMux I__8977 (
            .O(N__51532),
            .I(N__51529));
    Odrv4 I__8976 (
            .O(N__51529),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13577 ));
    CascadeMux I__8975 (
            .O(N__51526),
            .I(N__51522));
    InMux I__8974 (
            .O(N__51525),
            .I(N__51517));
    InMux I__8973 (
            .O(N__51522),
            .I(N__51517));
    LocalMux I__8972 (
            .O(N__51517),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_2 ));
    InMux I__8971 (
            .O(N__51514),
            .I(N__51511));
    LocalMux I__8970 (
            .O(N__51511),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14276 ));
    CascadeMux I__8969 (
            .O(N__51508),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12509_cascade_ ));
    InMux I__8968 (
            .O(N__51505),
            .I(N__51502));
    LocalMux I__8967 (
            .O(N__51502),
            .I(N__51499));
    Odrv4 I__8966 (
            .O(N__51499),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12508 ));
    InMux I__8965 (
            .O(N__51496),
            .I(N__51493));
    LocalMux I__8964 (
            .O(N__51493),
            .I(N__51490));
    Span12Mux_s8_v I__8963 (
            .O(N__51490),
            .I(N__51486));
    InMux I__8962 (
            .O(N__51489),
            .I(N__51483));
    Odrv12 I__8961 (
            .O(N__51486),
            .I(REG_mem_44_1));
    LocalMux I__8960 (
            .O(N__51483),
            .I(REG_mem_44_1));
    CascadeMux I__8959 (
            .O(N__51478),
            .I(N__51474));
    InMux I__8958 (
            .O(N__51477),
            .I(N__51469));
    InMux I__8957 (
            .O(N__51474),
            .I(N__51469));
    LocalMux I__8956 (
            .O(N__51469),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_5 ));
    InMux I__8955 (
            .O(N__51466),
            .I(N__51462));
    CascadeMux I__8954 (
            .O(N__51465),
            .I(N__51459));
    LocalMux I__8953 (
            .O(N__51462),
            .I(N__51456));
    InMux I__8952 (
            .O(N__51459),
            .I(N__51453));
    Odrv4 I__8951 (
            .O(N__51456),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_1 ));
    LocalMux I__8950 (
            .O(N__51453),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_1 ));
    InMux I__8949 (
            .O(N__51448),
            .I(N__51445));
    LocalMux I__8948 (
            .O(N__51445),
            .I(N__51442));
    Span4Mux_v I__8947 (
            .O(N__51442),
            .I(N__51438));
    CascadeMux I__8946 (
            .O(N__51441),
            .I(N__51435));
    Span4Mux_h I__8945 (
            .O(N__51438),
            .I(N__51432));
    InMux I__8944 (
            .O(N__51435),
            .I(N__51429));
    Odrv4 I__8943 (
            .O(N__51432),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_1 ));
    LocalMux I__8942 (
            .O(N__51429),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_1 ));
    CascadeMux I__8941 (
            .O(N__51424),
            .I(N__51421));
    InMux I__8940 (
            .O(N__51421),
            .I(N__51418));
    LocalMux I__8939 (
            .O(N__51418),
            .I(N__51415));
    Span4Mux_v I__8938 (
            .O(N__51415),
            .I(N__51411));
    InMux I__8937 (
            .O(N__51414),
            .I(N__51408));
    Odrv4 I__8936 (
            .O(N__51411),
            .I(REG_mem_40_1));
    LocalMux I__8935 (
            .O(N__51408),
            .I(REG_mem_40_1));
    InMux I__8934 (
            .O(N__51403),
            .I(N__51400));
    LocalMux I__8933 (
            .O(N__51400),
            .I(N__51397));
    Odrv4 I__8932 (
            .O(N__51397),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11704 ));
    CascadeMux I__8931 (
            .O(N__51394),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11489_cascade_ ));
    CascadeMux I__8930 (
            .O(N__51391),
            .I(N__51388));
    InMux I__8929 (
            .O(N__51388),
            .I(N__51385));
    LocalMux I__8928 (
            .O(N__51385),
            .I(N__51382));
    Span4Mux_v I__8927 (
            .O(N__51382),
            .I(N__51379));
    Odrv4 I__8926 (
            .O(N__51379),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13217 ));
    InMux I__8925 (
            .O(N__51376),
            .I(N__51373));
    LocalMux I__8924 (
            .O(N__51373),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14258 ));
    InMux I__8923 (
            .O(N__51370),
            .I(N__51366));
    InMux I__8922 (
            .O(N__51369),
            .I(N__51363));
    LocalMux I__8921 (
            .O(N__51366),
            .I(REG_mem_38_5));
    LocalMux I__8920 (
            .O(N__51363),
            .I(REG_mem_38_5));
    CascadeMux I__8919 (
            .O(N__51358),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12131_cascade_ ));
    InMux I__8918 (
            .O(N__51355),
            .I(N__51352));
    LocalMux I__8917 (
            .O(N__51352),
            .I(N__51349));
    Odrv4 I__8916 (
            .O(N__51349),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12130 ));
    InMux I__8915 (
            .O(N__51346),
            .I(N__51343));
    LocalMux I__8914 (
            .O(N__51343),
            .I(N__51340));
    Span4Mux_v I__8913 (
            .O(N__51340),
            .I(N__51337));
    Odrv4 I__8912 (
            .O(N__51337),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12088 ));
    CascadeMux I__8911 (
            .O(N__51334),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12818_cascade_ ));
    InMux I__8910 (
            .O(N__51331),
            .I(N__51328));
    LocalMux I__8909 (
            .O(N__51328),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12821 ));
    CascadeMux I__8908 (
            .O(N__51325),
            .I(N__51322));
    InMux I__8907 (
            .O(N__51322),
            .I(N__51319));
    LocalMux I__8906 (
            .O(N__51319),
            .I(N__51316));
    Span4Mux_v I__8905 (
            .O(N__51316),
            .I(N__51312));
    InMux I__8904 (
            .O(N__51315),
            .I(N__51309));
    Odrv4 I__8903 (
            .O(N__51312),
            .I(REG_mem_7_5));
    LocalMux I__8902 (
            .O(N__51309),
            .I(REG_mem_7_5));
    CascadeMux I__8901 (
            .O(N__51304),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11507_cascade_ ));
    InMux I__8900 (
            .O(N__51301),
            .I(N__51298));
    LocalMux I__8899 (
            .O(N__51298),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11506 ));
    InMux I__8898 (
            .O(N__51295),
            .I(N__51292));
    LocalMux I__8897 (
            .O(N__51292),
            .I(\spi0.n4409 ));
    CascadeMux I__8896 (
            .O(N__51289),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13844_cascade_ ));
    InMux I__8895 (
            .O(N__51286),
            .I(N__51283));
    LocalMux I__8894 (
            .O(N__51283),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11750 ));
    InMux I__8893 (
            .O(N__51280),
            .I(N__51277));
    LocalMux I__8892 (
            .O(N__51277),
            .I(N__51274));
    Sp12to4 I__8891 (
            .O(N__51274),
            .I(N__51271));
    Span12Mux_v I__8890 (
            .O(N__51271),
            .I(N__51268));
    Odrv12 I__8889 (
            .O(N__51268),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13847 ));
    CascadeMux I__8888 (
            .O(N__51265),
            .I(N__51262));
    InMux I__8887 (
            .O(N__51262),
            .I(N__51259));
    LocalMux I__8886 (
            .O(N__51259),
            .I(N__51256));
    Span4Mux_h I__8885 (
            .O(N__51256),
            .I(N__51253));
    Odrv4 I__8884 (
            .O(N__51253),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11713 ));
    InMux I__8883 (
            .O(N__51250),
            .I(N__51247));
    LocalMux I__8882 (
            .O(N__51247),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11714 ));
    CascadeMux I__8881 (
            .O(N__51244),
            .I(N__51241));
    InMux I__8880 (
            .O(N__51241),
            .I(N__51238));
    LocalMux I__8879 (
            .O(N__51238),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13970 ));
    InMux I__8878 (
            .O(N__51235),
            .I(N__51232));
    LocalMux I__8877 (
            .O(N__51232),
            .I(N__51229));
    Odrv12 I__8876 (
            .O(N__51229),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11698 ));
    CascadeMux I__8875 (
            .O(N__51226),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13358_cascade_ ));
    InMux I__8874 (
            .O(N__51223),
            .I(N__51220));
    LocalMux I__8873 (
            .O(N__51220),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13361 ));
    InMux I__8872 (
            .O(N__51217),
            .I(N__51214));
    LocalMux I__8871 (
            .O(N__51214),
            .I(N__51210));
    InMux I__8870 (
            .O(N__51213),
            .I(N__51207));
    Odrv4 I__8869 (
            .O(N__51210),
            .I(REG_mem_43_1));
    LocalMux I__8868 (
            .O(N__51207),
            .I(REG_mem_43_1));
    InMux I__8867 (
            .O(N__51202),
            .I(N__51199));
    LocalMux I__8866 (
            .O(N__51199),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11705 ));
    InMux I__8865 (
            .O(N__51196),
            .I(N__51193));
    LocalMux I__8864 (
            .O(N__51193),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13745 ));
    CascadeMux I__8863 (
            .O(N__51190),
            .I(\spi0.n19_cascade_ ));
    CascadeMux I__8862 (
            .O(N__51187),
            .I(N__51184));
    InMux I__8861 (
            .O(N__51184),
            .I(N__51181));
    LocalMux I__8860 (
            .O(N__51181),
            .I(\spi0.n88 ));
    InMux I__8859 (
            .O(N__51178),
            .I(N__51172));
    InMux I__8858 (
            .O(N__51177),
            .I(N__51172));
    LocalMux I__8857 (
            .O(N__51172),
            .I(\spi0.n8 ));
    InMux I__8856 (
            .O(N__51169),
            .I(N__51166));
    LocalMux I__8855 (
            .O(N__51166),
            .I(\spi0.n12566 ));
    CascadeMux I__8854 (
            .O(N__51163),
            .I(\spi0.n12567_cascade_ ));
    IoInMux I__8853 (
            .O(N__51160),
            .I(N__51157));
    LocalMux I__8852 (
            .O(N__51157),
            .I(N__51154));
    Span4Mux_s3_v I__8851 (
            .O(N__51154),
            .I(N__51151));
    Sp12to4 I__8850 (
            .O(N__51151),
            .I(N__51148));
    Span12Mux_h I__8849 (
            .O(N__51148),
            .I(N__51145));
    Odrv12 I__8848 (
            .O(N__51145),
            .I(\spi0.SCLK_N_977 ));
    InMux I__8847 (
            .O(N__51142),
            .I(N__51139));
    LocalMux I__8846 (
            .O(N__51139),
            .I(\spi0.n11351 ));
    CascadeMux I__8845 (
            .O(N__51136),
            .I(\spi0.n2_cascade_ ));
    CascadeMux I__8844 (
            .O(N__51133),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n4025_cascade_ ));
    InMux I__8843 (
            .O(N__51130),
            .I(N__51126));
    InMux I__8842 (
            .O(N__51129),
            .I(N__51123));
    LocalMux I__8841 (
            .O(N__51126),
            .I(N__51119));
    LocalMux I__8840 (
            .O(N__51123),
            .I(N__51116));
    InMux I__8839 (
            .O(N__51122),
            .I(N__51113));
    Span4Mux_v I__8838 (
            .O(N__51119),
            .I(N__51110));
    Span4Mux_v I__8837 (
            .O(N__51116),
            .I(N__51107));
    LocalMux I__8836 (
            .O(N__51113),
            .I(N__51104));
    Span4Mux_h I__8835 (
            .O(N__51110),
            .I(N__51097));
    Span4Mux_v I__8834 (
            .O(N__51107),
            .I(N__51097));
    Span4Mux_h I__8833 (
            .O(N__51104),
            .I(N__51097));
    Odrv4 I__8832 (
            .O(N__51097),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_0 ));
    InMux I__8831 (
            .O(N__51094),
            .I(N__51091));
    LocalMux I__8830 (
            .O(N__51091),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12_adj_1158 ));
    InMux I__8829 (
            .O(N__51088),
            .I(N__51085));
    LocalMux I__8828 (
            .O(N__51085),
            .I(N__51082));
    Span4Mux_v I__8827 (
            .O(N__51082),
            .I(N__51079));
    Span4Mux_h I__8826 (
            .O(N__51079),
            .I(N__51076));
    Sp12to4 I__8825 (
            .O(N__51076),
            .I(N__51073));
    Odrv12 I__8824 (
            .O(N__51073),
            .I(wr_grey_sync_r_0));
    InMux I__8823 (
            .O(N__51070),
            .I(N__51067));
    LocalMux I__8822 (
            .O(N__51067),
            .I(wp_sync1_r_0));
    InMux I__8821 (
            .O(N__51064),
            .I(N__51060));
    InMux I__8820 (
            .O(N__51063),
            .I(N__51057));
    LocalMux I__8819 (
            .O(N__51060),
            .I(\spi0.counter_5 ));
    LocalMux I__8818 (
            .O(N__51057),
            .I(\spi0.counter_5 ));
    InMux I__8817 (
            .O(N__51052),
            .I(N__51048));
    InMux I__8816 (
            .O(N__51051),
            .I(N__51045));
    LocalMux I__8815 (
            .O(N__51048),
            .I(\spi0.counter_9 ));
    LocalMux I__8814 (
            .O(N__51045),
            .I(\spi0.counter_9 ));
    CascadeMux I__8813 (
            .O(N__51040),
            .I(N__51037));
    InMux I__8812 (
            .O(N__51037),
            .I(N__51033));
    InMux I__8811 (
            .O(N__51036),
            .I(N__51030));
    LocalMux I__8810 (
            .O(N__51033),
            .I(\spi0.counter_8 ));
    LocalMux I__8809 (
            .O(N__51030),
            .I(\spi0.counter_8 ));
    InMux I__8808 (
            .O(N__51025),
            .I(N__51021));
    InMux I__8807 (
            .O(N__51024),
            .I(N__51018));
    LocalMux I__8806 (
            .O(N__51021),
            .I(\spi0.counter_6 ));
    LocalMux I__8805 (
            .O(N__51018),
            .I(\spi0.counter_6 ));
    InMux I__8804 (
            .O(N__51013),
            .I(N__51009));
    InMux I__8803 (
            .O(N__51012),
            .I(N__51006));
    LocalMux I__8802 (
            .O(N__51009),
            .I(\spi0.counter_7 ));
    LocalMux I__8801 (
            .O(N__51006),
            .I(\spi0.counter_7 ));
    InMux I__8800 (
            .O(N__51001),
            .I(N__50991));
    InMux I__8799 (
            .O(N__51000),
            .I(N__50991));
    InMux I__8798 (
            .O(N__50999),
            .I(N__50991));
    InMux I__8797 (
            .O(N__50998),
            .I(N__50988));
    LocalMux I__8796 (
            .O(N__50991),
            .I(\spi0.counter_3 ));
    LocalMux I__8795 (
            .O(N__50988),
            .I(\spi0.counter_3 ));
    InMux I__8794 (
            .O(N__50983),
            .I(N__50973));
    InMux I__8793 (
            .O(N__50982),
            .I(N__50973));
    InMux I__8792 (
            .O(N__50981),
            .I(N__50973));
    InMux I__8791 (
            .O(N__50980),
            .I(N__50970));
    LocalMux I__8790 (
            .O(N__50973),
            .I(\spi0.counter_1 ));
    LocalMux I__8789 (
            .O(N__50970),
            .I(\spi0.counter_1 ));
    CascadeMux I__8788 (
            .O(N__50965),
            .I(N__50960));
    InMux I__8787 (
            .O(N__50964),
            .I(N__50956));
    InMux I__8786 (
            .O(N__50963),
            .I(N__50951));
    InMux I__8785 (
            .O(N__50960),
            .I(N__50951));
    InMux I__8784 (
            .O(N__50959),
            .I(N__50948));
    LocalMux I__8783 (
            .O(N__50956),
            .I(\spi0.counter_2 ));
    LocalMux I__8782 (
            .O(N__50951),
            .I(\spi0.counter_2 ));
    LocalMux I__8781 (
            .O(N__50948),
            .I(\spi0.counter_2 ));
    CascadeMux I__8780 (
            .O(N__50941),
            .I(N__50937));
    InMux I__8779 (
            .O(N__50940),
            .I(N__50928));
    InMux I__8778 (
            .O(N__50937),
            .I(N__50928));
    InMux I__8777 (
            .O(N__50936),
            .I(N__50928));
    InMux I__8776 (
            .O(N__50935),
            .I(N__50925));
    LocalMux I__8775 (
            .O(N__50928),
            .I(\spi0.counter_0 ));
    LocalMux I__8774 (
            .O(N__50925),
            .I(\spi0.counter_0 ));
    InMux I__8773 (
            .O(N__50920),
            .I(N__50917));
    LocalMux I__8772 (
            .O(N__50917),
            .I(\spi0.n9 ));
    CascadeMux I__8771 (
            .O(N__50914),
            .I(\spi0.n3909_cascade_ ));
    InMux I__8770 (
            .O(N__50911),
            .I(N__50908));
    LocalMux I__8769 (
            .O(N__50908),
            .I(\spi0.n14 ));
    CascadeMux I__8768 (
            .O(N__50905),
            .I(N__50902));
    InMux I__8767 (
            .O(N__50902),
            .I(N__50899));
    LocalMux I__8766 (
            .O(N__50899),
            .I(N__50896));
    Span4Mux_v I__8765 (
            .O(N__50896),
            .I(N__50893));
    Odrv4 I__8764 (
            .O(N__50893),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n4 ));
    InMux I__8763 (
            .O(N__50890),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10622 ));
    InMux I__8762 (
            .O(N__50887),
            .I(N__50884));
    LocalMux I__8761 (
            .O(N__50884),
            .I(N__50881));
    Odrv12 I__8760 (
            .O(N__50881),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_sig_diff0_w_2 ));
    InMux I__8759 (
            .O(N__50878),
            .I(N__50875));
    LocalMux I__8758 (
            .O(N__50875),
            .I(N__50872));
    Span4Mux_v I__8757 (
            .O(N__50872),
            .I(N__50869));
    Sp12to4 I__8756 (
            .O(N__50869),
            .I(N__50866));
    Odrv12 I__8755 (
            .O(N__50866),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n3 ));
    CascadeMux I__8754 (
            .O(N__50863),
            .I(N__50860));
    InMux I__8753 (
            .O(N__50860),
            .I(N__50857));
    LocalMux I__8752 (
            .O(N__50857),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_5 ));
    InMux I__8751 (
            .O(N__50854),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10623 ));
    InMux I__8750 (
            .O(N__50851),
            .I(N__50848));
    LocalMux I__8749 (
            .O(N__50848),
            .I(N__50845));
    Span4Mux_v I__8748 (
            .O(N__50845),
            .I(N__50842));
    Odrv4 I__8747 (
            .O(N__50842),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n2_adj_1149 ));
    CascadeMux I__8746 (
            .O(N__50839),
            .I(N__50836));
    InMux I__8745 (
            .O(N__50836),
            .I(N__50833));
    LocalMux I__8744 (
            .O(N__50833),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_sig_diff0_w_4 ));
    InMux I__8743 (
            .O(N__50830),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10624 ));
    InMux I__8742 (
            .O(N__50827),
            .I(N__50824));
    LocalMux I__8741 (
            .O(N__50824),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n6 ));
    CascadeMux I__8740 (
            .O(N__50821),
            .I(N__50818));
    InMux I__8739 (
            .O(N__50818),
            .I(N__50815));
    LocalMux I__8738 (
            .O(N__50815),
            .I(N__50811));
    InMux I__8737 (
            .O(N__50814),
            .I(N__50808));
    Span4Mux_v I__8736 (
            .O(N__50811),
            .I(N__50805));
    LocalMux I__8735 (
            .O(N__50808),
            .I(N__50802));
    Span4Mux_h I__8734 (
            .O(N__50805),
            .I(N__50799));
    Span4Mux_v I__8733 (
            .O(N__50802),
            .I(N__50796));
    Odrv4 I__8732 (
            .O(N__50799),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_1 ));
    Odrv4 I__8731 (
            .O(N__50796),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_1 ));
    InMux I__8730 (
            .O(N__50791),
            .I(N__50787));
    InMux I__8729 (
            .O(N__50790),
            .I(N__50784));
    LocalMux I__8728 (
            .O(N__50787),
            .I(N__50781));
    LocalMux I__8727 (
            .O(N__50784),
            .I(N__50777));
    Span4Mux_v I__8726 (
            .O(N__50781),
            .I(N__50774));
    InMux I__8725 (
            .O(N__50780),
            .I(N__50771));
    Span4Mux_v I__8724 (
            .O(N__50777),
            .I(N__50768));
    Span4Mux_v I__8723 (
            .O(N__50774),
            .I(N__50763));
    LocalMux I__8722 (
            .O(N__50771),
            .I(N__50763));
    Sp12to4 I__8721 (
            .O(N__50768),
            .I(N__50758));
    Sp12to4 I__8720 (
            .O(N__50763),
            .I(N__50758));
    Odrv12 I__8719 (
            .O(N__50758),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_6 ));
    CascadeMux I__8718 (
            .O(N__50755),
            .I(N__50751));
    InMux I__8717 (
            .O(N__50754),
            .I(N__50747));
    InMux I__8716 (
            .O(N__50751),
            .I(N__50742));
    InMux I__8715 (
            .O(N__50750),
            .I(N__50742));
    LocalMux I__8714 (
            .O(N__50747),
            .I(N__50738));
    LocalMux I__8713 (
            .O(N__50742),
            .I(N__50735));
    InMux I__8712 (
            .O(N__50741),
            .I(N__50732));
    Span12Mux_h I__8711 (
            .O(N__50738),
            .I(N__50729));
    Span4Mux_v I__8710 (
            .O(N__50735),
            .I(N__50724));
    LocalMux I__8709 (
            .O(N__50732),
            .I(N__50724));
    Odrv12 I__8708 (
            .O(N__50729),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_2 ));
    Odrv4 I__8707 (
            .O(N__50724),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_2 ));
    CascadeMux I__8706 (
            .O(N__50719),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n8_adj_1157_cascade_ ));
    CascadeMux I__8705 (
            .O(N__50716),
            .I(N__50713));
    InMux I__8704 (
            .O(N__50713),
            .I(N__50710));
    LocalMux I__8703 (
            .O(N__50710),
            .I(N__50706));
    InMux I__8702 (
            .O(N__50709),
            .I(N__50703));
    Odrv4 I__8701 (
            .O(N__50706),
            .I(REG_mem_39_10));
    LocalMux I__8700 (
            .O(N__50703),
            .I(REG_mem_39_10));
    InMux I__8699 (
            .O(N__50698),
            .I(N__50695));
    LocalMux I__8698 (
            .O(N__50695),
            .I(N__50691));
    CascadeMux I__8697 (
            .O(N__50694),
            .I(N__50688));
    Span4Mux_v I__8696 (
            .O(N__50691),
            .I(N__50685));
    InMux I__8695 (
            .O(N__50688),
            .I(N__50682));
    Odrv4 I__8694 (
            .O(N__50685),
            .I(REG_mem_38_10));
    LocalMux I__8693 (
            .O(N__50682),
            .I(REG_mem_38_10));
    CascadeMux I__8692 (
            .O(N__50677),
            .I(N__50674));
    InMux I__8691 (
            .O(N__50674),
            .I(N__50671));
    LocalMux I__8690 (
            .O(N__50671),
            .I(N__50668));
    Span4Mux_v I__8689 (
            .O(N__50668),
            .I(N__50665));
    Span4Mux_h I__8688 (
            .O(N__50665),
            .I(N__50662));
    Span4Mux_h I__8687 (
            .O(N__50662),
            .I(N__50659));
    Odrv4 I__8686 (
            .O(N__50659),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11585 ));
    InMux I__8685 (
            .O(N__50656),
            .I(N__50650));
    InMux I__8684 (
            .O(N__50655),
            .I(N__50650));
    LocalMux I__8683 (
            .O(N__50650),
            .I(N__50646));
    InMux I__8682 (
            .O(N__50649),
            .I(N__50643));
    Odrv4 I__8681 (
            .O(N__50646),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_4 ));
    LocalMux I__8680 (
            .O(N__50643),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_4 ));
    InMux I__8679 (
            .O(N__50638),
            .I(N__50633));
    InMux I__8678 (
            .O(N__50637),
            .I(N__50628));
    InMux I__8677 (
            .O(N__50636),
            .I(N__50628));
    LocalMux I__8676 (
            .O(N__50633),
            .I(N__50625));
    LocalMux I__8675 (
            .O(N__50628),
            .I(N__50621));
    Span4Mux_v I__8674 (
            .O(N__50625),
            .I(N__50618));
    InMux I__8673 (
            .O(N__50624),
            .I(N__50615));
    Span4Mux_h I__8672 (
            .O(N__50621),
            .I(N__50612));
    Sp12to4 I__8671 (
            .O(N__50618),
            .I(N__50607));
    LocalMux I__8670 (
            .O(N__50615),
            .I(N__50607));
    Odrv4 I__8669 (
            .O(N__50612),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_4 ));
    Odrv12 I__8668 (
            .O(N__50607),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_4 ));
    InMux I__8667 (
            .O(N__50602),
            .I(N__50599));
    LocalMux I__8666 (
            .O(N__50599),
            .I(N__50596));
    Span4Mux_v I__8665 (
            .O(N__50596),
            .I(N__50593));
    Span4Mux_h I__8664 (
            .O(N__50593),
            .I(N__50590));
    Odrv4 I__8663 (
            .O(N__50590),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10 ));
    InMux I__8662 (
            .O(N__50587),
            .I(N__50584));
    LocalMux I__8661 (
            .O(N__50584),
            .I(wp_sync1_r_1));
    CascadeMux I__8660 (
            .O(N__50581),
            .I(N__50577));
    CascadeMux I__8659 (
            .O(N__50580),
            .I(N__50574));
    InMux I__8658 (
            .O(N__50577),
            .I(N__50571));
    InMux I__8657 (
            .O(N__50574),
            .I(N__50568));
    LocalMux I__8656 (
            .O(N__50571),
            .I(N__50565));
    LocalMux I__8655 (
            .O(N__50568),
            .I(N__50562));
    Span4Mux_v I__8654 (
            .O(N__50565),
            .I(N__50559));
    Span4Mux_v I__8653 (
            .O(N__50562),
            .I(N__50556));
    Span4Mux_h I__8652 (
            .O(N__50559),
            .I(N__50551));
    Span4Mux_h I__8651 (
            .O(N__50556),
            .I(N__50551));
    Odrv4 I__8650 (
            .O(N__50551),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n4027 ));
    InMux I__8649 (
            .O(N__50548),
            .I(N__50536));
    InMux I__8648 (
            .O(N__50547),
            .I(N__50536));
    InMux I__8647 (
            .O(N__50546),
            .I(N__50536));
    InMux I__8646 (
            .O(N__50545),
            .I(N__50536));
    LocalMux I__8645 (
            .O(N__50536),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_5 ));
    CascadeMux I__8644 (
            .O(N__50533),
            .I(N__50529));
    InMux I__8643 (
            .O(N__50532),
            .I(N__50526));
    InMux I__8642 (
            .O(N__50529),
            .I(N__50523));
    LocalMux I__8641 (
            .O(N__50526),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_4 ));
    LocalMux I__8640 (
            .O(N__50523),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_4 ));
    InMux I__8639 (
            .O(N__50518),
            .I(N__50512));
    InMux I__8638 (
            .O(N__50517),
            .I(N__50512));
    LocalMux I__8637 (
            .O(N__50512),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_3 ));
    InMux I__8636 (
            .O(N__50509),
            .I(N__50503));
    InMux I__8635 (
            .O(N__50508),
            .I(N__50503));
    LocalMux I__8634 (
            .O(N__50503),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_2 ));
    CascadeMux I__8633 (
            .O(N__50500),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_3_cascade_ ));
    InMux I__8632 (
            .O(N__50497),
            .I(N__50494));
    LocalMux I__8631 (
            .O(N__50494),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_1 ));
    CascadeMux I__8630 (
            .O(N__50491),
            .I(N__50488));
    InMux I__8629 (
            .O(N__50488),
            .I(N__50485));
    LocalMux I__8628 (
            .O(N__50485),
            .I(N__50482));
    Span4Mux_v I__8627 (
            .O(N__50482),
            .I(N__50479));
    Odrv4 I__8626 (
            .O(N__50479),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n8_adj_1152 ));
    InMux I__8625 (
            .O(N__50476),
            .I(bfn_12_16_0_));
    InMux I__8624 (
            .O(N__50473),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10619 ));
    CascadeMux I__8623 (
            .O(N__50470),
            .I(N__50467));
    InMux I__8622 (
            .O(N__50467),
            .I(N__50464));
    LocalMux I__8621 (
            .O(N__50464),
            .I(N__50461));
    Span4Mux_v I__8620 (
            .O(N__50461),
            .I(N__50458));
    Sp12to4 I__8619 (
            .O(N__50458),
            .I(N__50455));
    Odrv12 I__8618 (
            .O(N__50455),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n6_adj_1150 ));
    InMux I__8617 (
            .O(N__50452),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10620 ));
    InMux I__8616 (
            .O(N__50449),
            .I(N__50443));
    InMux I__8615 (
            .O(N__50448),
            .I(N__50443));
    LocalMux I__8614 (
            .O(N__50443),
            .I(N__50440));
    Span4Mux_v I__8613 (
            .O(N__50440),
            .I(N__50437));
    Span4Mux_h I__8612 (
            .O(N__50437),
            .I(N__50433));
    InMux I__8611 (
            .O(N__50436),
            .I(N__50430));
    Odrv4 I__8610 (
            .O(N__50433),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_3 ));
    LocalMux I__8609 (
            .O(N__50430),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_3 ));
    CascadeMux I__8608 (
            .O(N__50425),
            .I(N__50422));
    InMux I__8607 (
            .O(N__50422),
            .I(N__50419));
    LocalMux I__8606 (
            .O(N__50419),
            .I(N__50416));
    Span4Mux_v I__8605 (
            .O(N__50416),
            .I(N__50413));
    Span4Mux_h I__8604 (
            .O(N__50413),
            .I(N__50410));
    Odrv4 I__8603 (
            .O(N__50410),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n5 ));
    InMux I__8602 (
            .O(N__50407),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10621 ));
    InMux I__8601 (
            .O(N__50404),
            .I(N__50401));
    LocalMux I__8600 (
            .O(N__50401),
            .I(N__50398));
    Span4Mux_v I__8599 (
            .O(N__50398),
            .I(N__50395));
    Odrv4 I__8598 (
            .O(N__50395),
            .I(wr_grey_sync_r_4));
    InMux I__8597 (
            .O(N__50392),
            .I(N__50389));
    LocalMux I__8596 (
            .O(N__50389),
            .I(wp_sync1_r_4));
    InMux I__8595 (
            .O(N__50386),
            .I(N__50383));
    LocalMux I__8594 (
            .O(N__50383),
            .I(N__50380));
    Span4Mux_h I__8593 (
            .O(N__50380),
            .I(N__50377));
    Span4Mux_v I__8592 (
            .O(N__50377),
            .I(N__50374));
    Odrv4 I__8591 (
            .O(N__50374),
            .I(wr_grey_sync_r_3));
    InMux I__8590 (
            .O(N__50371),
            .I(N__50368));
    LocalMux I__8589 (
            .O(N__50368),
            .I(wp_sync1_r_3));
    InMux I__8588 (
            .O(N__50365),
            .I(N__50362));
    LocalMux I__8587 (
            .O(N__50362),
            .I(N__50359));
    Span4Mux_v I__8586 (
            .O(N__50359),
            .I(N__50356));
    Odrv4 I__8585 (
            .O(N__50356),
            .I(wr_grey_sync_r_5));
    InMux I__8584 (
            .O(N__50353),
            .I(N__50350));
    LocalMux I__8583 (
            .O(N__50350),
            .I(wp_sync1_r_5));
    CascadeMux I__8582 (
            .O(N__50347),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_4_cascade_ ));
    InMux I__8581 (
            .O(N__50344),
            .I(N__50341));
    LocalMux I__8580 (
            .O(N__50341),
            .I(N__50338));
    Span4Mux_v I__8579 (
            .O(N__50338),
            .I(N__50335));
    Sp12to4 I__8578 (
            .O(N__50335),
            .I(N__50332));
    Span12Mux_h I__8577 (
            .O(N__50332),
            .I(N__50329));
    Odrv12 I__8576 (
            .O(N__50329),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13157 ));
    CascadeMux I__8575 (
            .O(N__50326),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14318_cascade_ ));
    InMux I__8574 (
            .O(N__50323),
            .I(N__50320));
    LocalMux I__8573 (
            .O(N__50320),
            .I(N__50317));
    Span4Mux_v I__8572 (
            .O(N__50317),
            .I(N__50314));
    Span4Mux_v I__8571 (
            .O(N__50314),
            .I(N__50311));
    Odrv4 I__8570 (
            .O(N__50311),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12480 ));
    CascadeMux I__8569 (
            .O(N__50308),
            .I(N__50305));
    InMux I__8568 (
            .O(N__50305),
            .I(N__50302));
    LocalMux I__8567 (
            .O(N__50302),
            .I(N__50299));
    Span4Mux_v I__8566 (
            .O(N__50299),
            .I(N__50296));
    Span4Mux_v I__8565 (
            .O(N__50296),
            .I(N__50293));
    Span4Mux_v I__8564 (
            .O(N__50293),
            .I(N__50290));
    Odrv4 I__8563 (
            .O(N__50290),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14117 ));
    InMux I__8562 (
            .O(N__50287),
            .I(N__50284));
    LocalMux I__8561 (
            .O(N__50284),
            .I(N__50281));
    Span12Mux_v I__8560 (
            .O(N__50281),
            .I(N__50278));
    Odrv12 I__8559 (
            .O(N__50278),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13691 ));
    InMux I__8558 (
            .O(N__50275),
            .I(N__50272));
    LocalMux I__8557 (
            .O(N__50272),
            .I(N__50269));
    Span12Mux_v I__8556 (
            .O(N__50269),
            .I(N__50266));
    Odrv12 I__8555 (
            .O(N__50266),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13709 ));
    InMux I__8554 (
            .O(N__50263),
            .I(N__50260));
    LocalMux I__8553 (
            .O(N__50260),
            .I(N__50257));
    Span4Mux_v I__8552 (
            .O(N__50257),
            .I(N__50254));
    Span4Mux_v I__8551 (
            .O(N__50254),
            .I(N__50251));
    Odrv4 I__8550 (
            .O(N__50251),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14081 ));
    InMux I__8549 (
            .O(N__50248),
            .I(N__50245));
    LocalMux I__8548 (
            .O(N__50245),
            .I(N__50242));
    Span4Mux_h I__8547 (
            .O(N__50242),
            .I(N__50239));
    Span4Mux_h I__8546 (
            .O(N__50239),
            .I(N__50236));
    Span4Mux_v I__8545 (
            .O(N__50236),
            .I(N__50233));
    Odrv4 I__8544 (
            .O(N__50233),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14303 ));
    InMux I__8543 (
            .O(N__50230),
            .I(N__50227));
    LocalMux I__8542 (
            .O(N__50227),
            .I(N__50224));
    Span12Mux_h I__8541 (
            .O(N__50224),
            .I(N__50221));
    Odrv12 I__8540 (
            .O(N__50221),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13175 ));
    InMux I__8539 (
            .O(N__50218),
            .I(N__50215));
    LocalMux I__8538 (
            .O(N__50215),
            .I(N__50212));
    Span4Mux_v I__8537 (
            .O(N__50212),
            .I(N__50209));
    Span4Mux_h I__8536 (
            .O(N__50209),
            .I(N__50206));
    Span4Mux_h I__8535 (
            .O(N__50206),
            .I(N__50203));
    Odrv4 I__8534 (
            .O(N__50203),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13229 ));
    InMux I__8533 (
            .O(N__50200),
            .I(N__50197));
    LocalMux I__8532 (
            .O(N__50197),
            .I(N__50194));
    Span12Mux_h I__8531 (
            .O(N__50194),
            .I(N__50191));
    Odrv12 I__8530 (
            .O(N__50191),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13631 ));
    InMux I__8529 (
            .O(N__50188),
            .I(N__50185));
    LocalMux I__8528 (
            .O(N__50185),
            .I(N__50182));
    Sp12to4 I__8527 (
            .O(N__50182),
            .I(N__50179));
    Span12Mux_v I__8526 (
            .O(N__50179),
            .I(N__50176));
    Odrv12 I__8525 (
            .O(N__50176),
            .I(wr_grey_sync_r_1));
    InMux I__8524 (
            .O(N__50173),
            .I(N__50170));
    LocalMux I__8523 (
            .O(N__50170),
            .I(REG_out_raw_10));
    InMux I__8522 (
            .O(N__50167),
            .I(bfn_12_12_0_));
    InMux I__8521 (
            .O(N__50164),
            .I(N__50146));
    InMux I__8520 (
            .O(N__50163),
            .I(N__50146));
    InMux I__8519 (
            .O(N__50162),
            .I(N__50146));
    InMux I__8518 (
            .O(N__50161),
            .I(N__50146));
    CascadeMux I__8517 (
            .O(N__50160),
            .I(N__50143));
    InMux I__8516 (
            .O(N__50159),
            .I(N__50139));
    InMux I__8515 (
            .O(N__50158),
            .I(N__50134));
    InMux I__8514 (
            .O(N__50157),
            .I(N__50134));
    InMux I__8513 (
            .O(N__50156),
            .I(N__50131));
    InMux I__8512 (
            .O(N__50155),
            .I(N__50128));
    LocalMux I__8511 (
            .O(N__50146),
            .I(N__50125));
    InMux I__8510 (
            .O(N__50143),
            .I(N__50122));
    InMux I__8509 (
            .O(N__50142),
            .I(N__50119));
    LocalMux I__8508 (
            .O(N__50139),
            .I(N__50114));
    LocalMux I__8507 (
            .O(N__50134),
            .I(N__50114));
    LocalMux I__8506 (
            .O(N__50131),
            .I(N__50111));
    LocalMux I__8505 (
            .O(N__50128),
            .I(N__50104));
    Span4Mux_v I__8504 (
            .O(N__50125),
            .I(N__50104));
    LocalMux I__8503 (
            .O(N__50122),
            .I(N__50104));
    LocalMux I__8502 (
            .O(N__50119),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_1 ));
    Odrv4 I__8501 (
            .O(N__50114),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_1 ));
    Odrv4 I__8500 (
            .O(N__50111),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_1 ));
    Odrv4 I__8499 (
            .O(N__50104),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_1 ));
    CascadeMux I__8498 (
            .O(N__50095),
            .I(N__50092));
    InMux I__8497 (
            .O(N__50092),
            .I(N__50085));
    InMux I__8496 (
            .O(N__50091),
            .I(N__50085));
    CascadeMux I__8495 (
            .O(N__50090),
            .I(N__50081));
    LocalMux I__8494 (
            .O(N__50085),
            .I(N__50078));
    InMux I__8493 (
            .O(N__50084),
            .I(N__50075));
    InMux I__8492 (
            .O(N__50081),
            .I(N__50072));
    Span4Mux_h I__8491 (
            .O(N__50078),
            .I(N__50069));
    LocalMux I__8490 (
            .O(N__50075),
            .I(N__50064));
    LocalMux I__8489 (
            .O(N__50072),
            .I(N__50064));
    Odrv4 I__8488 (
            .O(N__50069),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_1 ));
    Odrv4 I__8487 (
            .O(N__50064),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_1 ));
    InMux I__8486 (
            .O(N__50059),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10631 ));
    CascadeMux I__8485 (
            .O(N__50056),
            .I(N__50050));
    CascadeMux I__8484 (
            .O(N__50055),
            .I(N__50047));
    CascadeMux I__8483 (
            .O(N__50054),
            .I(N__50044));
    CascadeMux I__8482 (
            .O(N__50053),
            .I(N__50030));
    InMux I__8481 (
            .O(N__50050),
            .I(N__50021));
    InMux I__8480 (
            .O(N__50047),
            .I(N__50018));
    InMux I__8479 (
            .O(N__50044),
            .I(N__50011));
    InMux I__8478 (
            .O(N__50043),
            .I(N__50011));
    InMux I__8477 (
            .O(N__50042),
            .I(N__50011));
    InMux I__8476 (
            .O(N__50041),
            .I(N__50002));
    InMux I__8475 (
            .O(N__50040),
            .I(N__50002));
    InMux I__8474 (
            .O(N__50039),
            .I(N__50002));
    InMux I__8473 (
            .O(N__50038),
            .I(N__50002));
    InMux I__8472 (
            .O(N__50037),
            .I(N__49993));
    InMux I__8471 (
            .O(N__50036),
            .I(N__49993));
    InMux I__8470 (
            .O(N__50035),
            .I(N__49993));
    InMux I__8469 (
            .O(N__50034),
            .I(N__49993));
    InMux I__8468 (
            .O(N__50033),
            .I(N__49986));
    InMux I__8467 (
            .O(N__50030),
            .I(N__49986));
    InMux I__8466 (
            .O(N__50029),
            .I(N__49986));
    InMux I__8465 (
            .O(N__50028),
            .I(N__49983));
    InMux I__8464 (
            .O(N__50027),
            .I(N__49978));
    InMux I__8463 (
            .O(N__50026),
            .I(N__49978));
    CascadeMux I__8462 (
            .O(N__50025),
            .I(N__49975));
    InMux I__8461 (
            .O(N__50024),
            .I(N__49972));
    LocalMux I__8460 (
            .O(N__50021),
            .I(N__49969));
    LocalMux I__8459 (
            .O(N__50018),
            .I(N__49958));
    LocalMux I__8458 (
            .O(N__50011),
            .I(N__49958));
    LocalMux I__8457 (
            .O(N__50002),
            .I(N__49958));
    LocalMux I__8456 (
            .O(N__49993),
            .I(N__49958));
    LocalMux I__8455 (
            .O(N__49986),
            .I(N__49958));
    LocalMux I__8454 (
            .O(N__49983),
            .I(N__49953));
    LocalMux I__8453 (
            .O(N__49978),
            .I(N__49953));
    InMux I__8452 (
            .O(N__49975),
            .I(N__49950));
    LocalMux I__8451 (
            .O(N__49972),
            .I(N__49947));
    Span4Mux_v I__8450 (
            .O(N__49969),
            .I(N__49942));
    Span4Mux_v I__8449 (
            .O(N__49958),
            .I(N__49942));
    Span4Mux_h I__8448 (
            .O(N__49953),
            .I(N__49938));
    LocalMux I__8447 (
            .O(N__49950),
            .I(N__49935));
    Span4Mux_h I__8446 (
            .O(N__49947),
            .I(N__49932));
    Span4Mux_h I__8445 (
            .O(N__49942),
            .I(N__49929));
    InMux I__8444 (
            .O(N__49941),
            .I(N__49926));
    Span4Mux_h I__8443 (
            .O(N__49938),
            .I(N__49921));
    Span4Mux_h I__8442 (
            .O(N__49935),
            .I(N__49921));
    Odrv4 I__8441 (
            .O(N__49932),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_2 ));
    Odrv4 I__8440 (
            .O(N__49929),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_2 ));
    LocalMux I__8439 (
            .O(N__49926),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_2 ));
    Odrv4 I__8438 (
            .O(N__49921),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_2 ));
    InMux I__8437 (
            .O(N__49912),
            .I(N__49908));
    CascadeMux I__8436 (
            .O(N__49911),
            .I(N__49905));
    LocalMux I__8435 (
            .O(N__49908),
            .I(N__49902));
    InMux I__8434 (
            .O(N__49905),
            .I(N__49899));
    Span4Mux_h I__8433 (
            .O(N__49902),
            .I(N__49896));
    LocalMux I__8432 (
            .O(N__49899),
            .I(N__49893));
    Odrv4 I__8431 (
            .O(N__49896),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_2 ));
    Odrv12 I__8430 (
            .O(N__49893),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_2 ));
    InMux I__8429 (
            .O(N__49888),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10632 ));
    CascadeMux I__8428 (
            .O(N__49885),
            .I(N__49879));
    InMux I__8427 (
            .O(N__49884),
            .I(N__49871));
    InMux I__8426 (
            .O(N__49883),
            .I(N__49871));
    InMux I__8425 (
            .O(N__49882),
            .I(N__49860));
    InMux I__8424 (
            .O(N__49879),
            .I(N__49860));
    InMux I__8423 (
            .O(N__49878),
            .I(N__49860));
    InMux I__8422 (
            .O(N__49877),
            .I(N__49860));
    InMux I__8421 (
            .O(N__49876),
            .I(N__49860));
    LocalMux I__8420 (
            .O(N__49871),
            .I(N__49851));
    LocalMux I__8419 (
            .O(N__49860),
            .I(N__49851));
    CascadeMux I__8418 (
            .O(N__49859),
            .I(N__49847));
    CascadeMux I__8417 (
            .O(N__49858),
            .I(N__49842));
    InMux I__8416 (
            .O(N__49857),
            .I(N__49832));
    InMux I__8415 (
            .O(N__49856),
            .I(N__49832));
    Span4Mux_v I__8414 (
            .O(N__49851),
            .I(N__49828));
    InMux I__8413 (
            .O(N__49850),
            .I(N__49817));
    InMux I__8412 (
            .O(N__49847),
            .I(N__49817));
    InMux I__8411 (
            .O(N__49846),
            .I(N__49817));
    InMux I__8410 (
            .O(N__49845),
            .I(N__49817));
    InMux I__8409 (
            .O(N__49842),
            .I(N__49817));
    CascadeMux I__8408 (
            .O(N__49841),
            .I(N__49812));
    CascadeMux I__8407 (
            .O(N__49840),
            .I(N__49801));
    CascadeMux I__8406 (
            .O(N__49839),
            .I(N__49789));
    CascadeMux I__8405 (
            .O(N__49838),
            .I(N__49786));
    CascadeMux I__8404 (
            .O(N__49837),
            .I(N__49779));
    LocalMux I__8403 (
            .O(N__49832),
            .I(N__49776));
    InMux I__8402 (
            .O(N__49831),
            .I(N__49773));
    Span4Mux_v I__8401 (
            .O(N__49828),
            .I(N__49768));
    LocalMux I__8400 (
            .O(N__49817),
            .I(N__49768));
    InMux I__8399 (
            .O(N__49816),
            .I(N__49765));
    InMux I__8398 (
            .O(N__49815),
            .I(N__49750));
    InMux I__8397 (
            .O(N__49812),
            .I(N__49750));
    InMux I__8396 (
            .O(N__49811),
            .I(N__49750));
    InMux I__8395 (
            .O(N__49810),
            .I(N__49750));
    InMux I__8394 (
            .O(N__49809),
            .I(N__49750));
    InMux I__8393 (
            .O(N__49808),
            .I(N__49750));
    InMux I__8392 (
            .O(N__49807),
            .I(N__49750));
    InMux I__8391 (
            .O(N__49806),
            .I(N__49743));
    InMux I__8390 (
            .O(N__49805),
            .I(N__49743));
    InMux I__8389 (
            .O(N__49804),
            .I(N__49743));
    InMux I__8388 (
            .O(N__49801),
            .I(N__49736));
    InMux I__8387 (
            .O(N__49800),
            .I(N__49736));
    InMux I__8386 (
            .O(N__49799),
            .I(N__49736));
    InMux I__8385 (
            .O(N__49798),
            .I(N__49733));
    InMux I__8384 (
            .O(N__49797),
            .I(N__49724));
    InMux I__8383 (
            .O(N__49796),
            .I(N__49724));
    InMux I__8382 (
            .O(N__49795),
            .I(N__49724));
    InMux I__8381 (
            .O(N__49794),
            .I(N__49724));
    InMux I__8380 (
            .O(N__49793),
            .I(N__49709));
    InMux I__8379 (
            .O(N__49792),
            .I(N__49709));
    InMux I__8378 (
            .O(N__49789),
            .I(N__49709));
    InMux I__8377 (
            .O(N__49786),
            .I(N__49709));
    InMux I__8376 (
            .O(N__49785),
            .I(N__49709));
    InMux I__8375 (
            .O(N__49784),
            .I(N__49709));
    InMux I__8374 (
            .O(N__49783),
            .I(N__49709));
    InMux I__8373 (
            .O(N__49782),
            .I(N__49706));
    InMux I__8372 (
            .O(N__49779),
            .I(N__49703));
    Span4Mux_h I__8371 (
            .O(N__49776),
            .I(N__49694));
    LocalMux I__8370 (
            .O(N__49773),
            .I(N__49694));
    Span4Mux_v I__8369 (
            .O(N__49768),
            .I(N__49694));
    LocalMux I__8368 (
            .O(N__49765),
            .I(N__49689));
    LocalMux I__8367 (
            .O(N__49750),
            .I(N__49689));
    LocalMux I__8366 (
            .O(N__49743),
            .I(N__49680));
    LocalMux I__8365 (
            .O(N__49736),
            .I(N__49680));
    LocalMux I__8364 (
            .O(N__49733),
            .I(N__49680));
    LocalMux I__8363 (
            .O(N__49724),
            .I(N__49680));
    LocalMux I__8362 (
            .O(N__49709),
            .I(N__49676));
    LocalMux I__8361 (
            .O(N__49706),
            .I(N__49671));
    LocalMux I__8360 (
            .O(N__49703),
            .I(N__49671));
    InMux I__8359 (
            .O(N__49702),
            .I(N__49668));
    InMux I__8358 (
            .O(N__49701),
            .I(N__49665));
    Span4Mux_h I__8357 (
            .O(N__49694),
            .I(N__49662));
    Span4Mux_v I__8356 (
            .O(N__49689),
            .I(N__49657));
    Span4Mux_v I__8355 (
            .O(N__49680),
            .I(N__49657));
    InMux I__8354 (
            .O(N__49679),
            .I(N__49654));
    Span4Mux_v I__8353 (
            .O(N__49676),
            .I(N__49649));
    Span4Mux_h I__8352 (
            .O(N__49671),
            .I(N__49649));
    LocalMux I__8351 (
            .O(N__49668),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_3 ));
    LocalMux I__8350 (
            .O(N__49665),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_3 ));
    Odrv4 I__8349 (
            .O(N__49662),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_3 ));
    Odrv4 I__8348 (
            .O(N__49657),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_3 ));
    LocalMux I__8347 (
            .O(N__49654),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_3 ));
    Odrv4 I__8346 (
            .O(N__49649),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_3 ));
    CascadeMux I__8345 (
            .O(N__49636),
            .I(N__49633));
    InMux I__8344 (
            .O(N__49633),
            .I(N__49626));
    InMux I__8343 (
            .O(N__49632),
            .I(N__49626));
    InMux I__8342 (
            .O(N__49631),
            .I(N__49623));
    LocalMux I__8341 (
            .O(N__49626),
            .I(N__49620));
    LocalMux I__8340 (
            .O(N__49623),
            .I(N__49616));
    Span4Mux_h I__8339 (
            .O(N__49620),
            .I(N__49613));
    InMux I__8338 (
            .O(N__49619),
            .I(N__49610));
    Span4Mux_h I__8337 (
            .O(N__49616),
            .I(N__49607));
    Odrv4 I__8336 (
            .O(N__49613),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_3 ));
    LocalMux I__8335 (
            .O(N__49610),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_3 ));
    Odrv4 I__8334 (
            .O(N__49607),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_3 ));
    InMux I__8333 (
            .O(N__49600),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10633 ));
    CascadeMux I__8332 (
            .O(N__49597),
            .I(N__49586));
    CascadeMux I__8331 (
            .O(N__49596),
            .I(N__49583));
    CascadeMux I__8330 (
            .O(N__49595),
            .I(N__49576));
    CascadeMux I__8329 (
            .O(N__49594),
            .I(N__49573));
    InMux I__8328 (
            .O(N__49593),
            .I(N__49565));
    InMux I__8327 (
            .O(N__49592),
            .I(N__49562));
    CascadeMux I__8326 (
            .O(N__49591),
            .I(N__49559));
    CascadeMux I__8325 (
            .O(N__49590),
            .I(N__49556));
    CascadeMux I__8324 (
            .O(N__49589),
            .I(N__49550));
    InMux I__8323 (
            .O(N__49586),
            .I(N__49528));
    InMux I__8322 (
            .O(N__49583),
            .I(N__49528));
    InMux I__8321 (
            .O(N__49582),
            .I(N__49528));
    InMux I__8320 (
            .O(N__49581),
            .I(N__49528));
    CascadeMux I__8319 (
            .O(N__49580),
            .I(N__49524));
    CascadeMux I__8318 (
            .O(N__49579),
            .I(N__49520));
    InMux I__8317 (
            .O(N__49576),
            .I(N__49516));
    InMux I__8316 (
            .O(N__49573),
            .I(N__49513));
    CascadeMux I__8315 (
            .O(N__49572),
            .I(N__49506));
    CascadeMux I__8314 (
            .O(N__49571),
            .I(N__49503));
    InMux I__8313 (
            .O(N__49570),
            .I(N__49493));
    InMux I__8312 (
            .O(N__49569),
            .I(N__49493));
    InMux I__8311 (
            .O(N__49568),
            .I(N__49493));
    LocalMux I__8310 (
            .O(N__49565),
            .I(N__49488));
    LocalMux I__8309 (
            .O(N__49562),
            .I(N__49488));
    InMux I__8308 (
            .O(N__49559),
            .I(N__49485));
    InMux I__8307 (
            .O(N__49556),
            .I(N__49482));
    InMux I__8306 (
            .O(N__49555),
            .I(N__49467));
    InMux I__8305 (
            .O(N__49554),
            .I(N__49467));
    InMux I__8304 (
            .O(N__49553),
            .I(N__49467));
    InMux I__8303 (
            .O(N__49550),
            .I(N__49467));
    InMux I__8302 (
            .O(N__49549),
            .I(N__49456));
    InMux I__8301 (
            .O(N__49548),
            .I(N__49456));
    InMux I__8300 (
            .O(N__49547),
            .I(N__49456));
    InMux I__8299 (
            .O(N__49546),
            .I(N__49456));
    InMux I__8298 (
            .O(N__49545),
            .I(N__49456));
    InMux I__8297 (
            .O(N__49544),
            .I(N__49449));
    InMux I__8296 (
            .O(N__49543),
            .I(N__49449));
    InMux I__8295 (
            .O(N__49542),
            .I(N__49449));
    InMux I__8294 (
            .O(N__49541),
            .I(N__49435));
    InMux I__8293 (
            .O(N__49540),
            .I(N__49435));
    InMux I__8292 (
            .O(N__49539),
            .I(N__49435));
    InMux I__8291 (
            .O(N__49538),
            .I(N__49435));
    InMux I__8290 (
            .O(N__49537),
            .I(N__49435));
    LocalMux I__8289 (
            .O(N__49528),
            .I(N__49432));
    InMux I__8288 (
            .O(N__49527),
            .I(N__49423));
    InMux I__8287 (
            .O(N__49524),
            .I(N__49423));
    InMux I__8286 (
            .O(N__49523),
            .I(N__49423));
    InMux I__8285 (
            .O(N__49520),
            .I(N__49423));
    InMux I__8284 (
            .O(N__49519),
            .I(N__49420));
    LocalMux I__8283 (
            .O(N__49516),
            .I(N__49415));
    LocalMux I__8282 (
            .O(N__49513),
            .I(N__49415));
    InMux I__8281 (
            .O(N__49512),
            .I(N__49408));
    InMux I__8280 (
            .O(N__49511),
            .I(N__49408));
    InMux I__8279 (
            .O(N__49510),
            .I(N__49408));
    InMux I__8278 (
            .O(N__49509),
            .I(N__49394));
    InMux I__8277 (
            .O(N__49506),
            .I(N__49394));
    InMux I__8276 (
            .O(N__49503),
            .I(N__49394));
    InMux I__8275 (
            .O(N__49502),
            .I(N__49394));
    InMux I__8274 (
            .O(N__49501),
            .I(N__49394));
    InMux I__8273 (
            .O(N__49500),
            .I(N__49394));
    LocalMux I__8272 (
            .O(N__49493),
            .I(N__49389));
    Span4Mux_h I__8271 (
            .O(N__49488),
            .I(N__49389));
    LocalMux I__8270 (
            .O(N__49485),
            .I(N__49384));
    LocalMux I__8269 (
            .O(N__49482),
            .I(N__49384));
    InMux I__8268 (
            .O(N__49481),
            .I(N__49371));
    InMux I__8267 (
            .O(N__49480),
            .I(N__49371));
    InMux I__8266 (
            .O(N__49479),
            .I(N__49371));
    InMux I__8265 (
            .O(N__49478),
            .I(N__49371));
    InMux I__8264 (
            .O(N__49477),
            .I(N__49371));
    InMux I__8263 (
            .O(N__49476),
            .I(N__49371));
    LocalMux I__8262 (
            .O(N__49467),
            .I(N__49366));
    LocalMux I__8261 (
            .O(N__49456),
            .I(N__49366));
    LocalMux I__8260 (
            .O(N__49449),
            .I(N__49363));
    InMux I__8259 (
            .O(N__49448),
            .I(N__49356));
    InMux I__8258 (
            .O(N__49447),
            .I(N__49356));
    InMux I__8257 (
            .O(N__49446),
            .I(N__49356));
    LocalMux I__8256 (
            .O(N__49435),
            .I(N__49349));
    Span4Mux_v I__8255 (
            .O(N__49432),
            .I(N__49349));
    LocalMux I__8254 (
            .O(N__49423),
            .I(N__49349));
    LocalMux I__8253 (
            .O(N__49420),
            .I(N__49342));
    Span4Mux_h I__8252 (
            .O(N__49415),
            .I(N__49342));
    LocalMux I__8251 (
            .O(N__49408),
            .I(N__49342));
    InMux I__8250 (
            .O(N__49407),
            .I(N__49338));
    LocalMux I__8249 (
            .O(N__49394),
            .I(N__49333));
    Span4Mux_v I__8248 (
            .O(N__49389),
            .I(N__49333));
    Span4Mux_h I__8247 (
            .O(N__49384),
            .I(N__49330));
    LocalMux I__8246 (
            .O(N__49371),
            .I(N__49323));
    Span4Mux_h I__8245 (
            .O(N__49366),
            .I(N__49323));
    Span4Mux_h I__8244 (
            .O(N__49363),
            .I(N__49323));
    LocalMux I__8243 (
            .O(N__49356),
            .I(N__49318));
    Span4Mux_h I__8242 (
            .O(N__49349),
            .I(N__49318));
    Span4Mux_h I__8241 (
            .O(N__49342),
            .I(N__49315));
    InMux I__8240 (
            .O(N__49341),
            .I(N__49312));
    LocalMux I__8239 (
            .O(N__49338),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_4 ));
    Odrv4 I__8238 (
            .O(N__49333),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_4 ));
    Odrv4 I__8237 (
            .O(N__49330),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_4 ));
    Odrv4 I__8236 (
            .O(N__49323),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_4 ));
    Odrv4 I__8235 (
            .O(N__49318),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_4 ));
    Odrv4 I__8234 (
            .O(N__49315),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_4 ));
    LocalMux I__8233 (
            .O(N__49312),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_4 ));
    InMux I__8232 (
            .O(N__49297),
            .I(N__49293));
    InMux I__8231 (
            .O(N__49296),
            .I(N__49290));
    LocalMux I__8230 (
            .O(N__49293),
            .I(N__49287));
    LocalMux I__8229 (
            .O(N__49290),
            .I(N__49284));
    Odrv4 I__8228 (
            .O(N__49287),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_4 ));
    Odrv4 I__8227 (
            .O(N__49284),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_4 ));
    InMux I__8226 (
            .O(N__49279),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10634 ));
    InMux I__8225 (
            .O(N__49276),
            .I(N__49271));
    InMux I__8224 (
            .O(N__49275),
            .I(N__49265));
    InMux I__8223 (
            .O(N__49274),
            .I(N__49265));
    LocalMux I__8222 (
            .O(N__49271),
            .I(N__49262));
    InMux I__8221 (
            .O(N__49270),
            .I(N__49259));
    LocalMux I__8220 (
            .O(N__49265),
            .I(N__49256));
    Span4Mux_h I__8219 (
            .O(N__49262),
            .I(N__49253));
    LocalMux I__8218 (
            .O(N__49259),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_5 ));
    Odrv4 I__8217 (
            .O(N__49256),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_5 ));
    Odrv4 I__8216 (
            .O(N__49253),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_5 ));
    InMux I__8215 (
            .O(N__49246),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10635 ));
    InMux I__8214 (
            .O(N__49243),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10636 ));
    InMux I__8213 (
            .O(N__49240),
            .I(N__49235));
    InMux I__8212 (
            .O(N__49239),
            .I(N__49230));
    InMux I__8211 (
            .O(N__49238),
            .I(N__49230));
    LocalMux I__8210 (
            .O(N__49235),
            .I(N__49225));
    LocalMux I__8209 (
            .O(N__49230),
            .I(N__49225));
    Odrv4 I__8208 (
            .O(N__49225),
            .I(wr_addr_p1_w_6));
    InMux I__8207 (
            .O(N__49222),
            .I(N__49219));
    LocalMux I__8206 (
            .O(N__49219),
            .I(N__49216));
    Span4Mux_v I__8205 (
            .O(N__49216),
            .I(N__49213));
    Sp12to4 I__8204 (
            .O(N__49213),
            .I(N__49210));
    Odrv12 I__8203 (
            .O(N__49210),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13301 ));
    InMux I__8202 (
            .O(N__49207),
            .I(N__49204));
    LocalMux I__8201 (
            .O(N__49204),
            .I(N__49201));
    Span4Mux_v I__8200 (
            .O(N__49201),
            .I(N__49198));
    Span4Mux_h I__8199 (
            .O(N__49198),
            .I(N__49195));
    Span4Mux_h I__8198 (
            .O(N__49195),
            .I(N__49192));
    Odrv4 I__8197 (
            .O(N__49192),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14231 ));
    InMux I__8196 (
            .O(N__49189),
            .I(N__49186));
    LocalMux I__8195 (
            .O(N__49186),
            .I(N__49183));
    Odrv12 I__8194 (
            .O(N__49183),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12486 ));
    CascadeMux I__8193 (
            .O(N__49180),
            .I(N__49177));
    InMux I__8192 (
            .O(N__49177),
            .I(N__49174));
    LocalMux I__8191 (
            .O(N__49174),
            .I(N__49171));
    Span4Mux_v I__8190 (
            .O(N__49171),
            .I(N__49168));
    Span4Mux_v I__8189 (
            .O(N__49168),
            .I(N__49165));
    Odrv4 I__8188 (
            .O(N__49165),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12498 ));
    InMux I__8187 (
            .O(N__49162),
            .I(N__49158));
    InMux I__8186 (
            .O(N__49161),
            .I(N__49155));
    LocalMux I__8185 (
            .O(N__49158),
            .I(REG_mem_15_3));
    LocalMux I__8184 (
            .O(N__49155),
            .I(REG_mem_15_3));
    InMux I__8183 (
            .O(N__49150),
            .I(N__49141));
    InMux I__8182 (
            .O(N__49149),
            .I(N__49141));
    InMux I__8181 (
            .O(N__49148),
            .I(N__49141));
    LocalMux I__8180 (
            .O(N__49141),
            .I(N__49135));
    InMux I__8179 (
            .O(N__49140),
            .I(N__49128));
    InMux I__8178 (
            .O(N__49139),
            .I(N__49128));
    InMux I__8177 (
            .O(N__49138),
            .I(N__49128));
    Span4Mux_v I__8176 (
            .O(N__49135),
            .I(N__49112));
    LocalMux I__8175 (
            .O(N__49128),
            .I(N__49112));
    InMux I__8174 (
            .O(N__49127),
            .I(N__49095));
    InMux I__8173 (
            .O(N__49126),
            .I(N__49095));
    InMux I__8172 (
            .O(N__49125),
            .I(N__49095));
    InMux I__8171 (
            .O(N__49124),
            .I(N__49095));
    InMux I__8170 (
            .O(N__49123),
            .I(N__49095));
    InMux I__8169 (
            .O(N__49122),
            .I(N__49095));
    InMux I__8168 (
            .O(N__49121),
            .I(N__49095));
    InMux I__8167 (
            .O(N__49120),
            .I(N__49095));
    InMux I__8166 (
            .O(N__49119),
            .I(N__49090));
    InMux I__8165 (
            .O(N__49118),
            .I(N__49090));
    InMux I__8164 (
            .O(N__49117),
            .I(N__49087));
    Span4Mux_h I__8163 (
            .O(N__49112),
            .I(N__49084));
    LocalMux I__8162 (
            .O(N__49095),
            .I(N__49081));
    LocalMux I__8161 (
            .O(N__49090),
            .I(n7596));
    LocalMux I__8160 (
            .O(N__49087),
            .I(n7596));
    Odrv4 I__8159 (
            .O(N__49084),
            .I(n7596));
    Odrv12 I__8158 (
            .O(N__49081),
            .I(n7596));
    InMux I__8157 (
            .O(N__49072),
            .I(N__49069));
    LocalMux I__8156 (
            .O(N__49069),
            .I(N__49065));
    InMux I__8155 (
            .O(N__49068),
            .I(N__49062));
    Span4Mux_h I__8154 (
            .O(N__49065),
            .I(N__49059));
    LocalMux I__8153 (
            .O(N__49062),
            .I(wr_addr_nxt_c_2));
    Odrv4 I__8152 (
            .O(N__49059),
            .I(wr_addr_nxt_c_2));
    InMux I__8151 (
            .O(N__49054),
            .I(N__49051));
    LocalMux I__8150 (
            .O(N__49051),
            .I(N__49048));
    Span12Mux_h I__8149 (
            .O(N__49048),
            .I(N__49044));
    InMux I__8148 (
            .O(N__49047),
            .I(N__49041));
    Odrv12 I__8147 (
            .O(N__49044),
            .I(wr_addr_nxt_c_4));
    LocalMux I__8146 (
            .O(N__49041),
            .I(wr_addr_nxt_c_4));
    CascadeMux I__8145 (
            .O(N__49036),
            .I(N__49031));
    InMux I__8144 (
            .O(N__49035),
            .I(N__49021));
    InMux I__8143 (
            .O(N__49034),
            .I(N__49021));
    InMux I__8142 (
            .O(N__49031),
            .I(N__49021));
    CascadeMux I__8141 (
            .O(N__49030),
            .I(N__49017));
    CascadeMux I__8140 (
            .O(N__49029),
            .I(N__49013));
    InMux I__8139 (
            .O(N__49028),
            .I(N__49010));
    LocalMux I__8138 (
            .O(N__49021),
            .I(N__49007));
    InMux I__8137 (
            .O(N__49020),
            .I(N__49003));
    InMux I__8136 (
            .O(N__49017),
            .I(N__48998));
    InMux I__8135 (
            .O(N__49016),
            .I(N__48998));
    InMux I__8134 (
            .O(N__49013),
            .I(N__48995));
    LocalMux I__8133 (
            .O(N__49010),
            .I(N__48992));
    Span4Mux_h I__8132 (
            .O(N__49007),
            .I(N__48989));
    InMux I__8131 (
            .O(N__49006),
            .I(N__48986));
    LocalMux I__8130 (
            .O(N__49003),
            .I(N__48983));
    LocalMux I__8129 (
            .O(N__48998),
            .I(N__48979));
    LocalMux I__8128 (
            .O(N__48995),
            .I(N__48976));
    Span4Mux_h I__8127 (
            .O(N__48992),
            .I(N__48971));
    Span4Mux_h I__8126 (
            .O(N__48989),
            .I(N__48971));
    LocalMux I__8125 (
            .O(N__48986),
            .I(N__48966));
    Span4Mux_v I__8124 (
            .O(N__48983),
            .I(N__48966));
    InMux I__8123 (
            .O(N__48982),
            .I(N__48963));
    Span4Mux_h I__8122 (
            .O(N__48979),
            .I(N__48958));
    Span4Mux_h I__8121 (
            .O(N__48976),
            .I(N__48958));
    Odrv4 I__8120 (
            .O(N__48971),
            .I(wr_addr_r_0));
    Odrv4 I__8119 (
            .O(N__48966),
            .I(wr_addr_r_0));
    LocalMux I__8118 (
            .O(N__48963),
            .I(wr_addr_r_0));
    Odrv4 I__8117 (
            .O(N__48958),
            .I(wr_addr_r_0));
    InMux I__8116 (
            .O(N__48949),
            .I(N__48946));
    LocalMux I__8115 (
            .O(N__48946),
            .I(N__48942));
    InMux I__8114 (
            .O(N__48945),
            .I(N__48939));
    Span4Mux_h I__8113 (
            .O(N__48942),
            .I(N__48935));
    LocalMux I__8112 (
            .O(N__48939),
            .I(N__48932));
    InMux I__8111 (
            .O(N__48938),
            .I(N__48929));
    Span4Mux_v I__8110 (
            .O(N__48935),
            .I(N__48924));
    Span4Mux_h I__8109 (
            .O(N__48932),
            .I(N__48924));
    LocalMux I__8108 (
            .O(N__48929),
            .I(wr_addr_p1_w_0));
    Odrv4 I__8107 (
            .O(N__48924),
            .I(wr_addr_p1_w_0));
    InMux I__8106 (
            .O(N__48919),
            .I(N__48916));
    LocalMux I__8105 (
            .O(N__48916),
            .I(N__48913));
    Span4Mux_v I__8104 (
            .O(N__48913),
            .I(N__48910));
    Span4Mux_h I__8103 (
            .O(N__48910),
            .I(N__48906));
    InMux I__8102 (
            .O(N__48909),
            .I(N__48903));
    Odrv4 I__8101 (
            .O(N__48906),
            .I(REG_mem_15_15));
    LocalMux I__8100 (
            .O(N__48903),
            .I(REG_mem_15_15));
    InMux I__8099 (
            .O(N__48898),
            .I(N__48886));
    InMux I__8098 (
            .O(N__48897),
            .I(N__48886));
    InMux I__8097 (
            .O(N__48896),
            .I(N__48883));
    InMux I__8096 (
            .O(N__48895),
            .I(N__48862));
    CascadeMux I__8095 (
            .O(N__48894),
            .I(N__48859));
    CascadeMux I__8094 (
            .O(N__48893),
            .I(N__48856));
    InMux I__8093 (
            .O(N__48892),
            .I(N__48847));
    InMux I__8092 (
            .O(N__48891),
            .I(N__48843));
    LocalMux I__8091 (
            .O(N__48886),
            .I(N__48837));
    LocalMux I__8090 (
            .O(N__48883),
            .I(N__48837));
    InMux I__8089 (
            .O(N__48882),
            .I(N__48832));
    InMux I__8088 (
            .O(N__48881),
            .I(N__48832));
    InMux I__8087 (
            .O(N__48880),
            .I(N__48823));
    InMux I__8086 (
            .O(N__48879),
            .I(N__48823));
    InMux I__8085 (
            .O(N__48878),
            .I(N__48823));
    InMux I__8084 (
            .O(N__48877),
            .I(N__48823));
    InMux I__8083 (
            .O(N__48876),
            .I(N__48814));
    InMux I__8082 (
            .O(N__48875),
            .I(N__48814));
    InMux I__8081 (
            .O(N__48874),
            .I(N__48814));
    InMux I__8080 (
            .O(N__48873),
            .I(N__48814));
    InMux I__8079 (
            .O(N__48872),
            .I(N__48799));
    InMux I__8078 (
            .O(N__48871),
            .I(N__48799));
    InMux I__8077 (
            .O(N__48870),
            .I(N__48799));
    InMux I__8076 (
            .O(N__48869),
            .I(N__48799));
    InMux I__8075 (
            .O(N__48868),
            .I(N__48799));
    InMux I__8074 (
            .O(N__48867),
            .I(N__48796));
    InMux I__8073 (
            .O(N__48866),
            .I(N__48791));
    InMux I__8072 (
            .O(N__48865),
            .I(N__48791));
    LocalMux I__8071 (
            .O(N__48862),
            .I(N__48788));
    InMux I__8070 (
            .O(N__48859),
            .I(N__48777));
    InMux I__8069 (
            .O(N__48856),
            .I(N__48777));
    InMux I__8068 (
            .O(N__48855),
            .I(N__48777));
    InMux I__8067 (
            .O(N__48854),
            .I(N__48777));
    InMux I__8066 (
            .O(N__48853),
            .I(N__48777));
    InMux I__8065 (
            .O(N__48852),
            .I(N__48770));
    InMux I__8064 (
            .O(N__48851),
            .I(N__48770));
    InMux I__8063 (
            .O(N__48850),
            .I(N__48770));
    LocalMux I__8062 (
            .O(N__48847),
            .I(N__48756));
    InMux I__8061 (
            .O(N__48846),
            .I(N__48752));
    LocalMux I__8060 (
            .O(N__48843),
            .I(N__48748));
    InMux I__8059 (
            .O(N__48842),
            .I(N__48745));
    Span4Mux_v I__8058 (
            .O(N__48837),
            .I(N__48735));
    LocalMux I__8057 (
            .O(N__48832),
            .I(N__48735));
    LocalMux I__8056 (
            .O(N__48823),
            .I(N__48735));
    LocalMux I__8055 (
            .O(N__48814),
            .I(N__48735));
    InMux I__8054 (
            .O(N__48813),
            .I(N__48726));
    InMux I__8053 (
            .O(N__48812),
            .I(N__48726));
    InMux I__8052 (
            .O(N__48811),
            .I(N__48722));
    InMux I__8051 (
            .O(N__48810),
            .I(N__48719));
    LocalMux I__8050 (
            .O(N__48799),
            .I(N__48712));
    LocalMux I__8049 (
            .O(N__48796),
            .I(N__48712));
    LocalMux I__8048 (
            .O(N__48791),
            .I(N__48712));
    Span4Mux_v I__8047 (
            .O(N__48788),
            .I(N__48705));
    LocalMux I__8046 (
            .O(N__48777),
            .I(N__48700));
    LocalMux I__8045 (
            .O(N__48770),
            .I(N__48700));
    InMux I__8044 (
            .O(N__48769),
            .I(N__48697));
    InMux I__8043 (
            .O(N__48768),
            .I(N__48694));
    InMux I__8042 (
            .O(N__48767),
            .I(N__48685));
    InMux I__8041 (
            .O(N__48766),
            .I(N__48685));
    InMux I__8040 (
            .O(N__48765),
            .I(N__48685));
    InMux I__8039 (
            .O(N__48764),
            .I(N__48676));
    InMux I__8038 (
            .O(N__48763),
            .I(N__48676));
    InMux I__8037 (
            .O(N__48762),
            .I(N__48676));
    InMux I__8036 (
            .O(N__48761),
            .I(N__48676));
    InMux I__8035 (
            .O(N__48760),
            .I(N__48673));
    InMux I__8034 (
            .O(N__48759),
            .I(N__48670));
    Span4Mux_h I__8033 (
            .O(N__48756),
            .I(N__48667));
    InMux I__8032 (
            .O(N__48755),
            .I(N__48664));
    LocalMux I__8031 (
            .O(N__48752),
            .I(N__48661));
    InMux I__8030 (
            .O(N__48751),
            .I(N__48658));
    Span4Mux_h I__8029 (
            .O(N__48748),
            .I(N__48655));
    LocalMux I__8028 (
            .O(N__48745),
            .I(N__48652));
    InMux I__8027 (
            .O(N__48744),
            .I(N__48649));
    Span4Mux_v I__8026 (
            .O(N__48735),
            .I(N__48645));
    InMux I__8025 (
            .O(N__48734),
            .I(N__48638));
    InMux I__8024 (
            .O(N__48733),
            .I(N__48638));
    InMux I__8023 (
            .O(N__48732),
            .I(N__48638));
    InMux I__8022 (
            .O(N__48731),
            .I(N__48635));
    LocalMux I__8021 (
            .O(N__48726),
            .I(N__48632));
    InMux I__8020 (
            .O(N__48725),
            .I(N__48629));
    LocalMux I__8019 (
            .O(N__48722),
            .I(N__48626));
    LocalMux I__8018 (
            .O(N__48719),
            .I(N__48621));
    Span4Mux_v I__8017 (
            .O(N__48712),
            .I(N__48621));
    InMux I__8016 (
            .O(N__48711),
            .I(N__48616));
    InMux I__8015 (
            .O(N__48710),
            .I(N__48616));
    InMux I__8014 (
            .O(N__48709),
            .I(N__48613));
    InMux I__8013 (
            .O(N__48708),
            .I(N__48610));
    Sp12to4 I__8012 (
            .O(N__48705),
            .I(N__48603));
    Span12Mux_h I__8011 (
            .O(N__48700),
            .I(N__48603));
    LocalMux I__8010 (
            .O(N__48697),
            .I(N__48603));
    LocalMux I__8009 (
            .O(N__48694),
            .I(N__48600));
    InMux I__8008 (
            .O(N__48693),
            .I(N__48597));
    InMux I__8007 (
            .O(N__48692),
            .I(N__48594));
    LocalMux I__8006 (
            .O(N__48685),
            .I(N__48589));
    LocalMux I__8005 (
            .O(N__48676),
            .I(N__48589));
    LocalMux I__8004 (
            .O(N__48673),
            .I(N__48584));
    LocalMux I__8003 (
            .O(N__48670),
            .I(N__48584));
    Span4Mux_v I__8002 (
            .O(N__48667),
            .I(N__48579));
    LocalMux I__8001 (
            .O(N__48664),
            .I(N__48579));
    Span4Mux_h I__8000 (
            .O(N__48661),
            .I(N__48568));
    LocalMux I__7999 (
            .O(N__48658),
            .I(N__48568));
    Span4Mux_h I__7998 (
            .O(N__48655),
            .I(N__48568));
    Span4Mux_h I__7997 (
            .O(N__48652),
            .I(N__48568));
    LocalMux I__7996 (
            .O(N__48649),
            .I(N__48568));
    InMux I__7995 (
            .O(N__48648),
            .I(N__48565));
    Span4Mux_h I__7994 (
            .O(N__48645),
            .I(N__48558));
    LocalMux I__7993 (
            .O(N__48638),
            .I(N__48558));
    LocalMux I__7992 (
            .O(N__48635),
            .I(N__48558));
    Span4Mux_v I__7991 (
            .O(N__48632),
            .I(N__48553));
    LocalMux I__7990 (
            .O(N__48629),
            .I(N__48553));
    Span4Mux_h I__7989 (
            .O(N__48626),
            .I(N__48542));
    Span4Mux_h I__7988 (
            .O(N__48621),
            .I(N__48542));
    LocalMux I__7987 (
            .O(N__48616),
            .I(N__48542));
    LocalMux I__7986 (
            .O(N__48613),
            .I(N__48542));
    LocalMux I__7985 (
            .O(N__48610),
            .I(N__48542));
    Span12Mux_v I__7984 (
            .O(N__48603),
            .I(N__48539));
    Span4Mux_v I__7983 (
            .O(N__48600),
            .I(N__48536));
    LocalMux I__7982 (
            .O(N__48597),
            .I(N__48521));
    LocalMux I__7981 (
            .O(N__48594),
            .I(N__48521));
    Span12Mux_v I__7980 (
            .O(N__48589),
            .I(N__48521));
    Span12Mux_h I__7979 (
            .O(N__48584),
            .I(N__48521));
    Sp12to4 I__7978 (
            .O(N__48579),
            .I(N__48521));
    Sp12to4 I__7977 (
            .O(N__48568),
            .I(N__48521));
    LocalMux I__7976 (
            .O(N__48565),
            .I(N__48521));
    Span4Mux_v I__7975 (
            .O(N__48558),
            .I(N__48518));
    Span4Mux_h I__7974 (
            .O(N__48553),
            .I(N__48513));
    Span4Mux_v I__7973 (
            .O(N__48542),
            .I(N__48513));
    Odrv12 I__7972 (
            .O(N__48539),
            .I(dc32_fifo_data_in_10));
    Odrv4 I__7971 (
            .O(N__48536),
            .I(dc32_fifo_data_in_10));
    Odrv12 I__7970 (
            .O(N__48521),
            .I(dc32_fifo_data_in_10));
    Odrv4 I__7969 (
            .O(N__48518),
            .I(dc32_fifo_data_in_10));
    Odrv4 I__7968 (
            .O(N__48513),
            .I(dc32_fifo_data_in_10));
    InMux I__7967 (
            .O(N__48502),
            .I(N__48499));
    LocalMux I__7966 (
            .O(N__48499),
            .I(N__48496));
    Span4Mux_v I__7965 (
            .O(N__48496),
            .I(N__48493));
    Span4Mux_h I__7964 (
            .O(N__48493),
            .I(N__48490));
    Span4Mux_v I__7963 (
            .O(N__48490),
            .I(N__48486));
    InMux I__7962 (
            .O(N__48489),
            .I(N__48483));
    Odrv4 I__7961 (
            .O(N__48486),
            .I(REG_mem_47_10));
    LocalMux I__7960 (
            .O(N__48483),
            .I(REG_mem_47_10));
    CascadeMux I__7959 (
            .O(N__48478),
            .I(N__48475));
    InMux I__7958 (
            .O(N__48475),
            .I(N__48472));
    LocalMux I__7957 (
            .O(N__48472),
            .I(N__48469));
    Span4Mux_v I__7956 (
            .O(N__48469),
            .I(N__48466));
    Sp12to4 I__7955 (
            .O(N__48466),
            .I(N__48463));
    Span12Mux_v I__7954 (
            .O(N__48463),
            .I(N__48459));
    InMux I__7953 (
            .O(N__48462),
            .I(N__48456));
    Odrv12 I__7952 (
            .O(N__48459),
            .I(REG_mem_9_7));
    LocalMux I__7951 (
            .O(N__48456),
            .I(REG_mem_9_7));
    InMux I__7950 (
            .O(N__48451),
            .I(N__48448));
    LocalMux I__7949 (
            .O(N__48448),
            .I(N__48444));
    InMux I__7948 (
            .O(N__48447),
            .I(N__48441));
    Odrv4 I__7947 (
            .O(N__48444),
            .I(REG_mem_13_9));
    LocalMux I__7946 (
            .O(N__48441),
            .I(REG_mem_13_9));
    InMux I__7945 (
            .O(N__48436),
            .I(N__48433));
    LocalMux I__7944 (
            .O(N__48433),
            .I(N__48430));
    Span4Mux_h I__7943 (
            .O(N__48430),
            .I(N__48426));
    InMux I__7942 (
            .O(N__48429),
            .I(N__48423));
    Odrv4 I__7941 (
            .O(N__48426),
            .I(REG_mem_18_9));
    LocalMux I__7940 (
            .O(N__48423),
            .I(REG_mem_18_9));
    CascadeMux I__7939 (
            .O(N__48418),
            .I(N__48414));
    InMux I__7938 (
            .O(N__48417),
            .I(N__48409));
    InMux I__7937 (
            .O(N__48414),
            .I(N__48409));
    LocalMux I__7936 (
            .O(N__48409),
            .I(REG_mem_37_7));
    CascadeMux I__7935 (
            .O(N__48406),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13862_cascade_ ));
    InMux I__7934 (
            .O(N__48403),
            .I(N__48399));
    InMux I__7933 (
            .O(N__48402),
            .I(N__48396));
    LocalMux I__7932 (
            .O(N__48399),
            .I(REG_mem_36_7));
    LocalMux I__7931 (
            .O(N__48396),
            .I(REG_mem_36_7));
    InMux I__7930 (
            .O(N__48391),
            .I(N__48388));
    LocalMux I__7929 (
            .O(N__48388),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11762 ));
    InMux I__7928 (
            .O(N__48385),
            .I(N__48382));
    LocalMux I__7927 (
            .O(N__48382),
            .I(N__48379));
    Span4Mux_v I__7926 (
            .O(N__48379),
            .I(N__48376));
    Odrv4 I__7925 (
            .O(N__48376),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13562 ));
    InMux I__7924 (
            .O(N__48373),
            .I(N__48369));
    InMux I__7923 (
            .O(N__48372),
            .I(N__48366));
    LocalMux I__7922 (
            .O(N__48369),
            .I(REG_mem_7_0));
    LocalMux I__7921 (
            .O(N__48366),
            .I(REG_mem_7_0));
    CascadeMux I__7920 (
            .O(N__48361),
            .I(N__48358));
    InMux I__7919 (
            .O(N__48358),
            .I(N__48354));
    InMux I__7918 (
            .O(N__48357),
            .I(N__48351));
    LocalMux I__7917 (
            .O(N__48354),
            .I(REG_mem_14_9));
    LocalMux I__7916 (
            .O(N__48351),
            .I(REG_mem_14_9));
    InMux I__7915 (
            .O(N__48346),
            .I(N__48342));
    InMux I__7914 (
            .O(N__48345),
            .I(N__48339));
    LocalMux I__7913 (
            .O(N__48342),
            .I(REG_mem_49_5));
    LocalMux I__7912 (
            .O(N__48339),
            .I(REG_mem_49_5));
    CascadeMux I__7911 (
            .O(N__48334),
            .I(N__48331));
    InMux I__7910 (
            .O(N__48331),
            .I(N__48328));
    LocalMux I__7909 (
            .O(N__48328),
            .I(N__48325));
    Odrv12 I__7908 (
            .O(N__48325),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12304 ));
    InMux I__7907 (
            .O(N__48322),
            .I(N__48319));
    LocalMux I__7906 (
            .O(N__48319),
            .I(N__48316));
    Odrv12 I__7905 (
            .O(N__48316),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12305 ));
    InMux I__7904 (
            .O(N__48313),
            .I(N__48310));
    LocalMux I__7903 (
            .O(N__48310),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12295 ));
    CascadeMux I__7902 (
            .O(N__48307),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13214_cascade_ ));
    CascadeMux I__7901 (
            .O(N__48304),
            .I(N__48301));
    InMux I__7900 (
            .O(N__48301),
            .I(N__48297));
    InMux I__7899 (
            .O(N__48300),
            .I(N__48294));
    LocalMux I__7898 (
            .O(N__48297),
            .I(REG_mem_50_5));
    LocalMux I__7897 (
            .O(N__48294),
            .I(REG_mem_50_5));
    InMux I__7896 (
            .O(N__48289),
            .I(N__48285));
    InMux I__7895 (
            .O(N__48288),
            .I(N__48282));
    LocalMux I__7894 (
            .O(N__48285),
            .I(REG_mem_51_5));
    LocalMux I__7893 (
            .O(N__48282),
            .I(REG_mem_51_5));
    InMux I__7892 (
            .O(N__48277),
            .I(N__48274));
    LocalMux I__7891 (
            .O(N__48274),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12296 ));
    InMux I__7890 (
            .O(N__48271),
            .I(N__48265));
    InMux I__7889 (
            .O(N__48270),
            .I(N__48265));
    LocalMux I__7888 (
            .O(N__48265),
            .I(REG_mem_48_5));
    CascadeMux I__7887 (
            .O(N__48262),
            .I(N__48259));
    InMux I__7886 (
            .O(N__48259),
            .I(N__48256));
    LocalMux I__7885 (
            .O(N__48256),
            .I(N__48252));
    InMux I__7884 (
            .O(N__48255),
            .I(N__48249));
    Odrv4 I__7883 (
            .O(N__48252),
            .I(REG_mem_39_7));
    LocalMux I__7882 (
            .O(N__48249),
            .I(REG_mem_39_7));
    CascadeMux I__7881 (
            .O(N__48244),
            .I(N__48241));
    InMux I__7880 (
            .O(N__48241),
            .I(N__48238));
    LocalMux I__7879 (
            .O(N__48238),
            .I(N__48235));
    Span4Mux_v I__7878 (
            .O(N__48235),
            .I(N__48231));
    InMux I__7877 (
            .O(N__48234),
            .I(N__48228));
    Odrv4 I__7876 (
            .O(N__48231),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_2 ));
    LocalMux I__7875 (
            .O(N__48228),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_2 ));
    InMux I__7874 (
            .O(N__48223),
            .I(N__48220));
    LocalMux I__7873 (
            .O(N__48220),
            .I(N__48217));
    Span4Mux_v I__7872 (
            .O(N__48217),
            .I(N__48213));
    CascadeMux I__7871 (
            .O(N__48216),
            .I(N__48210));
    Span4Mux_h I__7870 (
            .O(N__48213),
            .I(N__48207));
    InMux I__7869 (
            .O(N__48210),
            .I(N__48204));
    Odrv4 I__7868 (
            .O(N__48207),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_5 ));
    LocalMux I__7867 (
            .O(N__48204),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_5 ));
    CascadeMux I__7866 (
            .O(N__48199),
            .I(N__48195));
    InMux I__7865 (
            .O(N__48198),
            .I(N__48190));
    InMux I__7864 (
            .O(N__48195),
            .I(N__48190));
    LocalMux I__7863 (
            .O(N__48190),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_9 ));
    CascadeMux I__7862 (
            .O(N__48187),
            .I(N__48184));
    InMux I__7861 (
            .O(N__48184),
            .I(N__48181));
    LocalMux I__7860 (
            .O(N__48181),
            .I(N__48178));
    Span4Mux_h I__7859 (
            .O(N__48178),
            .I(N__48175));
    Odrv4 I__7858 (
            .O(N__48175),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12382 ));
    CascadeMux I__7857 (
            .O(N__48172),
            .I(N__48168));
    InMux I__7856 (
            .O(N__48171),
            .I(N__48163));
    InMux I__7855 (
            .O(N__48168),
            .I(N__48163));
    LocalMux I__7854 (
            .O(N__48163),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_9 ));
    InMux I__7853 (
            .O(N__48160),
            .I(N__48157));
    LocalMux I__7852 (
            .O(N__48157),
            .I(N__48153));
    CascadeMux I__7851 (
            .O(N__48156),
            .I(N__48150));
    Sp12to4 I__7850 (
            .O(N__48153),
            .I(N__48147));
    InMux I__7849 (
            .O(N__48150),
            .I(N__48144));
    Odrv12 I__7848 (
            .O(N__48147),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_5 ));
    LocalMux I__7847 (
            .O(N__48144),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_5 ));
    InMux I__7846 (
            .O(N__48139),
            .I(N__48136));
    LocalMux I__7845 (
            .O(N__48136),
            .I(N__48133));
    Span4Mux_h I__7844 (
            .O(N__48133),
            .I(N__48129));
    InMux I__7843 (
            .O(N__48132),
            .I(N__48126));
    Odrv4 I__7842 (
            .O(N__48129),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_5 ));
    LocalMux I__7841 (
            .O(N__48126),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_5 ));
    InMux I__7840 (
            .O(N__48121),
            .I(N__48118));
    LocalMux I__7839 (
            .O(N__48118),
            .I(N__48114));
    InMux I__7838 (
            .O(N__48117),
            .I(N__48111));
    Odrv12 I__7837 (
            .O(N__48114),
            .I(REG_mem_4_1));
    LocalMux I__7836 (
            .O(N__48111),
            .I(REG_mem_4_1));
    InMux I__7835 (
            .O(N__48106),
            .I(N__48100));
    InMux I__7834 (
            .O(N__48105),
            .I(N__48100));
    LocalMux I__7833 (
            .O(N__48100),
            .I(REG_mem_5_1));
    InMux I__7832 (
            .O(N__48097),
            .I(N__48094));
    LocalMux I__7831 (
            .O(N__48094),
            .I(N__48091));
    Span4Mux_v I__7830 (
            .O(N__48091),
            .I(N__48087));
    InMux I__7829 (
            .O(N__48090),
            .I(N__48084));
    Odrv4 I__7828 (
            .O(N__48087),
            .I(REG_mem_36_5));
    LocalMux I__7827 (
            .O(N__48084),
            .I(REG_mem_36_5));
    InMux I__7826 (
            .O(N__48079),
            .I(N__48076));
    LocalMux I__7825 (
            .O(N__48076),
            .I(N__48072));
    CascadeMux I__7824 (
            .O(N__48075),
            .I(N__48069));
    Span4Mux_v I__7823 (
            .O(N__48072),
            .I(N__48066));
    InMux I__7822 (
            .O(N__48069),
            .I(N__48063));
    Odrv4 I__7821 (
            .O(N__48066),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_0 ));
    LocalMux I__7820 (
            .O(N__48063),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_0 ));
    InMux I__7819 (
            .O(N__48058),
            .I(N__48054));
    InMux I__7818 (
            .O(N__48057),
            .I(N__48051));
    LocalMux I__7817 (
            .O(N__48054),
            .I(REG_mem_48_2));
    LocalMux I__7816 (
            .O(N__48051),
            .I(REG_mem_48_2));
    InMux I__7815 (
            .O(N__48046),
            .I(N__48043));
    LocalMux I__7814 (
            .O(N__48043),
            .I(N__48040));
    Span4Mux_v I__7813 (
            .O(N__48040),
            .I(N__48037));
    Span4Mux_h I__7812 (
            .O(N__48037),
            .I(N__48034));
    Odrv4 I__7811 (
            .O(N__48034),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13685 ));
    CascadeMux I__7810 (
            .O(N__48031),
            .I(N__48028));
    InMux I__7809 (
            .O(N__48028),
            .I(N__48025));
    LocalMux I__7808 (
            .O(N__48025),
            .I(N__48022));
    Span4Mux_v I__7807 (
            .O(N__48022),
            .I(N__48019));
    Odrv4 I__7806 (
            .O(N__48019),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12098 ));
    InMux I__7805 (
            .O(N__48016),
            .I(N__48013));
    LocalMux I__7804 (
            .O(N__48013),
            .I(N__48010));
    Span4Mux_v I__7803 (
            .O(N__48010),
            .I(N__48007));
    Span4Mux_h I__7802 (
            .O(N__48007),
            .I(N__48004));
    Odrv4 I__7801 (
            .O(N__48004),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14078 ));
    InMux I__7800 (
            .O(N__48001),
            .I(N__47997));
    InMux I__7799 (
            .O(N__48000),
            .I(N__47994));
    LocalMux I__7798 (
            .O(N__47997),
            .I(REG_mem_10_1));
    LocalMux I__7797 (
            .O(N__47994),
            .I(REG_mem_10_1));
    InMux I__7796 (
            .O(N__47989),
            .I(N__47985));
    InMux I__7795 (
            .O(N__47988),
            .I(N__47982));
    LocalMux I__7794 (
            .O(N__47985),
            .I(REG_mem_6_2));
    LocalMux I__7793 (
            .O(N__47982),
            .I(REG_mem_6_2));
    InMux I__7792 (
            .O(N__47977),
            .I(N__47974));
    LocalMux I__7791 (
            .O(N__47974),
            .I(N__47970));
    CascadeMux I__7790 (
            .O(N__47973),
            .I(N__47967));
    Span4Mux_h I__7789 (
            .O(N__47970),
            .I(N__47964));
    InMux I__7788 (
            .O(N__47967),
            .I(N__47961));
    Span4Mux_h I__7787 (
            .O(N__47964),
            .I(N__47958));
    LocalMux I__7786 (
            .O(N__47961),
            .I(N__47955));
    Odrv4 I__7785 (
            .O(N__47958),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_5 ));
    Odrv4 I__7784 (
            .O(N__47955),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_5 ));
    InMux I__7783 (
            .O(N__47950),
            .I(N__47946));
    InMux I__7782 (
            .O(N__47949),
            .I(N__47943));
    LocalMux I__7781 (
            .O(N__47946),
            .I(REG_mem_45_1));
    LocalMux I__7780 (
            .O(N__47943),
            .I(REG_mem_45_1));
    InMux I__7779 (
            .O(N__47938),
            .I(N__47935));
    LocalMux I__7778 (
            .O(N__47935),
            .I(N__47931));
    InMux I__7777 (
            .O(N__47934),
            .I(N__47928));
    Odrv4 I__7776 (
            .O(N__47931),
            .I(REG_mem_46_15));
    LocalMux I__7775 (
            .O(N__47928),
            .I(REG_mem_46_15));
    InMux I__7774 (
            .O(N__47923),
            .I(N__47919));
    InMux I__7773 (
            .O(N__47922),
            .I(N__47916));
    LocalMux I__7772 (
            .O(N__47919),
            .I(REG_mem_40_5));
    LocalMux I__7771 (
            .O(N__47916),
            .I(REG_mem_40_5));
    InMux I__7770 (
            .O(N__47911),
            .I(N__47907));
    InMux I__7769 (
            .O(N__47910),
            .I(N__47904));
    LocalMux I__7768 (
            .O(N__47907),
            .I(REG_mem_55_5));
    LocalMux I__7767 (
            .O(N__47904),
            .I(REG_mem_55_5));
    CascadeMux I__7766 (
            .O(N__47899),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14123_cascade_ ));
    InMux I__7765 (
            .O(N__47896),
            .I(N__47893));
    LocalMux I__7764 (
            .O(N__47893),
            .I(N__47890));
    Span4Mux_v I__7763 (
            .O(N__47890),
            .I(N__47886));
    InMux I__7762 (
            .O(N__47889),
            .I(N__47883));
    Odrv4 I__7761 (
            .O(N__47886),
            .I(REG_mem_7_2));
    LocalMux I__7760 (
            .O(N__47883),
            .I(REG_mem_7_2));
    CascadeMux I__7759 (
            .O(N__47878),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13886_cascade_ ));
    InMux I__7758 (
            .O(N__47875),
            .I(N__47872));
    LocalMux I__7757 (
            .O(N__47872),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13889 ));
    InMux I__7756 (
            .O(N__47869),
            .I(N__47866));
    LocalMux I__7755 (
            .O(N__47866),
            .I(N__47862));
    CascadeMux I__7754 (
            .O(N__47865),
            .I(N__47859));
    Span4Mux_v I__7753 (
            .O(N__47862),
            .I(N__47856));
    InMux I__7752 (
            .O(N__47859),
            .I(N__47853));
    Odrv4 I__7751 (
            .O(N__47856),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_2 ));
    LocalMux I__7750 (
            .O(N__47853),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_2 ));
    InMux I__7749 (
            .O(N__47848),
            .I(N__47845));
    LocalMux I__7748 (
            .O(N__47845),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14120 ));
    InMux I__7747 (
            .O(N__47842),
            .I(N__47836));
    InMux I__7746 (
            .O(N__47841),
            .I(N__47836));
    LocalMux I__7745 (
            .O(N__47836),
            .I(REG_mem_5_2));
    InMux I__7744 (
            .O(N__47833),
            .I(N__47827));
    InMux I__7743 (
            .O(N__47832),
            .I(N__47827));
    LocalMux I__7742 (
            .O(N__47827),
            .I(REG_mem_4_2));
    InMux I__7741 (
            .O(N__47824),
            .I(N__47820));
    InMux I__7740 (
            .O(N__47823),
            .I(N__47817));
    LocalMux I__7739 (
            .O(N__47820),
            .I(REG_mem_48_1));
    LocalMux I__7738 (
            .O(N__47817),
            .I(REG_mem_48_1));
    InMux I__7737 (
            .O(N__47812),
            .I(N__47808));
    InMux I__7736 (
            .O(N__47811),
            .I(N__47805));
    LocalMux I__7735 (
            .O(N__47808),
            .I(REG_mem_49_1));
    LocalMux I__7734 (
            .O(N__47805),
            .I(REG_mem_49_1));
    InMux I__7733 (
            .O(N__47800),
            .I(N__47796));
    InMux I__7732 (
            .O(N__47799),
            .I(N__47793));
    LocalMux I__7731 (
            .O(N__47796),
            .I(REG_mem_47_1));
    LocalMux I__7730 (
            .O(N__47793),
            .I(REG_mem_47_1));
    InMux I__7729 (
            .O(N__47788),
            .I(N__47784));
    InMux I__7728 (
            .O(N__47787),
            .I(N__47781));
    LocalMux I__7727 (
            .O(N__47784),
            .I(N__47778));
    LocalMux I__7726 (
            .O(N__47781),
            .I(REG_mem_46_1));
    Odrv4 I__7725 (
            .O(N__47778),
            .I(REG_mem_46_1));
    CascadeMux I__7724 (
            .O(N__47773),
            .I(N__47770));
    InMux I__7723 (
            .O(N__47770),
            .I(N__47767));
    LocalMux I__7722 (
            .O(N__47767),
            .I(N__47764));
    Span4Mux_h I__7721 (
            .O(N__47764),
            .I(N__47760));
    InMux I__7720 (
            .O(N__47763),
            .I(N__47757));
    Odrv4 I__7719 (
            .O(N__47760),
            .I(REG_mem_41_5));
    LocalMux I__7718 (
            .O(N__47757),
            .I(REG_mem_41_5));
    InMux I__7717 (
            .O(N__47752),
            .I(N__47749));
    LocalMux I__7716 (
            .O(N__47749),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13742 ));
    InMux I__7715 (
            .O(N__47746),
            .I(\spi0.n10702 ));
    InMux I__7714 (
            .O(N__47743),
            .I(N__47740));
    LocalMux I__7713 (
            .O(N__47740),
            .I(N__47737));
    Span4Mux_v I__7712 (
            .O(N__47737),
            .I(N__47733));
    InMux I__7711 (
            .O(N__47736),
            .I(N__47730));
    Odrv4 I__7710 (
            .O(N__47733),
            .I(REG_mem_58_11));
    LocalMux I__7709 (
            .O(N__47730),
            .I(REG_mem_58_11));
    CascadeMux I__7708 (
            .O(N__47725),
            .I(N__47722));
    InMux I__7707 (
            .O(N__47722),
            .I(N__47718));
    CascadeMux I__7706 (
            .O(N__47721),
            .I(N__47715));
    LocalMux I__7705 (
            .O(N__47718),
            .I(N__47712));
    InMux I__7704 (
            .O(N__47715),
            .I(N__47709));
    Odrv12 I__7703 (
            .O(N__47712),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_11 ));
    LocalMux I__7702 (
            .O(N__47709),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_11 ));
    InMux I__7701 (
            .O(N__47704),
            .I(N__47701));
    LocalMux I__7700 (
            .O(N__47701),
            .I(N__47698));
    Span4Mux_h I__7699 (
            .O(N__47698),
            .I(N__47694));
    CascadeMux I__7698 (
            .O(N__47697),
            .I(N__47691));
    Span4Mux_v I__7697 (
            .O(N__47694),
            .I(N__47688));
    InMux I__7696 (
            .O(N__47691),
            .I(N__47685));
    Odrv4 I__7695 (
            .O(N__47688),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_11 ));
    LocalMux I__7694 (
            .O(N__47685),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_11 ));
    CascadeMux I__7693 (
            .O(N__47680),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13748_cascade_ ));
    InMux I__7692 (
            .O(N__47677),
            .I(N__47673));
    InMux I__7691 (
            .O(N__47676),
            .I(N__47670));
    LocalMux I__7690 (
            .O(N__47673),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_11 ));
    LocalMux I__7689 (
            .O(N__47670),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_11 ));
    CascadeMux I__7688 (
            .O(N__47665),
            .I(N__47662));
    InMux I__7687 (
            .O(N__47662),
            .I(N__47659));
    LocalMux I__7686 (
            .O(N__47659),
            .I(N__47656));
    Span4Mux_v I__7685 (
            .O(N__47656),
            .I(N__47652));
    InMux I__7684 (
            .O(N__47655),
            .I(N__47649));
    Span4Mux_h I__7683 (
            .O(N__47652),
            .I(N__47646));
    LocalMux I__7682 (
            .O(N__47649),
            .I(N__47643));
    Odrv4 I__7681 (
            .O(N__47646),
            .I(REG_mem_63_11));
    Odrv4 I__7680 (
            .O(N__47643),
            .I(REG_mem_63_11));
    InMux I__7679 (
            .O(N__47638),
            .I(N__47634));
    CascadeMux I__7678 (
            .O(N__47637),
            .I(N__47631));
    LocalMux I__7677 (
            .O(N__47634),
            .I(N__47628));
    InMux I__7676 (
            .O(N__47631),
            .I(N__47625));
    Odrv4 I__7675 (
            .O(N__47628),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_11 ));
    LocalMux I__7674 (
            .O(N__47625),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_11 ));
    InMux I__7673 (
            .O(N__47620),
            .I(N__47617));
    LocalMux I__7672 (
            .O(N__47617),
            .I(N__47613));
    CascadeMux I__7671 (
            .O(N__47616),
            .I(N__47610));
    Span4Mux_v I__7670 (
            .O(N__47613),
            .I(N__47607));
    InMux I__7669 (
            .O(N__47610),
            .I(N__47604));
    Odrv4 I__7668 (
            .O(N__47607),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_11 ));
    LocalMux I__7667 (
            .O(N__47604),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_11 ));
    CascadeMux I__7666 (
            .O(N__47599),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13616_cascade_ ));
    InMux I__7665 (
            .O(N__47596),
            .I(N__47593));
    LocalMux I__7664 (
            .O(N__47593),
            .I(N__47590));
    Span4Mux_h I__7663 (
            .O(N__47590),
            .I(N__47586));
    CascadeMux I__7662 (
            .O(N__47589),
            .I(N__47583));
    Span4Mux_v I__7661 (
            .O(N__47586),
            .I(N__47580));
    InMux I__7660 (
            .O(N__47583),
            .I(N__47577));
    Odrv4 I__7659 (
            .O(N__47580),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_11 ));
    LocalMux I__7658 (
            .O(N__47577),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_11 ));
    CascadeMux I__7657 (
            .O(N__47572),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13619_cascade_ ));
    InMux I__7656 (
            .O(N__47569),
            .I(N__47566));
    LocalMux I__7655 (
            .O(N__47566),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13751 ));
    InMux I__7654 (
            .O(N__47563),
            .I(N__47560));
    LocalMux I__7653 (
            .O(N__47560),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14147 ));
    CascadeMux I__7652 (
            .O(N__47557),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14324_cascade_ ));
    InMux I__7651 (
            .O(N__47554),
            .I(N__47551));
    LocalMux I__7650 (
            .O(N__47551),
            .I(N__47548));
    Odrv12 I__7649 (
            .O(N__47548),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14207 ));
    InMux I__7648 (
            .O(N__47545),
            .I(bfn_11_18_0_));
    InMux I__7647 (
            .O(N__47542),
            .I(\spi0.n10694 ));
    InMux I__7646 (
            .O(N__47539),
            .I(\spi0.n10695 ));
    InMux I__7645 (
            .O(N__47536),
            .I(\spi0.n10696 ));
    InMux I__7644 (
            .O(N__47533),
            .I(\spi0.n10697 ));
    InMux I__7643 (
            .O(N__47530),
            .I(\spi0.n10698 ));
    InMux I__7642 (
            .O(N__47527),
            .I(\spi0.n10699 ));
    InMux I__7641 (
            .O(N__47524),
            .I(\spi0.n10700 ));
    InMux I__7640 (
            .O(N__47521),
            .I(bfn_11_19_0_));
    InMux I__7639 (
            .O(N__47518),
            .I(N__47515));
    LocalMux I__7638 (
            .O(N__47515),
            .I(N__47512));
    Odrv4 I__7637 (
            .O(N__47512),
            .I(rp_sync1_r_6));
    InMux I__7636 (
            .O(N__47509),
            .I(N__47503));
    InMux I__7635 (
            .O(N__47508),
            .I(N__47503));
    LocalMux I__7634 (
            .O(N__47503),
            .I(REG_mem_13_11));
    CascadeMux I__7633 (
            .O(N__47500),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14396_cascade_ ));
    InMux I__7632 (
            .O(N__47497),
            .I(N__47494));
    LocalMux I__7631 (
            .O(N__47494),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12456 ));
    InMux I__7630 (
            .O(N__47491),
            .I(N__47485));
    InMux I__7629 (
            .O(N__47490),
            .I(N__47485));
    LocalMux I__7628 (
            .O(N__47485),
            .I(REG_mem_12_11));
    InMux I__7627 (
            .O(N__47482),
            .I(N__47476));
    InMux I__7626 (
            .O(N__47481),
            .I(N__47476));
    LocalMux I__7625 (
            .O(N__47476),
            .I(REG_mem_14_11));
    CascadeMux I__7624 (
            .O(N__47473),
            .I(N__47470));
    InMux I__7623 (
            .O(N__47470),
            .I(N__47464));
    InMux I__7622 (
            .O(N__47469),
            .I(N__47464));
    LocalMux I__7621 (
            .O(N__47464),
            .I(REG_mem_15_11));
    CascadeMux I__7620 (
            .O(N__47461),
            .I(N__47455));
    CascadeMux I__7619 (
            .O(N__47460),
            .I(N__47448));
    InMux I__7618 (
            .O(N__47459),
            .I(N__47438));
    InMux I__7617 (
            .O(N__47458),
            .I(N__47438));
    InMux I__7616 (
            .O(N__47455),
            .I(N__47419));
    InMux I__7615 (
            .O(N__47454),
            .I(N__47419));
    InMux I__7614 (
            .O(N__47453),
            .I(N__47419));
    InMux I__7613 (
            .O(N__47452),
            .I(N__47419));
    CascadeMux I__7612 (
            .O(N__47451),
            .I(N__47413));
    InMux I__7611 (
            .O(N__47448),
            .I(N__47397));
    InMux I__7610 (
            .O(N__47447),
            .I(N__47397));
    InMux I__7609 (
            .O(N__47446),
            .I(N__47397));
    InMux I__7608 (
            .O(N__47445),
            .I(N__47397));
    InMux I__7607 (
            .O(N__47444),
            .I(N__47397));
    CascadeMux I__7606 (
            .O(N__47443),
            .I(N__47394));
    LocalMux I__7605 (
            .O(N__47438),
            .I(N__47379));
    InMux I__7604 (
            .O(N__47437),
            .I(N__47374));
    InMux I__7603 (
            .O(N__47436),
            .I(N__47374));
    InMux I__7602 (
            .O(N__47435),
            .I(N__47364));
    InMux I__7601 (
            .O(N__47434),
            .I(N__47364));
    InMux I__7600 (
            .O(N__47433),
            .I(N__47364));
    InMux I__7599 (
            .O(N__47432),
            .I(N__47364));
    InMux I__7598 (
            .O(N__47431),
            .I(N__47361));
    InMux I__7597 (
            .O(N__47430),
            .I(N__47356));
    InMux I__7596 (
            .O(N__47429),
            .I(N__47356));
    InMux I__7595 (
            .O(N__47428),
            .I(N__47353));
    LocalMux I__7594 (
            .O(N__47419),
            .I(N__47350));
    InMux I__7593 (
            .O(N__47418),
            .I(N__47343));
    InMux I__7592 (
            .O(N__47417),
            .I(N__47343));
    InMux I__7591 (
            .O(N__47416),
            .I(N__47343));
    InMux I__7590 (
            .O(N__47413),
            .I(N__47334));
    InMux I__7589 (
            .O(N__47412),
            .I(N__47331));
    InMux I__7588 (
            .O(N__47411),
            .I(N__47326));
    InMux I__7587 (
            .O(N__47410),
            .I(N__47326));
    InMux I__7586 (
            .O(N__47409),
            .I(N__47321));
    InMux I__7585 (
            .O(N__47408),
            .I(N__47321));
    LocalMux I__7584 (
            .O(N__47397),
            .I(N__47318));
    InMux I__7583 (
            .O(N__47394),
            .I(N__47297));
    InMux I__7582 (
            .O(N__47393),
            .I(N__47297));
    InMux I__7581 (
            .O(N__47392),
            .I(N__47297));
    InMux I__7580 (
            .O(N__47391),
            .I(N__47297));
    InMux I__7579 (
            .O(N__47390),
            .I(N__47297));
    InMux I__7578 (
            .O(N__47389),
            .I(N__47297));
    CascadeMux I__7577 (
            .O(N__47388),
            .I(N__47293));
    CascadeMux I__7576 (
            .O(N__47387),
            .I(N__47290));
    InMux I__7575 (
            .O(N__47386),
            .I(N__47279));
    InMux I__7574 (
            .O(N__47385),
            .I(N__47279));
    InMux I__7573 (
            .O(N__47384),
            .I(N__47279));
    InMux I__7572 (
            .O(N__47383),
            .I(N__47279));
    InMux I__7571 (
            .O(N__47382),
            .I(N__47279));
    Span4Mux_v I__7570 (
            .O(N__47379),
            .I(N__47274));
    LocalMux I__7569 (
            .O(N__47374),
            .I(N__47274));
    InMux I__7568 (
            .O(N__47373),
            .I(N__47271));
    LocalMux I__7567 (
            .O(N__47364),
            .I(N__47268));
    LocalMux I__7566 (
            .O(N__47361),
            .I(N__47257));
    LocalMux I__7565 (
            .O(N__47356),
            .I(N__47257));
    LocalMux I__7564 (
            .O(N__47353),
            .I(N__47257));
    Span4Mux_v I__7563 (
            .O(N__47350),
            .I(N__47257));
    LocalMux I__7562 (
            .O(N__47343),
            .I(N__47257));
    InMux I__7561 (
            .O(N__47342),
            .I(N__47252));
    InMux I__7560 (
            .O(N__47341),
            .I(N__47252));
    InMux I__7559 (
            .O(N__47340),
            .I(N__47247));
    InMux I__7558 (
            .O(N__47339),
            .I(N__47247));
    InMux I__7557 (
            .O(N__47338),
            .I(N__47244));
    InMux I__7556 (
            .O(N__47337),
            .I(N__47241));
    LocalMux I__7555 (
            .O(N__47334),
            .I(N__47230));
    LocalMux I__7554 (
            .O(N__47331),
            .I(N__47230));
    LocalMux I__7553 (
            .O(N__47326),
            .I(N__47230));
    LocalMux I__7552 (
            .O(N__47321),
            .I(N__47230));
    Span4Mux_v I__7551 (
            .O(N__47318),
            .I(N__47230));
    InMux I__7550 (
            .O(N__47317),
            .I(N__47223));
    InMux I__7549 (
            .O(N__47316),
            .I(N__47223));
    InMux I__7548 (
            .O(N__47315),
            .I(N__47223));
    InMux I__7547 (
            .O(N__47314),
            .I(N__47214));
    InMux I__7546 (
            .O(N__47313),
            .I(N__47214));
    InMux I__7545 (
            .O(N__47312),
            .I(N__47214));
    InMux I__7544 (
            .O(N__47311),
            .I(N__47214));
    InMux I__7543 (
            .O(N__47310),
            .I(N__47210));
    LocalMux I__7542 (
            .O(N__47297),
            .I(N__47207));
    CascadeMux I__7541 (
            .O(N__47296),
            .I(N__47204));
    InMux I__7540 (
            .O(N__47293),
            .I(N__47199));
    InMux I__7539 (
            .O(N__47290),
            .I(N__47199));
    LocalMux I__7538 (
            .O(N__47279),
            .I(N__47196));
    Span4Mux_v I__7537 (
            .O(N__47274),
            .I(N__47193));
    LocalMux I__7536 (
            .O(N__47271),
            .I(N__47184));
    Span4Mux_h I__7535 (
            .O(N__47268),
            .I(N__47184));
    Span4Mux_v I__7534 (
            .O(N__47257),
            .I(N__47184));
    LocalMux I__7533 (
            .O(N__47252),
            .I(N__47184));
    LocalMux I__7532 (
            .O(N__47247),
            .I(N__47181));
    LocalMux I__7531 (
            .O(N__47244),
            .I(N__47177));
    LocalMux I__7530 (
            .O(N__47241),
            .I(N__47174));
    Span4Mux_v I__7529 (
            .O(N__47230),
            .I(N__47169));
    LocalMux I__7528 (
            .O(N__47223),
            .I(N__47169));
    LocalMux I__7527 (
            .O(N__47214),
            .I(N__47166));
    InMux I__7526 (
            .O(N__47213),
            .I(N__47163));
    LocalMux I__7525 (
            .O(N__47210),
            .I(N__47158));
    Span4Mux_v I__7524 (
            .O(N__47207),
            .I(N__47158));
    InMux I__7523 (
            .O(N__47204),
            .I(N__47152));
    LocalMux I__7522 (
            .O(N__47199),
            .I(N__47143));
    Span4Mux_v I__7521 (
            .O(N__47196),
            .I(N__47143));
    Span4Mux_h I__7520 (
            .O(N__47193),
            .I(N__47143));
    Span4Mux_v I__7519 (
            .O(N__47184),
            .I(N__47143));
    Span4Mux_h I__7518 (
            .O(N__47181),
            .I(N__47140));
    InMux I__7517 (
            .O(N__47180),
            .I(N__47137));
    Span4Mux_v I__7516 (
            .O(N__47177),
            .I(N__47134));
    Span4Mux_v I__7515 (
            .O(N__47174),
            .I(N__47127));
    Span4Mux_h I__7514 (
            .O(N__47169),
            .I(N__47127));
    Span4Mux_v I__7513 (
            .O(N__47166),
            .I(N__47127));
    LocalMux I__7512 (
            .O(N__47163),
            .I(N__47122));
    Span4Mux_v I__7511 (
            .O(N__47158),
            .I(N__47122));
    InMux I__7510 (
            .O(N__47157),
            .I(N__47119));
    InMux I__7509 (
            .O(N__47156),
            .I(N__47116));
    InMux I__7508 (
            .O(N__47155),
            .I(N__47113));
    LocalMux I__7507 (
            .O(N__47152),
            .I(N__47110));
    Span4Mux_h I__7506 (
            .O(N__47143),
            .I(N__47107));
    Sp12to4 I__7505 (
            .O(N__47140),
            .I(N__47104));
    LocalMux I__7504 (
            .O(N__47137),
            .I(N__47101));
    Span4Mux_h I__7503 (
            .O(N__47134),
            .I(N__47096));
    Span4Mux_v I__7502 (
            .O(N__47127),
            .I(N__47096));
    Span4Mux_v I__7501 (
            .O(N__47122),
            .I(N__47093));
    LocalMux I__7500 (
            .O(N__47119),
            .I(N__47080));
    LocalMux I__7499 (
            .O(N__47116),
            .I(N__47080));
    LocalMux I__7498 (
            .O(N__47113),
            .I(N__47080));
    Sp12to4 I__7497 (
            .O(N__47110),
            .I(N__47080));
    Sp12to4 I__7496 (
            .O(N__47107),
            .I(N__47080));
    Span12Mux_s8_v I__7495 (
            .O(N__47104),
            .I(N__47080));
    Span4Mux_h I__7494 (
            .O(N__47101),
            .I(N__47073));
    Span4Mux_h I__7493 (
            .O(N__47096),
            .I(N__47073));
    Span4Mux_v I__7492 (
            .O(N__47093),
            .I(N__47073));
    Span12Mux_v I__7491 (
            .O(N__47080),
            .I(N__47070));
    Span4Mux_v I__7490 (
            .O(N__47073),
            .I(N__47067));
    Odrv12 I__7489 (
            .O(N__47070),
            .I(dc32_fifo_data_in_11));
    Odrv4 I__7488 (
            .O(N__47067),
            .I(dc32_fifo_data_in_11));
    CascadeMux I__7487 (
            .O(N__47062),
            .I(N__47059));
    InMux I__7486 (
            .O(N__47059),
            .I(N__47056));
    LocalMux I__7485 (
            .O(N__47056),
            .I(N__47053));
    Span4Mux_v I__7484 (
            .O(N__47053),
            .I(N__47049));
    InMux I__7483 (
            .O(N__47052),
            .I(N__47046));
    Odrv4 I__7482 (
            .O(N__47049),
            .I(REG_mem_6_11));
    LocalMux I__7481 (
            .O(N__47046),
            .I(REG_mem_6_11));
    CascadeMux I__7480 (
            .O(N__47041),
            .I(N__47035));
    InMux I__7479 (
            .O(N__47040),
            .I(N__47032));
    CascadeMux I__7478 (
            .O(N__47039),
            .I(N__47027));
    CascadeMux I__7477 (
            .O(N__47038),
            .I(N__47017));
    InMux I__7476 (
            .O(N__47035),
            .I(N__47006));
    LocalMux I__7475 (
            .O(N__47032),
            .I(N__47001));
    CascadeMux I__7474 (
            .O(N__47031),
            .I(N__46991));
    InMux I__7473 (
            .O(N__47030),
            .I(N__46977));
    InMux I__7472 (
            .O(N__47027),
            .I(N__46977));
    InMux I__7471 (
            .O(N__47026),
            .I(N__46977));
    InMux I__7470 (
            .O(N__47025),
            .I(N__46966));
    InMux I__7469 (
            .O(N__47024),
            .I(N__46966));
    InMux I__7468 (
            .O(N__47023),
            .I(N__46966));
    InMux I__7467 (
            .O(N__47022),
            .I(N__46957));
    InMux I__7466 (
            .O(N__47021),
            .I(N__46957));
    InMux I__7465 (
            .O(N__47020),
            .I(N__46952));
    InMux I__7464 (
            .O(N__47017),
            .I(N__46952));
    InMux I__7463 (
            .O(N__47016),
            .I(N__46949));
    InMux I__7462 (
            .O(N__47015),
            .I(N__46942));
    InMux I__7461 (
            .O(N__47014),
            .I(N__46942));
    InMux I__7460 (
            .O(N__47013),
            .I(N__46942));
    InMux I__7459 (
            .O(N__47012),
            .I(N__46939));
    InMux I__7458 (
            .O(N__47011),
            .I(N__46936));
    InMux I__7457 (
            .O(N__47010),
            .I(N__46930));
    InMux I__7456 (
            .O(N__47009),
            .I(N__46930));
    LocalMux I__7455 (
            .O(N__47006),
            .I(N__46926));
    InMux I__7454 (
            .O(N__47005),
            .I(N__46921));
    InMux I__7453 (
            .O(N__47004),
            .I(N__46921));
    Span4Mux_v I__7452 (
            .O(N__47001),
            .I(N__46918));
    InMux I__7451 (
            .O(N__47000),
            .I(N__46915));
    InMux I__7450 (
            .O(N__46999),
            .I(N__46910));
    InMux I__7449 (
            .O(N__46998),
            .I(N__46910));
    InMux I__7448 (
            .O(N__46997),
            .I(N__46903));
    InMux I__7447 (
            .O(N__46996),
            .I(N__46903));
    InMux I__7446 (
            .O(N__46995),
            .I(N__46903));
    InMux I__7445 (
            .O(N__46994),
            .I(N__46896));
    InMux I__7444 (
            .O(N__46991),
            .I(N__46891));
    InMux I__7443 (
            .O(N__46990),
            .I(N__46891));
    InMux I__7442 (
            .O(N__46989),
            .I(N__46888));
    InMux I__7441 (
            .O(N__46988),
            .I(N__46885));
    InMux I__7440 (
            .O(N__46987),
            .I(N__46876));
    InMux I__7439 (
            .O(N__46986),
            .I(N__46876));
    InMux I__7438 (
            .O(N__46985),
            .I(N__46876));
    InMux I__7437 (
            .O(N__46984),
            .I(N__46876));
    LocalMux I__7436 (
            .O(N__46977),
            .I(N__46873));
    InMux I__7435 (
            .O(N__46976),
            .I(N__46864));
    InMux I__7434 (
            .O(N__46975),
            .I(N__46864));
    InMux I__7433 (
            .O(N__46974),
            .I(N__46864));
    InMux I__7432 (
            .O(N__46973),
            .I(N__46864));
    LocalMux I__7431 (
            .O(N__46966),
            .I(N__46861));
    InMux I__7430 (
            .O(N__46965),
            .I(N__46847));
    InMux I__7429 (
            .O(N__46964),
            .I(N__46847));
    InMux I__7428 (
            .O(N__46963),
            .I(N__46847));
    InMux I__7427 (
            .O(N__46962),
            .I(N__46844));
    LocalMux I__7426 (
            .O(N__46957),
            .I(N__46839));
    LocalMux I__7425 (
            .O(N__46952),
            .I(N__46839));
    LocalMux I__7424 (
            .O(N__46949),
            .I(N__46836));
    LocalMux I__7423 (
            .O(N__46942),
            .I(N__46831));
    LocalMux I__7422 (
            .O(N__46939),
            .I(N__46831));
    LocalMux I__7421 (
            .O(N__46936),
            .I(N__46828));
    InMux I__7420 (
            .O(N__46935),
            .I(N__46825));
    LocalMux I__7419 (
            .O(N__46930),
            .I(N__46822));
    InMux I__7418 (
            .O(N__46929),
            .I(N__46819));
    Span4Mux_v I__7417 (
            .O(N__46926),
            .I(N__46806));
    LocalMux I__7416 (
            .O(N__46921),
            .I(N__46806));
    Span4Mux_h I__7415 (
            .O(N__46918),
            .I(N__46806));
    LocalMux I__7414 (
            .O(N__46915),
            .I(N__46806));
    LocalMux I__7413 (
            .O(N__46910),
            .I(N__46806));
    LocalMux I__7412 (
            .O(N__46903),
            .I(N__46806));
    InMux I__7411 (
            .O(N__46902),
            .I(N__46803));
    InMux I__7410 (
            .O(N__46901),
            .I(N__46798));
    InMux I__7409 (
            .O(N__46900),
            .I(N__46798));
    InMux I__7408 (
            .O(N__46899),
            .I(N__46795));
    LocalMux I__7407 (
            .O(N__46896),
            .I(N__46792));
    LocalMux I__7406 (
            .O(N__46891),
            .I(N__46789));
    LocalMux I__7405 (
            .O(N__46888),
            .I(N__46782));
    LocalMux I__7404 (
            .O(N__46885),
            .I(N__46782));
    LocalMux I__7403 (
            .O(N__46876),
            .I(N__46782));
    Span4Mux_v I__7402 (
            .O(N__46873),
            .I(N__46779));
    LocalMux I__7401 (
            .O(N__46864),
            .I(N__46776));
    Span4Mux_h I__7400 (
            .O(N__46861),
            .I(N__46769));
    InMux I__7399 (
            .O(N__46860),
            .I(N__46762));
    InMux I__7398 (
            .O(N__46859),
            .I(N__46762));
    InMux I__7397 (
            .O(N__46858),
            .I(N__46762));
    InMux I__7396 (
            .O(N__46857),
            .I(N__46759));
    InMux I__7395 (
            .O(N__46856),
            .I(N__46756));
    InMux I__7394 (
            .O(N__46855),
            .I(N__46751));
    InMux I__7393 (
            .O(N__46854),
            .I(N__46751));
    LocalMux I__7392 (
            .O(N__46847),
            .I(N__46742));
    LocalMux I__7391 (
            .O(N__46844),
            .I(N__46742));
    Span4Mux_h I__7390 (
            .O(N__46839),
            .I(N__46742));
    Span4Mux_h I__7389 (
            .O(N__46836),
            .I(N__46742));
    Span4Mux_h I__7388 (
            .O(N__46831),
            .I(N__46733));
    Span4Mux_h I__7387 (
            .O(N__46828),
            .I(N__46733));
    LocalMux I__7386 (
            .O(N__46825),
            .I(N__46733));
    Span4Mux_h I__7385 (
            .O(N__46822),
            .I(N__46733));
    LocalMux I__7384 (
            .O(N__46819),
            .I(N__46722));
    Span4Mux_v I__7383 (
            .O(N__46806),
            .I(N__46722));
    LocalMux I__7382 (
            .O(N__46803),
            .I(N__46722));
    LocalMux I__7381 (
            .O(N__46798),
            .I(N__46722));
    LocalMux I__7380 (
            .O(N__46795),
            .I(N__46719));
    Span4Mux_v I__7379 (
            .O(N__46792),
            .I(N__46710));
    Span4Mux_h I__7378 (
            .O(N__46789),
            .I(N__46710));
    Span4Mux_v I__7377 (
            .O(N__46782),
            .I(N__46710));
    Span4Mux_h I__7376 (
            .O(N__46779),
            .I(N__46710));
    Span4Mux_v I__7375 (
            .O(N__46776),
            .I(N__46707));
    InMux I__7374 (
            .O(N__46775),
            .I(N__46704));
    InMux I__7373 (
            .O(N__46774),
            .I(N__46701));
    InMux I__7372 (
            .O(N__46773),
            .I(N__46696));
    InMux I__7371 (
            .O(N__46772),
            .I(N__46696));
    Span4Mux_v I__7370 (
            .O(N__46769),
            .I(N__46693));
    LocalMux I__7369 (
            .O(N__46762),
            .I(N__46690));
    LocalMux I__7368 (
            .O(N__46759),
            .I(N__46679));
    LocalMux I__7367 (
            .O(N__46756),
            .I(N__46679));
    LocalMux I__7366 (
            .O(N__46751),
            .I(N__46679));
    Sp12to4 I__7365 (
            .O(N__46742),
            .I(N__46679));
    Sp12to4 I__7364 (
            .O(N__46733),
            .I(N__46679));
    InMux I__7363 (
            .O(N__46732),
            .I(N__46676));
    InMux I__7362 (
            .O(N__46731),
            .I(N__46673));
    Span4Mux_v I__7361 (
            .O(N__46722),
            .I(N__46670));
    Span4Mux_v I__7360 (
            .O(N__46719),
            .I(N__46663));
    Span4Mux_v I__7359 (
            .O(N__46710),
            .I(N__46663));
    Span4Mux_h I__7358 (
            .O(N__46707),
            .I(N__46663));
    LocalMux I__7357 (
            .O(N__46704),
            .I(N__46650));
    LocalMux I__7356 (
            .O(N__46701),
            .I(N__46650));
    LocalMux I__7355 (
            .O(N__46696),
            .I(N__46650));
    Sp12to4 I__7354 (
            .O(N__46693),
            .I(N__46650));
    Span12Mux_s11_h I__7353 (
            .O(N__46690),
            .I(N__46650));
    Span12Mux_v I__7352 (
            .O(N__46679),
            .I(N__46650));
    LocalMux I__7351 (
            .O(N__46676),
            .I(N__46643));
    LocalMux I__7350 (
            .O(N__46673),
            .I(N__46643));
    Span4Mux_h I__7349 (
            .O(N__46670),
            .I(N__46643));
    Span4Mux_v I__7348 (
            .O(N__46663),
            .I(N__46640));
    Span12Mux_v I__7347 (
            .O(N__46650),
            .I(N__46637));
    Span4Mux_v I__7346 (
            .O(N__46643),
            .I(N__46634));
    Odrv4 I__7345 (
            .O(N__46640),
            .I(dc32_fifo_data_in_13));
    Odrv12 I__7344 (
            .O(N__46637),
            .I(dc32_fifo_data_in_13));
    Odrv4 I__7343 (
            .O(N__46634),
            .I(dc32_fifo_data_in_13));
    InMux I__7342 (
            .O(N__46627),
            .I(N__46624));
    LocalMux I__7341 (
            .O(N__46624),
            .I(N__46621));
    Span4Mux_v I__7340 (
            .O(N__46621),
            .I(N__46617));
    InMux I__7339 (
            .O(N__46620),
            .I(N__46614));
    Odrv4 I__7338 (
            .O(N__46617),
            .I(REG_mem_45_13));
    LocalMux I__7337 (
            .O(N__46614),
            .I(REG_mem_45_13));
    InMux I__7336 (
            .O(N__46609),
            .I(N__46606));
    LocalMux I__7335 (
            .O(N__46606),
            .I(N__46603));
    Span4Mux_v I__7334 (
            .O(N__46603),
            .I(N__46600));
    Span4Mux_h I__7333 (
            .O(N__46600),
            .I(N__46596));
    InMux I__7332 (
            .O(N__46599),
            .I(N__46593));
    Odrv4 I__7331 (
            .O(N__46596),
            .I(REG_mem_50_12));
    LocalMux I__7330 (
            .O(N__46593),
            .I(REG_mem_50_12));
    InMux I__7329 (
            .O(N__46588),
            .I(N__46576));
    CascadeMux I__7328 (
            .O(N__46587),
            .I(N__46573));
    CascadeMux I__7327 (
            .O(N__46586),
            .I(N__46570));
    InMux I__7326 (
            .O(N__46585),
            .I(N__46562));
    InMux I__7325 (
            .O(N__46584),
            .I(N__46555));
    InMux I__7324 (
            .O(N__46583),
            .I(N__46555));
    InMux I__7323 (
            .O(N__46582),
            .I(N__46555));
    InMux I__7322 (
            .O(N__46581),
            .I(N__46549));
    InMux I__7321 (
            .O(N__46580),
            .I(N__46545));
    InMux I__7320 (
            .O(N__46579),
            .I(N__46542));
    LocalMux I__7319 (
            .O(N__46576),
            .I(N__46534));
    InMux I__7318 (
            .O(N__46573),
            .I(N__46531));
    InMux I__7317 (
            .O(N__46570),
            .I(N__46526));
    InMux I__7316 (
            .O(N__46569),
            .I(N__46526));
    InMux I__7315 (
            .O(N__46568),
            .I(N__46521));
    InMux I__7314 (
            .O(N__46567),
            .I(N__46521));
    InMux I__7313 (
            .O(N__46566),
            .I(N__46516));
    InMux I__7312 (
            .O(N__46565),
            .I(N__46516));
    LocalMux I__7311 (
            .O(N__46562),
            .I(N__46513));
    LocalMux I__7310 (
            .O(N__46555),
            .I(N__46510));
    InMux I__7309 (
            .O(N__46554),
            .I(N__46501));
    InMux I__7308 (
            .O(N__46553),
            .I(N__46501));
    InMux I__7307 (
            .O(N__46552),
            .I(N__46501));
    LocalMux I__7306 (
            .O(N__46549),
            .I(N__46498));
    CascadeMux I__7305 (
            .O(N__46548),
            .I(N__46494));
    LocalMux I__7304 (
            .O(N__46545),
            .I(N__46488));
    LocalMux I__7303 (
            .O(N__46542),
            .I(N__46484));
    InMux I__7302 (
            .O(N__46541),
            .I(N__46473));
    InMux I__7301 (
            .O(N__46540),
            .I(N__46473));
    InMux I__7300 (
            .O(N__46539),
            .I(N__46473));
    InMux I__7299 (
            .O(N__46538),
            .I(N__46473));
    CascadeMux I__7298 (
            .O(N__46537),
            .I(N__46465));
    Span4Mux_h I__7297 (
            .O(N__46534),
            .I(N__46457));
    LocalMux I__7296 (
            .O(N__46531),
            .I(N__46457));
    LocalMux I__7295 (
            .O(N__46526),
            .I(N__46448));
    LocalMux I__7294 (
            .O(N__46521),
            .I(N__46443));
    LocalMux I__7293 (
            .O(N__46516),
            .I(N__46443));
    Span4Mux_h I__7292 (
            .O(N__46513),
            .I(N__46438));
    Span4Mux_v I__7291 (
            .O(N__46510),
            .I(N__46438));
    InMux I__7290 (
            .O(N__46509),
            .I(N__46433));
    InMux I__7289 (
            .O(N__46508),
            .I(N__46433));
    LocalMux I__7288 (
            .O(N__46501),
            .I(N__46430));
    Span4Mux_v I__7287 (
            .O(N__46498),
            .I(N__46427));
    InMux I__7286 (
            .O(N__46497),
            .I(N__46416));
    InMux I__7285 (
            .O(N__46494),
            .I(N__46416));
    InMux I__7284 (
            .O(N__46493),
            .I(N__46416));
    InMux I__7283 (
            .O(N__46492),
            .I(N__46416));
    InMux I__7282 (
            .O(N__46491),
            .I(N__46416));
    Span4Mux_v I__7281 (
            .O(N__46488),
            .I(N__46413));
    InMux I__7280 (
            .O(N__46487),
            .I(N__46410));
    Span4Mux_h I__7279 (
            .O(N__46484),
            .I(N__46403));
    InMux I__7278 (
            .O(N__46483),
            .I(N__46398));
    InMux I__7277 (
            .O(N__46482),
            .I(N__46398));
    LocalMux I__7276 (
            .O(N__46473),
            .I(N__46391));
    CascadeMux I__7275 (
            .O(N__46472),
            .I(N__46388));
    InMux I__7274 (
            .O(N__46471),
            .I(N__46381));
    InMux I__7273 (
            .O(N__46470),
            .I(N__46373));
    InMux I__7272 (
            .O(N__46469),
            .I(N__46373));
    InMux I__7271 (
            .O(N__46468),
            .I(N__46373));
    InMux I__7270 (
            .O(N__46465),
            .I(N__46370));
    InMux I__7269 (
            .O(N__46464),
            .I(N__46363));
    InMux I__7268 (
            .O(N__46463),
            .I(N__46363));
    InMux I__7267 (
            .O(N__46462),
            .I(N__46363));
    Span4Mux_v I__7266 (
            .O(N__46457),
            .I(N__46360));
    InMux I__7265 (
            .O(N__46456),
            .I(N__46357));
    InMux I__7264 (
            .O(N__46455),
            .I(N__46350));
    InMux I__7263 (
            .O(N__46454),
            .I(N__46350));
    InMux I__7262 (
            .O(N__46453),
            .I(N__46350));
    InMux I__7261 (
            .O(N__46452),
            .I(N__46344));
    InMux I__7260 (
            .O(N__46451),
            .I(N__46341));
    Span4Mux_v I__7259 (
            .O(N__46448),
            .I(N__46336));
    Span4Mux_v I__7258 (
            .O(N__46443),
            .I(N__46336));
    Span4Mux_h I__7257 (
            .O(N__46438),
            .I(N__46327));
    LocalMux I__7256 (
            .O(N__46433),
            .I(N__46327));
    Span4Mux_h I__7255 (
            .O(N__46430),
            .I(N__46327));
    Span4Mux_h I__7254 (
            .O(N__46427),
            .I(N__46327));
    LocalMux I__7253 (
            .O(N__46416),
            .I(N__46320));
    Span4Mux_h I__7252 (
            .O(N__46413),
            .I(N__46320));
    LocalMux I__7251 (
            .O(N__46410),
            .I(N__46320));
    InMux I__7250 (
            .O(N__46409),
            .I(N__46317));
    InMux I__7249 (
            .O(N__46408),
            .I(N__46312));
    InMux I__7248 (
            .O(N__46407),
            .I(N__46312));
    InMux I__7247 (
            .O(N__46406),
            .I(N__46309));
    Span4Mux_v I__7246 (
            .O(N__46403),
            .I(N__46303));
    LocalMux I__7245 (
            .O(N__46398),
            .I(N__46303));
    InMux I__7244 (
            .O(N__46397),
            .I(N__46300));
    InMux I__7243 (
            .O(N__46396),
            .I(N__46293));
    InMux I__7242 (
            .O(N__46395),
            .I(N__46293));
    InMux I__7241 (
            .O(N__46394),
            .I(N__46293));
    Span4Mux_v I__7240 (
            .O(N__46391),
            .I(N__46290));
    InMux I__7239 (
            .O(N__46388),
            .I(N__46287));
    InMux I__7238 (
            .O(N__46387),
            .I(N__46278));
    InMux I__7237 (
            .O(N__46386),
            .I(N__46278));
    InMux I__7236 (
            .O(N__46385),
            .I(N__46278));
    InMux I__7235 (
            .O(N__46384),
            .I(N__46278));
    LocalMux I__7234 (
            .O(N__46381),
            .I(N__46275));
    InMux I__7233 (
            .O(N__46380),
            .I(N__46272));
    LocalMux I__7232 (
            .O(N__46373),
            .I(N__46269));
    LocalMux I__7231 (
            .O(N__46370),
            .I(N__46264));
    LocalMux I__7230 (
            .O(N__46363),
            .I(N__46264));
    Sp12to4 I__7229 (
            .O(N__46360),
            .I(N__46261));
    LocalMux I__7228 (
            .O(N__46357),
            .I(N__46256));
    LocalMux I__7227 (
            .O(N__46350),
            .I(N__46256));
    InMux I__7226 (
            .O(N__46349),
            .I(N__46253));
    InMux I__7225 (
            .O(N__46348),
            .I(N__46248));
    InMux I__7224 (
            .O(N__46347),
            .I(N__46248));
    LocalMux I__7223 (
            .O(N__46344),
            .I(N__46245));
    LocalMux I__7222 (
            .O(N__46341),
            .I(N__46236));
    Span4Mux_h I__7221 (
            .O(N__46336),
            .I(N__46236));
    Span4Mux_v I__7220 (
            .O(N__46327),
            .I(N__46236));
    Span4Mux_v I__7219 (
            .O(N__46320),
            .I(N__46236));
    LocalMux I__7218 (
            .O(N__46317),
            .I(N__46229));
    LocalMux I__7217 (
            .O(N__46312),
            .I(N__46229));
    LocalMux I__7216 (
            .O(N__46309),
            .I(N__46229));
    InMux I__7215 (
            .O(N__46308),
            .I(N__46226));
    Sp12to4 I__7214 (
            .O(N__46303),
            .I(N__46211));
    LocalMux I__7213 (
            .O(N__46300),
            .I(N__46211));
    LocalMux I__7212 (
            .O(N__46293),
            .I(N__46211));
    Sp12to4 I__7211 (
            .O(N__46290),
            .I(N__46211));
    LocalMux I__7210 (
            .O(N__46287),
            .I(N__46211));
    LocalMux I__7209 (
            .O(N__46278),
            .I(N__46211));
    Span12Mux_h I__7208 (
            .O(N__46275),
            .I(N__46211));
    LocalMux I__7207 (
            .O(N__46272),
            .I(N__46198));
    Span12Mux_h I__7206 (
            .O(N__46269),
            .I(N__46198));
    Span12Mux_h I__7205 (
            .O(N__46264),
            .I(N__46198));
    Span12Mux_v I__7204 (
            .O(N__46261),
            .I(N__46198));
    Sp12to4 I__7203 (
            .O(N__46256),
            .I(N__46198));
    LocalMux I__7202 (
            .O(N__46253),
            .I(N__46198));
    LocalMux I__7201 (
            .O(N__46248),
            .I(N__46191));
    Span4Mux_h I__7200 (
            .O(N__46245),
            .I(N__46191));
    Span4Mux_v I__7199 (
            .O(N__46236),
            .I(N__46191));
    Span12Mux_v I__7198 (
            .O(N__46229),
            .I(N__46188));
    LocalMux I__7197 (
            .O(N__46226),
            .I(N__46183));
    Span12Mux_v I__7196 (
            .O(N__46211),
            .I(N__46183));
    Span12Mux_v I__7195 (
            .O(N__46198),
            .I(N__46180));
    Span4Mux_v I__7194 (
            .O(N__46191),
            .I(N__46177));
    Odrv12 I__7193 (
            .O(N__46188),
            .I(dc32_fifo_data_in_12));
    Odrv12 I__7192 (
            .O(N__46183),
            .I(dc32_fifo_data_in_12));
    Odrv12 I__7191 (
            .O(N__46180),
            .I(dc32_fifo_data_in_12));
    Odrv4 I__7190 (
            .O(N__46177),
            .I(dc32_fifo_data_in_12));
    InMux I__7189 (
            .O(N__46168),
            .I(N__46164));
    InMux I__7188 (
            .O(N__46167),
            .I(N__46161));
    LocalMux I__7187 (
            .O(N__46164),
            .I(REG_mem_6_12));
    LocalMux I__7186 (
            .O(N__46161),
            .I(REG_mem_6_12));
    CascadeMux I__7185 (
            .O(N__46156),
            .I(N__46153));
    InMux I__7184 (
            .O(N__46153),
            .I(N__46149));
    InMux I__7183 (
            .O(N__46152),
            .I(N__46146));
    LocalMux I__7182 (
            .O(N__46149),
            .I(REG_mem_5_13));
    LocalMux I__7181 (
            .O(N__46146),
            .I(REG_mem_5_13));
    InMux I__7180 (
            .O(N__46141),
            .I(N__46138));
    LocalMux I__7179 (
            .O(N__46138),
            .I(N__46135));
    Span4Mux_v I__7178 (
            .O(N__46135),
            .I(N__46132));
    Odrv4 I__7177 (
            .O(N__46132),
            .I(rd_grey_sync_r_4));
    InMux I__7176 (
            .O(N__46129),
            .I(N__46126));
    LocalMux I__7175 (
            .O(N__46126),
            .I(rp_sync1_r_4));
    InMux I__7174 (
            .O(N__46123),
            .I(N__46120));
    LocalMux I__7173 (
            .O(N__46120),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_4 ));
    InMux I__7172 (
            .O(N__46117),
            .I(N__46113));
    InMux I__7171 (
            .O(N__46116),
            .I(N__46110));
    LocalMux I__7170 (
            .O(N__46113),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_5 ));
    LocalMux I__7169 (
            .O(N__46110),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_5 ));
    CascadeMux I__7168 (
            .O(N__46105),
            .I(N__46102));
    InMux I__7167 (
            .O(N__46102),
            .I(N__46099));
    LocalMux I__7166 (
            .O(N__46099),
            .I(N__46095));
    CascadeMux I__7165 (
            .O(N__46098),
            .I(N__46092));
    Span4Mux_h I__7164 (
            .O(N__46095),
            .I(N__46088));
    InMux I__7163 (
            .O(N__46092),
            .I(N__46083));
    InMux I__7162 (
            .O(N__46091),
            .I(N__46083));
    Odrv4 I__7161 (
            .O(N__46088),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_5 ));
    LocalMux I__7160 (
            .O(N__46083),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_5 ));
    InMux I__7159 (
            .O(N__46078),
            .I(N__46075));
    LocalMux I__7158 (
            .O(N__46075),
            .I(N__46072));
    Span4Mux_h I__7157 (
            .O(N__46072),
            .I(N__46069));
    Odrv4 I__7156 (
            .O(N__46069),
            .I(rd_grey_sync_r_5));
    InMux I__7155 (
            .O(N__46066),
            .I(N__46063));
    LocalMux I__7154 (
            .O(N__46063),
            .I(rp_sync1_r_5));
    CascadeMux I__7153 (
            .O(N__46060),
            .I(N__46057));
    InMux I__7152 (
            .O(N__46057),
            .I(N__46054));
    LocalMux I__7151 (
            .O(N__46054),
            .I(N__46050));
    InMux I__7150 (
            .O(N__46053),
            .I(N__46047));
    Odrv4 I__7149 (
            .O(N__46050),
            .I(REG_mem_6_13));
    LocalMux I__7148 (
            .O(N__46047),
            .I(REG_mem_6_13));
    InMux I__7147 (
            .O(N__46042),
            .I(N__46036));
    InMux I__7146 (
            .O(N__46041),
            .I(N__46036));
    LocalMux I__7145 (
            .O(N__46036),
            .I(REG_mem_51_11));
    CascadeMux I__7144 (
            .O(N__46033),
            .I(N__46030));
    InMux I__7143 (
            .O(N__46030),
            .I(N__46027));
    LocalMux I__7142 (
            .O(N__46027),
            .I(N__46023));
    CascadeMux I__7141 (
            .O(N__46026),
            .I(N__46020));
    Span4Mux_h I__7140 (
            .O(N__46023),
            .I(N__46017));
    InMux I__7139 (
            .O(N__46020),
            .I(N__46014));
    Odrv4 I__7138 (
            .O(N__46017),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_11 ));
    LocalMux I__7137 (
            .O(N__46014),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_11 ));
    InMux I__7136 (
            .O(N__46009),
            .I(N__46006));
    LocalMux I__7135 (
            .O(N__46006),
            .I(N__46003));
    Span4Mux_v I__7134 (
            .O(N__46003),
            .I(N__45999));
    InMux I__7133 (
            .O(N__46002),
            .I(N__45996));
    Odrv4 I__7132 (
            .O(N__45999),
            .I(REG_mem_5_11));
    LocalMux I__7131 (
            .O(N__45996),
            .I(REG_mem_5_11));
    InMux I__7130 (
            .O(N__45991),
            .I(N__45985));
    InMux I__7129 (
            .O(N__45990),
            .I(N__45985));
    LocalMux I__7128 (
            .O(N__45985),
            .I(REG_mem_37_13));
    CascadeMux I__7127 (
            .O(N__45982),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13838_cascade_ ));
    InMux I__7126 (
            .O(N__45979),
            .I(N__45976));
    LocalMux I__7125 (
            .O(N__45976),
            .I(N__45972));
    InMux I__7124 (
            .O(N__45975),
            .I(N__45969));
    Span4Mux_v I__7123 (
            .O(N__45972),
            .I(N__45964));
    LocalMux I__7122 (
            .O(N__45969),
            .I(N__45964));
    Odrv4 I__7121 (
            .O(N__45964),
            .I(REG_mem_36_13));
    CascadeMux I__7120 (
            .O(N__45961),
            .I(N__45958));
    InMux I__7119 (
            .O(N__45958),
            .I(N__45955));
    LocalMux I__7118 (
            .O(N__45955),
            .I(N__45952));
    Span4Mux_v I__7117 (
            .O(N__45952),
            .I(N__45949));
    Odrv4 I__7116 (
            .O(N__45949),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12189 ));
    InMux I__7115 (
            .O(N__45946),
            .I(N__45943));
    LocalMux I__7114 (
            .O(N__45943),
            .I(N__45939));
    InMux I__7113 (
            .O(N__45942),
            .I(N__45936));
    Span4Mux_h I__7112 (
            .O(N__45939),
            .I(N__45930));
    LocalMux I__7111 (
            .O(N__45936),
            .I(N__45927));
    InMux I__7110 (
            .O(N__45935),
            .I(N__45924));
    InMux I__7109 (
            .O(N__45934),
            .I(N__45919));
    InMux I__7108 (
            .O(N__45933),
            .I(N__45919));
    Odrv4 I__7107 (
            .O(N__45930),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_4 ));
    Odrv4 I__7106 (
            .O(N__45927),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_4 ));
    LocalMux I__7105 (
            .O(N__45924),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_4 ));
    LocalMux I__7104 (
            .O(N__45919),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_4 ));
    InMux I__7103 (
            .O(N__45910),
            .I(N__45904));
    InMux I__7102 (
            .O(N__45909),
            .I(N__45904));
    LocalMux I__7101 (
            .O(N__45904),
            .I(REG_mem_38_13));
    CascadeMux I__7100 (
            .O(N__45901),
            .I(N__45898));
    InMux I__7099 (
            .O(N__45898),
            .I(N__45892));
    InMux I__7098 (
            .O(N__45897),
            .I(N__45892));
    LocalMux I__7097 (
            .O(N__45892),
            .I(N__45889));
    Odrv4 I__7096 (
            .O(N__45889),
            .I(REG_mem_39_13));
    InMux I__7095 (
            .O(N__45886),
            .I(N__45880));
    InMux I__7094 (
            .O(N__45885),
            .I(N__45880));
    LocalMux I__7093 (
            .O(N__45880),
            .I(REG_mem_14_12));
    InMux I__7092 (
            .O(N__45877),
            .I(N__45871));
    InMux I__7091 (
            .O(N__45876),
            .I(N__45871));
    LocalMux I__7090 (
            .O(N__45871),
            .I(REG_mem_15_12));
    InMux I__7089 (
            .O(N__45868),
            .I(N__45865));
    LocalMux I__7088 (
            .O(N__45865),
            .I(N__45861));
    InMux I__7087 (
            .O(N__45864),
            .I(N__45858));
    Odrv12 I__7086 (
            .O(N__45861),
            .I(REG_mem_50_11));
    LocalMux I__7085 (
            .O(N__45858),
            .I(REG_mem_50_11));
    InMux I__7084 (
            .O(N__45853),
            .I(N__45847));
    InMux I__7083 (
            .O(N__45852),
            .I(N__45847));
    LocalMux I__7082 (
            .O(N__45847),
            .I(REG_mem_49_11));
    CascadeMux I__7081 (
            .O(N__45844),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14204_cascade_ ));
    InMux I__7080 (
            .O(N__45841),
            .I(N__45837));
    InMux I__7079 (
            .O(N__45840),
            .I(N__45834));
    LocalMux I__7078 (
            .O(N__45837),
            .I(N__45829));
    LocalMux I__7077 (
            .O(N__45834),
            .I(N__45829));
    Odrv4 I__7076 (
            .O(N__45829),
            .I(REG_mem_48_11));
    InMux I__7075 (
            .O(N__45826),
            .I(N__45823));
    LocalMux I__7074 (
            .O(N__45823),
            .I(N__45820));
    Span4Mux_v I__7073 (
            .O(N__45820),
            .I(N__45816));
    InMux I__7072 (
            .O(N__45819),
            .I(N__45813));
    Odrv4 I__7071 (
            .O(N__45816),
            .I(REG_mem_50_13));
    LocalMux I__7070 (
            .O(N__45813),
            .I(REG_mem_50_13));
    InMux I__7069 (
            .O(N__45808),
            .I(N__45805));
    LocalMux I__7068 (
            .O(N__45805),
            .I(N__45802));
    Span4Mux_v I__7067 (
            .O(N__45802),
            .I(N__45798));
    InMux I__7066 (
            .O(N__45801),
            .I(N__45795));
    Odrv4 I__7065 (
            .O(N__45798),
            .I(REG_mem_47_13));
    LocalMux I__7064 (
            .O(N__45795),
            .I(REG_mem_47_13));
    InMux I__7063 (
            .O(N__45790),
            .I(N__45787));
    LocalMux I__7062 (
            .O(N__45787),
            .I(N__45784));
    Span4Mux_v I__7061 (
            .O(N__45784),
            .I(N__45781));
    Span4Mux_h I__7060 (
            .O(N__45781),
            .I(N__45778));
    Span4Mux_h I__7059 (
            .O(N__45778),
            .I(N__45774));
    InMux I__7058 (
            .O(N__45777),
            .I(N__45771));
    Odrv4 I__7057 (
            .O(N__45774),
            .I(REG_mem_14_7));
    LocalMux I__7056 (
            .O(N__45771),
            .I(REG_mem_14_7));
    InMux I__7055 (
            .O(N__45766),
            .I(N__45763));
    LocalMux I__7054 (
            .O(N__45763),
            .I(N__45760));
    Span4Mux_v I__7053 (
            .O(N__45760),
            .I(N__45756));
    InMux I__7052 (
            .O(N__45759),
            .I(N__45753));
    Span4Mux_h I__7051 (
            .O(N__45756),
            .I(N__45748));
    LocalMux I__7050 (
            .O(N__45753),
            .I(N__45748));
    Odrv4 I__7049 (
            .O(N__45748),
            .I(REG_mem_46_12));
    CascadeMux I__7048 (
            .O(N__45745),
            .I(N__45741));
    InMux I__7047 (
            .O(N__45744),
            .I(N__45736));
    InMux I__7046 (
            .O(N__45741),
            .I(N__45736));
    LocalMux I__7045 (
            .O(N__45736),
            .I(N__45733));
    Odrv4 I__7044 (
            .O(N__45733),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_11 ));
    InMux I__7043 (
            .O(N__45730),
            .I(N__45727));
    LocalMux I__7042 (
            .O(N__45727),
            .I(N__45724));
    Span4Mux_h I__7041 (
            .O(N__45724),
            .I(N__45721));
    Span4Mux_h I__7040 (
            .O(N__45721),
            .I(N__45717));
    InMux I__7039 (
            .O(N__45720),
            .I(N__45714));
    Odrv4 I__7038 (
            .O(N__45717),
            .I(REG_mem_58_3));
    LocalMux I__7037 (
            .O(N__45714),
            .I(REG_mem_58_3));
    InMux I__7036 (
            .O(N__45709),
            .I(N__45706));
    LocalMux I__7035 (
            .O(N__45706),
            .I(N__45703));
    Span4Mux_v I__7034 (
            .O(N__45703),
            .I(N__45700));
    Span4Mux_h I__7033 (
            .O(N__45700),
            .I(N__45696));
    InMux I__7032 (
            .O(N__45699),
            .I(N__45693));
    Odrv4 I__7031 (
            .O(N__45696),
            .I(REG_mem_31_13));
    LocalMux I__7030 (
            .O(N__45693),
            .I(REG_mem_31_13));
    CascadeMux I__7029 (
            .O(N__45688),
            .I(N__45685));
    InMux I__7028 (
            .O(N__45685),
            .I(N__45682));
    LocalMux I__7027 (
            .O(N__45682),
            .I(N__45678));
    InMux I__7026 (
            .O(N__45681),
            .I(N__45675));
    Odrv12 I__7025 (
            .O(N__45678),
            .I(REG_mem_46_11));
    LocalMux I__7024 (
            .O(N__45675),
            .I(REG_mem_46_11));
    InMux I__7023 (
            .O(N__45670),
            .I(N__45664));
    InMux I__7022 (
            .O(N__45669),
            .I(N__45664));
    LocalMux I__7021 (
            .O(N__45664),
            .I(REG_mem_13_12));
    CascadeMux I__7020 (
            .O(N__45661),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13412_cascade_ ));
    InMux I__7019 (
            .O(N__45658),
            .I(N__45655));
    LocalMux I__7018 (
            .O(N__45655),
            .I(N__45652));
    Span4Mux_h I__7017 (
            .O(N__45652),
            .I(N__45649));
    Span4Mux_h I__7016 (
            .O(N__45649),
            .I(N__45646));
    Odrv4 I__7015 (
            .O(N__45646),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13415 ));
    InMux I__7014 (
            .O(N__45643),
            .I(N__45637));
    InMux I__7013 (
            .O(N__45642),
            .I(N__45637));
    LocalMux I__7012 (
            .O(N__45637),
            .I(REG_mem_12_12));
    CascadeMux I__7011 (
            .O(N__45634),
            .I(N__45631));
    InMux I__7010 (
            .O(N__45631),
            .I(N__45627));
    InMux I__7009 (
            .O(N__45630),
            .I(N__45624));
    LocalMux I__7008 (
            .O(N__45627),
            .I(REG_mem_14_3));
    LocalMux I__7007 (
            .O(N__45624),
            .I(REG_mem_14_3));
    InMux I__7006 (
            .O(N__45619),
            .I(N__45616));
    LocalMux I__7005 (
            .O(N__45616),
            .I(N__45612));
    InMux I__7004 (
            .O(N__45615),
            .I(N__45609));
    Odrv12 I__7003 (
            .O(N__45612),
            .I(REG_mem_13_3));
    LocalMux I__7002 (
            .O(N__45609),
            .I(REG_mem_13_3));
    InMux I__7001 (
            .O(N__45604),
            .I(N__45601));
    LocalMux I__7000 (
            .O(N__45601),
            .I(N__45598));
    Span4Mux_v I__6999 (
            .O(N__45598),
            .I(N__45595));
    Span4Mux_v I__6998 (
            .O(N__45595),
            .I(N__45591));
    InMux I__6997 (
            .O(N__45594),
            .I(N__45588));
    Odrv4 I__6996 (
            .O(N__45591),
            .I(REG_mem_15_13));
    LocalMux I__6995 (
            .O(N__45588),
            .I(REG_mem_15_13));
    InMux I__6994 (
            .O(N__45583),
            .I(N__45580));
    LocalMux I__6993 (
            .O(N__45580),
            .I(N__45577));
    Span4Mux_h I__6992 (
            .O(N__45577),
            .I(N__45574));
    Span4Mux_v I__6991 (
            .O(N__45574),
            .I(N__45570));
    InMux I__6990 (
            .O(N__45573),
            .I(N__45567));
    Odrv4 I__6989 (
            .O(N__45570),
            .I(REG_mem_43_13));
    LocalMux I__6988 (
            .O(N__45567),
            .I(REG_mem_43_13));
    InMux I__6987 (
            .O(N__45562),
            .I(N__45556));
    InMux I__6986 (
            .O(N__45561),
            .I(N__45549));
    InMux I__6985 (
            .O(N__45560),
            .I(N__45549));
    InMux I__6984 (
            .O(N__45559),
            .I(N__45549));
    LocalMux I__6983 (
            .O(N__45556),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n17 ));
    LocalMux I__6982 (
            .O(N__45549),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n17 ));
    InMux I__6981 (
            .O(N__45544),
            .I(N__45541));
    LocalMux I__6980 (
            .O(N__45541),
            .I(N__45538));
    Span4Mux_v I__6979 (
            .O(N__45538),
            .I(N__45535));
    Span4Mux_h I__6978 (
            .O(N__45535),
            .I(N__45531));
    InMux I__6977 (
            .O(N__45534),
            .I(N__45528));
    Odrv4 I__6976 (
            .O(N__45531),
            .I(REG_mem_47_11));
    LocalMux I__6975 (
            .O(N__45528),
            .I(REG_mem_47_11));
    InMux I__6974 (
            .O(N__45523),
            .I(N__45520));
    LocalMux I__6973 (
            .O(N__45520),
            .I(N__45517));
    Span4Mux_v I__6972 (
            .O(N__45517),
            .I(N__45514));
    Span4Mux_h I__6971 (
            .O(N__45514),
            .I(N__45510));
    InMux I__6970 (
            .O(N__45513),
            .I(N__45507));
    Odrv4 I__6969 (
            .O(N__45510),
            .I(REG_mem_38_3));
    LocalMux I__6968 (
            .O(N__45507),
            .I(REG_mem_38_3));
    InMux I__6967 (
            .O(N__45502),
            .I(N__45499));
    LocalMux I__6966 (
            .O(N__45499),
            .I(N__45496));
    Span4Mux_h I__6965 (
            .O(N__45496),
            .I(N__45493));
    Odrv4 I__6964 (
            .O(N__45493),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13754 ));
    InMux I__6963 (
            .O(N__45490),
            .I(N__45487));
    LocalMux I__6962 (
            .O(N__45487),
            .I(N__45484));
    Span4Mux_h I__6961 (
            .O(N__45484),
            .I(N__45481));
    Odrv4 I__6960 (
            .O(N__45481),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_w_6 ));
    CascadeMux I__6959 (
            .O(N__45478),
            .I(wr_addr_nxt_c_4_cascade_));
    InMux I__6958 (
            .O(N__45475),
            .I(N__45463));
    InMux I__6957 (
            .O(N__45474),
            .I(N__45463));
    InMux I__6956 (
            .O(N__45473),
            .I(N__45463));
    InMux I__6955 (
            .O(N__45472),
            .I(N__45463));
    LocalMux I__6954 (
            .O(N__45463),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n35 ));
    InMux I__6953 (
            .O(N__45460),
            .I(N__45455));
    InMux I__6952 (
            .O(N__45459),
            .I(N__45450));
    InMux I__6951 (
            .O(N__45458),
            .I(N__45450));
    LocalMux I__6950 (
            .O(N__45455),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n26_adj_1146 ));
    LocalMux I__6949 (
            .O(N__45450),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n26_adj_1146 ));
    CascadeMux I__6948 (
            .O(N__45445),
            .I(N__45442));
    InMux I__6947 (
            .O(N__45442),
            .I(N__45439));
    LocalMux I__6946 (
            .O(N__45439),
            .I(N__45436));
    Span4Mux_h I__6945 (
            .O(N__45436),
            .I(N__45433));
    Odrv4 I__6944 (
            .O(N__45433),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14306 ));
    InMux I__6943 (
            .O(N__45430),
            .I(N__45427));
    LocalMux I__6942 (
            .O(N__45427),
            .I(N__45424));
    Span4Mux_v I__6941 (
            .O(N__45424),
            .I(N__45421));
    Span4Mux_h I__6940 (
            .O(N__45421),
            .I(N__45417));
    InMux I__6939 (
            .O(N__45420),
            .I(N__45414));
    Odrv4 I__6938 (
            .O(N__45417),
            .I(REG_mem_5_9));
    LocalMux I__6937 (
            .O(N__45414),
            .I(REG_mem_5_9));
    InMux I__6936 (
            .O(N__45409),
            .I(N__45397));
    InMux I__6935 (
            .O(N__45408),
            .I(N__45397));
    InMux I__6934 (
            .O(N__45407),
            .I(N__45397));
    InMux I__6933 (
            .O(N__45406),
            .I(N__45397));
    LocalMux I__6932 (
            .O(N__45397),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n15 ));
    CascadeMux I__6931 (
            .O(N__45394),
            .I(N__45391));
    InMux I__6930 (
            .O(N__45391),
            .I(N__45388));
    LocalMux I__6929 (
            .O(N__45388),
            .I(N__45385));
    Span12Mux_v I__6928 (
            .O(N__45385),
            .I(N__45381));
    InMux I__6927 (
            .O(N__45384),
            .I(N__45378));
    Odrv12 I__6926 (
            .O(N__45381),
            .I(REG_mem_63_10));
    LocalMux I__6925 (
            .O(N__45378),
            .I(REG_mem_63_10));
    InMux I__6924 (
            .O(N__45373),
            .I(N__45369));
    InMux I__6923 (
            .O(N__45372),
            .I(N__45366));
    LocalMux I__6922 (
            .O(N__45369),
            .I(REG_mem_37_15));
    LocalMux I__6921 (
            .O(N__45366),
            .I(REG_mem_37_15));
    CascadeMux I__6920 (
            .O(N__45361),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13202_cascade_ ));
    InMux I__6919 (
            .O(N__45358),
            .I(N__45355));
    LocalMux I__6918 (
            .O(N__45355),
            .I(N__45352));
    Span4Mux_h I__6917 (
            .O(N__45352),
            .I(N__45349));
    Span4Mux_v I__6916 (
            .O(N__45349),
            .I(N__45346));
    Odrv4 I__6915 (
            .O(N__45346),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13205 ));
    InMux I__6914 (
            .O(N__45343),
            .I(N__45337));
    InMux I__6913 (
            .O(N__45342),
            .I(N__45337));
    LocalMux I__6912 (
            .O(N__45337),
            .I(REG_mem_12_9));
    InMux I__6911 (
            .O(N__45334),
            .I(N__45331));
    LocalMux I__6910 (
            .O(N__45331),
            .I(N__45327));
    InMux I__6909 (
            .O(N__45330),
            .I(N__45324));
    Odrv12 I__6908 (
            .O(N__45327),
            .I(REG_mem_7_15));
    LocalMux I__6907 (
            .O(N__45324),
            .I(REG_mem_7_15));
    InMux I__6906 (
            .O(N__45319),
            .I(N__45313));
    InMux I__6905 (
            .O(N__45318),
            .I(N__45313));
    LocalMux I__6904 (
            .O(N__45313),
            .I(REG_mem_51_2));
    InMux I__6903 (
            .O(N__45310),
            .I(N__45307));
    LocalMux I__6902 (
            .O(N__45307),
            .I(N__45304));
    Span4Mux_h I__6901 (
            .O(N__45304),
            .I(N__45301));
    Span4Mux_v I__6900 (
            .O(N__45301),
            .I(N__45297));
    InMux I__6899 (
            .O(N__45300),
            .I(N__45294));
    Odrv4 I__6898 (
            .O(N__45297),
            .I(REG_mem_38_9));
    LocalMux I__6897 (
            .O(N__45294),
            .I(REG_mem_38_9));
    CascadeMux I__6896 (
            .O(N__45289),
            .I(N__45286));
    InMux I__6895 (
            .O(N__45286),
            .I(N__45283));
    LocalMux I__6894 (
            .O(N__45283),
            .I(N__45279));
    InMux I__6893 (
            .O(N__45282),
            .I(N__45276));
    Odrv12 I__6892 (
            .O(N__45279),
            .I(REG_mem_41_9));
    LocalMux I__6891 (
            .O(N__45276),
            .I(REG_mem_41_9));
    InMux I__6890 (
            .O(N__45271),
            .I(N__45268));
    LocalMux I__6889 (
            .O(N__45268),
            .I(N__45264));
    InMux I__6888 (
            .O(N__45267),
            .I(N__45261));
    Odrv4 I__6887 (
            .O(N__45264),
            .I(REG_mem_49_15));
    LocalMux I__6886 (
            .O(N__45261),
            .I(REG_mem_49_15));
    InMux I__6885 (
            .O(N__45256),
            .I(N__45253));
    LocalMux I__6884 (
            .O(N__45253),
            .I(N__45249));
    InMux I__6883 (
            .O(N__45252),
            .I(N__45246));
    Odrv4 I__6882 (
            .O(N__45249),
            .I(REG_mem_48_15));
    LocalMux I__6881 (
            .O(N__45246),
            .I(REG_mem_48_15));
    InMux I__6880 (
            .O(N__45241),
            .I(N__45238));
    LocalMux I__6879 (
            .O(N__45238),
            .I(N__45235));
    Span4Mux_v I__6878 (
            .O(N__45235),
            .I(N__45232));
    Span4Mux_v I__6877 (
            .O(N__45232),
            .I(N__45229));
    Span4Mux_h I__6876 (
            .O(N__45229),
            .I(N__45225));
    InMux I__6875 (
            .O(N__45228),
            .I(N__45222));
    Odrv4 I__6874 (
            .O(N__45225),
            .I(REG_mem_45_11));
    LocalMux I__6873 (
            .O(N__45222),
            .I(REG_mem_45_11));
    CascadeMux I__6872 (
            .O(N__45217),
            .I(N__45214));
    InMux I__6871 (
            .O(N__45214),
            .I(N__45210));
    InMux I__6870 (
            .O(N__45213),
            .I(N__45207));
    LocalMux I__6869 (
            .O(N__45210),
            .I(N__45204));
    LocalMux I__6868 (
            .O(N__45207),
            .I(N__45201));
    Odrv12 I__6867 (
            .O(N__45204),
            .I(REG_mem_50_2));
    Odrv4 I__6866 (
            .O(N__45201),
            .I(REG_mem_50_2));
    InMux I__6865 (
            .O(N__45196),
            .I(N__45193));
    LocalMux I__6864 (
            .O(N__45193),
            .I(N__45190));
    Odrv4 I__6863 (
            .O(N__45190),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13976 ));
    CascadeMux I__6862 (
            .O(N__45187),
            .I(N__45184));
    InMux I__6861 (
            .O(N__45184),
            .I(N__45181));
    LocalMux I__6860 (
            .O(N__45181),
            .I(N__45178));
    Span4Mux_v I__6859 (
            .O(N__45178),
            .I(N__45175));
    Odrv4 I__6858 (
            .O(N__45175),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12014 ));
    InMux I__6857 (
            .O(N__45172),
            .I(N__45166));
    InMux I__6856 (
            .O(N__45171),
            .I(N__45166));
    LocalMux I__6855 (
            .O(N__45166),
            .I(REG_mem_47_15));
    InMux I__6854 (
            .O(N__45163),
            .I(N__45160));
    LocalMux I__6853 (
            .O(N__45160),
            .I(N__45157));
    Span4Mux_v I__6852 (
            .O(N__45157),
            .I(N__45153));
    InMux I__6851 (
            .O(N__45156),
            .I(N__45150));
    Odrv4 I__6850 (
            .O(N__45153),
            .I(REG_mem_45_15));
    LocalMux I__6849 (
            .O(N__45150),
            .I(REG_mem_45_15));
    CascadeMux I__6848 (
            .O(N__45145),
            .I(N__45142));
    InMux I__6847 (
            .O(N__45142),
            .I(N__45138));
    InMux I__6846 (
            .O(N__45141),
            .I(N__45135));
    LocalMux I__6845 (
            .O(N__45138),
            .I(REG_mem_15_0));
    LocalMux I__6844 (
            .O(N__45135),
            .I(REG_mem_15_0));
    CascadeMux I__6843 (
            .O(N__45130),
            .I(N__45127));
    InMux I__6842 (
            .O(N__45127),
            .I(N__45124));
    LocalMux I__6841 (
            .O(N__45124),
            .I(N__45121));
    Span4Mux_v I__6840 (
            .O(N__45121),
            .I(N__45117));
    InMux I__6839 (
            .O(N__45120),
            .I(N__45114));
    Odrv4 I__6838 (
            .O(N__45117),
            .I(REG_mem_49_2));
    LocalMux I__6837 (
            .O(N__45114),
            .I(REG_mem_49_2));
    InMux I__6836 (
            .O(N__45109),
            .I(N__45106));
    LocalMux I__6835 (
            .O(N__45106),
            .I(N__45103));
    Span4Mux_h I__6834 (
            .O(N__45103),
            .I(N__45099));
    InMux I__6833 (
            .O(N__45102),
            .I(N__45096));
    Odrv4 I__6832 (
            .O(N__45099),
            .I(REG_mem_10_15));
    LocalMux I__6831 (
            .O(N__45096),
            .I(REG_mem_10_15));
    InMux I__6830 (
            .O(N__45091),
            .I(N__45088));
    LocalMux I__6829 (
            .O(N__45088),
            .I(N__45085));
    Span4Mux_v I__6828 (
            .O(N__45085),
            .I(N__45082));
    Span4Mux_v I__6827 (
            .O(N__45082),
            .I(N__45078));
    CascadeMux I__6826 (
            .O(N__45081),
            .I(N__45075));
    Span4Mux_h I__6825 (
            .O(N__45078),
            .I(N__45072));
    InMux I__6824 (
            .O(N__45075),
            .I(N__45069));
    Odrv4 I__6823 (
            .O(N__45072),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_7 ));
    LocalMux I__6822 (
            .O(N__45069),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_7 ));
    InMux I__6821 (
            .O(N__45064),
            .I(N__45061));
    LocalMux I__6820 (
            .O(N__45061),
            .I(N__45057));
    InMux I__6819 (
            .O(N__45060),
            .I(N__45054));
    Odrv4 I__6818 (
            .O(N__45057),
            .I(REG_mem_12_0));
    LocalMux I__6817 (
            .O(N__45054),
            .I(REG_mem_12_0));
    CascadeMux I__6816 (
            .O(N__45049),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13835_cascade_ ));
    InMux I__6815 (
            .O(N__45046),
            .I(N__45043));
    LocalMux I__6814 (
            .O(N__45043),
            .I(N__45040));
    Odrv4 I__6813 (
            .O(N__45040),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12038 ));
    InMux I__6812 (
            .O(N__45037),
            .I(N__45034));
    LocalMux I__6811 (
            .O(N__45034),
            .I(N__45031));
    Span4Mux_v I__6810 (
            .O(N__45031),
            .I(N__45028));
    Sp12to4 I__6809 (
            .O(N__45028),
            .I(N__45025));
    Odrv12 I__6808 (
            .O(N__45025),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12019 ));
    CascadeMux I__6807 (
            .O(N__45022),
            .I(N__45019));
    InMux I__6806 (
            .O(N__45019),
            .I(N__45016));
    LocalMux I__6805 (
            .O(N__45016),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13832 ));
    InMux I__6804 (
            .O(N__45013),
            .I(N__45007));
    InMux I__6803 (
            .O(N__45012),
            .I(N__45007));
    LocalMux I__6802 (
            .O(N__45007),
            .I(REG_mem_13_0));
    InMux I__6801 (
            .O(N__45004),
            .I(N__44998));
    InMux I__6800 (
            .O(N__45003),
            .I(N__44998));
    LocalMux I__6799 (
            .O(N__44998),
            .I(REG_mem_14_0));
    CascadeMux I__6798 (
            .O(N__44995),
            .I(N__44992));
    InMux I__6797 (
            .O(N__44992),
            .I(N__44988));
    CascadeMux I__6796 (
            .O(N__44991),
            .I(N__44985));
    LocalMux I__6795 (
            .O(N__44988),
            .I(N__44982));
    InMux I__6794 (
            .O(N__44985),
            .I(N__44979));
    Odrv4 I__6793 (
            .O(N__44982),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_15 ));
    LocalMux I__6792 (
            .O(N__44979),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_15 ));
    CascadeMux I__6791 (
            .O(N__44974),
            .I(N__44971));
    InMux I__6790 (
            .O(N__44971),
            .I(N__44968));
    LocalMux I__6789 (
            .O(N__44968),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13040 ));
    InMux I__6788 (
            .O(N__44965),
            .I(N__44959));
    InMux I__6787 (
            .O(N__44964),
            .I(N__44959));
    LocalMux I__6786 (
            .O(N__44959),
            .I(REG_mem_5_15));
    InMux I__6785 (
            .O(N__44956),
            .I(N__44952));
    InMux I__6784 (
            .O(N__44955),
            .I(N__44949));
    LocalMux I__6783 (
            .O(N__44952),
            .I(REG_mem_42_5));
    LocalMux I__6782 (
            .O(N__44949),
            .I(REG_mem_42_5));
    InMux I__6781 (
            .O(N__44944),
            .I(N__44938));
    InMux I__6780 (
            .O(N__44943),
            .I(N__44938));
    LocalMux I__6779 (
            .O(N__44938),
            .I(REG_mem_6_15));
    InMux I__6778 (
            .O(N__44935),
            .I(N__44931));
    InMux I__6777 (
            .O(N__44934),
            .I(N__44928));
    LocalMux I__6776 (
            .O(N__44931),
            .I(N__44923));
    LocalMux I__6775 (
            .O(N__44928),
            .I(N__44923));
    Odrv4 I__6774 (
            .O(N__44923),
            .I(REG_mem_50_0));
    InMux I__6773 (
            .O(N__44920),
            .I(N__44917));
    LocalMux I__6772 (
            .O(N__44917),
            .I(N__44913));
    IoInMux I__6771 (
            .O(N__44916),
            .I(N__44910));
    Sp12to4 I__6770 (
            .O(N__44913),
            .I(N__44907));
    LocalMux I__6769 (
            .O(N__44910),
            .I(N__44904));
    Span12Mux_v I__6768 (
            .O(N__44907),
            .I(N__44901));
    IoSpan4Mux I__6767 (
            .O(N__44904),
            .I(N__44898));
    Span12Mux_h I__6766 (
            .O(N__44901),
            .I(N__44895));
    IoSpan4Mux I__6765 (
            .O(N__44898),
            .I(N__44892));
    Odrv12 I__6764 (
            .O(N__44895),
            .I(DEBUG_1_c_0_c));
    Odrv4 I__6763 (
            .O(N__44892),
            .I(DEBUG_1_c_0_c));
    InMux I__6762 (
            .O(N__44887),
            .I(N__44884));
    LocalMux I__6761 (
            .O(N__44884),
            .I(N__44881));
    Odrv12 I__6760 (
            .O(N__44881),
            .I(\usb3_if_inst.usb3_data_in_latched_0 ));
    InMux I__6759 (
            .O(N__44878),
            .I(N__44875));
    LocalMux I__6758 (
            .O(N__44875),
            .I(N__44871));
    InMux I__6757 (
            .O(N__44874),
            .I(N__44868));
    Odrv4 I__6756 (
            .O(N__44871),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_13 ));
    LocalMux I__6755 (
            .O(N__44868),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_13 ));
    InMux I__6754 (
            .O(N__44863),
            .I(N__44860));
    LocalMux I__6753 (
            .O(N__44860),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14144 ));
    CascadeMux I__6752 (
            .O(N__44857),
            .I(N__44854));
    InMux I__6751 (
            .O(N__44854),
            .I(N__44851));
    LocalMux I__6750 (
            .O(N__44851),
            .I(N__44847));
    CascadeMux I__6749 (
            .O(N__44850),
            .I(N__44844));
    Span4Mux_v I__6748 (
            .O(N__44847),
            .I(N__44841));
    InMux I__6747 (
            .O(N__44844),
            .I(N__44838));
    Odrv4 I__6746 (
            .O(N__44841),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_11 ));
    LocalMux I__6745 (
            .O(N__44838),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_11 ));
    InMux I__6744 (
            .O(N__44833),
            .I(N__44829));
    CascadeMux I__6743 (
            .O(N__44832),
            .I(N__44826));
    LocalMux I__6742 (
            .O(N__44829),
            .I(N__44823));
    InMux I__6741 (
            .O(N__44826),
            .I(N__44820));
    Odrv12 I__6740 (
            .O(N__44823),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_11 ));
    LocalMux I__6739 (
            .O(N__44820),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_11 ));
    InMux I__6738 (
            .O(N__44815),
            .I(N__44812));
    LocalMux I__6737 (
            .O(N__44812),
            .I(N__44808));
    CascadeMux I__6736 (
            .O(N__44811),
            .I(N__44805));
    Span4Mux_v I__6735 (
            .O(N__44808),
            .I(N__44802));
    InMux I__6734 (
            .O(N__44805),
            .I(N__44799));
    Odrv4 I__6733 (
            .O(N__44802),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_13 ));
    LocalMux I__6732 (
            .O(N__44799),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_13 ));
    InMux I__6731 (
            .O(N__44794),
            .I(N__44791));
    LocalMux I__6730 (
            .O(N__44791),
            .I(N__44788));
    Span4Mux_v I__6729 (
            .O(N__44788),
            .I(N__44784));
    CascadeMux I__6728 (
            .O(N__44787),
            .I(N__44781));
    Span4Mux_v I__6727 (
            .O(N__44784),
            .I(N__44778));
    InMux I__6726 (
            .O(N__44781),
            .I(N__44775));
    Odrv4 I__6725 (
            .O(N__44778),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_11 ));
    LocalMux I__6724 (
            .O(N__44775),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_11 ));
    CascadeMux I__6723 (
            .O(N__44770),
            .I(N__44767));
    InMux I__6722 (
            .O(N__44767),
            .I(N__44764));
    LocalMux I__6721 (
            .O(N__44764),
            .I(N__44760));
    InMux I__6720 (
            .O(N__44763),
            .I(N__44757));
    Odrv4 I__6719 (
            .O(N__44760),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_11 ));
    LocalMux I__6718 (
            .O(N__44757),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_11 ));
    InMux I__6717 (
            .O(N__44752),
            .I(N__44749));
    LocalMux I__6716 (
            .O(N__44749),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13874 ));
    InMux I__6715 (
            .O(N__44746),
            .I(N__44743));
    LocalMux I__6714 (
            .O(N__44743),
            .I(N__44740));
    Odrv4 I__6713 (
            .O(N__44740),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13877 ));
    InMux I__6712 (
            .O(N__44737),
            .I(N__44734));
    LocalMux I__6711 (
            .O(N__44734),
            .I(N__44730));
    CascadeMux I__6710 (
            .O(N__44733),
            .I(N__44727));
    Span4Mux_v I__6709 (
            .O(N__44730),
            .I(N__44724));
    InMux I__6708 (
            .O(N__44727),
            .I(N__44721));
    Odrv4 I__6707 (
            .O(N__44724),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_15 ));
    LocalMux I__6706 (
            .O(N__44721),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_15 ));
    InMux I__6705 (
            .O(N__44716),
            .I(N__44713));
    LocalMux I__6704 (
            .O(N__44713),
            .I(N__44709));
    InMux I__6703 (
            .O(N__44712),
            .I(N__44706));
    Odrv4 I__6702 (
            .O(N__44709),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_15 ));
    LocalMux I__6701 (
            .O(N__44706),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_15 ));
    CascadeMux I__6700 (
            .O(N__44701),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13043_cascade_ ));
    InMux I__6699 (
            .O(N__44698),
            .I(N__44695));
    LocalMux I__6698 (
            .O(N__44695),
            .I(N__44692));
    Span4Mux_h I__6697 (
            .O(N__44692),
            .I(N__44689));
    Span4Mux_h I__6696 (
            .O(N__44689),
            .I(N__44686));
    Span4Mux_v I__6695 (
            .O(N__44686),
            .I(N__44683));
    Odrv4 I__6694 (
            .O(N__44683),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12058 ));
    CascadeMux I__6693 (
            .O(N__44680),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12926_cascade_ ));
    InMux I__6692 (
            .O(N__44677),
            .I(N__44674));
    LocalMux I__6691 (
            .O(N__44674),
            .I(N__44670));
    InMux I__6690 (
            .O(N__44673),
            .I(N__44667));
    Odrv4 I__6689 (
            .O(N__44670),
            .I(REG_mem_4_15));
    LocalMux I__6688 (
            .O(N__44667),
            .I(REG_mem_4_15));
    InMux I__6687 (
            .O(N__44662),
            .I(N__44659));
    LocalMux I__6686 (
            .O(N__44659),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12929 ));
    InMux I__6685 (
            .O(N__44656),
            .I(N__44650));
    InMux I__6684 (
            .O(N__44655),
            .I(N__44650));
    LocalMux I__6683 (
            .O(N__44650),
            .I(REG_mem_49_13));
    CascadeMux I__6682 (
            .O(N__44647),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13592_cascade_ ));
    InMux I__6681 (
            .O(N__44644),
            .I(N__44641));
    LocalMux I__6680 (
            .O(N__44641),
            .I(N__44637));
    InMux I__6679 (
            .O(N__44640),
            .I(N__44634));
    Odrv4 I__6678 (
            .O(N__44637),
            .I(REG_mem_48_13));
    LocalMux I__6677 (
            .O(N__44634),
            .I(REG_mem_48_13));
    InMux I__6676 (
            .O(N__44629),
            .I(N__44626));
    LocalMux I__6675 (
            .O(N__44626),
            .I(N__44623));
    Span4Mux_v I__6674 (
            .O(N__44623),
            .I(N__44620));
    Odrv4 I__6673 (
            .O(N__44620),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12255 ));
    CascadeMux I__6672 (
            .O(N__44617),
            .I(N__44614));
    InMux I__6671 (
            .O(N__44614),
            .I(N__44611));
    LocalMux I__6670 (
            .O(N__44611),
            .I(N__44608));
    Odrv4 I__6669 (
            .O(N__44608),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12453 ));
    InMux I__6668 (
            .O(N__44605),
            .I(N__44602));
    LocalMux I__6667 (
            .O(N__44602),
            .I(N__44599));
    Odrv4 I__6666 (
            .O(N__44599),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13154 ));
    InMux I__6665 (
            .O(N__44596),
            .I(N__44593));
    LocalMux I__6664 (
            .O(N__44593),
            .I(N__44589));
    CascadeMux I__6663 (
            .O(N__44592),
            .I(N__44586));
    Span4Mux_v I__6662 (
            .O(N__44589),
            .I(N__44583));
    InMux I__6661 (
            .O(N__44586),
            .I(N__44580));
    Odrv4 I__6660 (
            .O(N__44583),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_11 ));
    LocalMux I__6659 (
            .O(N__44580),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_11 ));
    InMux I__6658 (
            .O(N__44575),
            .I(N__44571));
    InMux I__6657 (
            .O(N__44574),
            .I(N__44568));
    LocalMux I__6656 (
            .O(N__44571),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_13 ));
    LocalMux I__6655 (
            .O(N__44568),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_13 ));
    InMux I__6654 (
            .O(N__44563),
            .I(N__44560));
    LocalMux I__6653 (
            .O(N__44560),
            .I(N__44557));
    Span4Mux_h I__6652 (
            .O(N__44557),
            .I(N__44554));
    Span4Mux_v I__6651 (
            .O(N__44554),
            .I(N__44550));
    InMux I__6650 (
            .O(N__44553),
            .I(N__44547));
    Odrv4 I__6649 (
            .O(N__44550),
            .I(REG_mem_18_12));
    LocalMux I__6648 (
            .O(N__44547),
            .I(REG_mem_18_12));
    CascadeMux I__6647 (
            .O(N__44542),
            .I(N__44539));
    InMux I__6646 (
            .O(N__44539),
            .I(N__44536));
    LocalMux I__6645 (
            .O(N__44536),
            .I(N__44533));
    Span4Mux_v I__6644 (
            .O(N__44533),
            .I(N__44529));
    InMux I__6643 (
            .O(N__44532),
            .I(N__44526));
    Odrv4 I__6642 (
            .O(N__44529),
            .I(REG_mem_26_11));
    LocalMux I__6641 (
            .O(N__44526),
            .I(REG_mem_26_11));
    InMux I__6640 (
            .O(N__44521),
            .I(N__44517));
    CascadeMux I__6639 (
            .O(N__44520),
            .I(N__44514));
    LocalMux I__6638 (
            .O(N__44517),
            .I(N__44511));
    InMux I__6637 (
            .O(N__44514),
            .I(N__44508));
    Odrv4 I__6636 (
            .O(N__44511),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_11 ));
    LocalMux I__6635 (
            .O(N__44508),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_11 ));
    InMux I__6634 (
            .O(N__44503),
            .I(N__44500));
    LocalMux I__6633 (
            .O(N__44500),
            .I(N__44497));
    Span4Mux_h I__6632 (
            .O(N__44497),
            .I(N__44493));
    InMux I__6631 (
            .O(N__44496),
            .I(N__44490));
    Odrv4 I__6630 (
            .O(N__44493),
            .I(REG_mem_19_11));
    LocalMux I__6629 (
            .O(N__44490),
            .I(REG_mem_19_11));
    InMux I__6628 (
            .O(N__44485),
            .I(N__44479));
    InMux I__6627 (
            .O(N__44484),
            .I(N__44479));
    LocalMux I__6626 (
            .O(N__44479),
            .I(REG_mem_4_13));
    CascadeMux I__6625 (
            .O(N__44476),
            .I(N__44473));
    InMux I__6624 (
            .O(N__44473),
            .I(N__44470));
    LocalMux I__6623 (
            .O(N__44470),
            .I(N__44467));
    Span4Mux_h I__6622 (
            .O(N__44467),
            .I(N__44464));
    Odrv4 I__6621 (
            .O(N__44464),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12051 ));
    InMux I__6620 (
            .O(N__44461),
            .I(N__44458));
    LocalMux I__6619 (
            .O(N__44458),
            .I(N__44455));
    Span4Mux_v I__6618 (
            .O(N__44455),
            .I(N__44452));
    Span4Mux_v I__6617 (
            .O(N__44452),
            .I(N__44448));
    InMux I__6616 (
            .O(N__44451),
            .I(N__44445));
    Odrv4 I__6615 (
            .O(N__44448),
            .I(REG_mem_38_11));
    LocalMux I__6614 (
            .O(N__44445),
            .I(REG_mem_38_11));
    CascadeMux I__6613 (
            .O(N__44440),
            .I(N__44437));
    InMux I__6612 (
            .O(N__44437),
            .I(N__44434));
    LocalMux I__6611 (
            .O(N__44434),
            .I(N__44431));
    Span4Mux_h I__6610 (
            .O(N__44431),
            .I(N__44428));
    Odrv4 I__6609 (
            .O(N__44428),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13424 ));
    InMux I__6608 (
            .O(N__44425),
            .I(N__44422));
    LocalMux I__6607 (
            .O(N__44422),
            .I(N__44418));
    InMux I__6606 (
            .O(N__44421),
            .I(N__44415));
    Odrv12 I__6605 (
            .O(N__44418),
            .I(REG_mem_7_13));
    LocalMux I__6604 (
            .O(N__44415),
            .I(REG_mem_7_13));
    InMux I__6603 (
            .O(N__44410),
            .I(N__44407));
    LocalMux I__6602 (
            .O(N__44407),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14222 ));
    InMux I__6601 (
            .O(N__44404),
            .I(N__44400));
    InMux I__6600 (
            .O(N__44403),
            .I(N__44397));
    LocalMux I__6599 (
            .O(N__44400),
            .I(REG_mem_39_11));
    LocalMux I__6598 (
            .O(N__44397),
            .I(REG_mem_39_11));
    InMux I__6597 (
            .O(N__44392),
            .I(N__44387));
    CascadeMux I__6596 (
            .O(N__44391),
            .I(N__44382));
    InMux I__6595 (
            .O(N__44390),
            .I(N__44379));
    LocalMux I__6594 (
            .O(N__44387),
            .I(N__44376));
    InMux I__6593 (
            .O(N__44386),
            .I(N__44373));
    InMux I__6592 (
            .O(N__44385),
            .I(N__44368));
    InMux I__6591 (
            .O(N__44382),
            .I(N__44368));
    LocalMux I__6590 (
            .O(N__44379),
            .I(rd_addr_r_6));
    Odrv4 I__6589 (
            .O(N__44376),
            .I(rd_addr_r_6));
    LocalMux I__6588 (
            .O(N__44373),
            .I(rd_addr_r_6));
    LocalMux I__6587 (
            .O(N__44368),
            .I(rd_addr_r_6));
    CascadeMux I__6586 (
            .O(N__44359),
            .I(N__44356));
    InMux I__6585 (
            .O(N__44356),
            .I(N__44352));
    InMux I__6584 (
            .O(N__44355),
            .I(N__44349));
    LocalMux I__6583 (
            .O(N__44352),
            .I(REG_mem_51_13));
    LocalMux I__6582 (
            .O(N__44349),
            .I(REG_mem_51_13));
    InMux I__6581 (
            .O(N__44344),
            .I(N__44338));
    InMux I__6580 (
            .O(N__44343),
            .I(N__44338));
    LocalMux I__6579 (
            .O(N__44338),
            .I(REG_mem_8_12));
    InMux I__6578 (
            .O(N__44335),
            .I(N__44329));
    InMux I__6577 (
            .O(N__44334),
            .I(N__44329));
    LocalMux I__6576 (
            .O(N__44329),
            .I(REG_mem_10_12));
    InMux I__6575 (
            .O(N__44326),
            .I(N__44323));
    LocalMux I__6574 (
            .O(N__44323),
            .I(N__44320));
    Span4Mux_h I__6573 (
            .O(N__44320),
            .I(N__44316));
    InMux I__6572 (
            .O(N__44319),
            .I(N__44313));
    Odrv4 I__6571 (
            .O(N__44316),
            .I(REG_mem_41_13));
    LocalMux I__6570 (
            .O(N__44313),
            .I(REG_mem_41_13));
    CascadeMux I__6569 (
            .O(N__44308),
            .I(N__44305));
    InMux I__6568 (
            .O(N__44305),
            .I(N__44301));
    InMux I__6567 (
            .O(N__44304),
            .I(N__44298));
    LocalMux I__6566 (
            .O(N__44301),
            .I(REG_mem_7_12));
    LocalMux I__6565 (
            .O(N__44298),
            .I(REG_mem_7_12));
    InMux I__6564 (
            .O(N__44293),
            .I(N__44290));
    LocalMux I__6563 (
            .O(N__44290),
            .I(N__44287));
    Odrv12 I__6562 (
            .O(N__44287),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12299 ));
    InMux I__6561 (
            .O(N__44284),
            .I(N__44281));
    LocalMux I__6560 (
            .O(N__44281),
            .I(N__44278));
    Odrv4 I__6559 (
            .O(N__44278),
            .I(rp_sync1_r_3));
    InMux I__6558 (
            .O(N__44275),
            .I(N__44270));
    InMux I__6557 (
            .O(N__44274),
            .I(N__44265));
    InMux I__6556 (
            .O(N__44273),
            .I(N__44265));
    LocalMux I__6555 (
            .O(N__44270),
            .I(N__44262));
    LocalMux I__6554 (
            .O(N__44265),
            .I(N__44259));
    Odrv4 I__6553 (
            .O(N__44262),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_3 ));
    Odrv4 I__6552 (
            .O(N__44259),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_3 ));
    CascadeMux I__6551 (
            .O(N__44254),
            .I(N__44251));
    InMux I__6550 (
            .O(N__44251),
            .I(N__44248));
    LocalMux I__6549 (
            .O(N__44248),
            .I(N__44244));
    InMux I__6548 (
            .O(N__44247),
            .I(N__44241));
    Odrv4 I__6547 (
            .O(N__44244),
            .I(REG_mem_11_12));
    LocalMux I__6546 (
            .O(N__44241),
            .I(REG_mem_11_12));
    CascadeMux I__6545 (
            .O(N__44236),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_3_cascade_ ));
    InMux I__6544 (
            .O(N__44233),
            .I(N__44230));
    LocalMux I__6543 (
            .O(N__44230),
            .I(N__44227));
    Odrv4 I__6542 (
            .O(N__44227),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11384 ));
    InMux I__6541 (
            .O(N__44224),
            .I(N__44221));
    LocalMux I__6540 (
            .O(N__44221),
            .I(N__44218));
    Span4Mux_v I__6539 (
            .O(N__44218),
            .I(N__44215));
    Odrv4 I__6538 (
            .O(N__44215),
            .I(rd_grey_sync_r_2));
    InMux I__6537 (
            .O(N__44212),
            .I(N__44209));
    LocalMux I__6536 (
            .O(N__44209),
            .I(N__44205));
    InMux I__6535 (
            .O(N__44208),
            .I(N__44201));
    Span4Mux_h I__6534 (
            .O(N__44205),
            .I(N__44198));
    InMux I__6533 (
            .O(N__44204),
            .I(N__44195));
    LocalMux I__6532 (
            .O(N__44201),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_1 ));
    Odrv4 I__6531 (
            .O(N__44198),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_1 ));
    LocalMux I__6530 (
            .O(N__44195),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_1 ));
    InMux I__6529 (
            .O(N__44188),
            .I(N__44185));
    LocalMux I__6528 (
            .O(N__44185),
            .I(N__44182));
    Sp12to4 I__6527 (
            .O(N__44182),
            .I(N__44179));
    Odrv12 I__6526 (
            .O(N__44179),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11402 ));
    InMux I__6525 (
            .O(N__44176),
            .I(N__44173));
    LocalMux I__6524 (
            .O(N__44173),
            .I(rp_sync1_r_2));
    InMux I__6523 (
            .O(N__44170),
            .I(N__44167));
    LocalMux I__6522 (
            .O(N__44167),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_2 ));
    InMux I__6521 (
            .O(N__44164),
            .I(N__44161));
    LocalMux I__6520 (
            .O(N__44161),
            .I(N__44158));
    Span4Mux_h I__6519 (
            .O(N__44158),
            .I(N__44155));
    Odrv4 I__6518 (
            .O(N__44155),
            .I(rd_grey_sync_r_3));
    InMux I__6517 (
            .O(N__44152),
            .I(N__44148));
    InMux I__6516 (
            .O(N__44151),
            .I(N__44145));
    LocalMux I__6515 (
            .O(N__44148),
            .I(REG_mem_9_12));
    LocalMux I__6514 (
            .O(N__44145),
            .I(REG_mem_9_12));
    CascadeMux I__6513 (
            .O(N__44140),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13430_cascade_ ));
    InMux I__6512 (
            .O(N__44137),
            .I(N__44134));
    LocalMux I__6511 (
            .O(N__44134),
            .I(N__44131));
    Odrv12 I__6510 (
            .O(N__44131),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13433 ));
    CascadeMux I__6509 (
            .O(N__44128),
            .I(N__44125));
    InMux I__6508 (
            .O(N__44125),
            .I(N__44119));
    InMux I__6507 (
            .O(N__44124),
            .I(N__44119));
    LocalMux I__6506 (
            .O(N__44119),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_sig_diff0_w_1 ));
    InMux I__6505 (
            .O(N__44116),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10625 ));
    InMux I__6504 (
            .O(N__44113),
            .I(N__44107));
    InMux I__6503 (
            .O(N__44112),
            .I(N__44107));
    LocalMux I__6502 (
            .O(N__44107),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_sig_diff0_w_2 ));
    InMux I__6501 (
            .O(N__44104),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10626 ));
    InMux I__6500 (
            .O(N__44101),
            .I(N__44095));
    InMux I__6499 (
            .O(N__44100),
            .I(N__44095));
    LocalMux I__6498 (
            .O(N__44095),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_sig_diff0_w_3 ));
    InMux I__6497 (
            .O(N__44092),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10627 ));
    InMux I__6496 (
            .O(N__44089),
            .I(N__44086));
    LocalMux I__6495 (
            .O(N__44086),
            .I(N__44083));
    Odrv4 I__6494 (
            .O(N__44083),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n3_adj_1166 ));
    InMux I__6493 (
            .O(N__44080),
            .I(N__44077));
    LocalMux I__6492 (
            .O(N__44077),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11436 ));
    InMux I__6491 (
            .O(N__44074),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10628 ));
    InMux I__6490 (
            .O(N__44071),
            .I(N__44068));
    LocalMux I__6489 (
            .O(N__44068),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11463 ));
    InMux I__6488 (
            .O(N__44065),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10629 ));
    InMux I__6487 (
            .O(N__44062),
            .I(N__44059));
    LocalMux I__6486 (
            .O(N__44059),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11475 ));
    InMux I__6485 (
            .O(N__44056),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10630 ));
    InMux I__6484 (
            .O(N__44053),
            .I(N__44047));
    InMux I__6483 (
            .O(N__44052),
            .I(N__44047));
    LocalMux I__6482 (
            .O(N__44047),
            .I(N__44041));
    InMux I__6481 (
            .O(N__44046),
            .I(N__44038));
    InMux I__6480 (
            .O(N__44045),
            .I(N__44033));
    InMux I__6479 (
            .O(N__44044),
            .I(N__44033));
    Odrv4 I__6478 (
            .O(N__44041),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_2 ));
    LocalMux I__6477 (
            .O(N__44038),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_2 ));
    LocalMux I__6476 (
            .O(N__44033),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_2 ));
    InMux I__6475 (
            .O(N__44026),
            .I(N__44023));
    LocalMux I__6474 (
            .O(N__44023),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_3 ));
    CascadeMux I__6473 (
            .O(N__44020),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10784_cascade_ ));
    IoInMux I__6472 (
            .O(N__44017),
            .I(N__44014));
    LocalMux I__6471 (
            .O(N__44014),
            .I(N__44010));
    IoInMux I__6470 (
            .O(N__44013),
            .I(N__44007));
    IoSpan4Mux I__6469 (
            .O(N__44010),
            .I(N__44004));
    LocalMux I__6468 (
            .O(N__44007),
            .I(N__44001));
    Span4Mux_s0_h I__6467 (
            .O(N__44004),
            .I(N__43998));
    IoSpan4Mux I__6466 (
            .O(N__44001),
            .I(N__43995));
    Span4Mux_v I__6465 (
            .O(N__43998),
            .I(N__43992));
    Span4Mux_s3_h I__6464 (
            .O(N__43995),
            .I(N__43989));
    Span4Mux_h I__6463 (
            .O(N__43992),
            .I(N__43986));
    Span4Mux_h I__6462 (
            .O(N__43989),
            .I(N__43983));
    Span4Mux_h I__6461 (
            .O(N__43986),
            .I(N__43980));
    Span4Mux_h I__6460 (
            .O(N__43983),
            .I(N__43977));
    Span4Mux_h I__6459 (
            .O(N__43980),
            .I(N__43974));
    Span4Mux_v I__6458 (
            .O(N__43977),
            .I(N__43971));
    Span4Mux_h I__6457 (
            .O(N__43974),
            .I(N__43965));
    Span4Mux_v I__6456 (
            .O(N__43971),
            .I(N__43965));
    InMux I__6455 (
            .O(N__43970),
            .I(N__43962));
    Odrv4 I__6454 (
            .O(N__43965),
            .I(DEBUG_3_c));
    LocalMux I__6453 (
            .O(N__43962),
            .I(DEBUG_3_c));
    IoInMux I__6452 (
            .O(N__43957),
            .I(N__43954));
    LocalMux I__6451 (
            .O(N__43954),
            .I(N__43951));
    Span4Mux_s2_v I__6450 (
            .O(N__43951),
            .I(N__43948));
    Span4Mux_v I__6449 (
            .O(N__43948),
            .I(N__43945));
    Sp12to4 I__6448 (
            .O(N__43945),
            .I(N__43942));
    Span12Mux_h I__6447 (
            .O(N__43942),
            .I(N__43936));
    InMux I__6446 (
            .O(N__43941),
            .I(N__43933));
    InMux I__6445 (
            .O(N__43940),
            .I(N__43928));
    InMux I__6444 (
            .O(N__43939),
            .I(N__43928));
    Span12Mux_v I__6443 (
            .O(N__43936),
            .I(N__43924));
    LocalMux I__6442 (
            .O(N__43933),
            .I(N__43921));
    LocalMux I__6441 (
            .O(N__43928),
            .I(N__43918));
    InMux I__6440 (
            .O(N__43927),
            .I(N__43915));
    Odrv12 I__6439 (
            .O(N__43924),
            .I(afull_flag_impl_af_flag_p_w_N_603_3));
    Odrv12 I__6438 (
            .O(N__43921),
            .I(afull_flag_impl_af_flag_p_w_N_603_3));
    Odrv4 I__6437 (
            .O(N__43918),
            .I(afull_flag_impl_af_flag_p_w_N_603_3));
    LocalMux I__6436 (
            .O(N__43915),
            .I(afull_flag_impl_af_flag_p_w_N_603_3));
    CascadeMux I__6435 (
            .O(N__43906),
            .I(afull_flag_impl_af_flag_p_w_N_603_3_cascade_));
    InMux I__6434 (
            .O(N__43903),
            .I(N__43900));
    LocalMux I__6433 (
            .O(N__43900),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n6_adj_1172 ));
    IoInMux I__6432 (
            .O(N__43897),
            .I(N__43894));
    LocalMux I__6431 (
            .O(N__43894),
            .I(N__43891));
    IoSpan4Mux I__6430 (
            .O(N__43891),
            .I(N__43888));
    Span4Mux_s3_h I__6429 (
            .O(N__43888),
            .I(N__43885));
    Sp12to4 I__6428 (
            .O(N__43885),
            .I(N__43882));
    Span12Mux_v I__6427 (
            .O(N__43882),
            .I(N__43878));
    InMux I__6426 (
            .O(N__43881),
            .I(N__43875));
    Odrv12 I__6425 (
            .O(N__43878),
            .I(FT_OE_c));
    LocalMux I__6424 (
            .O(N__43875),
            .I(FT_OE_c));
    InMux I__6423 (
            .O(N__43870),
            .I(N__43861));
    InMux I__6422 (
            .O(N__43869),
            .I(N__43861));
    InMux I__6421 (
            .O(N__43868),
            .I(N__43861));
    LocalMux I__6420 (
            .O(N__43861),
            .I(N__43858));
    Span4Mux_v I__6419 (
            .O(N__43858),
            .I(N__43855));
    Span4Mux_h I__6418 (
            .O(N__43855),
            .I(N__43852));
    Span4Mux_v I__6417 (
            .O(N__43852),
            .I(N__43849));
    Span4Mux_v I__6416 (
            .O(N__43849),
            .I(N__43846));
    Odrv4 I__6415 (
            .O(N__43846),
            .I(\usb3_if_inst.n551 ));
    InMux I__6414 (
            .O(N__43843),
            .I(N__43837));
    InMux I__6413 (
            .O(N__43842),
            .I(N__43837));
    LocalMux I__6412 (
            .O(N__43837),
            .I(N__43833));
    InMux I__6411 (
            .O(N__43836),
            .I(N__43830));
    Odrv4 I__6410 (
            .O(N__43833),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_0 ));
    LocalMux I__6409 (
            .O(N__43830),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_0 ));
    InMux I__6408 (
            .O(N__43825),
            .I(N__43819));
    InMux I__6407 (
            .O(N__43824),
            .I(N__43819));
    LocalMux I__6406 (
            .O(N__43819),
            .I(N__43816));
    Odrv4 I__6405 (
            .O(N__43816),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_sig_diff0_w_0 ));
    InMux I__6404 (
            .O(N__43813),
            .I(bfn_10_14_0_));
    InMux I__6403 (
            .O(N__43810),
            .I(N__43798));
    InMux I__6402 (
            .O(N__43809),
            .I(N__43798));
    InMux I__6401 (
            .O(N__43808),
            .I(N__43798));
    InMux I__6400 (
            .O(N__43807),
            .I(N__43798));
    LocalMux I__6399 (
            .O(N__43798),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n25 ));
    InMux I__6398 (
            .O(N__43795),
            .I(N__43792));
    LocalMux I__6397 (
            .O(N__43792),
            .I(N__43788));
    CascadeMux I__6396 (
            .O(N__43791),
            .I(N__43785));
    Span4Mux_v I__6395 (
            .O(N__43788),
            .I(N__43782));
    InMux I__6394 (
            .O(N__43785),
            .I(N__43779));
    Odrv4 I__6393 (
            .O(N__43782),
            .I(REG_mem_47_7));
    LocalMux I__6392 (
            .O(N__43779),
            .I(REG_mem_47_7));
    CascadeMux I__6391 (
            .O(N__43774),
            .I(N__43771));
    InMux I__6390 (
            .O(N__43771),
            .I(N__43768));
    LocalMux I__6389 (
            .O(N__43768),
            .I(N__43765));
    Sp12to4 I__6388 (
            .O(N__43765),
            .I(N__43761));
    InMux I__6387 (
            .O(N__43764),
            .I(N__43758));
    Odrv12 I__6386 (
            .O(N__43761),
            .I(REG_mem_55_11));
    LocalMux I__6385 (
            .O(N__43758),
            .I(REG_mem_55_11));
    CascadeMux I__6384 (
            .O(N__43753),
            .I(N__43750));
    InMux I__6383 (
            .O(N__43750),
            .I(N__43747));
    LocalMux I__6382 (
            .O(N__43747),
            .I(N__43744));
    Span4Mux_v I__6381 (
            .O(N__43744),
            .I(N__43741));
    Span4Mux_h I__6380 (
            .O(N__43741),
            .I(N__43737));
    InMux I__6379 (
            .O(N__43740),
            .I(N__43734));
    Odrv4 I__6378 (
            .O(N__43737),
            .I(REG_mem_47_9));
    LocalMux I__6377 (
            .O(N__43734),
            .I(REG_mem_47_9));
    InMux I__6376 (
            .O(N__43729),
            .I(N__43726));
    LocalMux I__6375 (
            .O(N__43726),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11447 ));
    InMux I__6374 (
            .O(N__43723),
            .I(N__43720));
    LocalMux I__6373 (
            .O(N__43720),
            .I(N__43717));
    Span4Mux_h I__6372 (
            .O(N__43717),
            .I(N__43710));
    InMux I__6371 (
            .O(N__43716),
            .I(N__43707));
    InMux I__6370 (
            .O(N__43715),
            .I(N__43700));
    InMux I__6369 (
            .O(N__43714),
            .I(N__43700));
    InMux I__6368 (
            .O(N__43713),
            .I(N__43700));
    Odrv4 I__6367 (
            .O(N__43710),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12_adj_1156 ));
    LocalMux I__6366 (
            .O(N__43707),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12_adj_1156 ));
    LocalMux I__6365 (
            .O(N__43700),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12_adj_1156 ));
    CascadeMux I__6364 (
            .O(N__43693),
            .I(N__43690));
    InMux I__6363 (
            .O(N__43690),
            .I(N__43686));
    CascadeMux I__6362 (
            .O(N__43689),
            .I(N__43682));
    LocalMux I__6361 (
            .O(N__43686),
            .I(N__43679));
    InMux I__6360 (
            .O(N__43685),
            .I(N__43674));
    InMux I__6359 (
            .O(N__43682),
            .I(N__43674));
    Span4Mux_v I__6358 (
            .O(N__43679),
            .I(N__43667));
    LocalMux I__6357 (
            .O(N__43674),
            .I(N__43667));
    InMux I__6356 (
            .O(N__43673),
            .I(N__43662));
    InMux I__6355 (
            .O(N__43672),
            .I(N__43662));
    Odrv4 I__6354 (
            .O(N__43667),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.full_o ));
    LocalMux I__6353 (
            .O(N__43662),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.full_o ));
    CascadeMux I__6352 (
            .O(N__43657),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n9_cascade_ ));
    InMux I__6351 (
            .O(N__43654),
            .I(N__43651));
    LocalMux I__6350 (
            .O(N__43651),
            .I(N__43645));
    InMux I__6349 (
            .O(N__43650),
            .I(N__43642));
    InMux I__6348 (
            .O(N__43649),
            .I(N__43637));
    InMux I__6347 (
            .O(N__43648),
            .I(N__43637));
    Odrv4 I__6346 (
            .O(N__43645),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n9 ));
    LocalMux I__6345 (
            .O(N__43642),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n9 ));
    LocalMux I__6344 (
            .O(N__43637),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n9 ));
    CascadeMux I__6343 (
            .O(N__43630),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12_adj_1156_cascade_ ));
    InMux I__6342 (
            .O(N__43627),
            .I(N__43622));
    InMux I__6341 (
            .O(N__43626),
            .I(N__43617));
    InMux I__6340 (
            .O(N__43625),
            .I(N__43617));
    LocalMux I__6339 (
            .O(N__43622),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n20_adj_1160 ));
    LocalMux I__6338 (
            .O(N__43617),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n20_adj_1160 ));
    InMux I__6337 (
            .O(N__43612),
            .I(N__43604));
    InMux I__6336 (
            .O(N__43611),
            .I(N__43604));
    InMux I__6335 (
            .O(N__43610),
            .I(N__43599));
    InMux I__6334 (
            .O(N__43609),
            .I(N__43599));
    LocalMux I__6333 (
            .O(N__43604),
            .I(N__43596));
    LocalMux I__6332 (
            .O(N__43599),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n36 ));
    Odrv4 I__6331 (
            .O(N__43596),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n36 ));
    CascadeMux I__6330 (
            .O(N__43591),
            .I(N__43588));
    InMux I__6329 (
            .O(N__43588),
            .I(N__43582));
    InMux I__6328 (
            .O(N__43587),
            .I(N__43575));
    InMux I__6327 (
            .O(N__43586),
            .I(N__43575));
    InMux I__6326 (
            .O(N__43585),
            .I(N__43575));
    LocalMux I__6325 (
            .O(N__43582),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11 ));
    LocalMux I__6324 (
            .O(N__43575),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11 ));
    CascadeMux I__6323 (
            .O(N__43570),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11_cascade_ ));
    CascadeMux I__6322 (
            .O(N__43567),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n16_cascade_ ));
    InMux I__6321 (
            .O(N__43564),
            .I(N__43555));
    InMux I__6320 (
            .O(N__43563),
            .I(N__43555));
    InMux I__6319 (
            .O(N__43562),
            .I(N__43555));
    LocalMux I__6318 (
            .O(N__43555),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n16 ));
    CascadeMux I__6317 (
            .O(N__43552),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n20_adj_1160_cascade_ ));
    InMux I__6316 (
            .O(N__43549),
            .I(N__43546));
    LocalMux I__6315 (
            .O(N__43546),
            .I(N__43543));
    Span4Mux_v I__6314 (
            .O(N__43543),
            .I(N__43539));
    InMux I__6313 (
            .O(N__43542),
            .I(N__43536));
    Odrv4 I__6312 (
            .O(N__43539),
            .I(REG_mem_11_15));
    LocalMux I__6311 (
            .O(N__43536),
            .I(REG_mem_11_15));
    CascadeMux I__6310 (
            .O(N__43531),
            .I(n26_cascade_));
    InMux I__6309 (
            .O(N__43528),
            .I(N__43525));
    LocalMux I__6308 (
            .O(N__43525),
            .I(N__43522));
    Span4Mux_v I__6307 (
            .O(N__43522),
            .I(N__43519));
    Span4Mux_v I__6306 (
            .O(N__43519),
            .I(N__43515));
    InMux I__6305 (
            .O(N__43518),
            .I(N__43512));
    Span4Mux_h I__6304 (
            .O(N__43515),
            .I(N__43509));
    LocalMux I__6303 (
            .O(N__43512),
            .I(N__43506));
    Odrv4 I__6302 (
            .O(N__43509),
            .I(REG_mem_39_3));
    Odrv4 I__6301 (
            .O(N__43506),
            .I(REG_mem_39_3));
    InMux I__6300 (
            .O(N__43501),
            .I(N__43498));
    LocalMux I__6299 (
            .O(N__43498),
            .I(N__43495));
    Span4Mux_v I__6298 (
            .O(N__43495),
            .I(N__43491));
    InMux I__6297 (
            .O(N__43494),
            .I(N__43488));
    Odrv4 I__6296 (
            .O(N__43491),
            .I(REG_mem_17_9));
    LocalMux I__6295 (
            .O(N__43488),
            .I(REG_mem_17_9));
    InMux I__6294 (
            .O(N__43483),
            .I(N__43480));
    LocalMux I__6293 (
            .O(N__43480),
            .I(N__43477));
    Span4Mux_h I__6292 (
            .O(N__43477),
            .I(N__43473));
    InMux I__6291 (
            .O(N__43476),
            .I(N__43470));
    Odrv4 I__6290 (
            .O(N__43473),
            .I(REG_mem_9_9));
    LocalMux I__6289 (
            .O(N__43470),
            .I(REG_mem_9_9));
    InMux I__6288 (
            .O(N__43465),
            .I(N__43462));
    LocalMux I__6287 (
            .O(N__43462),
            .I(N__43459));
    Span4Mux_v I__6286 (
            .O(N__43459),
            .I(N__43456));
    Sp12to4 I__6285 (
            .O(N__43456),
            .I(N__43453));
    Span12Mux_s9_h I__6284 (
            .O(N__43453),
            .I(N__43449));
    InMux I__6283 (
            .O(N__43452),
            .I(N__43446));
    Odrv12 I__6282 (
            .O(N__43449),
            .I(REG_mem_43_9));
    LocalMux I__6281 (
            .O(N__43446),
            .I(REG_mem_43_9));
    InMux I__6280 (
            .O(N__43441),
            .I(N__43438));
    LocalMux I__6279 (
            .O(N__43438),
            .I(N__43435));
    Span4Mux_h I__6278 (
            .O(N__43435),
            .I(N__43431));
    InMux I__6277 (
            .O(N__43434),
            .I(N__43428));
    Odrv4 I__6276 (
            .O(N__43431),
            .I(REG_mem_51_15));
    LocalMux I__6275 (
            .O(N__43428),
            .I(REG_mem_51_15));
    InMux I__6274 (
            .O(N__43423),
            .I(N__43420));
    LocalMux I__6273 (
            .O(N__43420),
            .I(N__43417));
    Span4Mux_v I__6272 (
            .O(N__43417),
            .I(N__43414));
    Span4Mux_v I__6271 (
            .O(N__43414),
            .I(N__43411));
    Span4Mux_h I__6270 (
            .O(N__43411),
            .I(N__43408));
    Span4Mux_h I__6269 (
            .O(N__43408),
            .I(N__43404));
    InMux I__6268 (
            .O(N__43407),
            .I(N__43401));
    Odrv4 I__6267 (
            .O(N__43404),
            .I(REG_mem_7_10));
    LocalMux I__6266 (
            .O(N__43401),
            .I(REG_mem_7_10));
    InMux I__6265 (
            .O(N__43396),
            .I(N__43390));
    InMux I__6264 (
            .O(N__43395),
            .I(N__43390));
    LocalMux I__6263 (
            .O(N__43390),
            .I(REG_mem_36_15));
    InMux I__6262 (
            .O(N__43387),
            .I(N__43384));
    LocalMux I__6261 (
            .O(N__43384),
            .I(N__43381));
    Sp12to4 I__6260 (
            .O(N__43381),
            .I(N__43378));
    Odrv12 I__6259 (
            .O(N__43378),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11995 ));
    InMux I__6258 (
            .O(N__43375),
            .I(N__43372));
    LocalMux I__6257 (
            .O(N__43372),
            .I(N__43369));
    Span4Mux_v I__6256 (
            .O(N__43369),
            .I(N__43365));
    InMux I__6255 (
            .O(N__43368),
            .I(N__43362));
    Odrv4 I__6254 (
            .O(N__43365),
            .I(REG_mem_9_15));
    LocalMux I__6253 (
            .O(N__43362),
            .I(REG_mem_9_15));
    InMux I__6252 (
            .O(N__43357),
            .I(N__43354));
    LocalMux I__6251 (
            .O(N__43354),
            .I(N__43350));
    InMux I__6250 (
            .O(N__43353),
            .I(N__43347));
    Odrv4 I__6249 (
            .O(N__43350),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_7 ));
    LocalMux I__6248 (
            .O(N__43347),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_7 ));
    InMux I__6247 (
            .O(N__43342),
            .I(N__43339));
    LocalMux I__6246 (
            .O(N__43339),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12383 ));
    InMux I__6245 (
            .O(N__43336),
            .I(N__43332));
    CascadeMux I__6244 (
            .O(N__43335),
            .I(N__43329));
    LocalMux I__6243 (
            .O(N__43332),
            .I(N__43326));
    InMux I__6242 (
            .O(N__43329),
            .I(N__43323));
    Odrv4 I__6241 (
            .O(N__43326),
            .I(REG_mem_31_0));
    LocalMux I__6240 (
            .O(N__43323),
            .I(REG_mem_31_0));
    CascadeMux I__6239 (
            .O(N__43318),
            .I(N__43315));
    InMux I__6238 (
            .O(N__43315),
            .I(N__43312));
    LocalMux I__6237 (
            .O(N__43312),
            .I(N__43309));
    Sp12to4 I__6236 (
            .O(N__43309),
            .I(N__43306));
    Span12Mux_s9_v I__6235 (
            .O(N__43306),
            .I(N__43302));
    InMux I__6234 (
            .O(N__43305),
            .I(N__43299));
    Odrv12 I__6233 (
            .O(N__43302),
            .I(REG_mem_18_15));
    LocalMux I__6232 (
            .O(N__43299),
            .I(REG_mem_18_15));
    InMux I__6231 (
            .O(N__43294),
            .I(N__43291));
    LocalMux I__6230 (
            .O(N__43291),
            .I(N__43288));
    Span4Mux_v I__6229 (
            .O(N__43288),
            .I(N__43284));
    InMux I__6228 (
            .O(N__43287),
            .I(N__43281));
    Odrv4 I__6227 (
            .O(N__43284),
            .I(REG_mem_16_9));
    LocalMux I__6226 (
            .O(N__43281),
            .I(REG_mem_16_9));
    InMux I__6225 (
            .O(N__43276),
            .I(N__43273));
    LocalMux I__6224 (
            .O(N__43273),
            .I(N__43270));
    Span4Mux_h I__6223 (
            .O(N__43270),
            .I(N__43266));
    InMux I__6222 (
            .O(N__43269),
            .I(N__43263));
    Odrv4 I__6221 (
            .O(N__43266),
            .I(REG_mem_26_0));
    LocalMux I__6220 (
            .O(N__43263),
            .I(REG_mem_26_0));
    InMux I__6219 (
            .O(N__43258),
            .I(N__43255));
    LocalMux I__6218 (
            .O(N__43255),
            .I(N__43251));
    InMux I__6217 (
            .O(N__43254),
            .I(N__43248));
    Odrv4 I__6216 (
            .O(N__43251),
            .I(REG_mem_49_9));
    LocalMux I__6215 (
            .O(N__43248),
            .I(REG_mem_49_9));
    InMux I__6214 (
            .O(N__43243),
            .I(N__43240));
    LocalMux I__6213 (
            .O(N__43240),
            .I(N__43237));
    Span12Mux_v I__6212 (
            .O(N__43237),
            .I(N__43233));
    InMux I__6211 (
            .O(N__43236),
            .I(N__43230));
    Odrv12 I__6210 (
            .O(N__43233),
            .I(REG_mem_19_9));
    LocalMux I__6209 (
            .O(N__43230),
            .I(REG_mem_19_9));
    InMux I__6208 (
            .O(N__43225),
            .I(N__43222));
    LocalMux I__6207 (
            .O(N__43222),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12908 ));
    InMux I__6206 (
            .O(N__43219),
            .I(N__43216));
    LocalMux I__6205 (
            .O(N__43216),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12361 ));
    CascadeMux I__6204 (
            .O(N__43213),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12362_cascade_ ));
    CascadeMux I__6203 (
            .O(N__43210),
            .I(N__43207));
    InMux I__6202 (
            .O(N__43207),
            .I(N__43204));
    LocalMux I__6201 (
            .O(N__43204),
            .I(N__43201));
    Span4Mux_h I__6200 (
            .O(N__43201),
            .I(N__43198));
    Sp12to4 I__6199 (
            .O(N__43198),
            .I(N__43195));
    Odrv12 I__6198 (
            .O(N__43195),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12911 ));
    InMux I__6197 (
            .O(N__43192),
            .I(N__43189));
    LocalMux I__6196 (
            .O(N__43189),
            .I(N__43186));
    Span4Mux_h I__6195 (
            .O(N__43186),
            .I(N__43182));
    InMux I__6194 (
            .O(N__43185),
            .I(N__43179));
    Odrv4 I__6193 (
            .O(N__43182),
            .I(REG_mem_19_0));
    LocalMux I__6192 (
            .O(N__43179),
            .I(REG_mem_19_0));
    InMux I__6191 (
            .O(N__43174),
            .I(N__43171));
    LocalMux I__6190 (
            .O(N__43171),
            .I(N__43167));
    InMux I__6189 (
            .O(N__43170),
            .I(N__43164));
    Odrv4 I__6188 (
            .O(N__43167),
            .I(REG_mem_11_9));
    LocalMux I__6187 (
            .O(N__43164),
            .I(REG_mem_11_9));
    InMux I__6186 (
            .O(N__43159),
            .I(N__43156));
    LocalMux I__6185 (
            .O(N__43156),
            .I(N__43153));
    Odrv12 I__6184 (
            .O(N__43153),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13232 ));
    CascadeMux I__6183 (
            .O(N__43150),
            .I(N__43147));
    InMux I__6182 (
            .O(N__43147),
            .I(N__43143));
    InMux I__6181 (
            .O(N__43146),
            .I(N__43140));
    LocalMux I__6180 (
            .O(N__43143),
            .I(N__43137));
    LocalMux I__6179 (
            .O(N__43140),
            .I(N__43134));
    Odrv4 I__6178 (
            .O(N__43137),
            .I(REG_mem_18_0));
    Odrv4 I__6177 (
            .O(N__43134),
            .I(REG_mem_18_0));
    CascadeMux I__6176 (
            .O(N__43129),
            .I(N__43126));
    InMux I__6175 (
            .O(N__43126),
            .I(N__43120));
    InMux I__6174 (
            .O(N__43125),
            .I(N__43120));
    LocalMux I__6173 (
            .O(N__43120),
            .I(REG_mem_10_9));
    InMux I__6172 (
            .O(N__43117),
            .I(N__43114));
    LocalMux I__6171 (
            .O(N__43114),
            .I(N__43111));
    Odrv4 I__6170 (
            .O(N__43111),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11971 ));
    CascadeMux I__6169 (
            .O(N__43108),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13682_cascade_ ));
    CascadeMux I__6168 (
            .O(N__43105),
            .I(N__43102));
    InMux I__6167 (
            .O(N__43102),
            .I(N__43099));
    LocalMux I__6166 (
            .O(N__43099),
            .I(N__43096));
    Span4Mux_h I__6165 (
            .O(N__43096),
            .I(N__43093));
    Span4Mux_h I__6164 (
            .O(N__43093),
            .I(N__43090));
    Odrv4 I__6163 (
            .O(N__43090),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14132 ));
    InMux I__6162 (
            .O(N__43087),
            .I(N__43084));
    LocalMux I__6161 (
            .O(N__43084),
            .I(N__43081));
    Span4Mux_v I__6160 (
            .O(N__43081),
            .I(N__43078));
    Odrv4 I__6159 (
            .O(N__43078),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12007 ));
    InMux I__6158 (
            .O(N__43075),
            .I(N__43072));
    LocalMux I__6157 (
            .O(N__43072),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11972 ));
    InMux I__6156 (
            .O(N__43069),
            .I(N__43063));
    InMux I__6155 (
            .O(N__43068),
            .I(N__43063));
    LocalMux I__6154 (
            .O(N__43063),
            .I(REG_mem_51_0));
    InMux I__6153 (
            .O(N__43060),
            .I(N__43054));
    InMux I__6152 (
            .O(N__43059),
            .I(N__43054));
    LocalMux I__6151 (
            .O(N__43054),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_5 ));
    CascadeMux I__6150 (
            .O(N__43051),
            .I(N__43047));
    InMux I__6149 (
            .O(N__43050),
            .I(N__43042));
    InMux I__6148 (
            .O(N__43047),
            .I(N__43042));
    LocalMux I__6147 (
            .O(N__43042),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_5 ));
    InMux I__6146 (
            .O(N__43039),
            .I(N__43035));
    CascadeMux I__6145 (
            .O(N__43038),
            .I(N__43032));
    LocalMux I__6144 (
            .O(N__43035),
            .I(N__43029));
    InMux I__6143 (
            .O(N__43032),
            .I(N__43026));
    Odrv4 I__6142 (
            .O(N__43029),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_0 ));
    LocalMux I__6141 (
            .O(N__43026),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_0 ));
    InMux I__6140 (
            .O(N__43021),
            .I(N__43018));
    LocalMux I__6139 (
            .O(N__43018),
            .I(N__43015));
    Span4Mux_v I__6138 (
            .O(N__43015),
            .I(N__43012));
    Span4Mux_v I__6137 (
            .O(N__43012),
            .I(N__43008));
    InMux I__6136 (
            .O(N__43011),
            .I(N__43005));
    Odrv4 I__6135 (
            .O(N__43008),
            .I(REG_mem_19_3));
    LocalMux I__6134 (
            .O(N__43005),
            .I(REG_mem_19_3));
    CascadeMux I__6133 (
            .O(N__43000),
            .I(N__42997));
    InMux I__6132 (
            .O(N__42997),
            .I(N__42991));
    InMux I__6131 (
            .O(N__42996),
            .I(N__42991));
    LocalMux I__6130 (
            .O(N__42991),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_9 ));
    InMux I__6129 (
            .O(N__42988),
            .I(N__42985));
    LocalMux I__6128 (
            .O(N__42985),
            .I(N__42981));
    InMux I__6127 (
            .O(N__42984),
            .I(N__42978));
    Odrv4 I__6126 (
            .O(N__42981),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_9 ));
    LocalMux I__6125 (
            .O(N__42978),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_9 ));
    InMux I__6124 (
            .O(N__42973),
            .I(N__42970));
    LocalMux I__6123 (
            .O(N__42970),
            .I(N__42967));
    Span4Mux_h I__6122 (
            .O(N__42967),
            .I(N__42964));
    Odrv4 I__6121 (
            .O(N__42964),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12341 ));
    InMux I__6120 (
            .O(N__42961),
            .I(N__42955));
    InMux I__6119 (
            .O(N__42960),
            .I(N__42955));
    LocalMux I__6118 (
            .O(N__42955),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_15 ));
    InMux I__6117 (
            .O(N__42952),
            .I(N__42946));
    InMux I__6116 (
            .O(N__42951),
            .I(N__42946));
    LocalMux I__6115 (
            .O(N__42946),
            .I(N__42943));
    Odrv4 I__6114 (
            .O(N__42943),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_15 ));
    InMux I__6113 (
            .O(N__42940),
            .I(N__42937));
    LocalMux I__6112 (
            .O(N__42937),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11987 ));
    CascadeMux I__6111 (
            .O(N__42934),
            .I(N__42931));
    InMux I__6110 (
            .O(N__42931),
            .I(N__42928));
    LocalMux I__6109 (
            .O(N__42928),
            .I(N__42925));
    Span4Mux_h I__6108 (
            .O(N__42925),
            .I(N__42922));
    Odrv4 I__6107 (
            .O(N__42922),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11984 ));
    InMux I__6106 (
            .O(N__42919),
            .I(N__42916));
    LocalMux I__6105 (
            .O(N__42916),
            .I(N__42913));
    Span4Mux_h I__6104 (
            .O(N__42913),
            .I(N__42910));
    Odrv4 I__6103 (
            .O(N__42910),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11983 ));
    InMux I__6102 (
            .O(N__42907),
            .I(N__42904));
    LocalMux I__6101 (
            .O(N__42904),
            .I(N__42900));
    InMux I__6100 (
            .O(N__42903),
            .I(N__42897));
    Odrv4 I__6099 (
            .O(N__42900),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_11 ));
    LocalMux I__6098 (
            .O(N__42897),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_11 ));
    InMux I__6097 (
            .O(N__42892),
            .I(N__42889));
    LocalMux I__6096 (
            .O(N__42889),
            .I(N__42885));
    CascadeMux I__6095 (
            .O(N__42888),
            .I(N__42882));
    Span4Mux_v I__6094 (
            .O(N__42885),
            .I(N__42879));
    InMux I__6093 (
            .O(N__42882),
            .I(N__42876));
    Odrv4 I__6092 (
            .O(N__42879),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_13 ));
    LocalMux I__6091 (
            .O(N__42876),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_13 ));
    CascadeMux I__6090 (
            .O(N__42871),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13904_cascade_ ));
    InMux I__6089 (
            .O(N__42868),
            .I(N__42865));
    LocalMux I__6088 (
            .O(N__42865),
            .I(N__42862));
    Span4Mux_v I__6087 (
            .O(N__42862),
            .I(N__42859));
    Odrv4 I__6086 (
            .O(N__42859),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12174 ));
    CascadeMux I__6085 (
            .O(N__42856),
            .I(N__42852));
    InMux I__6084 (
            .O(N__42855),
            .I(N__42847));
    InMux I__6083 (
            .O(N__42852),
            .I(N__42847));
    LocalMux I__6082 (
            .O(N__42847),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_13 ));
    CascadeMux I__6081 (
            .O(N__42844),
            .I(N__42840));
    InMux I__6080 (
            .O(N__42843),
            .I(N__42835));
    InMux I__6079 (
            .O(N__42840),
            .I(N__42835));
    LocalMux I__6078 (
            .O(N__42835),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_13 ));
    InMux I__6077 (
            .O(N__42832),
            .I(N__42829));
    LocalMux I__6076 (
            .O(N__42829),
            .I(N__42826));
    Odrv4 I__6075 (
            .O(N__42826),
            .I(rd_grey_sync_r_0));
    InMux I__6074 (
            .O(N__42823),
            .I(N__42820));
    LocalMux I__6073 (
            .O(N__42820),
            .I(N__42817));
    Span4Mux_v I__6072 (
            .O(N__42817),
            .I(N__42814));
    Odrv4 I__6071 (
            .O(N__42814),
            .I(rp_sync1_r_0));
    CascadeMux I__6070 (
            .O(N__42811),
            .I(N__42808));
    InMux I__6069 (
            .O(N__42808),
            .I(N__42802));
    InMux I__6068 (
            .O(N__42807),
            .I(N__42802));
    LocalMux I__6067 (
            .O(N__42802),
            .I(N__42799));
    Odrv4 I__6066 (
            .O(N__42799),
            .I(rd_addr_nxt_c_6_N_465_5));
    CascadeMux I__6065 (
            .O(N__42796),
            .I(rd_addr_nxt_c_6_N_465_1_cascade_));
    CascadeMux I__6064 (
            .O(N__42793),
            .I(N__42789));
    CascadeMux I__6063 (
            .O(N__42792),
            .I(N__42786));
    InMux I__6062 (
            .O(N__42789),
            .I(N__42783));
    InMux I__6061 (
            .O(N__42786),
            .I(N__42780));
    LocalMux I__6060 (
            .O(N__42783),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_13 ));
    LocalMux I__6059 (
            .O(N__42780),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_13 ));
    CascadeMux I__6058 (
            .O(N__42775),
            .I(N__42772));
    InMux I__6057 (
            .O(N__42772),
            .I(N__42769));
    LocalMux I__6056 (
            .O(N__42769),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14240 ));
    CascadeMux I__6055 (
            .O(N__42766),
            .I(N__42762));
    InMux I__6054 (
            .O(N__42765),
            .I(N__42757));
    InMux I__6053 (
            .O(N__42762),
            .I(N__42757));
    LocalMux I__6052 (
            .O(N__42757),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_11 ));
    CascadeMux I__6051 (
            .O(N__42754),
            .I(N__42750));
    CascadeMux I__6050 (
            .O(N__42753),
            .I(N__42747));
    InMux I__6049 (
            .O(N__42750),
            .I(N__42742));
    InMux I__6048 (
            .O(N__42747),
            .I(N__42742));
    LocalMux I__6047 (
            .O(N__42742),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_11 ));
    InMux I__6046 (
            .O(N__42739),
            .I(N__42735));
    InMux I__6045 (
            .O(N__42738),
            .I(N__42732));
    LocalMux I__6044 (
            .O(N__42735),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_11 ));
    LocalMux I__6043 (
            .O(N__42732),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_11 ));
    InMux I__6042 (
            .O(N__42727),
            .I(N__42724));
    LocalMux I__6041 (
            .O(N__42724),
            .I(N__42721));
    Odrv4 I__6040 (
            .O(N__42721),
            .I(rd_grey_sync_r_1));
    CascadeMux I__6039 (
            .O(N__42718),
            .I(N__42714));
    InMux I__6038 (
            .O(N__42717),
            .I(N__42710));
    InMux I__6037 (
            .O(N__42714),
            .I(N__42705));
    InMux I__6036 (
            .O(N__42713),
            .I(N__42705));
    LocalMux I__6035 (
            .O(N__42710),
            .I(N__42702));
    LocalMux I__6034 (
            .O(N__42705),
            .I(N__42699));
    Odrv4 I__6033 (
            .O(N__42702),
            .I(rd_addr_nxt_c_6_N_465_3));
    Odrv4 I__6032 (
            .O(N__42699),
            .I(rd_addr_nxt_c_6_N_465_3));
    InMux I__6031 (
            .O(N__42694),
            .I(N__42691));
    LocalMux I__6030 (
            .O(N__42691),
            .I(N__42687));
    CascadeMux I__6029 (
            .O(N__42690),
            .I(N__42684));
    Span4Mux_v I__6028 (
            .O(N__42687),
            .I(N__42681));
    InMux I__6027 (
            .O(N__42684),
            .I(N__42678));
    Odrv4 I__6026 (
            .O(N__42681),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_13 ));
    LocalMux I__6025 (
            .O(N__42678),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_13 ));
    InMux I__6024 (
            .O(N__42673),
            .I(N__42670));
    LocalMux I__6023 (
            .O(N__42670),
            .I(N__42667));
    Span4Mux_v I__6022 (
            .O(N__42667),
            .I(N__42664));
    Odrv4 I__6021 (
            .O(N__42664),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12042 ));
    CascadeMux I__6020 (
            .O(N__42661),
            .I(N__42657));
    InMux I__6019 (
            .O(N__42660),
            .I(N__42652));
    InMux I__6018 (
            .O(N__42657),
            .I(N__42652));
    LocalMux I__6017 (
            .O(N__42652),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_13 ));
    InMux I__6016 (
            .O(N__42649),
            .I(N__42643));
    InMux I__6015 (
            .O(N__42648),
            .I(N__42643));
    LocalMux I__6014 (
            .O(N__42643),
            .I(REG_mem_31_11));
    CascadeMux I__6013 (
            .O(N__42640),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13940_cascade_ ));
    CascadeMux I__6012 (
            .O(N__42637),
            .I(N__42633));
    InMux I__6011 (
            .O(N__42636),
            .I(N__42630));
    InMux I__6010 (
            .O(N__42633),
            .I(N__42627));
    LocalMux I__6009 (
            .O(N__42630),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_11 ));
    LocalMux I__6008 (
            .O(N__42627),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_11 ));
    InMux I__6007 (
            .O(N__42622),
            .I(N__42619));
    LocalMux I__6006 (
            .O(N__42619),
            .I(N__42616));
    Odrv4 I__6005 (
            .O(N__42616),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13943 ));
    CascadeMux I__6004 (
            .O(N__42613),
            .I(N__42610));
    InMux I__6003 (
            .O(N__42610),
            .I(N__42607));
    LocalMux I__6002 (
            .O(N__42607),
            .I(N__42604));
    Span4Mux_v I__6001 (
            .O(N__42604),
            .I(N__42600));
    InMux I__6000 (
            .O(N__42603),
            .I(N__42597));
    Odrv4 I__5999 (
            .O(N__42600),
            .I(REG_mem_23_11));
    LocalMux I__5998 (
            .O(N__42597),
            .I(REG_mem_23_11));
    InMux I__5997 (
            .O(N__42592),
            .I(N__42589));
    LocalMux I__5996 (
            .O(N__42589),
            .I(rp_sync1_r_1));
    InMux I__5995 (
            .O(N__42586),
            .I(N__42583));
    LocalMux I__5994 (
            .O(N__42583),
            .I(N__42579));
    CascadeMux I__5993 (
            .O(N__42582),
            .I(N__42576));
    Span4Mux_v I__5992 (
            .O(N__42579),
            .I(N__42573));
    InMux I__5991 (
            .O(N__42576),
            .I(N__42570));
    Odrv4 I__5990 (
            .O(N__42573),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_11 ));
    LocalMux I__5989 (
            .O(N__42570),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_11 ));
    InMux I__5988 (
            .O(N__42565),
            .I(N__42562));
    LocalMux I__5987 (
            .O(N__42562),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_0 ));
    InMux I__5986 (
            .O(N__42559),
            .I(N__42553));
    InMux I__5985 (
            .O(N__42558),
            .I(N__42553));
    LocalMux I__5984 (
            .O(N__42553),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_1 ));
    CascadeMux I__5983 (
            .O(N__42550),
            .I(N__42547));
    InMux I__5982 (
            .O(N__42547),
            .I(N__42543));
    InMux I__5981 (
            .O(N__42546),
            .I(N__42540));
    LocalMux I__5980 (
            .O(N__42543),
            .I(REG_mem_9_11));
    LocalMux I__5979 (
            .O(N__42540),
            .I(REG_mem_9_11));
    InMux I__5978 (
            .O(N__42535),
            .I(N__42532));
    LocalMux I__5977 (
            .O(N__42532),
            .I(N__42528));
    InMux I__5976 (
            .O(N__42531),
            .I(N__42525));
    Odrv4 I__5975 (
            .O(N__42528),
            .I(REG_mem_8_11));
    LocalMux I__5974 (
            .O(N__42525),
            .I(REG_mem_8_11));
    CascadeMux I__5973 (
            .O(N__42520),
            .I(N__42517));
    InMux I__5972 (
            .O(N__42517),
            .I(N__42514));
    LocalMux I__5971 (
            .O(N__42514),
            .I(N__42511));
    Span12Mux_v I__5970 (
            .O(N__42511),
            .I(N__42507));
    InMux I__5969 (
            .O(N__42510),
            .I(N__42504));
    Odrv12 I__5968 (
            .O(N__42507),
            .I(REG_mem_11_11));
    LocalMux I__5967 (
            .O(N__42504),
            .I(REG_mem_11_11));
    InMux I__5966 (
            .O(N__42499),
            .I(N__42496));
    LocalMux I__5965 (
            .O(N__42496),
            .I(N__42493));
    Odrv4 I__5964 (
            .O(N__42493),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14402 ));
    InMux I__5963 (
            .O(N__42490),
            .I(N__42484));
    InMux I__5962 (
            .O(N__42489),
            .I(N__42484));
    LocalMux I__5961 (
            .O(N__42484),
            .I(REG_mem_10_11));
    InMux I__5960 (
            .O(N__42481),
            .I(N__42478));
    LocalMux I__5959 (
            .O(N__42478),
            .I(N__42474));
    InMux I__5958 (
            .O(N__42477),
            .I(N__42471));
    Odrv4 I__5957 (
            .O(N__42474),
            .I(REG_mem_47_3));
    LocalMux I__5956 (
            .O(N__42471),
            .I(REG_mem_47_3));
    CascadeMux I__5955 (
            .O(N__42466),
            .I(N__42462));
    InMux I__5954 (
            .O(N__42465),
            .I(N__42459));
    InMux I__5953 (
            .O(N__42462),
            .I(N__42456));
    LocalMux I__5952 (
            .O(N__42459),
            .I(N__42453));
    LocalMux I__5951 (
            .O(N__42456),
            .I(REG_mem_19_12));
    Odrv4 I__5950 (
            .O(N__42453),
            .I(REG_mem_19_12));
    InMux I__5949 (
            .O(N__42448),
            .I(N__42445));
    LocalMux I__5948 (
            .O(N__42445),
            .I(N__42442));
    Span4Mux_v I__5947 (
            .O(N__42442),
            .I(N__42439));
    Span4Mux_h I__5946 (
            .O(N__42439),
            .I(N__42435));
    InMux I__5945 (
            .O(N__42438),
            .I(N__42432));
    Odrv4 I__5944 (
            .O(N__42435),
            .I(REG_mem_41_12));
    LocalMux I__5943 (
            .O(N__42432),
            .I(REG_mem_41_12));
    InMux I__5942 (
            .O(N__42427),
            .I(N__42424));
    LocalMux I__5941 (
            .O(N__42424),
            .I(N__42421));
    Span4Mux_v I__5940 (
            .O(N__42421),
            .I(N__42417));
    InMux I__5939 (
            .O(N__42420),
            .I(N__42414));
    Odrv4 I__5938 (
            .O(N__42417),
            .I(REG_mem_11_13));
    LocalMux I__5937 (
            .O(N__42414),
            .I(REG_mem_11_13));
    InMux I__5936 (
            .O(N__42409),
            .I(N__42406));
    LocalMux I__5935 (
            .O(N__42406),
            .I(N__42402));
    InMux I__5934 (
            .O(N__42405),
            .I(N__42399));
    Odrv4 I__5933 (
            .O(N__42402),
            .I(REG_mem_9_13));
    LocalMux I__5932 (
            .O(N__42399),
            .I(REG_mem_9_13));
    InMux I__5931 (
            .O(N__42394),
            .I(N__42391));
    LocalMux I__5930 (
            .O(N__42391),
            .I(N__42388));
    Span4Mux_h I__5929 (
            .O(N__42388),
            .I(N__42384));
    InMux I__5928 (
            .O(N__42387),
            .I(N__42381));
    Odrv4 I__5927 (
            .O(N__42384),
            .I(REG_mem_51_12));
    LocalMux I__5926 (
            .O(N__42381),
            .I(REG_mem_51_12));
    InMux I__5925 (
            .O(N__42376),
            .I(N__42373));
    LocalMux I__5924 (
            .O(N__42373),
            .I(N__42370));
    Odrv4 I__5923 (
            .O(N__42370),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11400 ));
    CascadeMux I__5922 (
            .O(N__42367),
            .I(n7596_cascade_));
    InMux I__5921 (
            .O(N__42364),
            .I(N__42361));
    LocalMux I__5920 (
            .O(N__42361),
            .I(N__42358));
    Span4Mux_v I__5919 (
            .O(N__42358),
            .I(N__42355));
    Span4Mux_h I__5918 (
            .O(N__42355),
            .I(N__42352));
    Odrv4 I__5917 (
            .O(N__42352),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11831 ));
    CascadeMux I__5916 (
            .O(N__42349),
            .I(N__42346));
    InMux I__5915 (
            .O(N__42346),
            .I(N__42342));
    CascadeMux I__5914 (
            .O(N__42345),
            .I(N__42339));
    LocalMux I__5913 (
            .O(N__42342),
            .I(N__42336));
    InMux I__5912 (
            .O(N__42339),
            .I(N__42333));
    Span4Mux_v I__5911 (
            .O(N__42336),
            .I(N__42328));
    LocalMux I__5910 (
            .O(N__42333),
            .I(N__42328));
    Odrv4 I__5909 (
            .O(N__42328),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_13 ));
    CascadeMux I__5908 (
            .O(N__42325),
            .I(N__42322));
    InMux I__5907 (
            .O(N__42322),
            .I(N__42319));
    LocalMux I__5906 (
            .O(N__42319),
            .I(N__42316));
    Span4Mux_v I__5905 (
            .O(N__42316),
            .I(N__42312));
    InMux I__5904 (
            .O(N__42315),
            .I(N__42309));
    Odrv4 I__5903 (
            .O(N__42312),
            .I(REG_mem_42_13));
    LocalMux I__5902 (
            .O(N__42309),
            .I(REG_mem_42_13));
    InMux I__5901 (
            .O(N__42304),
            .I(N__42301));
    LocalMux I__5900 (
            .O(N__42301),
            .I(N__42298));
    Span4Mux_v I__5899 (
            .O(N__42298),
            .I(N__42294));
    InMux I__5898 (
            .O(N__42297),
            .I(N__42291));
    Odrv4 I__5897 (
            .O(N__42294),
            .I(REG_mem_40_12));
    LocalMux I__5896 (
            .O(N__42291),
            .I(REG_mem_40_12));
    InMux I__5895 (
            .O(N__42286),
            .I(N__42283));
    LocalMux I__5894 (
            .O(N__42283),
            .I(N__42280));
    Span4Mux_h I__5893 (
            .O(N__42280),
            .I(N__42277));
    Span4Mux_v I__5892 (
            .O(N__42277),
            .I(N__42273));
    InMux I__5891 (
            .O(N__42276),
            .I(N__42270));
    Odrv4 I__5890 (
            .O(N__42273),
            .I(REG_mem_17_11));
    LocalMux I__5889 (
            .O(N__42270),
            .I(REG_mem_17_11));
    InMux I__5888 (
            .O(N__42265),
            .I(N__42259));
    InMux I__5887 (
            .O(N__42264),
            .I(N__42259));
    LocalMux I__5886 (
            .O(N__42259),
            .I(REG_mem_18_13));
    CascadeMux I__5885 (
            .O(N__42256),
            .I(N__42253));
    InMux I__5884 (
            .O(N__42253),
            .I(N__42247));
    InMux I__5883 (
            .O(N__42252),
            .I(N__42247));
    LocalMux I__5882 (
            .O(N__42247),
            .I(REG_mem_19_13));
    InMux I__5881 (
            .O(N__42244),
            .I(N__42241));
    LocalMux I__5880 (
            .O(N__42241),
            .I(N__42238));
    Span4Mux_h I__5879 (
            .O(N__42238),
            .I(N__42235));
    Span4Mux_v I__5878 (
            .O(N__42235),
            .I(N__42231));
    InMux I__5877 (
            .O(N__42234),
            .I(N__42228));
    Odrv4 I__5876 (
            .O(N__42231),
            .I(REG_mem_4_11));
    LocalMux I__5875 (
            .O(N__42228),
            .I(REG_mem_4_11));
    CascadeMux I__5874 (
            .O(N__42223),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11481_cascade_ ));
    InMux I__5873 (
            .O(N__42220),
            .I(N__42217));
    LocalMux I__5872 (
            .O(N__42217),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11420 ));
    InMux I__5871 (
            .O(N__42214),
            .I(N__42211));
    LocalMux I__5870 (
            .O(N__42211),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12527 ));
    CascadeMux I__5869 (
            .O(N__42208),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.full_max_w_cascade_ ));
    InMux I__5868 (
            .O(N__42205),
            .I(N__42202));
    LocalMux I__5867 (
            .O(N__42202),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12 ));
    CascadeMux I__5866 (
            .O(N__42199),
            .I(N__42196));
    InMux I__5865 (
            .O(N__42196),
            .I(N__42193));
    LocalMux I__5864 (
            .O(N__42193),
            .I(N__42190));
    Span4Mux_v I__5863 (
            .O(N__42190),
            .I(N__42186));
    CascadeMux I__5862 (
            .O(N__42189),
            .I(N__42183));
    Span4Mux_v I__5861 (
            .O(N__42186),
            .I(N__42180));
    InMux I__5860 (
            .O(N__42183),
            .I(N__42177));
    Odrv4 I__5859 (
            .O(N__42180),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_11 ));
    LocalMux I__5858 (
            .O(N__42177),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_11 ));
    InMux I__5857 (
            .O(N__42172),
            .I(N__42169));
    LocalMux I__5856 (
            .O(N__42169),
            .I(N__42166));
    Span4Mux_h I__5855 (
            .O(N__42166),
            .I(N__42162));
    InMux I__5854 (
            .O(N__42165),
            .I(N__42159));
    Odrv4 I__5853 (
            .O(N__42162),
            .I(REG_mem_41_11));
    LocalMux I__5852 (
            .O(N__42159),
            .I(REG_mem_41_11));
    InMux I__5851 (
            .O(N__42154),
            .I(N__42148));
    InMux I__5850 (
            .O(N__42153),
            .I(N__42148));
    LocalMux I__5849 (
            .O(N__42148),
            .I(REG_mem_17_13));
    CascadeMux I__5848 (
            .O(N__42145),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14102_cascade_ ));
    CascadeMux I__5847 (
            .O(N__42142),
            .I(N__42139));
    InMux I__5846 (
            .O(N__42139),
            .I(N__42136));
    LocalMux I__5845 (
            .O(N__42136),
            .I(N__42133));
    Span4Mux_h I__5844 (
            .O(N__42133),
            .I(N__42130));
    Sp12to4 I__5843 (
            .O(N__42130),
            .I(N__42127));
    Odrv12 I__5842 (
            .O(N__42127),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12108 ));
    InMux I__5841 (
            .O(N__42124),
            .I(N__42118));
    InMux I__5840 (
            .O(N__42123),
            .I(N__42118));
    LocalMux I__5839 (
            .O(N__42118),
            .I(REG_mem_16_13));
    InMux I__5838 (
            .O(N__42115),
            .I(N__42107));
    InMux I__5837 (
            .O(N__42114),
            .I(N__42096));
    InMux I__5836 (
            .O(N__42113),
            .I(N__42096));
    InMux I__5835 (
            .O(N__42112),
            .I(N__42096));
    InMux I__5834 (
            .O(N__42111),
            .I(N__42096));
    InMux I__5833 (
            .O(N__42110),
            .I(N__42096));
    LocalMux I__5832 (
            .O(N__42107),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7612 ));
    LocalMux I__5831 (
            .O(N__42096),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7612 ));
    CascadeMux I__5830 (
            .O(N__42091),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616_cascade_ ));
    InMux I__5829 (
            .O(N__42088),
            .I(N__42085));
    LocalMux I__5828 (
            .O(N__42085),
            .I(N__42081));
    InMux I__5827 (
            .O(N__42084),
            .I(N__42078));
    Odrv12 I__5826 (
            .O(N__42081),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_0 ));
    LocalMux I__5825 (
            .O(N__42078),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_0 ));
    InMux I__5824 (
            .O(N__42073),
            .I(N__42070));
    LocalMux I__5823 (
            .O(N__42070),
            .I(N__42066));
    CascadeMux I__5822 (
            .O(N__42069),
            .I(N__42063));
    Sp12to4 I__5821 (
            .O(N__42066),
            .I(N__42060));
    InMux I__5820 (
            .O(N__42063),
            .I(N__42057));
    Odrv12 I__5819 (
            .O(N__42060),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_0 ));
    LocalMux I__5818 (
            .O(N__42057),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_0 ));
    InMux I__5817 (
            .O(N__42052),
            .I(N__42049));
    LocalMux I__5816 (
            .O(N__42049),
            .I(N__42046));
    Span4Mux_v I__5815 (
            .O(N__42046),
            .I(N__42042));
    InMux I__5814 (
            .O(N__42045),
            .I(N__42039));
    Odrv4 I__5813 (
            .O(N__42042),
            .I(REG_mem_39_12));
    LocalMux I__5812 (
            .O(N__42039),
            .I(REG_mem_39_12));
    InMux I__5811 (
            .O(N__42034),
            .I(N__42031));
    LocalMux I__5810 (
            .O(N__42031),
            .I(N__42028));
    Span12Mux_s9_v I__5809 (
            .O(N__42028),
            .I(N__42024));
    InMux I__5808 (
            .O(N__42027),
            .I(N__42021));
    Odrv12 I__5807 (
            .O(N__42024),
            .I(REG_mem_41_15));
    LocalMux I__5806 (
            .O(N__42021),
            .I(REG_mem_41_15));
    CascadeMux I__5805 (
            .O(N__42016),
            .I(n10_cascade_));
    CascadeMux I__5804 (
            .O(N__42013),
            .I(N__42010));
    InMux I__5803 (
            .O(N__42010),
            .I(N__42007));
    LocalMux I__5802 (
            .O(N__42007),
            .I(N__42003));
    InMux I__5801 (
            .O(N__42006),
            .I(N__42000));
    Odrv12 I__5800 (
            .O(N__42003),
            .I(REG_mem_55_3));
    LocalMux I__5799 (
            .O(N__42000),
            .I(REG_mem_55_3));
    CascadeMux I__5798 (
            .O(N__41995),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_nxt_c_0_cascade_ ));
    CascadeMux I__5797 (
            .O(N__41992),
            .I(wr_addr_nxt_c_2_cascade_));
    InMux I__5796 (
            .O(N__41989),
            .I(N__41986));
    LocalMux I__5795 (
            .O(N__41986),
            .I(N__41983));
    Span4Mux_v I__5794 (
            .O(N__41983),
            .I(N__41980));
    Span4Mux_v I__5793 (
            .O(N__41980),
            .I(N__41976));
    InMux I__5792 (
            .O(N__41979),
            .I(N__41973));
    Odrv4 I__5791 (
            .O(N__41976),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_0 ));
    LocalMux I__5790 (
            .O(N__41973),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_0 ));
    InMux I__5789 (
            .O(N__41968),
            .I(N__41952));
    InMux I__5788 (
            .O(N__41967),
            .I(N__41952));
    InMux I__5787 (
            .O(N__41966),
            .I(N__41952));
    InMux I__5786 (
            .O(N__41965),
            .I(N__41952));
    InMux I__5785 (
            .O(N__41964),
            .I(N__41952));
    InMux I__5784 (
            .O(N__41963),
            .I(N__41949));
    LocalMux I__5783 (
            .O(N__41952),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13 ));
    LocalMux I__5782 (
            .O(N__41949),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13 ));
    InMux I__5781 (
            .O(N__41944),
            .I(N__41941));
    LocalMux I__5780 (
            .O(N__41941),
            .I(N__41937));
    CascadeMux I__5779 (
            .O(N__41940),
            .I(N__41934));
    Span4Mux_h I__5778 (
            .O(N__41937),
            .I(N__41931));
    InMux I__5777 (
            .O(N__41934),
            .I(N__41928));
    Odrv4 I__5776 (
            .O(N__41931),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_15 ));
    LocalMux I__5775 (
            .O(N__41928),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_15 ));
    InMux I__5774 (
            .O(N__41923),
            .I(N__41920));
    LocalMux I__5773 (
            .O(N__41920),
            .I(N__41917));
    Span4Mux_h I__5772 (
            .O(N__41917),
            .I(N__41913));
    InMux I__5771 (
            .O(N__41916),
            .I(N__41910));
    Odrv4 I__5770 (
            .O(N__41913),
            .I(REG_mem_38_14));
    LocalMux I__5769 (
            .O(N__41910),
            .I(REG_mem_38_14));
    InMux I__5768 (
            .O(N__41905),
            .I(N__41902));
    LocalMux I__5767 (
            .O(N__41902),
            .I(N__41899));
    Span4Mux_v I__5766 (
            .O(N__41899),
            .I(N__41896));
    Span4Mux_h I__5765 (
            .O(N__41896),
            .I(N__41893));
    Span4Mux_v I__5764 (
            .O(N__41893),
            .I(N__41890));
    Odrv4 I__5763 (
            .O(N__41890),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12356 ));
    InMux I__5762 (
            .O(N__41887),
            .I(N__41884));
    LocalMux I__5761 (
            .O(N__41884),
            .I(N__41880));
    InMux I__5760 (
            .O(N__41883),
            .I(N__41877));
    Odrv4 I__5759 (
            .O(N__41880),
            .I(REG_mem_16_0));
    LocalMux I__5758 (
            .O(N__41877),
            .I(REG_mem_16_0));
    InMux I__5757 (
            .O(N__41872),
            .I(N__41866));
    InMux I__5756 (
            .O(N__41871),
            .I(N__41866));
    LocalMux I__5755 (
            .O(N__41866),
            .I(REG_mem_39_14));
    CascadeMux I__5754 (
            .O(N__41863),
            .I(N__41860));
    InMux I__5753 (
            .O(N__41860),
            .I(N__41857));
    LocalMux I__5752 (
            .O(N__41857),
            .I(N__41853));
    InMux I__5751 (
            .O(N__41856),
            .I(N__41850));
    Odrv12 I__5750 (
            .O(N__41853),
            .I(REG_mem_43_0));
    LocalMux I__5749 (
            .O(N__41850),
            .I(REG_mem_43_0));
    InMux I__5748 (
            .O(N__41845),
            .I(N__41842));
    LocalMux I__5747 (
            .O(N__41842),
            .I(N__41839));
    Span4Mux_h I__5746 (
            .O(N__41839),
            .I(N__41835));
    InMux I__5745 (
            .O(N__41838),
            .I(N__41832));
    Odrv4 I__5744 (
            .O(N__41835),
            .I(REG_mem_43_14));
    LocalMux I__5743 (
            .O(N__41832),
            .I(REG_mem_43_14));
    CascadeMux I__5742 (
            .O(N__41827),
            .I(N__41824));
    InMux I__5741 (
            .O(N__41824),
            .I(N__41821));
    LocalMux I__5740 (
            .O(N__41821),
            .I(N__41818));
    Span4Mux_v I__5739 (
            .O(N__41818),
            .I(N__41815));
    Span4Mux_h I__5738 (
            .O(N__41815),
            .I(N__41811));
    InMux I__5737 (
            .O(N__41814),
            .I(N__41808));
    Odrv4 I__5736 (
            .O(N__41811),
            .I(REG_mem_8_14));
    LocalMux I__5735 (
            .O(N__41808),
            .I(REG_mem_8_14));
    InMux I__5734 (
            .O(N__41803),
            .I(N__41798));
    InMux I__5733 (
            .O(N__41802),
            .I(N__41794));
    InMux I__5732 (
            .O(N__41801),
            .I(N__41787));
    LocalMux I__5731 (
            .O(N__41798),
            .I(N__41779));
    InMux I__5730 (
            .O(N__41797),
            .I(N__41776));
    LocalMux I__5729 (
            .O(N__41794),
            .I(N__41762));
    InMux I__5728 (
            .O(N__41793),
            .I(N__41759));
    InMux I__5727 (
            .O(N__41792),
            .I(N__41752));
    InMux I__5726 (
            .O(N__41791),
            .I(N__41752));
    InMux I__5725 (
            .O(N__41790),
            .I(N__41752));
    LocalMux I__5724 (
            .O(N__41787),
            .I(N__41741));
    InMux I__5723 (
            .O(N__41786),
            .I(N__41738));
    InMux I__5722 (
            .O(N__41785),
            .I(N__41735));
    InMux I__5721 (
            .O(N__41784),
            .I(N__41732));
    InMux I__5720 (
            .O(N__41783),
            .I(N__41727));
    InMux I__5719 (
            .O(N__41782),
            .I(N__41727));
    Span4Mux_v I__5718 (
            .O(N__41779),
            .I(N__41714));
    LocalMux I__5717 (
            .O(N__41776),
            .I(N__41714));
    InMux I__5716 (
            .O(N__41775),
            .I(N__41711));
    InMux I__5715 (
            .O(N__41774),
            .I(N__41704));
    InMux I__5714 (
            .O(N__41773),
            .I(N__41704));
    InMux I__5713 (
            .O(N__41772),
            .I(N__41704));
    InMux I__5712 (
            .O(N__41771),
            .I(N__41701));
    InMux I__5711 (
            .O(N__41770),
            .I(N__41690));
    InMux I__5710 (
            .O(N__41769),
            .I(N__41690));
    InMux I__5709 (
            .O(N__41768),
            .I(N__41690));
    InMux I__5708 (
            .O(N__41767),
            .I(N__41690));
    InMux I__5707 (
            .O(N__41766),
            .I(N__41690));
    InMux I__5706 (
            .O(N__41765),
            .I(N__41682));
    Span4Mux_h I__5705 (
            .O(N__41762),
            .I(N__41675));
    LocalMux I__5704 (
            .O(N__41759),
            .I(N__41675));
    LocalMux I__5703 (
            .O(N__41752),
            .I(N__41675));
    InMux I__5702 (
            .O(N__41751),
            .I(N__41672));
    InMux I__5701 (
            .O(N__41750),
            .I(N__41660));
    InMux I__5700 (
            .O(N__41749),
            .I(N__41660));
    InMux I__5699 (
            .O(N__41748),
            .I(N__41660));
    InMux I__5698 (
            .O(N__41747),
            .I(N__41651));
    InMux I__5697 (
            .O(N__41746),
            .I(N__41651));
    InMux I__5696 (
            .O(N__41745),
            .I(N__41651));
    InMux I__5695 (
            .O(N__41744),
            .I(N__41651));
    Span4Mux_h I__5694 (
            .O(N__41741),
            .I(N__41639));
    LocalMux I__5693 (
            .O(N__41738),
            .I(N__41639));
    LocalMux I__5692 (
            .O(N__41735),
            .I(N__41639));
    LocalMux I__5691 (
            .O(N__41732),
            .I(N__41636));
    LocalMux I__5690 (
            .O(N__41727),
            .I(N__41633));
    InMux I__5689 (
            .O(N__41726),
            .I(N__41630));
    InMux I__5688 (
            .O(N__41725),
            .I(N__41623));
    InMux I__5687 (
            .O(N__41724),
            .I(N__41623));
    InMux I__5686 (
            .O(N__41723),
            .I(N__41623));
    InMux I__5685 (
            .O(N__41722),
            .I(N__41614));
    InMux I__5684 (
            .O(N__41721),
            .I(N__41614));
    InMux I__5683 (
            .O(N__41720),
            .I(N__41614));
    InMux I__5682 (
            .O(N__41719),
            .I(N__41614));
    Span4Mux_v I__5681 (
            .O(N__41714),
            .I(N__41603));
    LocalMux I__5680 (
            .O(N__41711),
            .I(N__41603));
    LocalMux I__5679 (
            .O(N__41704),
            .I(N__41603));
    LocalMux I__5678 (
            .O(N__41701),
            .I(N__41603));
    LocalMux I__5677 (
            .O(N__41690),
            .I(N__41600));
    InMux I__5676 (
            .O(N__41689),
            .I(N__41589));
    InMux I__5675 (
            .O(N__41688),
            .I(N__41589));
    InMux I__5674 (
            .O(N__41687),
            .I(N__41589));
    InMux I__5673 (
            .O(N__41686),
            .I(N__41589));
    InMux I__5672 (
            .O(N__41685),
            .I(N__41589));
    LocalMux I__5671 (
            .O(N__41682),
            .I(N__41586));
    Span4Mux_v I__5670 (
            .O(N__41675),
            .I(N__41581));
    LocalMux I__5669 (
            .O(N__41672),
            .I(N__41581));
    InMux I__5668 (
            .O(N__41671),
            .I(N__41578));
    InMux I__5667 (
            .O(N__41670),
            .I(N__41575));
    InMux I__5666 (
            .O(N__41669),
            .I(N__41572));
    InMux I__5665 (
            .O(N__41668),
            .I(N__41567));
    InMux I__5664 (
            .O(N__41667),
            .I(N__41567));
    LocalMux I__5663 (
            .O(N__41660),
            .I(N__41562));
    LocalMux I__5662 (
            .O(N__41651),
            .I(N__41562));
    InMux I__5661 (
            .O(N__41650),
            .I(N__41547));
    InMux I__5660 (
            .O(N__41649),
            .I(N__41547));
    InMux I__5659 (
            .O(N__41648),
            .I(N__41547));
    InMux I__5658 (
            .O(N__41647),
            .I(N__41547));
    InMux I__5657 (
            .O(N__41646),
            .I(N__41547));
    Span4Mux_v I__5656 (
            .O(N__41639),
            .I(N__41542));
    Span4Mux_h I__5655 (
            .O(N__41636),
            .I(N__41542));
    Span4Mux_v I__5654 (
            .O(N__41633),
            .I(N__41533));
    LocalMux I__5653 (
            .O(N__41630),
            .I(N__41533));
    LocalMux I__5652 (
            .O(N__41623),
            .I(N__41533));
    LocalMux I__5651 (
            .O(N__41614),
            .I(N__41533));
    InMux I__5650 (
            .O(N__41613),
            .I(N__41530));
    InMux I__5649 (
            .O(N__41612),
            .I(N__41524));
    Span4Mux_v I__5648 (
            .O(N__41603),
            .I(N__41521));
    Span4Mux_h I__5647 (
            .O(N__41600),
            .I(N__41512));
    LocalMux I__5646 (
            .O(N__41589),
            .I(N__41512));
    Span4Mux_v I__5645 (
            .O(N__41586),
            .I(N__41512));
    Span4Mux_h I__5644 (
            .O(N__41581),
            .I(N__41512));
    LocalMux I__5643 (
            .O(N__41578),
            .I(N__41509));
    LocalMux I__5642 (
            .O(N__41575),
            .I(N__41504));
    LocalMux I__5641 (
            .O(N__41572),
            .I(N__41504));
    LocalMux I__5640 (
            .O(N__41567),
            .I(N__41499));
    Span4Mux_h I__5639 (
            .O(N__41562),
            .I(N__41499));
    InMux I__5638 (
            .O(N__41561),
            .I(N__41496));
    InMux I__5637 (
            .O(N__41560),
            .I(N__41489));
    InMux I__5636 (
            .O(N__41559),
            .I(N__41489));
    InMux I__5635 (
            .O(N__41558),
            .I(N__41489));
    LocalMux I__5634 (
            .O(N__41547),
            .I(N__41480));
    Span4Mux_h I__5633 (
            .O(N__41542),
            .I(N__41480));
    Span4Mux_v I__5632 (
            .O(N__41533),
            .I(N__41480));
    LocalMux I__5631 (
            .O(N__41530),
            .I(N__41480));
    InMux I__5630 (
            .O(N__41529),
            .I(N__41473));
    InMux I__5629 (
            .O(N__41528),
            .I(N__41473));
    InMux I__5628 (
            .O(N__41527),
            .I(N__41473));
    LocalMux I__5627 (
            .O(N__41524),
            .I(N__41470));
    Span4Mux_h I__5626 (
            .O(N__41521),
            .I(N__41467));
    Span4Mux_v I__5625 (
            .O(N__41512),
            .I(N__41464));
    Span12Mux_v I__5624 (
            .O(N__41509),
            .I(N__41449));
    Span12Mux_h I__5623 (
            .O(N__41504),
            .I(N__41449));
    Sp12to4 I__5622 (
            .O(N__41499),
            .I(N__41449));
    LocalMux I__5621 (
            .O(N__41496),
            .I(N__41449));
    LocalMux I__5620 (
            .O(N__41489),
            .I(N__41449));
    Sp12to4 I__5619 (
            .O(N__41480),
            .I(N__41449));
    LocalMux I__5618 (
            .O(N__41473),
            .I(N__41449));
    Odrv12 I__5617 (
            .O(N__41470),
            .I(dc32_fifo_data_in_14));
    Odrv4 I__5616 (
            .O(N__41467),
            .I(dc32_fifo_data_in_14));
    Odrv4 I__5615 (
            .O(N__41464),
            .I(dc32_fifo_data_in_14));
    Odrv12 I__5614 (
            .O(N__41449),
            .I(dc32_fifo_data_in_14));
    InMux I__5613 (
            .O(N__41440),
            .I(N__41437));
    LocalMux I__5612 (
            .O(N__41437),
            .I(N__41433));
    InMux I__5611 (
            .O(N__41436),
            .I(N__41430));
    Odrv12 I__5610 (
            .O(N__41433),
            .I(REG_mem_42_14));
    LocalMux I__5609 (
            .O(N__41430),
            .I(REG_mem_42_14));
    InMux I__5608 (
            .O(N__41425),
            .I(N__41422));
    LocalMux I__5607 (
            .O(N__41422),
            .I(N__41419));
    Span4Mux_v I__5606 (
            .O(N__41419),
            .I(N__41416));
    Span4Mux_h I__5605 (
            .O(N__41416),
            .I(N__41413));
    Span4Mux_v I__5604 (
            .O(N__41413),
            .I(N__41409));
    InMux I__5603 (
            .O(N__41412),
            .I(N__41406));
    Odrv4 I__5602 (
            .O(N__41409),
            .I(REG_mem_7_3));
    LocalMux I__5601 (
            .O(N__41406),
            .I(REG_mem_7_3));
    CascadeMux I__5600 (
            .O(N__41401),
            .I(N__41398));
    InMux I__5599 (
            .O(N__41398),
            .I(N__41395));
    LocalMux I__5598 (
            .O(N__41395),
            .I(N__41391));
    InMux I__5597 (
            .O(N__41394),
            .I(N__41388));
    Odrv4 I__5596 (
            .O(N__41391),
            .I(REG_mem_23_15));
    LocalMux I__5595 (
            .O(N__41388),
            .I(REG_mem_23_15));
    InMux I__5594 (
            .O(N__41383),
            .I(N__41380));
    LocalMux I__5593 (
            .O(N__41380),
            .I(N__41376));
    CascadeMux I__5592 (
            .O(N__41379),
            .I(N__41373));
    Span4Mux_v I__5591 (
            .O(N__41376),
            .I(N__41370));
    InMux I__5590 (
            .O(N__41373),
            .I(N__41367));
    Odrv4 I__5589 (
            .O(N__41370),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_0 ));
    LocalMux I__5588 (
            .O(N__41367),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_0 ));
    InMux I__5587 (
            .O(N__41362),
            .I(N__41356));
    InMux I__5586 (
            .O(N__41361),
            .I(N__41356));
    LocalMux I__5585 (
            .O(N__41356),
            .I(REG_mem_55_0));
    CascadeMux I__5584 (
            .O(N__41353),
            .I(N__41350));
    InMux I__5583 (
            .O(N__41350),
            .I(N__41346));
    InMux I__5582 (
            .O(N__41349),
            .I(N__41343));
    LocalMux I__5581 (
            .O(N__41346),
            .I(REG_mem_41_0));
    LocalMux I__5580 (
            .O(N__41343),
            .I(REG_mem_41_0));
    InMux I__5579 (
            .O(N__41338),
            .I(N__41334));
    InMux I__5578 (
            .O(N__41337),
            .I(N__41331));
    LocalMux I__5577 (
            .O(N__41334),
            .I(REG_mem_42_0));
    LocalMux I__5576 (
            .O(N__41331),
            .I(REG_mem_42_0));
    InMux I__5575 (
            .O(N__41326),
            .I(N__41323));
    LocalMux I__5574 (
            .O(N__41323),
            .I(N__41319));
    InMux I__5573 (
            .O(N__41322),
            .I(N__41316));
    Odrv12 I__5572 (
            .O(N__41319),
            .I(REG_mem_9_14));
    LocalMux I__5571 (
            .O(N__41316),
            .I(REG_mem_9_14));
    InMux I__5570 (
            .O(N__41311),
            .I(N__41307));
    CascadeMux I__5569 (
            .O(N__41310),
            .I(N__41304));
    LocalMux I__5568 (
            .O(N__41307),
            .I(N__41301));
    InMux I__5567 (
            .O(N__41304),
            .I(N__41298));
    Odrv12 I__5566 (
            .O(N__41301),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_7 ));
    LocalMux I__5565 (
            .O(N__41298),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_7 ));
    InMux I__5564 (
            .O(N__41293),
            .I(N__41289));
    CascadeMux I__5563 (
            .O(N__41292),
            .I(N__41286));
    LocalMux I__5562 (
            .O(N__41289),
            .I(N__41283));
    InMux I__5561 (
            .O(N__41286),
            .I(N__41280));
    Odrv12 I__5560 (
            .O(N__41283),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_7 ));
    LocalMux I__5559 (
            .O(N__41280),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_7 ));
    InMux I__5558 (
            .O(N__41275),
            .I(N__41271));
    InMux I__5557 (
            .O(N__41274),
            .I(N__41268));
    LocalMux I__5556 (
            .O(N__41271),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_0 ));
    LocalMux I__5555 (
            .O(N__41268),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_0 ));
    InMux I__5554 (
            .O(N__41263),
            .I(N__41259));
    CascadeMux I__5553 (
            .O(N__41262),
            .I(N__41256));
    LocalMux I__5552 (
            .O(N__41259),
            .I(N__41253));
    InMux I__5551 (
            .O(N__41256),
            .I(N__41250));
    Odrv4 I__5550 (
            .O(N__41253),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_9 ));
    LocalMux I__5549 (
            .O(N__41250),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_9 ));
    InMux I__5548 (
            .O(N__41245),
            .I(N__41239));
    InMux I__5547 (
            .O(N__41244),
            .I(N__41239));
    LocalMux I__5546 (
            .O(N__41239),
            .I(REG_mem_23_9));
    InMux I__5545 (
            .O(N__41236),
            .I(N__41233));
    LocalMux I__5544 (
            .O(N__41233),
            .I(N__41230));
    Span4Mux_h I__5543 (
            .O(N__41230),
            .I(N__41226));
    InMux I__5542 (
            .O(N__41229),
            .I(N__41223));
    Odrv4 I__5541 (
            .O(N__41226),
            .I(REG_mem_55_1));
    LocalMux I__5540 (
            .O(N__41223),
            .I(REG_mem_55_1));
    InMux I__5539 (
            .O(N__41218),
            .I(N__41215));
    LocalMux I__5538 (
            .O(N__41215),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12938 ));
    CascadeMux I__5537 (
            .O(N__41212),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13112_cascade_ ));
    InMux I__5536 (
            .O(N__41209),
            .I(N__41206));
    LocalMux I__5535 (
            .O(N__41206),
            .I(N__41203));
    Odrv4 I__5534 (
            .O(N__41203),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13115 ));
    InMux I__5533 (
            .O(N__41200),
            .I(N__41196));
    CascadeMux I__5532 (
            .O(N__41199),
            .I(N__41193));
    LocalMux I__5531 (
            .O(N__41196),
            .I(N__41190));
    InMux I__5530 (
            .O(N__41193),
            .I(N__41187));
    Odrv4 I__5529 (
            .O(N__41190),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_0 ));
    LocalMux I__5528 (
            .O(N__41187),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_0 ));
    CascadeMux I__5527 (
            .O(N__41182),
            .I(N__41178));
    InMux I__5526 (
            .O(N__41181),
            .I(N__41173));
    InMux I__5525 (
            .O(N__41178),
            .I(N__41173));
    LocalMux I__5524 (
            .O(N__41173),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_0 ));
    CascadeMux I__5523 (
            .O(N__41170),
            .I(N__41166));
    InMux I__5522 (
            .O(N__41169),
            .I(N__41163));
    InMux I__5521 (
            .O(N__41166),
            .I(N__41160));
    LocalMux I__5520 (
            .O(N__41163),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_0 ));
    LocalMux I__5519 (
            .O(N__41160),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_0 ));
    InMux I__5518 (
            .O(N__41155),
            .I(N__41149));
    InMux I__5517 (
            .O(N__41154),
            .I(N__41149));
    LocalMux I__5516 (
            .O(N__41149),
            .I(REG_mem_7_9));
    CascadeMux I__5515 (
            .O(N__41146),
            .I(N__41143));
    InMux I__5514 (
            .O(N__41143),
            .I(N__41140));
    LocalMux I__5513 (
            .O(N__41140),
            .I(N__41137));
    Span4Mux_v I__5512 (
            .O(N__41137),
            .I(N__41134));
    Odrv4 I__5511 (
            .O(N__41134),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12344 ));
    CascadeMux I__5510 (
            .O(N__41131),
            .I(N__41128));
    InMux I__5509 (
            .O(N__41128),
            .I(N__41125));
    LocalMux I__5508 (
            .O(N__41125),
            .I(N__41122));
    Span4Mux_h I__5507 (
            .O(N__41122),
            .I(N__41119));
    Odrv4 I__5506 (
            .O(N__41119),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13706 ));
    InMux I__5505 (
            .O(N__41116),
            .I(N__41113));
    LocalMux I__5504 (
            .O(N__41113),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14156 ));
    CascadeMux I__5503 (
            .O(N__41110),
            .I(N__41107));
    InMux I__5502 (
            .O(N__41107),
            .I(N__41104));
    LocalMux I__5501 (
            .O(N__41104),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11998 ));
    InMux I__5500 (
            .O(N__41101),
            .I(N__41098));
    LocalMux I__5499 (
            .O(N__41098),
            .I(N__41095));
    Odrv4 I__5498 (
            .O(N__41095),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11999 ));
    InMux I__5497 (
            .O(N__41092),
            .I(N__41089));
    LocalMux I__5496 (
            .O(N__41089),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13673 ));
    CascadeMux I__5495 (
            .O(N__41086),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12080_cascade_ ));
    InMux I__5494 (
            .O(N__41083),
            .I(N__41080));
    LocalMux I__5493 (
            .O(N__41080),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14114 ));
    CascadeMux I__5492 (
            .O(N__41077),
            .I(N__41074));
    InMux I__5491 (
            .O(N__41074),
            .I(N__41071));
    LocalMux I__5490 (
            .O(N__41071),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11732 ));
    InMux I__5489 (
            .O(N__41068),
            .I(N__41065));
    LocalMux I__5488 (
            .O(N__41065),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11731 ));
    InMux I__5487 (
            .O(N__41062),
            .I(N__41059));
    LocalMux I__5486 (
            .O(N__41059),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13565 ));
    InMux I__5485 (
            .O(N__41056),
            .I(N__41053));
    LocalMux I__5484 (
            .O(N__41053),
            .I(N__41050));
    Span4Mux_v I__5483 (
            .O(N__41050),
            .I(N__41047));
    Span4Mux_h I__5482 (
            .O(N__41047),
            .I(N__41043));
    CascadeMux I__5481 (
            .O(N__41046),
            .I(N__41040));
    Span4Mux_v I__5480 (
            .O(N__41043),
            .I(N__41037));
    InMux I__5479 (
            .O(N__41040),
            .I(N__41034));
    Odrv4 I__5478 (
            .O(N__41037),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_14 ));
    LocalMux I__5477 (
            .O(N__41034),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_14 ));
    InMux I__5476 (
            .O(N__41029),
            .I(N__41026));
    LocalMux I__5475 (
            .O(N__41026),
            .I(N__41022));
    CascadeMux I__5474 (
            .O(N__41025),
            .I(N__41019));
    Span12Mux_v I__5473 (
            .O(N__41022),
            .I(N__41016));
    InMux I__5472 (
            .O(N__41019),
            .I(N__41013));
    Odrv12 I__5471 (
            .O(N__41016),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_14 ));
    LocalMux I__5470 (
            .O(N__41013),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_14 ));
    InMux I__5469 (
            .O(N__41008),
            .I(N__41005));
    LocalMux I__5468 (
            .O(N__41005),
            .I(N__41002));
    Span4Mux_v I__5467 (
            .O(N__41002),
            .I(N__40999));
    Span4Mux_h I__5466 (
            .O(N__40999),
            .I(N__40996));
    Odrv4 I__5465 (
            .O(N__40996),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12184 ));
    InMux I__5464 (
            .O(N__40993),
            .I(N__40989));
    CascadeMux I__5463 (
            .O(N__40992),
            .I(N__40986));
    LocalMux I__5462 (
            .O(N__40989),
            .I(N__40983));
    InMux I__5461 (
            .O(N__40986),
            .I(N__40980));
    Odrv12 I__5460 (
            .O(N__40983),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_0 ));
    LocalMux I__5459 (
            .O(N__40980),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_0 ));
    CascadeMux I__5458 (
            .O(N__40975),
            .I(N__40972));
    InMux I__5457 (
            .O(N__40972),
            .I(N__40969));
    LocalMux I__5456 (
            .O(N__40969),
            .I(N__40965));
    InMux I__5455 (
            .O(N__40968),
            .I(N__40962));
    Odrv4 I__5454 (
            .O(N__40965),
            .I(REG_mem_49_0));
    LocalMux I__5453 (
            .O(N__40962),
            .I(REG_mem_49_0));
    InMux I__5452 (
            .O(N__40957),
            .I(N__40954));
    LocalMux I__5451 (
            .O(N__40954),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11986 ));
    CascadeMux I__5450 (
            .O(N__40951),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13670_cascade_ ));
    InMux I__5449 (
            .O(N__40948),
            .I(N__40945));
    LocalMux I__5448 (
            .O(N__40945),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12013 ));
    InMux I__5447 (
            .O(N__40942),
            .I(N__40939));
    LocalMux I__5446 (
            .O(N__40939),
            .I(N__40936));
    Span4Mux_v I__5445 (
            .O(N__40936),
            .I(N__40933));
    Odrv4 I__5444 (
            .O(N__40933),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12020 ));
    CascadeMux I__5443 (
            .O(N__40930),
            .I(N__40927));
    InMux I__5442 (
            .O(N__40927),
            .I(N__40924));
    LocalMux I__5441 (
            .O(N__40924),
            .I(N__40921));
    Span4Mux_v I__5440 (
            .O(N__40921),
            .I(N__40918));
    Span4Mux_h I__5439 (
            .O(N__40918),
            .I(N__40915));
    Odrv4 I__5438 (
            .O(N__40915),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13676 ));
    CascadeMux I__5437 (
            .O(N__40912),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13679_cascade_ ));
    InMux I__5436 (
            .O(N__40909),
            .I(N__40906));
    LocalMux I__5435 (
            .O(N__40906),
            .I(N__40903));
    Span4Mux_v I__5434 (
            .O(N__40903),
            .I(N__40900));
    Odrv4 I__5433 (
            .O(N__40900),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12083 ));
    InMux I__5432 (
            .O(N__40897),
            .I(N__40893));
    InMux I__5431 (
            .O(N__40896),
            .I(N__40890));
    LocalMux I__5430 (
            .O(N__40893),
            .I(REG_mem_40_15));
    LocalMux I__5429 (
            .O(N__40890),
            .I(REG_mem_40_15));
    CascadeMux I__5428 (
            .O(N__40885),
            .I(N__40881));
    InMux I__5427 (
            .O(N__40884),
            .I(N__40876));
    InMux I__5426 (
            .O(N__40881),
            .I(N__40876));
    LocalMux I__5425 (
            .O(N__40876),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_1 ));
    CascadeMux I__5424 (
            .O(N__40873),
            .I(N__40869));
    InMux I__5423 (
            .O(N__40872),
            .I(N__40864));
    InMux I__5422 (
            .O(N__40869),
            .I(N__40864));
    LocalMux I__5421 (
            .O(N__40864),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_1 ));
    CascadeMux I__5420 (
            .O(N__40861),
            .I(N__40857));
    InMux I__5419 (
            .O(N__40860),
            .I(N__40854));
    InMux I__5418 (
            .O(N__40857),
            .I(N__40851));
    LocalMux I__5417 (
            .O(N__40854),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_15 ));
    LocalMux I__5416 (
            .O(N__40851),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_15 ));
    CascadeMux I__5415 (
            .O(N__40846),
            .I(N__40842));
    InMux I__5414 (
            .O(N__40845),
            .I(N__40837));
    InMux I__5413 (
            .O(N__40842),
            .I(N__40837));
    LocalMux I__5412 (
            .O(N__40837),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_15 ));
    CascadeMux I__5411 (
            .O(N__40834),
            .I(N__40830));
    InMux I__5410 (
            .O(N__40833),
            .I(N__40827));
    InMux I__5409 (
            .O(N__40830),
            .I(N__40824));
    LocalMux I__5408 (
            .O(N__40827),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_1 ));
    LocalMux I__5407 (
            .O(N__40824),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_1 ));
    CascadeMux I__5406 (
            .O(N__40819),
            .I(N__40815));
    InMux I__5405 (
            .O(N__40818),
            .I(N__40812));
    InMux I__5404 (
            .O(N__40815),
            .I(N__40809));
    LocalMux I__5403 (
            .O(N__40812),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_1 ));
    LocalMux I__5402 (
            .O(N__40809),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_1 ));
    CascadeMux I__5401 (
            .O(N__40804),
            .I(N__40800));
    InMux I__5400 (
            .O(N__40803),
            .I(N__40797));
    InMux I__5399 (
            .O(N__40800),
            .I(N__40794));
    LocalMux I__5398 (
            .O(N__40797),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_11 ));
    LocalMux I__5397 (
            .O(N__40794),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_11 ));
    CascadeMux I__5396 (
            .O(N__40789),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14366_cascade_ ));
    CascadeMux I__5395 (
            .O(N__40786),
            .I(N__40783));
    InMux I__5394 (
            .O(N__40783),
            .I(N__40779));
    InMux I__5393 (
            .O(N__40782),
            .I(N__40776));
    LocalMux I__5392 (
            .O(N__40779),
            .I(REG_mem_18_11));
    LocalMux I__5391 (
            .O(N__40776),
            .I(REG_mem_18_11));
    CascadeMux I__5390 (
            .O(N__40771),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14378_cascade_ ));
    InMux I__5389 (
            .O(N__40768),
            .I(N__40765));
    LocalMux I__5388 (
            .O(N__40765),
            .I(N__40761));
    InMux I__5387 (
            .O(N__40764),
            .I(N__40758));
    Odrv12 I__5386 (
            .O(N__40761),
            .I(REG_mem_16_11));
    LocalMux I__5385 (
            .O(N__40758),
            .I(REG_mem_16_11));
    InMux I__5384 (
            .O(N__40753),
            .I(N__40750));
    LocalMux I__5383 (
            .O(N__40750),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12471 ));
    CascadeMux I__5382 (
            .O(N__40747),
            .I(N__40744));
    InMux I__5381 (
            .O(N__40744),
            .I(N__40741));
    LocalMux I__5380 (
            .O(N__40741),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13436 ));
    CascadeMux I__5379 (
            .O(N__40738),
            .I(N__40734));
    InMux I__5378 (
            .O(N__40737),
            .I(N__40731));
    InMux I__5377 (
            .O(N__40734),
            .I(N__40728));
    LocalMux I__5376 (
            .O(N__40731),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_11 ));
    LocalMux I__5375 (
            .O(N__40728),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_11 ));
    InMux I__5374 (
            .O(N__40723),
            .I(N__40720));
    LocalMux I__5373 (
            .O(N__40720),
            .I(N__40717));
    Odrv4 I__5372 (
            .O(N__40717),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13439 ));
    InMux I__5371 (
            .O(N__40714),
            .I(N__40711));
    LocalMux I__5370 (
            .O(N__40711),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12953 ));
    CascadeMux I__5369 (
            .O(N__40708),
            .I(N__40705));
    InMux I__5368 (
            .O(N__40705),
            .I(N__40702));
    LocalMux I__5367 (
            .O(N__40702),
            .I(N__40698));
    InMux I__5366 (
            .O(N__40701),
            .I(N__40695));
    Odrv4 I__5365 (
            .O(N__40698),
            .I(REG_mem_23_13));
    LocalMux I__5364 (
            .O(N__40695),
            .I(REG_mem_23_13));
    InMux I__5363 (
            .O(N__40690),
            .I(N__40687));
    LocalMux I__5362 (
            .O(N__40687),
            .I(N__40684));
    Odrv12 I__5361 (
            .O(N__40684),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14066 ));
    CascadeMux I__5360 (
            .O(N__40681),
            .I(N__40677));
    CascadeMux I__5359 (
            .O(N__40680),
            .I(N__40674));
    InMux I__5358 (
            .O(N__40677),
            .I(N__40671));
    InMux I__5357 (
            .O(N__40674),
            .I(N__40668));
    LocalMux I__5356 (
            .O(N__40671),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_11 ));
    LocalMux I__5355 (
            .O(N__40668),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_11 ));
    InMux I__5354 (
            .O(N__40663),
            .I(N__40660));
    LocalMux I__5353 (
            .O(N__40660),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12950 ));
    CascadeMux I__5352 (
            .O(N__40657),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12075_cascade_ ));
    InMux I__5351 (
            .O(N__40654),
            .I(N__40651));
    LocalMux I__5350 (
            .O(N__40651),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13076 ));
    CascadeMux I__5349 (
            .O(N__40648),
            .I(N__40645));
    InMux I__5348 (
            .O(N__40645),
            .I(N__40642));
    LocalMux I__5347 (
            .O(N__40642),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14126 ));
    InMux I__5346 (
            .O(N__40639),
            .I(N__40636));
    LocalMux I__5345 (
            .O(N__40636),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12102 ));
    InMux I__5344 (
            .O(N__40633),
            .I(N__40630));
    LocalMux I__5343 (
            .O(N__40630),
            .I(N__40627));
    Span4Mux_h I__5342 (
            .O(N__40627),
            .I(N__40623));
    InMux I__5341 (
            .O(N__40626),
            .I(N__40620));
    Odrv4 I__5340 (
            .O(N__40623),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_12 ));
    LocalMux I__5339 (
            .O(N__40620),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_12 ));
    InMux I__5338 (
            .O(N__40615),
            .I(N__40609));
    InMux I__5337 (
            .O(N__40614),
            .I(N__40609));
    LocalMux I__5336 (
            .O(N__40609),
            .I(REG_mem_13_13));
    InMux I__5335 (
            .O(N__40606),
            .I(N__40600));
    InMux I__5334 (
            .O(N__40605),
            .I(N__40600));
    LocalMux I__5333 (
            .O(N__40600),
            .I(REG_mem_12_13));
    InMux I__5332 (
            .O(N__40597),
            .I(N__40591));
    InMux I__5331 (
            .O(N__40596),
            .I(N__40591));
    LocalMux I__5330 (
            .O(N__40591),
            .I(REG_mem_14_13));
    InMux I__5329 (
            .O(N__40588),
            .I(N__40585));
    LocalMux I__5328 (
            .O(N__40585),
            .I(N__40582));
    Span4Mux_v I__5327 (
            .O(N__40582),
            .I(N__40579));
    Span4Mux_h I__5326 (
            .O(N__40579),
            .I(N__40575));
    InMux I__5325 (
            .O(N__40578),
            .I(N__40572));
    Odrv4 I__5324 (
            .O(N__40575),
            .I(REG_mem_7_11));
    LocalMux I__5323 (
            .O(N__40572),
            .I(REG_mem_7_11));
    CascadeMux I__5322 (
            .O(N__40567),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12884_cascade_ ));
    CascadeMux I__5321 (
            .O(N__40564),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12887_cascade_ ));
    InMux I__5320 (
            .O(N__40561),
            .I(N__40555));
    InMux I__5319 (
            .O(N__40560),
            .I(N__40555));
    LocalMux I__5318 (
            .O(N__40555),
            .I(REG_mem_55_13));
    CascadeMux I__5317 (
            .O(N__40552),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13508_cascade_ ));
    InMux I__5316 (
            .O(N__40549),
            .I(N__40545));
    CascadeMux I__5315 (
            .O(N__40548),
            .I(N__40542));
    LocalMux I__5314 (
            .O(N__40545),
            .I(N__40539));
    InMux I__5313 (
            .O(N__40542),
            .I(N__40536));
    Odrv4 I__5312 (
            .O(N__40539),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_13 ));
    LocalMux I__5311 (
            .O(N__40536),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_13 ));
    InMux I__5310 (
            .O(N__40531),
            .I(N__40528));
    LocalMux I__5309 (
            .O(N__40528),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12276 ));
    CascadeMux I__5308 (
            .O(N__40525),
            .I(N__40522));
    InMux I__5307 (
            .O(N__40522),
            .I(N__40519));
    LocalMux I__5306 (
            .O(N__40519),
            .I(N__40515));
    InMux I__5305 (
            .O(N__40518),
            .I(N__40512));
    Span4Mux_h I__5304 (
            .O(N__40515),
            .I(N__40509));
    LocalMux I__5303 (
            .O(N__40512),
            .I(N__40506));
    Odrv4 I__5302 (
            .O(N__40509),
            .I(REG_mem_40_10));
    Odrv4 I__5301 (
            .O(N__40506),
            .I(REG_mem_40_10));
    CascadeMux I__5300 (
            .O(N__40501),
            .I(N__40497));
    InMux I__5299 (
            .O(N__40500),
            .I(N__40492));
    InMux I__5298 (
            .O(N__40497),
            .I(N__40492));
    LocalMux I__5297 (
            .O(N__40492),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_13 ));
    CascadeMux I__5296 (
            .O(N__40489),
            .I(N__40485));
    CascadeMux I__5295 (
            .O(N__40488),
            .I(N__40482));
    InMux I__5294 (
            .O(N__40485),
            .I(N__40477));
    InMux I__5293 (
            .O(N__40482),
            .I(N__40477));
    LocalMux I__5292 (
            .O(N__40477),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_13 ));
    CascadeMux I__5291 (
            .O(N__40474),
            .I(N__40470));
    InMux I__5290 (
            .O(N__40473),
            .I(N__40465));
    InMux I__5289 (
            .O(N__40470),
            .I(N__40465));
    LocalMux I__5288 (
            .O(N__40465),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_13 ));
    InMux I__5287 (
            .O(N__40462),
            .I(N__40459));
    LocalMux I__5286 (
            .O(N__40459),
            .I(N__40456));
    Span4Mux_h I__5285 (
            .O(N__40456),
            .I(N__40453));
    Odrv4 I__5284 (
            .O(N__40453),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12123 ));
    CascadeMux I__5283 (
            .O(N__40450),
            .I(N__40447));
    InMux I__5282 (
            .O(N__40447),
            .I(N__40444));
    LocalMux I__5281 (
            .O(N__40444),
            .I(N__40441));
    Span4Mux_v I__5280 (
            .O(N__40441),
            .I(N__40438));
    Odrv4 I__5279 (
            .O(N__40438),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14174 ));
    InMux I__5278 (
            .O(N__40435),
            .I(N__40432));
    LocalMux I__5277 (
            .O(N__40432),
            .I(N__40428));
    InMux I__5276 (
            .O(N__40431),
            .I(N__40425));
    Odrv4 I__5275 (
            .O(N__40428),
            .I(REG_mem_8_13));
    LocalMux I__5274 (
            .O(N__40425),
            .I(REG_mem_8_13));
    InMux I__5273 (
            .O(N__40420),
            .I(N__40417));
    LocalMux I__5272 (
            .O(N__40417),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13427 ));
    InMux I__5271 (
            .O(N__40414),
            .I(N__40411));
    LocalMux I__5270 (
            .O(N__40411),
            .I(N__40407));
    InMux I__5269 (
            .O(N__40410),
            .I(N__40404));
    Odrv4 I__5268 (
            .O(N__40407),
            .I(REG_mem_40_13));
    LocalMux I__5267 (
            .O(N__40404),
            .I(REG_mem_40_13));
    CascadeMux I__5266 (
            .O(N__40399),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13802_cascade_ ));
    CascadeMux I__5265 (
            .O(N__40396),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12204_cascade_ ));
    InMux I__5264 (
            .O(N__40393),
            .I(N__40390));
    LocalMux I__5263 (
            .O(N__40390),
            .I(N__40387));
    Odrv4 I__5262 (
            .O(N__40387),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12968 ));
    InMux I__5261 (
            .O(N__40384),
            .I(N__40381));
    LocalMux I__5260 (
            .O(N__40381),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12225 ));
    CascadeMux I__5259 (
            .O(N__40378),
            .I(N__40375));
    InMux I__5258 (
            .O(N__40375),
            .I(N__40372));
    LocalMux I__5257 (
            .O(N__40372),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13712 ));
    InMux I__5256 (
            .O(N__40369),
            .I(N__40363));
    InMux I__5255 (
            .O(N__40368),
            .I(N__40363));
    LocalMux I__5254 (
            .O(N__40363),
            .I(REG_mem_44_13));
    InMux I__5253 (
            .O(N__40360),
            .I(N__40354));
    InMux I__5252 (
            .O(N__40359),
            .I(N__40354));
    LocalMux I__5251 (
            .O(N__40354),
            .I(REG_mem_46_13));
    InMux I__5250 (
            .O(N__40351),
            .I(N__40347));
    CascadeMux I__5249 (
            .O(N__40350),
            .I(N__40344));
    LocalMux I__5248 (
            .O(N__40347),
            .I(N__40341));
    InMux I__5247 (
            .O(N__40344),
            .I(N__40338));
    Odrv12 I__5246 (
            .O(N__40341),
            .I(REG_mem_37_12));
    LocalMux I__5245 (
            .O(N__40338),
            .I(REG_mem_37_12));
    InMux I__5244 (
            .O(N__40333),
            .I(N__40327));
    InMux I__5243 (
            .O(N__40332),
            .I(N__40327));
    LocalMux I__5242 (
            .O(N__40327),
            .I(REG_mem_17_12));
    CascadeMux I__5241 (
            .O(N__40324),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13406_cascade_ ));
    InMux I__5240 (
            .O(N__40321),
            .I(N__40318));
    LocalMux I__5239 (
            .O(N__40318),
            .I(N__40315));
    Span4Mux_v I__5238 (
            .O(N__40315),
            .I(N__40312));
    Odrv4 I__5237 (
            .O(N__40312),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12312 ));
    InMux I__5236 (
            .O(N__40309),
            .I(N__40303));
    InMux I__5235 (
            .O(N__40308),
            .I(N__40303));
    LocalMux I__5234 (
            .O(N__40303),
            .I(REG_mem_16_12));
    InMux I__5233 (
            .O(N__40300),
            .I(N__40296));
    InMux I__5232 (
            .O(N__40299),
            .I(N__40293));
    LocalMux I__5231 (
            .O(N__40296),
            .I(REG_mem_38_12));
    LocalMux I__5230 (
            .O(N__40293),
            .I(REG_mem_38_12));
    InMux I__5229 (
            .O(N__40288),
            .I(N__40285));
    LocalMux I__5228 (
            .O(N__40285),
            .I(N__40282));
    Odrv12 I__5227 (
            .O(N__40282),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12482 ));
    InMux I__5226 (
            .O(N__40279),
            .I(N__40276));
    LocalMux I__5225 (
            .O(N__40276),
            .I(N__40273));
    Span4Mux_v I__5224 (
            .O(N__40273),
            .I(N__40269));
    InMux I__5223 (
            .O(N__40272),
            .I(N__40266));
    Odrv4 I__5222 (
            .O(N__40269),
            .I(REG_mem_4_12));
    LocalMux I__5221 (
            .O(N__40266),
            .I(REG_mem_4_12));
    InMux I__5220 (
            .O(N__40261),
            .I(N__40258));
    LocalMux I__5219 (
            .O(N__40258),
            .I(N__40254));
    InMux I__5218 (
            .O(N__40257),
            .I(N__40251));
    Odrv12 I__5217 (
            .O(N__40254),
            .I(REG_mem_37_11));
    LocalMux I__5216 (
            .O(N__40251),
            .I(REG_mem_37_11));
    InMux I__5215 (
            .O(N__40246),
            .I(N__40243));
    LocalMux I__5214 (
            .O(N__40243),
            .I(N__40239));
    InMux I__5213 (
            .O(N__40242),
            .I(N__40236));
    Odrv4 I__5212 (
            .O(N__40239),
            .I(REG_mem_36_11));
    LocalMux I__5211 (
            .O(N__40236),
            .I(REG_mem_36_11));
    InMux I__5210 (
            .O(N__40231),
            .I(N__40228));
    LocalMux I__5209 (
            .O(N__40228),
            .I(N__40225));
    Span4Mux_v I__5208 (
            .O(N__40225),
            .I(N__40222));
    Span4Mux_h I__5207 (
            .O(N__40222),
            .I(N__40218));
    InMux I__5206 (
            .O(N__40221),
            .I(N__40215));
    Odrv4 I__5205 (
            .O(N__40218),
            .I(REG_mem_47_14));
    LocalMux I__5204 (
            .O(N__40215),
            .I(REG_mem_47_14));
    InMux I__5203 (
            .O(N__40210),
            .I(N__40206));
    CascadeMux I__5202 (
            .O(N__40209),
            .I(N__40203));
    LocalMux I__5201 (
            .O(N__40206),
            .I(N__40200));
    InMux I__5200 (
            .O(N__40203),
            .I(N__40197));
    Odrv12 I__5199 (
            .O(N__40200),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_11 ));
    LocalMux I__5198 (
            .O(N__40197),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_11 ));
    InMux I__5197 (
            .O(N__40192),
            .I(N__40189));
    LocalMux I__5196 (
            .O(N__40189),
            .I(N__40185));
    CascadeMux I__5195 (
            .O(N__40188),
            .I(N__40182));
    Span12Mux_v I__5194 (
            .O(N__40185),
            .I(N__40179));
    InMux I__5193 (
            .O(N__40182),
            .I(N__40176));
    Odrv12 I__5192 (
            .O(N__40179),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_3 ));
    LocalMux I__5191 (
            .O(N__40176),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_3 ));
    InMux I__5190 (
            .O(N__40171),
            .I(N__40167));
    InMux I__5189 (
            .O(N__40170),
            .I(N__40164));
    LocalMux I__5188 (
            .O(N__40167),
            .I(REG_mem_44_3));
    LocalMux I__5187 (
            .O(N__40164),
            .I(REG_mem_44_3));
    InMux I__5186 (
            .O(N__40159),
            .I(N__40156));
    LocalMux I__5185 (
            .O(N__40156),
            .I(N__40152));
    InMux I__5184 (
            .O(N__40155),
            .I(N__40149));
    Odrv4 I__5183 (
            .O(N__40152),
            .I(REG_mem_36_12));
    LocalMux I__5182 (
            .O(N__40149),
            .I(REG_mem_36_12));
    CascadeMux I__5181 (
            .O(N__40144),
            .I(N__40140));
    InMux I__5180 (
            .O(N__40143),
            .I(N__40135));
    InMux I__5179 (
            .O(N__40140),
            .I(N__40135));
    LocalMux I__5178 (
            .O(N__40135),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_9 ));
    InMux I__5177 (
            .O(N__40132),
            .I(N__40129));
    LocalMux I__5176 (
            .O(N__40129),
            .I(N__40126));
    Span4Mux_v I__5175 (
            .O(N__40126),
            .I(N__40122));
    CascadeMux I__5174 (
            .O(N__40125),
            .I(N__40119));
    Span4Mux_h I__5173 (
            .O(N__40122),
            .I(N__40116));
    InMux I__5172 (
            .O(N__40119),
            .I(N__40113));
    Odrv4 I__5171 (
            .O(N__40116),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_9 ));
    LocalMux I__5170 (
            .O(N__40113),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_9 ));
    InMux I__5169 (
            .O(N__40108),
            .I(N__40105));
    LocalMux I__5168 (
            .O(N__40105),
            .I(N__40102));
    Span4Mux_v I__5167 (
            .O(N__40102),
            .I(N__40099));
    Span4Mux_v I__5166 (
            .O(N__40099),
            .I(N__40096));
    Odrv4 I__5165 (
            .O(N__40096),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12340 ));
    InMux I__5164 (
            .O(N__40093),
            .I(N__40090));
    LocalMux I__5163 (
            .O(N__40090),
            .I(N__40087));
    Span4Mux_v I__5162 (
            .O(N__40087),
            .I(N__40083));
    CascadeMux I__5161 (
            .O(N__40086),
            .I(N__40080));
    Span4Mux_v I__5160 (
            .O(N__40083),
            .I(N__40077));
    InMux I__5159 (
            .O(N__40080),
            .I(N__40074));
    Odrv4 I__5158 (
            .O(N__40077),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_12 ));
    LocalMux I__5157 (
            .O(N__40074),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_12 ));
    InMux I__5156 (
            .O(N__40069),
            .I(N__40066));
    LocalMux I__5155 (
            .O(N__40066),
            .I(N__40062));
    InMux I__5154 (
            .O(N__40065),
            .I(N__40059));
    Odrv4 I__5153 (
            .O(N__40062),
            .I(REG_mem_46_9));
    LocalMux I__5152 (
            .O(N__40059),
            .I(REG_mem_46_9));
    InMux I__5151 (
            .O(N__40054),
            .I(N__40050));
    InMux I__5150 (
            .O(N__40053),
            .I(N__40047));
    LocalMux I__5149 (
            .O(N__40050),
            .I(REG_mem_8_3));
    LocalMux I__5148 (
            .O(N__40047),
            .I(REG_mem_8_3));
    InMux I__5147 (
            .O(N__40042),
            .I(N__40039));
    LocalMux I__5146 (
            .O(N__40039),
            .I(N__40035));
    InMux I__5145 (
            .O(N__40038),
            .I(N__40032));
    Odrv12 I__5144 (
            .O(N__40035),
            .I(REG_mem_40_11));
    LocalMux I__5143 (
            .O(N__40032),
            .I(REG_mem_40_11));
    CascadeMux I__5142 (
            .O(N__40027),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n63_cascade_ ));
    CascadeMux I__5141 (
            .O(N__40024),
            .I(N__40021));
    InMux I__5140 (
            .O(N__40021),
            .I(N__40018));
    LocalMux I__5139 (
            .O(N__40018),
            .I(N__40014));
    InMux I__5138 (
            .O(N__40017),
            .I(N__40011));
    Span12Mux_v I__5137 (
            .O(N__40014),
            .I(N__40008));
    LocalMux I__5136 (
            .O(N__40011),
            .I(N__40005));
    Odrv12 I__5135 (
            .O(N__40008),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_0 ));
    Odrv4 I__5134 (
            .O(N__40005),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_0 ));
    CascadeMux I__5133 (
            .O(N__40000),
            .I(N__39997));
    InMux I__5132 (
            .O(N__39997),
            .I(N__39994));
    LocalMux I__5131 (
            .O(N__39994),
            .I(N__39991));
    Span4Mux_v I__5130 (
            .O(N__39991),
            .I(N__39988));
    Span4Mux_h I__5129 (
            .O(N__39988),
            .I(N__39984));
    InMux I__5128 (
            .O(N__39987),
            .I(N__39981));
    Odrv4 I__5127 (
            .O(N__39984),
            .I(REG_mem_50_14));
    LocalMux I__5126 (
            .O(N__39981),
            .I(REG_mem_50_14));
    InMux I__5125 (
            .O(N__39976),
            .I(N__39973));
    LocalMux I__5124 (
            .O(N__39973),
            .I(N__39970));
    Span4Mux_v I__5123 (
            .O(N__39970),
            .I(N__39966));
    InMux I__5122 (
            .O(N__39969),
            .I(N__39963));
    Odrv4 I__5121 (
            .O(N__39966),
            .I(REG_mem_44_11));
    LocalMux I__5120 (
            .O(N__39963),
            .I(REG_mem_44_11));
    CascadeMux I__5119 (
            .O(N__39958),
            .I(N__39954));
    InMux I__5118 (
            .O(N__39957),
            .I(N__39951));
    InMux I__5117 (
            .O(N__39954),
            .I(N__39948));
    LocalMux I__5116 (
            .O(N__39951),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_7 ));
    LocalMux I__5115 (
            .O(N__39948),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_7 ));
    InMux I__5114 (
            .O(N__39943),
            .I(N__39939));
    CascadeMux I__5113 (
            .O(N__39942),
            .I(N__39936));
    LocalMux I__5112 (
            .O(N__39939),
            .I(N__39933));
    InMux I__5111 (
            .O(N__39936),
            .I(N__39930));
    Odrv4 I__5110 (
            .O(N__39933),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_7 ));
    LocalMux I__5109 (
            .O(N__39930),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_7 ));
    InMux I__5108 (
            .O(N__39925),
            .I(N__39922));
    LocalMux I__5107 (
            .O(N__39922),
            .I(N__39919));
    Span4Mux_v I__5106 (
            .O(N__39919),
            .I(N__39915));
    CascadeMux I__5105 (
            .O(N__39918),
            .I(N__39912));
    Span4Mux_h I__5104 (
            .O(N__39915),
            .I(N__39909));
    InMux I__5103 (
            .O(N__39912),
            .I(N__39906));
    Odrv4 I__5102 (
            .O(N__39909),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_13 ));
    LocalMux I__5101 (
            .O(N__39906),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_13 ));
    CascadeMux I__5100 (
            .O(N__39901),
            .I(N__39898));
    InMux I__5099 (
            .O(N__39898),
            .I(N__39895));
    LocalMux I__5098 (
            .O(N__39895),
            .I(N__39891));
    CascadeMux I__5097 (
            .O(N__39894),
            .I(N__39888));
    Span4Mux_v I__5096 (
            .O(N__39891),
            .I(N__39885));
    InMux I__5095 (
            .O(N__39888),
            .I(N__39882));
    Odrv4 I__5094 (
            .O(N__39885),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_13 ));
    LocalMux I__5093 (
            .O(N__39882),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_13 ));
    CascadeMux I__5092 (
            .O(N__39877),
            .I(n53_cascade_));
    InMux I__5091 (
            .O(N__39874),
            .I(N__39871));
    LocalMux I__5090 (
            .O(N__39871),
            .I(N__39868));
    Span4Mux_h I__5089 (
            .O(N__39868),
            .I(N__39864));
    InMux I__5088 (
            .O(N__39867),
            .I(N__39861));
    Odrv4 I__5087 (
            .O(N__39864),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_0 ));
    LocalMux I__5086 (
            .O(N__39861),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_0 ));
    InMux I__5085 (
            .O(N__39856),
            .I(N__39853));
    LocalMux I__5084 (
            .O(N__39853),
            .I(N__39849));
    CascadeMux I__5083 (
            .O(N__39852),
            .I(N__39846));
    Span4Mux_v I__5082 (
            .O(N__39849),
            .I(N__39843));
    InMux I__5081 (
            .O(N__39846),
            .I(N__39840));
    Odrv4 I__5080 (
            .O(N__39843),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_5 ));
    LocalMux I__5079 (
            .O(N__39840),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_5 ));
    InMux I__5078 (
            .O(N__39835),
            .I(N__39832));
    LocalMux I__5077 (
            .O(N__39832),
            .I(N__39828));
    CascadeMux I__5076 (
            .O(N__39831),
            .I(N__39825));
    Span4Mux_v I__5075 (
            .O(N__39828),
            .I(N__39822));
    InMux I__5074 (
            .O(N__39825),
            .I(N__39819));
    Odrv4 I__5073 (
            .O(N__39822),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_0 ));
    LocalMux I__5072 (
            .O(N__39819),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_0 ));
    CascadeMux I__5071 (
            .O(N__39814),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53_cascade_ ));
    InMux I__5070 (
            .O(N__39811),
            .I(N__39808));
    LocalMux I__5069 (
            .O(N__39808),
            .I(N__39805));
    Span4Mux_v I__5068 (
            .O(N__39805),
            .I(N__39801));
    InMux I__5067 (
            .O(N__39804),
            .I(N__39798));
    Odrv4 I__5066 (
            .O(N__39801),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_0 ));
    LocalMux I__5065 (
            .O(N__39798),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_0 ));
    InMux I__5064 (
            .O(N__39793),
            .I(N__39790));
    LocalMux I__5063 (
            .O(N__39790),
            .I(N__39787));
    Span4Mux_h I__5062 (
            .O(N__39787),
            .I(N__39784));
    Span4Mux_h I__5061 (
            .O(N__39784),
            .I(N__39780));
    InMux I__5060 (
            .O(N__39783),
            .I(N__39777));
    Odrv4 I__5059 (
            .O(N__39780),
            .I(REG_mem_41_14));
    LocalMux I__5058 (
            .O(N__39777),
            .I(REG_mem_41_14));
    CascadeMux I__5057 (
            .O(N__39772),
            .I(N__39768));
    InMux I__5056 (
            .O(N__39771),
            .I(N__39765));
    InMux I__5055 (
            .O(N__39768),
            .I(N__39762));
    LocalMux I__5054 (
            .O(N__39765),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_12 ));
    LocalMux I__5053 (
            .O(N__39762),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_12 ));
    InMux I__5052 (
            .O(N__39757),
            .I(N__39754));
    LocalMux I__5051 (
            .O(N__39754),
            .I(N__39751));
    Span4Mux_v I__5050 (
            .O(N__39751),
            .I(N__39747));
    InMux I__5049 (
            .O(N__39750),
            .I(N__39744));
    Odrv4 I__5048 (
            .O(N__39747),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_15 ));
    LocalMux I__5047 (
            .O(N__39744),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_15 ));
    InMux I__5046 (
            .O(N__39739),
            .I(N__39736));
    LocalMux I__5045 (
            .O(N__39736),
            .I(N__39733));
    Span4Mux_v I__5044 (
            .O(N__39733),
            .I(N__39730));
    Span4Mux_h I__5043 (
            .O(N__39730),
            .I(N__39726));
    InMux I__5042 (
            .O(N__39729),
            .I(N__39723));
    Odrv4 I__5041 (
            .O(N__39726),
            .I(REG_mem_12_15));
    LocalMux I__5040 (
            .O(N__39723),
            .I(REG_mem_12_15));
    CascadeMux I__5039 (
            .O(N__39718),
            .I(N__39715));
    InMux I__5038 (
            .O(N__39715),
            .I(N__39711));
    CascadeMux I__5037 (
            .O(N__39714),
            .I(N__39708));
    LocalMux I__5036 (
            .O(N__39711),
            .I(N__39705));
    InMux I__5035 (
            .O(N__39708),
            .I(N__39702));
    Odrv4 I__5034 (
            .O(N__39705),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_0 ));
    LocalMux I__5033 (
            .O(N__39702),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_0 ));
    InMux I__5032 (
            .O(N__39697),
            .I(N__39694));
    LocalMux I__5031 (
            .O(N__39694),
            .I(N__39691));
    Span4Mux_v I__5030 (
            .O(N__39691),
            .I(N__39688));
    Span4Mux_h I__5029 (
            .O(N__39688),
            .I(N__39685));
    Span4Mux_h I__5028 (
            .O(N__39685),
            .I(N__39681));
    InMux I__5027 (
            .O(N__39684),
            .I(N__39678));
    Odrv4 I__5026 (
            .O(N__39681),
            .I(REG_mem_7_14));
    LocalMux I__5025 (
            .O(N__39678),
            .I(REG_mem_7_14));
    InMux I__5024 (
            .O(N__39673),
            .I(N__39670));
    LocalMux I__5023 (
            .O(N__39670),
            .I(N__39666));
    InMux I__5022 (
            .O(N__39669),
            .I(N__39663));
    Odrv12 I__5021 (
            .O(N__39666),
            .I(REG_mem_40_9));
    LocalMux I__5020 (
            .O(N__39663),
            .I(REG_mem_40_9));
    InMux I__5019 (
            .O(N__39658),
            .I(N__39655));
    LocalMux I__5018 (
            .O(N__39655),
            .I(N__39651));
    InMux I__5017 (
            .O(N__39654),
            .I(N__39648));
    Odrv4 I__5016 (
            .O(N__39651),
            .I(REG_mem_48_9));
    LocalMux I__5015 (
            .O(N__39648),
            .I(REG_mem_48_9));
    InMux I__5014 (
            .O(N__39643),
            .I(N__39640));
    LocalMux I__5013 (
            .O(N__39640),
            .I(N__39637));
    Span4Mux_v I__5012 (
            .O(N__39637),
            .I(N__39633));
    InMux I__5011 (
            .O(N__39636),
            .I(N__39630));
    Odrv4 I__5010 (
            .O(N__39633),
            .I(REG_mem_40_0));
    LocalMux I__5009 (
            .O(N__39630),
            .I(REG_mem_40_0));
    CascadeMux I__5008 (
            .O(N__39625),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12941_cascade_ ));
    InMux I__5007 (
            .O(N__39622),
            .I(N__39619));
    LocalMux I__5006 (
            .O(N__39619),
            .I(N__39616));
    Odrv4 I__5005 (
            .O(N__39616),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12815 ));
    CascadeMux I__5004 (
            .O(N__39613),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12095_cascade_ ));
    InMux I__5003 (
            .O(N__39610),
            .I(N__39607));
    LocalMux I__5002 (
            .O(N__39607),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12094 ));
    CascadeMux I__5001 (
            .O(N__39604),
            .I(N__39601));
    InMux I__5000 (
            .O(N__39601),
            .I(N__39597));
    InMux I__4999 (
            .O(N__39600),
            .I(N__39594));
    LocalMux I__4998 (
            .O(N__39597),
            .I(REG_mem_45_0));
    LocalMux I__4997 (
            .O(N__39594),
            .I(REG_mem_45_0));
    CascadeMux I__4996 (
            .O(N__39589),
            .I(N__39585));
    InMux I__4995 (
            .O(N__39588),
            .I(N__39582));
    InMux I__4994 (
            .O(N__39585),
            .I(N__39579));
    LocalMux I__4993 (
            .O(N__39582),
            .I(N__39576));
    LocalMux I__4992 (
            .O(N__39579),
            .I(N__39573));
    Odrv12 I__4991 (
            .O(N__39576),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_3 ));
    Odrv12 I__4990 (
            .O(N__39573),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_3 ));
    InMux I__4989 (
            .O(N__39568),
            .I(N__39564));
    CascadeMux I__4988 (
            .O(N__39567),
            .I(N__39561));
    LocalMux I__4987 (
            .O(N__39564),
            .I(N__39558));
    InMux I__4986 (
            .O(N__39561),
            .I(N__39555));
    Odrv12 I__4985 (
            .O(N__39558),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_12 ));
    LocalMux I__4984 (
            .O(N__39555),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_12 ));
    CascadeMux I__4983 (
            .O(N__39550),
            .I(N__39547));
    InMux I__4982 (
            .O(N__39547),
            .I(N__39544));
    LocalMux I__4981 (
            .O(N__39544),
            .I(N__39540));
    InMux I__4980 (
            .O(N__39543),
            .I(N__39537));
    Odrv4 I__4979 (
            .O(N__39540),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_0 ));
    LocalMux I__4978 (
            .O(N__39537),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_0 ));
    CascadeMux I__4977 (
            .O(N__39532),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13586_cascade_ ));
    InMux I__4976 (
            .O(N__39529),
            .I(N__39526));
    LocalMux I__4975 (
            .O(N__39526),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13589 ));
    InMux I__4974 (
            .O(N__39523),
            .I(N__39519));
    CascadeMux I__4973 (
            .O(N__39522),
            .I(N__39516));
    LocalMux I__4972 (
            .O(N__39519),
            .I(N__39513));
    InMux I__4971 (
            .O(N__39516),
            .I(N__39510));
    Odrv12 I__4970 (
            .O(N__39513),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_0 ));
    LocalMux I__4969 (
            .O(N__39510),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_0 ));
    InMux I__4968 (
            .O(N__39505),
            .I(N__39502));
    LocalMux I__4967 (
            .O(N__39502),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13502 ));
    CascadeMux I__4966 (
            .O(N__39499),
            .I(N__39496));
    InMux I__4965 (
            .O(N__39496),
            .I(N__39490));
    InMux I__4964 (
            .O(N__39495),
            .I(N__39490));
    LocalMux I__4963 (
            .O(N__39490),
            .I(REG_mem_23_0));
    InMux I__4962 (
            .O(N__39487),
            .I(N__39481));
    InMux I__4961 (
            .O(N__39486),
            .I(N__39481));
    LocalMux I__4960 (
            .O(N__39481),
            .I(REG_mem_17_0));
    InMux I__4959 (
            .O(N__39478),
            .I(N__39475));
    LocalMux I__4958 (
            .O(N__39475),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12920 ));
    InMux I__4957 (
            .O(N__39472),
            .I(N__39469));
    LocalMux I__4956 (
            .O(N__39469),
            .I(N__39466));
    Span4Mux_h I__4955 (
            .O(N__39466),
            .I(N__39463));
    Odrv4 I__4954 (
            .O(N__39463),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12445 ));
    InMux I__4953 (
            .O(N__39460),
            .I(N__39457));
    LocalMux I__4952 (
            .O(N__39457),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11495 ));
    InMux I__4951 (
            .O(N__39454),
            .I(N__39451));
    LocalMux I__4950 (
            .O(N__39451),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11492 ));
    CascadeMux I__4949 (
            .O(N__39448),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13172_cascade_ ));
    InMux I__4948 (
            .O(N__39445),
            .I(N__39442));
    LocalMux I__4947 (
            .O(N__39442),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12863 ));
    InMux I__4946 (
            .O(N__39439),
            .I(N__39436));
    LocalMux I__4945 (
            .O(N__39436),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13505 ));
    InMux I__4944 (
            .O(N__39433),
            .I(N__39430));
    LocalMux I__4943 (
            .O(N__39430),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12067 ));
    InMux I__4942 (
            .O(N__39427),
            .I(N__39424));
    LocalMux I__4941 (
            .O(N__39424),
            .I(N__39420));
    CascadeMux I__4940 (
            .O(N__39423),
            .I(N__39417));
    Span4Mux_v I__4939 (
            .O(N__39420),
            .I(N__39414));
    InMux I__4938 (
            .O(N__39417),
            .I(N__39411));
    Odrv4 I__4937 (
            .O(N__39414),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_0 ));
    LocalMux I__4936 (
            .O(N__39411),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_0 ));
    InMux I__4935 (
            .O(N__39406),
            .I(N__39402));
    InMux I__4934 (
            .O(N__39405),
            .I(N__39399));
    LocalMux I__4933 (
            .O(N__39402),
            .I(REG_mem_39_9));
    LocalMux I__4932 (
            .O(N__39399),
            .I(REG_mem_39_9));
    InMux I__4931 (
            .O(N__39394),
            .I(N__39391));
    LocalMux I__4930 (
            .O(N__39391),
            .I(N__39388));
    Odrv4 I__4929 (
            .O(N__39388),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12932 ));
    InMux I__4928 (
            .O(N__39385),
            .I(N__39382));
    LocalMux I__4927 (
            .O(N__39382),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13151 ));
    InMux I__4926 (
            .O(N__39379),
            .I(N__39376));
    LocalMux I__4925 (
            .O(N__39376),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13148 ));
    CascadeMux I__4924 (
            .O(N__39373),
            .I(N__39370));
    InMux I__4923 (
            .O(N__39370),
            .I(N__39366));
    InMux I__4922 (
            .O(N__39369),
            .I(N__39363));
    LocalMux I__4921 (
            .O(N__39366),
            .I(REG_mem_8_9));
    LocalMux I__4920 (
            .O(N__39363),
            .I(REG_mem_8_9));
    InMux I__4919 (
            .O(N__39358),
            .I(N__39355));
    LocalMux I__4918 (
            .O(N__39355),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11722 ));
    CascadeMux I__4917 (
            .O(N__39352),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11723_cascade_ ));
    InMux I__4916 (
            .O(N__39349),
            .I(N__39346));
    LocalMux I__4915 (
            .O(N__39346),
            .I(N__39343));
    Span4Mux_v I__4914 (
            .O(N__39343),
            .I(N__39339));
    InMux I__4913 (
            .O(N__39342),
            .I(N__39336));
    Odrv4 I__4912 (
            .O(N__39339),
            .I(REG_mem_48_0));
    LocalMux I__4911 (
            .O(N__39336),
            .I(REG_mem_48_0));
    InMux I__4910 (
            .O(N__39331),
            .I(N__39327));
    InMux I__4909 (
            .O(N__39330),
            .I(N__39324));
    LocalMux I__4908 (
            .O(N__39327),
            .I(REG_mem_50_15));
    LocalMux I__4907 (
            .O(N__39324),
            .I(REG_mem_50_15));
    InMux I__4906 (
            .O(N__39319),
            .I(N__39315));
    InMux I__4905 (
            .O(N__39318),
            .I(N__39312));
    LocalMux I__4904 (
            .O(N__39315),
            .I(REG_mem_44_15));
    LocalMux I__4903 (
            .O(N__39312),
            .I(REG_mem_44_15));
    InMux I__4902 (
            .O(N__39307),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10640 ));
    InMux I__4901 (
            .O(N__39304),
            .I(N__39300));
    InMux I__4900 (
            .O(N__39303),
            .I(N__39297));
    LocalMux I__4899 (
            .O(N__39300),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_5 ));
    LocalMux I__4898 (
            .O(N__39297),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_5 ));
    InMux I__4897 (
            .O(N__39292),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10641 ));
    InMux I__4896 (
            .O(N__39289),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10642 ));
    InMux I__4895 (
            .O(N__39286),
            .I(N__39283));
    LocalMux I__4894 (
            .O(N__39283),
            .I(N__39279));
    InMux I__4893 (
            .O(N__39282),
            .I(N__39276));
    Odrv4 I__4892 (
            .O(N__39279),
            .I(REG_mem_36_9));
    LocalMux I__4891 (
            .O(N__39276),
            .I(REG_mem_36_9));
    CascadeMux I__4890 (
            .O(N__39271),
            .I(N__39267));
    InMux I__4889 (
            .O(N__39270),
            .I(N__39262));
    InMux I__4888 (
            .O(N__39267),
            .I(N__39262));
    LocalMux I__4887 (
            .O(N__39262),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_1 ));
    CascadeMux I__4886 (
            .O(N__39259),
            .I(N__39255));
    InMux I__4885 (
            .O(N__39258),
            .I(N__39250));
    InMux I__4884 (
            .O(N__39255),
            .I(N__39250));
    LocalMux I__4883 (
            .O(N__39250),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_1 ));
    CascadeMux I__4882 (
            .O(N__39247),
            .I(rd_addr_nxt_c_6_N_465_5_cascade_));
    InMux I__4881 (
            .O(N__39244),
            .I(N__39241));
    LocalMux I__4880 (
            .O(N__39241),
            .I(N__39238));
    Odrv4 I__4879 (
            .O(N__39238),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12153 ));
    InMux I__4878 (
            .O(N__39235),
            .I(N__39232));
    LocalMux I__4877 (
            .O(N__39232),
            .I(N__39229));
    Span4Mux_h I__4876 (
            .O(N__39229),
            .I(N__39226));
    Span4Mux_v I__4875 (
            .O(N__39226),
            .I(N__39223));
    Odrv4 I__4874 (
            .O(N__39223),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12138 ));
    InMux I__4873 (
            .O(N__39220),
            .I(N__39217));
    LocalMux I__4872 (
            .O(N__39217),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13034 ));
    InMux I__4871 (
            .O(N__39214),
            .I(bfn_7_19_0_));
    InMux I__4870 (
            .O(N__39211),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10637 ));
    InMux I__4869 (
            .O(N__39208),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10638 ));
    InMux I__4868 (
            .O(N__39205),
            .I(N__39199));
    InMux I__4867 (
            .O(N__39204),
            .I(N__39199));
    LocalMux I__4866 (
            .O(N__39199),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_3 ));
    InMux I__4865 (
            .O(N__39196),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10639 ));
    CascadeMux I__4864 (
            .O(N__39193),
            .I(N__39190));
    InMux I__4863 (
            .O(N__39190),
            .I(N__39187));
    LocalMux I__4862 (
            .O(N__39187),
            .I(N__39184));
    Span4Mux_h I__4861 (
            .O(N__39184),
            .I(N__39181));
    Odrv4 I__4860 (
            .O(N__39181),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12902 ));
    InMux I__4859 (
            .O(N__39178),
            .I(N__39175));
    LocalMux I__4858 (
            .O(N__39175),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12420 ));
    CascadeMux I__4857 (
            .O(N__39172),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12405_cascade_ ));
    InMux I__4856 (
            .O(N__39169),
            .I(N__39166));
    LocalMux I__4855 (
            .O(N__39166),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12387 ));
    CascadeMux I__4854 (
            .O(N__39163),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12375_cascade_ ));
    InMux I__4853 (
            .O(N__39160),
            .I(N__39157));
    LocalMux I__4852 (
            .O(N__39157),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12794 ));
    CascadeMux I__4851 (
            .O(N__39154),
            .I(N__39151));
    InMux I__4850 (
            .O(N__39151),
            .I(N__39145));
    InMux I__4849 (
            .O(N__39150),
            .I(N__39145));
    LocalMux I__4848 (
            .O(N__39145),
            .I(REG_mem_46_7));
    InMux I__4847 (
            .O(N__39142),
            .I(N__39139));
    LocalMux I__4846 (
            .O(N__39139),
            .I(N__39136));
    Span4Mux_v I__4845 (
            .O(N__39136),
            .I(N__39133));
    Span4Mux_v I__4844 (
            .O(N__39133),
            .I(N__39130));
    Odrv4 I__4843 (
            .O(N__39130),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12517 ));
    InMux I__4842 (
            .O(N__39127),
            .I(N__39124));
    LocalMux I__4841 (
            .O(N__39124),
            .I(N__39121));
    Span4Mux_h I__4840 (
            .O(N__39121),
            .I(N__39118));
    Odrv4 I__4839 (
            .O(N__39118),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12518 ));
    InMux I__4838 (
            .O(N__39115),
            .I(N__39112));
    LocalMux I__4837 (
            .O(N__39112),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12506 ));
    CascadeMux I__4836 (
            .O(N__39109),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13310_cascade_ ));
    InMux I__4835 (
            .O(N__39106),
            .I(N__39103));
    LocalMux I__4834 (
            .O(N__39103),
            .I(N__39100));
    Odrv4 I__4833 (
            .O(N__39100),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13313 ));
    InMux I__4832 (
            .O(N__39097),
            .I(N__39094));
    LocalMux I__4831 (
            .O(N__39094),
            .I(N__39091));
    Odrv4 I__4830 (
            .O(N__39091),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13958 ));
    InMux I__4829 (
            .O(N__39088),
            .I(N__39085));
    LocalMux I__4828 (
            .O(N__39085),
            .I(N__39081));
    InMux I__4827 (
            .O(N__39084),
            .I(N__39078));
    Odrv12 I__4826 (
            .O(N__39081),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_13 ));
    LocalMux I__4825 (
            .O(N__39078),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_13 ));
    InMux I__4824 (
            .O(N__39073),
            .I(N__39070));
    LocalMux I__4823 (
            .O(N__39070),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12505 ));
    InMux I__4822 (
            .O(N__39067),
            .I(N__39061));
    InMux I__4821 (
            .O(N__39066),
            .I(N__39061));
    LocalMux I__4820 (
            .O(N__39061),
            .I(REG_mem_48_12));
    InMux I__4819 (
            .O(N__39058),
            .I(N__39052));
    InMux I__4818 (
            .O(N__39057),
            .I(N__39052));
    LocalMux I__4817 (
            .O(N__39052),
            .I(REG_mem_49_12));
    InMux I__4816 (
            .O(N__39049),
            .I(N__39046));
    LocalMux I__4815 (
            .O(N__39046),
            .I(N__39042));
    CascadeMux I__4814 (
            .O(N__39045),
            .I(N__39039));
    Span12Mux_v I__4813 (
            .O(N__39042),
            .I(N__39036));
    InMux I__4812 (
            .O(N__39039),
            .I(N__39033));
    Odrv12 I__4811 (
            .O(N__39036),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_12 ));
    LocalMux I__4810 (
            .O(N__39033),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_12 ));
    CascadeMux I__4809 (
            .O(N__39028),
            .I(N__39025));
    InMux I__4808 (
            .O(N__39025),
            .I(N__39022));
    LocalMux I__4807 (
            .O(N__39022),
            .I(N__39018));
    InMux I__4806 (
            .O(N__39021),
            .I(N__39015));
    Odrv4 I__4805 (
            .O(N__39018),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_13 ));
    LocalMux I__4804 (
            .O(N__39015),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_13 ));
    CascadeMux I__4803 (
            .O(N__39010),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13820_cascade_ ));
    CascadeMux I__4802 (
            .O(N__39007),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12198_cascade_ ));
    InMux I__4801 (
            .O(N__39004),
            .I(N__39001));
    LocalMux I__4800 (
            .O(N__39001),
            .I(N__38997));
    InMux I__4799 (
            .O(N__39000),
            .I(N__38994));
    Odrv12 I__4798 (
            .O(N__38997),
            .I(REG_mem_40_7));
    LocalMux I__4797 (
            .O(N__38994),
            .I(REG_mem_40_7));
    CascadeMux I__4796 (
            .O(N__38989),
            .I(N__38986));
    InMux I__4795 (
            .O(N__38986),
            .I(N__38983));
    LocalMux I__4794 (
            .O(N__38983),
            .I(N__38980));
    Odrv4 I__4793 (
            .O(N__38980),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13826 ));
    InMux I__4792 (
            .O(N__38977),
            .I(N__38974));
    LocalMux I__4791 (
            .O(N__38974),
            .I(N__38970));
    InMux I__4790 (
            .O(N__38973),
            .I(N__38967));
    Odrv12 I__4789 (
            .O(N__38970),
            .I(REG_mem_41_7));
    LocalMux I__4788 (
            .O(N__38967),
            .I(REG_mem_41_7));
    InMux I__4787 (
            .O(N__38962),
            .I(N__38959));
    LocalMux I__4786 (
            .O(N__38959),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12195 ));
    CascadeMux I__4785 (
            .O(N__38956),
            .I(N__38952));
    InMux I__4784 (
            .O(N__38955),
            .I(N__38949));
    InMux I__4783 (
            .O(N__38952),
            .I(N__38946));
    LocalMux I__4782 (
            .O(N__38949),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_12 ));
    LocalMux I__4781 (
            .O(N__38946),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_12 ));
    InMux I__4780 (
            .O(N__38941),
            .I(N__38937));
    InMux I__4779 (
            .O(N__38940),
            .I(N__38934));
    LocalMux I__4778 (
            .O(N__38937),
            .I(REG_mem_45_7));
    LocalMux I__4777 (
            .O(N__38934),
            .I(REG_mem_45_7));
    InMux I__4776 (
            .O(N__38929),
            .I(N__38923));
    InMux I__4775 (
            .O(N__38928),
            .I(N__38923));
    LocalMux I__4774 (
            .O(N__38923),
            .I(REG_mem_44_7));
    InMux I__4773 (
            .O(N__38920),
            .I(N__38914));
    InMux I__4772 (
            .O(N__38919),
            .I(N__38914));
    LocalMux I__4771 (
            .O(N__38914),
            .I(REG_mem_46_3));
    InMux I__4770 (
            .O(N__38911),
            .I(N__38908));
    LocalMux I__4769 (
            .O(N__38908),
            .I(N__38905));
    Span4Mux_v I__4768 (
            .O(N__38905),
            .I(N__38902));
    Span4Mux_h I__4767 (
            .O(N__38902),
            .I(N__38898));
    InMux I__4766 (
            .O(N__38901),
            .I(N__38895));
    Odrv4 I__4765 (
            .O(N__38898),
            .I(REG_mem_23_10));
    LocalMux I__4764 (
            .O(N__38895),
            .I(REG_mem_23_10));
    CascadeMux I__4763 (
            .O(N__38890),
            .I(N__38887));
    InMux I__4762 (
            .O(N__38887),
            .I(N__38884));
    LocalMux I__4761 (
            .O(N__38884),
            .I(N__38880));
    InMux I__4760 (
            .O(N__38883),
            .I(N__38877));
    Odrv12 I__4759 (
            .O(N__38880),
            .I(REG_mem_10_7));
    LocalMux I__4758 (
            .O(N__38877),
            .I(REG_mem_10_7));
    InMux I__4757 (
            .O(N__38872),
            .I(N__38869));
    LocalMux I__4756 (
            .O(N__38869),
            .I(N__38866));
    Span4Mux_v I__4755 (
            .O(N__38866),
            .I(N__38863));
    Odrv4 I__4754 (
            .O(N__38863),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14354 ));
    CascadeMux I__4753 (
            .O(N__38860),
            .I(N__38857));
    InMux I__4752 (
            .O(N__38857),
            .I(N__38854));
    LocalMux I__4751 (
            .O(N__38854),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13757 ));
    InMux I__4750 (
            .O(N__38851),
            .I(N__38848));
    LocalMux I__4749 (
            .O(N__38848),
            .I(N__38845));
    Span4Mux_v I__4748 (
            .O(N__38845),
            .I(N__38841));
    InMux I__4747 (
            .O(N__38844),
            .I(N__38838));
    Odrv4 I__4746 (
            .O(N__38841),
            .I(REG_mem_23_12));
    LocalMux I__4745 (
            .O(N__38838),
            .I(REG_mem_23_12));
    InMux I__4744 (
            .O(N__38833),
            .I(N__38830));
    LocalMux I__4743 (
            .O(N__38830),
            .I(N__38826));
    CascadeMux I__4742 (
            .O(N__38829),
            .I(N__38823));
    Span12Mux_s10_h I__4741 (
            .O(N__38826),
            .I(N__38820));
    InMux I__4740 (
            .O(N__38823),
            .I(N__38817));
    Odrv12 I__4739 (
            .O(N__38820),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_3 ));
    LocalMux I__4738 (
            .O(N__38817),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_3 ));
    InMux I__4737 (
            .O(N__38812),
            .I(N__38808));
    InMux I__4736 (
            .O(N__38811),
            .I(N__38805));
    LocalMux I__4735 (
            .O(N__38808),
            .I(REG_mem_47_12));
    LocalMux I__4734 (
            .O(N__38805),
            .I(REG_mem_47_12));
    InMux I__4733 (
            .O(N__38800),
            .I(N__38797));
    LocalMux I__4732 (
            .O(N__38797),
            .I(N__38794));
    Span4Mux_v I__4731 (
            .O(N__38794),
            .I(N__38790));
    InMux I__4730 (
            .O(N__38793),
            .I(N__38787));
    Odrv4 I__4729 (
            .O(N__38790),
            .I(REG_mem_63_12));
    LocalMux I__4728 (
            .O(N__38787),
            .I(REG_mem_63_12));
    InMux I__4727 (
            .O(N__38782),
            .I(N__38779));
    LocalMux I__4726 (
            .O(N__38779),
            .I(N__38775));
    InMux I__4725 (
            .O(N__38778),
            .I(N__38772));
    Span4Mux_v I__4724 (
            .O(N__38775),
            .I(N__38769));
    LocalMux I__4723 (
            .O(N__38772),
            .I(N__38766));
    Odrv4 I__4722 (
            .O(N__38769),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_12 ));
    Odrv4 I__4721 (
            .O(N__38766),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_12 ));
    CascadeMux I__4720 (
            .O(N__38761),
            .I(N__38758));
    InMux I__4719 (
            .O(N__38758),
            .I(N__38755));
    LocalMux I__4718 (
            .O(N__38755),
            .I(N__38752));
    Span4Mux_v I__4717 (
            .O(N__38752),
            .I(N__38749));
    Span4Mux_h I__4716 (
            .O(N__38749),
            .I(N__38745));
    InMux I__4715 (
            .O(N__38748),
            .I(N__38742));
    Odrv4 I__4714 (
            .O(N__38745),
            .I(REG_mem_15_7));
    LocalMux I__4713 (
            .O(N__38742),
            .I(REG_mem_15_7));
    InMux I__4712 (
            .O(N__38737),
            .I(N__38731));
    InMux I__4711 (
            .O(N__38736),
            .I(N__38731));
    LocalMux I__4710 (
            .O(N__38731),
            .I(REG_mem_9_3));
    CascadeMux I__4709 (
            .O(N__38728),
            .I(N__38725));
    InMux I__4708 (
            .O(N__38725),
            .I(N__38722));
    LocalMux I__4707 (
            .O(N__38722),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13088 ));
    InMux I__4706 (
            .O(N__38719),
            .I(N__38716));
    LocalMux I__4705 (
            .O(N__38716),
            .I(N__38713));
    Span4Mux_v I__4704 (
            .O(N__38713),
            .I(N__38710));
    Odrv4 I__4703 (
            .O(N__38710),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11598 ));
    InMux I__4702 (
            .O(N__38707),
            .I(N__38704));
    LocalMux I__4701 (
            .O(N__38704),
            .I(N__38701));
    Span4Mux_h I__4700 (
            .O(N__38701),
            .I(N__38697));
    InMux I__4699 (
            .O(N__38700),
            .I(N__38694));
    Odrv4 I__4698 (
            .O(N__38697),
            .I(REG_mem_11_7));
    LocalMux I__4697 (
            .O(N__38694),
            .I(REG_mem_11_7));
    CascadeMux I__4696 (
            .O(N__38689),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13334_cascade_ ));
    InMux I__4695 (
            .O(N__38686),
            .I(N__38683));
    LocalMux I__4694 (
            .O(N__38683),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13337 ));
    InMux I__4693 (
            .O(N__38680),
            .I(N__38674));
    InMux I__4692 (
            .O(N__38679),
            .I(N__38674));
    LocalMux I__4691 (
            .O(N__38674),
            .I(REG_mem_45_3));
    InMux I__4690 (
            .O(N__38671),
            .I(N__38667));
    CascadeMux I__4689 (
            .O(N__38670),
            .I(N__38664));
    LocalMux I__4688 (
            .O(N__38667),
            .I(N__38661));
    InMux I__4687 (
            .O(N__38664),
            .I(N__38658));
    Odrv12 I__4686 (
            .O(N__38661),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_7 ));
    LocalMux I__4685 (
            .O(N__38658),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_7 ));
    CascadeMux I__4684 (
            .O(N__38653),
            .I(N__38650));
    InMux I__4683 (
            .O(N__38650),
            .I(N__38647));
    LocalMux I__4682 (
            .O(N__38647),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13700 ));
    InMux I__4681 (
            .O(N__38644),
            .I(N__38641));
    LocalMux I__4680 (
            .O(N__38641),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13652 ));
    CascadeMux I__4679 (
            .O(N__38638),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12237_cascade_ ));
    InMux I__4678 (
            .O(N__38635),
            .I(N__38632));
    LocalMux I__4677 (
            .O(N__38632),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12228 ));
    InMux I__4676 (
            .O(N__38629),
            .I(N__38626));
    LocalMux I__4675 (
            .O(N__38626),
            .I(N__38623));
    Span4Mux_v I__4674 (
            .O(N__38623),
            .I(N__38619));
    CascadeMux I__4673 (
            .O(N__38622),
            .I(N__38616));
    Span4Mux_h I__4672 (
            .O(N__38619),
            .I(N__38613));
    InMux I__4671 (
            .O(N__38616),
            .I(N__38610));
    Odrv4 I__4670 (
            .O(N__38613),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_3 ));
    LocalMux I__4669 (
            .O(N__38610),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_3 ));
    InMux I__4668 (
            .O(N__38605),
            .I(N__38599));
    InMux I__4667 (
            .O(N__38604),
            .I(N__38599));
    LocalMux I__4666 (
            .O(N__38599),
            .I(REG_mem_58_7));
    CascadeMux I__4665 (
            .O(N__38596),
            .I(N__38592));
    CascadeMux I__4664 (
            .O(N__38595),
            .I(N__38589));
    InMux I__4663 (
            .O(N__38592),
            .I(N__38584));
    InMux I__4662 (
            .O(N__38589),
            .I(N__38584));
    LocalMux I__4661 (
            .O(N__38584),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_7 ));
    InMux I__4660 (
            .O(N__38581),
            .I(N__38578));
    LocalMux I__4659 (
            .O(N__38578),
            .I(N__38575));
    Span4Mux_v I__4658 (
            .O(N__38575),
            .I(N__38572));
    Span4Mux_h I__4657 (
            .O(N__38572),
            .I(N__38568));
    InMux I__4656 (
            .O(N__38571),
            .I(N__38565));
    Odrv4 I__4655 (
            .O(N__38568),
            .I(REG_mem_8_7));
    LocalMux I__4654 (
            .O(N__38565),
            .I(REG_mem_8_7));
    InMux I__4653 (
            .O(N__38560),
            .I(N__38557));
    LocalMux I__4652 (
            .O(N__38557),
            .I(N__38554));
    Span4Mux_h I__4651 (
            .O(N__38554),
            .I(N__38550));
    InMux I__4650 (
            .O(N__38553),
            .I(N__38547));
    Odrv4 I__4649 (
            .O(N__38550),
            .I(REG_mem_4_3));
    LocalMux I__4648 (
            .O(N__38547),
            .I(REG_mem_4_3));
    InMux I__4647 (
            .O(N__38542),
            .I(N__38538));
    InMux I__4646 (
            .O(N__38541),
            .I(N__38535));
    LocalMux I__4645 (
            .O(N__38538),
            .I(REG_mem_40_3));
    LocalMux I__4644 (
            .O(N__38535),
            .I(REG_mem_40_3));
    InMux I__4643 (
            .O(N__38530),
            .I(N__38527));
    LocalMux I__4642 (
            .O(N__38527),
            .I(N__38524));
    Span4Mux_h I__4641 (
            .O(N__38524),
            .I(N__38520));
    InMux I__4640 (
            .O(N__38523),
            .I(N__38517));
    Odrv4 I__4639 (
            .O(N__38520),
            .I(REG_mem_51_14));
    LocalMux I__4638 (
            .O(N__38517),
            .I(REG_mem_51_14));
    InMux I__4637 (
            .O(N__38512),
            .I(N__38509));
    LocalMux I__4636 (
            .O(N__38509),
            .I(N__38505));
    InMux I__4635 (
            .O(N__38508),
            .I(N__38502));
    Odrv12 I__4634 (
            .O(N__38505),
            .I(REG_mem_17_10));
    LocalMux I__4633 (
            .O(N__38502),
            .I(REG_mem_17_10));
    InMux I__4632 (
            .O(N__38497),
            .I(N__38494));
    LocalMux I__4631 (
            .O(N__38494),
            .I(N__38490));
    InMux I__4630 (
            .O(N__38493),
            .I(N__38487));
    Span4Mux_h I__4629 (
            .O(N__38490),
            .I(N__38484));
    LocalMux I__4628 (
            .O(N__38487),
            .I(N__38481));
    Odrv4 I__4627 (
            .O(N__38484),
            .I(REG_mem_63_7));
    Odrv4 I__4626 (
            .O(N__38481),
            .I(REG_mem_63_7));
    InMux I__4625 (
            .O(N__38476),
            .I(N__38473));
    LocalMux I__4624 (
            .O(N__38473),
            .I(N__38470));
    Span4Mux_v I__4623 (
            .O(N__38470),
            .I(N__38466));
    InMux I__4622 (
            .O(N__38469),
            .I(N__38463));
    Odrv4 I__4621 (
            .O(N__38466),
            .I(REG_mem_5_3));
    LocalMux I__4620 (
            .O(N__38463),
            .I(REG_mem_5_3));
    CascadeMux I__4619 (
            .O(N__38458),
            .I(N__38455));
    InMux I__4618 (
            .O(N__38455),
            .I(N__38452));
    LocalMux I__4617 (
            .O(N__38452),
            .I(N__38448));
    InMux I__4616 (
            .O(N__38451),
            .I(N__38445));
    Odrv12 I__4615 (
            .O(N__38448),
            .I(REG_mem_50_3));
    LocalMux I__4614 (
            .O(N__38445),
            .I(REG_mem_50_3));
    InMux I__4613 (
            .O(N__38440),
            .I(N__38437));
    LocalMux I__4612 (
            .O(N__38437),
            .I(N__38434));
    Span4Mux_v I__4611 (
            .O(N__38434),
            .I(N__38430));
    CascadeMux I__4610 (
            .O(N__38433),
            .I(N__38427));
    Span4Mux_v I__4609 (
            .O(N__38430),
            .I(N__38424));
    InMux I__4608 (
            .O(N__38427),
            .I(N__38421));
    Odrv4 I__4607 (
            .O(N__38424),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_12 ));
    LocalMux I__4606 (
            .O(N__38421),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_12 ));
    InMux I__4605 (
            .O(N__38416),
            .I(N__38413));
    LocalMux I__4604 (
            .O(N__38413),
            .I(N__38410));
    Span4Mux_v I__4603 (
            .O(N__38410),
            .I(N__38407));
    Span4Mux_h I__4602 (
            .O(N__38407),
            .I(N__38403));
    InMux I__4601 (
            .O(N__38406),
            .I(N__38400));
    Odrv4 I__4600 (
            .O(N__38403),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_7 ));
    LocalMux I__4599 (
            .O(N__38400),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_7 ));
    InMux I__4598 (
            .O(N__38395),
            .I(N__38392));
    LocalMux I__4597 (
            .O(N__38392),
            .I(N__38389));
    Span4Mux_h I__4596 (
            .O(N__38389),
            .I(N__38385));
    InMux I__4595 (
            .O(N__38388),
            .I(N__38382));
    Odrv4 I__4594 (
            .O(N__38385),
            .I(REG_mem_15_10));
    LocalMux I__4593 (
            .O(N__38382),
            .I(REG_mem_15_10));
    InMux I__4592 (
            .O(N__38377),
            .I(N__38373));
    InMux I__4591 (
            .O(N__38376),
            .I(N__38370));
    LocalMux I__4590 (
            .O(N__38373),
            .I(REG_mem_13_10));
    LocalMux I__4589 (
            .O(N__38370),
            .I(REG_mem_13_10));
    CascadeMux I__4588 (
            .O(N__38365),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14162_cascade_ ));
    InMux I__4587 (
            .O(N__38362),
            .I(N__38359));
    LocalMux I__4586 (
            .O(N__38359),
            .I(N__38356));
    Span12Mux_s10_h I__4585 (
            .O(N__38356),
            .I(N__38353));
    Odrv12 I__4584 (
            .O(N__38353),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14165 ));
    InMux I__4583 (
            .O(N__38350),
            .I(N__38344));
    InMux I__4582 (
            .O(N__38349),
            .I(N__38344));
    LocalMux I__4581 (
            .O(N__38344),
            .I(REG_mem_12_10));
    InMux I__4580 (
            .O(N__38341),
            .I(N__38335));
    InMux I__4579 (
            .O(N__38340),
            .I(N__38335));
    LocalMux I__4578 (
            .O(N__38335),
            .I(REG_mem_14_10));
    InMux I__4577 (
            .O(N__38332),
            .I(N__38329));
    LocalMux I__4576 (
            .O(N__38329),
            .I(N__38326));
    Span4Mux_v I__4575 (
            .O(N__38326),
            .I(N__38322));
    InMux I__4574 (
            .O(N__38325),
            .I(N__38319));
    Odrv4 I__4573 (
            .O(N__38322),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_13 ));
    LocalMux I__4572 (
            .O(N__38319),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_13 ));
    InMux I__4571 (
            .O(N__38314),
            .I(N__38311));
    LocalMux I__4570 (
            .O(N__38311),
            .I(N__38308));
    Span4Mux_v I__4569 (
            .O(N__38308),
            .I(N__38305));
    Span4Mux_h I__4568 (
            .O(N__38305),
            .I(N__38301));
    InMux I__4567 (
            .O(N__38304),
            .I(N__38298));
    Odrv4 I__4566 (
            .O(N__38301),
            .I(REG_mem_4_10));
    LocalMux I__4565 (
            .O(N__38298),
            .I(REG_mem_4_10));
    InMux I__4564 (
            .O(N__38293),
            .I(N__38290));
    LocalMux I__4563 (
            .O(N__38290),
            .I(N__38286));
    InMux I__4562 (
            .O(N__38289),
            .I(N__38283));
    Span4Mux_v I__4561 (
            .O(N__38286),
            .I(N__38280));
    LocalMux I__4560 (
            .O(N__38283),
            .I(N__38277));
    Odrv4 I__4559 (
            .O(N__38280),
            .I(REG_mem_4_14));
    Odrv4 I__4558 (
            .O(N__38277),
            .I(REG_mem_4_14));
    InMux I__4557 (
            .O(N__38272),
            .I(N__38268));
    InMux I__4556 (
            .O(N__38271),
            .I(N__38265));
    LocalMux I__4555 (
            .O(N__38268),
            .I(REG_mem_48_3));
    LocalMux I__4554 (
            .O(N__38265),
            .I(REG_mem_48_3));
    InMux I__4553 (
            .O(N__38260),
            .I(N__38257));
    LocalMux I__4552 (
            .O(N__38257),
            .I(N__38253));
    InMux I__4551 (
            .O(N__38256),
            .I(N__38250));
    Odrv12 I__4550 (
            .O(N__38253),
            .I(REG_mem_45_14));
    LocalMux I__4549 (
            .O(N__38250),
            .I(REG_mem_45_14));
    InMux I__4548 (
            .O(N__38245),
            .I(N__38241));
    InMux I__4547 (
            .O(N__38244),
            .I(N__38238));
    LocalMux I__4546 (
            .O(N__38241),
            .I(REG_mem_50_10));
    LocalMux I__4545 (
            .O(N__38238),
            .I(REG_mem_50_10));
    InMux I__4544 (
            .O(N__38233),
            .I(N__38230));
    LocalMux I__4543 (
            .O(N__38230),
            .I(N__38227));
    Span4Mux_v I__4542 (
            .O(N__38227),
            .I(N__38224));
    Span4Mux_v I__4541 (
            .O(N__38224),
            .I(N__38220));
    InMux I__4540 (
            .O(N__38223),
            .I(N__38217));
    Odrv4 I__4539 (
            .O(N__38220),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_9 ));
    LocalMux I__4538 (
            .O(N__38217),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_9 ));
    InMux I__4537 (
            .O(N__38212),
            .I(N__38208));
    CascadeMux I__4536 (
            .O(N__38211),
            .I(N__38205));
    LocalMux I__4535 (
            .O(N__38208),
            .I(N__38202));
    InMux I__4534 (
            .O(N__38205),
            .I(N__38199));
    Odrv4 I__4533 (
            .O(N__38202),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_3 ));
    LocalMux I__4532 (
            .O(N__38199),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_3 ));
    InMux I__4531 (
            .O(N__38194),
            .I(N__38191));
    LocalMux I__4530 (
            .O(N__38191),
            .I(N__38188));
    Span4Mux_v I__4529 (
            .O(N__38188),
            .I(N__38184));
    CascadeMux I__4528 (
            .O(N__38187),
            .I(N__38181));
    Span4Mux_v I__4527 (
            .O(N__38184),
            .I(N__38178));
    InMux I__4526 (
            .O(N__38181),
            .I(N__38175));
    Odrv4 I__4525 (
            .O(N__38178),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_12 ));
    LocalMux I__4524 (
            .O(N__38175),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_12 ));
    InMux I__4523 (
            .O(N__38170),
            .I(N__38166));
    InMux I__4522 (
            .O(N__38169),
            .I(N__38163));
    LocalMux I__4521 (
            .O(N__38166),
            .I(N__38160));
    LocalMux I__4520 (
            .O(N__38163),
            .I(REG_mem_16_14));
    Odrv4 I__4519 (
            .O(N__38160),
            .I(REG_mem_16_14));
    CascadeMux I__4518 (
            .O(N__38155),
            .I(N__38152));
    InMux I__4517 (
            .O(N__38152),
            .I(N__38146));
    InMux I__4516 (
            .O(N__38151),
            .I(N__38146));
    LocalMux I__4515 (
            .O(N__38146),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_12 ));
    InMux I__4514 (
            .O(N__38143),
            .I(N__38140));
    LocalMux I__4513 (
            .O(N__38140),
            .I(N__38137));
    Span4Mux_h I__4512 (
            .O(N__38137),
            .I(N__38134));
    Span4Mux_v I__4511 (
            .O(N__38134),
            .I(N__38130));
    InMux I__4510 (
            .O(N__38133),
            .I(N__38127));
    Odrv4 I__4509 (
            .O(N__38130),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_9 ));
    LocalMux I__4508 (
            .O(N__38127),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_9 ));
    InMux I__4507 (
            .O(N__38122),
            .I(N__38116));
    InMux I__4506 (
            .O(N__38121),
            .I(N__38116));
    LocalMux I__4505 (
            .O(N__38116),
            .I(REG_mem_31_7));
    CascadeMux I__4504 (
            .O(N__38113),
            .I(N__38110));
    InMux I__4503 (
            .O(N__38110),
            .I(N__38106));
    InMux I__4502 (
            .O(N__38109),
            .I(N__38103));
    LocalMux I__4501 (
            .O(N__38106),
            .I(REG_mem_26_7));
    LocalMux I__4500 (
            .O(N__38103),
            .I(REG_mem_26_7));
    InMux I__4499 (
            .O(N__38098),
            .I(N__38094));
    InMux I__4498 (
            .O(N__38097),
            .I(N__38091));
    LocalMux I__4497 (
            .O(N__38094),
            .I(REG_mem_14_15));
    LocalMux I__4496 (
            .O(N__38091),
            .I(REG_mem_14_15));
    InMux I__4495 (
            .O(N__38086),
            .I(N__38082));
    CascadeMux I__4494 (
            .O(N__38085),
            .I(N__38079));
    LocalMux I__4493 (
            .O(N__38082),
            .I(N__38076));
    InMux I__4492 (
            .O(N__38079),
            .I(N__38073));
    Odrv12 I__4491 (
            .O(N__38076),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_7 ));
    LocalMux I__4490 (
            .O(N__38073),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_7 ));
    InMux I__4489 (
            .O(N__38068),
            .I(N__38065));
    LocalMux I__4488 (
            .O(N__38065),
            .I(N__38062));
    Span4Mux_h I__4487 (
            .O(N__38062),
            .I(N__38058));
    InMux I__4486 (
            .O(N__38061),
            .I(N__38055));
    Odrv4 I__4485 (
            .O(N__38058),
            .I(REG_mem_40_14));
    LocalMux I__4484 (
            .O(N__38055),
            .I(REG_mem_40_14));
    CascadeMux I__4483 (
            .O(N__38050),
            .I(N__38047));
    InMux I__4482 (
            .O(N__38047),
            .I(N__38043));
    InMux I__4481 (
            .O(N__38046),
            .I(N__38040));
    LocalMux I__4480 (
            .O(N__38043),
            .I(N__38037));
    LocalMux I__4479 (
            .O(N__38040),
            .I(N__38034));
    Odrv4 I__4478 (
            .O(N__38037),
            .I(REG_mem_8_15));
    Odrv4 I__4477 (
            .O(N__38034),
            .I(REG_mem_8_15));
    CascadeMux I__4476 (
            .O(N__38029),
            .I(N__38026));
    InMux I__4475 (
            .O(N__38026),
            .I(N__38023));
    LocalMux I__4474 (
            .O(N__38023),
            .I(N__38020));
    Span4Mux_h I__4473 (
            .O(N__38020),
            .I(N__38016));
    CascadeMux I__4472 (
            .O(N__38019),
            .I(N__38013));
    Span4Mux_v I__4471 (
            .O(N__38016),
            .I(N__38010));
    InMux I__4470 (
            .O(N__38013),
            .I(N__38007));
    Odrv4 I__4469 (
            .O(N__38010),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_13 ));
    LocalMux I__4468 (
            .O(N__38007),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_13 ));
    CascadeMux I__4467 (
            .O(N__38002),
            .I(N__37998));
    InMux I__4466 (
            .O(N__38001),
            .I(N__37995));
    InMux I__4465 (
            .O(N__37998),
            .I(N__37992));
    LocalMux I__4464 (
            .O(N__37995),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_7 ));
    LocalMux I__4463 (
            .O(N__37992),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_7 ));
    InMux I__4462 (
            .O(N__37987),
            .I(N__37984));
    LocalMux I__4461 (
            .O(N__37984),
            .I(N__37980));
    CascadeMux I__4460 (
            .O(N__37983),
            .I(N__37977));
    Span4Mux_v I__4459 (
            .O(N__37980),
            .I(N__37974));
    InMux I__4458 (
            .O(N__37977),
            .I(N__37971));
    Odrv4 I__4457 (
            .O(N__37974),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_0 ));
    LocalMux I__4456 (
            .O(N__37971),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_0 ));
    InMux I__4455 (
            .O(N__37966),
            .I(N__37963));
    LocalMux I__4454 (
            .O(N__37963),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12812 ));
    InMux I__4453 (
            .O(N__37960),
            .I(N__37954));
    InMux I__4452 (
            .O(N__37959),
            .I(N__37954));
    LocalMux I__4451 (
            .O(N__37954),
            .I(N__37951));
    Odrv4 I__4450 (
            .O(N__37951),
            .I(REG_mem_13_15));
    InMux I__4449 (
            .O(N__37948),
            .I(N__37942));
    InMux I__4448 (
            .O(N__37947),
            .I(N__37942));
    LocalMux I__4447 (
            .O(N__37942),
            .I(N__37939));
    Odrv4 I__4446 (
            .O(N__37939),
            .I(REG_mem_44_0));
    InMux I__4445 (
            .O(N__37936),
            .I(N__37933));
    LocalMux I__4444 (
            .O(N__37933),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12830 ));
    CascadeMux I__4443 (
            .O(N__37930),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13916_cascade_ ));
    CascadeMux I__4442 (
            .O(N__37927),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12168_cascade_ ));
    InMux I__4441 (
            .O(N__37924),
            .I(N__37921));
    LocalMux I__4440 (
            .O(N__37921),
            .I(N__37917));
    CascadeMux I__4439 (
            .O(N__37920),
            .I(N__37914));
    Span4Mux_v I__4438 (
            .O(N__37917),
            .I(N__37911));
    InMux I__4437 (
            .O(N__37914),
            .I(N__37908));
    Odrv4 I__4436 (
            .O(N__37911),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_7 ));
    LocalMux I__4435 (
            .O(N__37908),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_7 ));
    CascadeMux I__4434 (
            .O(N__37903),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13922_cascade_ ));
    InMux I__4433 (
            .O(N__37900),
            .I(N__37897));
    LocalMux I__4432 (
            .O(N__37897),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12165 ));
    CascadeMux I__4431 (
            .O(N__37894),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13235_cascade_ ));
    InMux I__4430 (
            .O(N__37891),
            .I(N__37887));
    InMux I__4429 (
            .O(N__37890),
            .I(N__37884));
    LocalMux I__4428 (
            .O(N__37887),
            .I(REG_mem_47_0));
    LocalMux I__4427 (
            .O(N__37884),
            .I(REG_mem_47_0));
    InMux I__4426 (
            .O(N__37879),
            .I(N__37876));
    LocalMux I__4425 (
            .O(N__37876),
            .I(N__37873));
    Span4Mux_v I__4424 (
            .O(N__37873),
            .I(N__37869));
    InMux I__4423 (
            .O(N__37872),
            .I(N__37866));
    Odrv4 I__4422 (
            .O(N__37869),
            .I(REG_mem_4_9));
    LocalMux I__4421 (
            .O(N__37866),
            .I(REG_mem_4_9));
    InMux I__4420 (
            .O(N__37861),
            .I(N__37858));
    LocalMux I__4419 (
            .O(N__37858),
            .I(N__37855));
    Odrv4 I__4418 (
            .O(N__37855),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12343 ));
    CascadeMux I__4417 (
            .O(N__37852),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12923_cascade_ ));
    InMux I__4416 (
            .O(N__37849),
            .I(N__37846));
    LocalMux I__4415 (
            .O(N__37846),
            .I(N__37843));
    Span4Mux_h I__4414 (
            .O(N__37843),
            .I(N__37840));
    Odrv4 I__4413 (
            .O(N__37840),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12059 ));
    CascadeMux I__4412 (
            .O(N__37837),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12896_cascade_ ));
    InMux I__4411 (
            .O(N__37834),
            .I(N__37831));
    LocalMux I__4410 (
            .O(N__37831),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12899 ));
    InMux I__4409 (
            .O(N__37828),
            .I(N__37824));
    InMux I__4408 (
            .O(N__37827),
            .I(N__37821));
    LocalMux I__4407 (
            .O(N__37824),
            .I(REG_mem_42_15));
    LocalMux I__4406 (
            .O(N__37821),
            .I(REG_mem_42_15));
    InMux I__4405 (
            .O(N__37816),
            .I(N__37812));
    InMux I__4404 (
            .O(N__37815),
            .I(N__37809));
    LocalMux I__4403 (
            .O(N__37812),
            .I(REG_mem_43_15));
    LocalMux I__4402 (
            .O(N__37809),
            .I(REG_mem_43_15));
    CascadeMux I__4401 (
            .O(N__37804),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13400_cascade_ ));
    CascadeMux I__4400 (
            .O(N__37801),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13403_cascade_ ));
    CascadeMux I__4399 (
            .O(N__37798),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12068_cascade_ ));
    CascadeMux I__4398 (
            .O(N__37795),
            .I(N__37792));
    InMux I__4397 (
            .O(N__37792),
            .I(N__37789));
    LocalMux I__4396 (
            .O(N__37789),
            .I(N__37786));
    Span4Mux_h I__4395 (
            .O(N__37786),
            .I(N__37783));
    Span4Mux_v I__4394 (
            .O(N__37783),
            .I(N__37780));
    Odrv4 I__4393 (
            .O(N__37780),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12017 ));
    InMux I__4392 (
            .O(N__37777),
            .I(N__37774));
    LocalMux I__4391 (
            .O(N__37774),
            .I(N__37771));
    Span4Mux_v I__4390 (
            .O(N__37771),
            .I(N__37768));
    Odrv4 I__4389 (
            .O(N__37768),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12016 ));
    InMux I__4388 (
            .O(N__37765),
            .I(N__37762));
    LocalMux I__4387 (
            .O(N__37762),
            .I(N__37759));
    Span4Mux_v I__4386 (
            .O(N__37759),
            .I(N__37756));
    Odrv4 I__4385 (
            .O(N__37756),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12935 ));
    InMux I__4384 (
            .O(N__37753),
            .I(N__37750));
    LocalMux I__4383 (
            .O(N__37750),
            .I(N__37747));
    Span4Mux_v I__4382 (
            .O(N__37747),
            .I(N__37744));
    Odrv4 I__4381 (
            .O(N__37744),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12983 ));
    InMux I__4380 (
            .O(N__37741),
            .I(N__37738));
    LocalMux I__4379 (
            .O(N__37738),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13031 ));
    CascadeMux I__4378 (
            .O(N__37735),
            .I(N__37732));
    InMux I__4377 (
            .O(N__37732),
            .I(N__37726));
    InMux I__4376 (
            .O(N__37731),
            .I(N__37726));
    LocalMux I__4375 (
            .O(N__37726),
            .I(REG_mem_37_9));
    InMux I__4374 (
            .O(N__37723),
            .I(N__37720));
    LocalMux I__4373 (
            .O(N__37720),
            .I(N__37717));
    Span4Mux_v I__4372 (
            .O(N__37717),
            .I(N__37714));
    Odrv4 I__4371 (
            .O(N__37714),
            .I(FIFO_D9_c_9));
    InMux I__4370 (
            .O(N__37711),
            .I(N__37708));
    LocalMux I__4369 (
            .O(N__37708),
            .I(\usb3_if_inst.usb3_data_in_latched_9 ));
    CascadeMux I__4368 (
            .O(N__37705),
            .I(N__37702));
    InMux I__4367 (
            .O(N__37702),
            .I(N__37696));
    InMux I__4366 (
            .O(N__37701),
            .I(N__37696));
    LocalMux I__4365 (
            .O(N__37696),
            .I(REG_mem_63_15));
    InMux I__4364 (
            .O(N__37693),
            .I(N__37690));
    LocalMux I__4363 (
            .O(N__37690),
            .I(N__37687));
    Span12Mux_s10_h I__4362 (
            .O(N__37687),
            .I(N__37684));
    Odrv12 I__4361 (
            .O(N__37684),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12044 ));
    CascadeMux I__4360 (
            .O(N__37681),
            .I(N__37677));
    InMux I__4359 (
            .O(N__37680),
            .I(N__37672));
    InMux I__4358 (
            .O(N__37677),
            .I(N__37672));
    LocalMux I__4357 (
            .O(N__37672),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_15 ));
    CascadeMux I__4356 (
            .O(N__37669),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12860_cascade_ ));
    CascadeMux I__4355 (
            .O(N__37666),
            .I(N__37662));
    InMux I__4354 (
            .O(N__37665),
            .I(N__37659));
    InMux I__4353 (
            .O(N__37662),
            .I(N__37656));
    LocalMux I__4352 (
            .O(N__37659),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_0 ));
    LocalMux I__4351 (
            .O(N__37656),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_0 ));
    CascadeMux I__4350 (
            .O(N__37651),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13142_cascade_ ));
    InMux I__4349 (
            .O(N__37648),
            .I(N__37645));
    LocalMux I__4348 (
            .O(N__37645),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13145 ));
    InMux I__4347 (
            .O(N__37642),
            .I(N__37638));
    InMux I__4346 (
            .O(N__37641),
            .I(N__37635));
    LocalMux I__4345 (
            .O(N__37638),
            .I(REG_mem_42_10));
    LocalMux I__4344 (
            .O(N__37635),
            .I(REG_mem_42_10));
    InMux I__4343 (
            .O(N__37630),
            .I(N__37627));
    LocalMux I__4342 (
            .O(N__37627),
            .I(N__37623));
    InMux I__4341 (
            .O(N__37626),
            .I(N__37620));
    Odrv4 I__4340 (
            .O(N__37623),
            .I(REG_mem_43_10));
    LocalMux I__4339 (
            .O(N__37620),
            .I(REG_mem_43_10));
    InMux I__4338 (
            .O(N__37615),
            .I(N__37612));
    LocalMux I__4337 (
            .O(N__37612),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13394 ));
    InMux I__4336 (
            .O(N__37609),
            .I(N__37603));
    InMux I__4335 (
            .O(N__37608),
            .I(N__37603));
    LocalMux I__4334 (
            .O(N__37603),
            .I(REG_mem_45_10));
    InMux I__4333 (
            .O(N__37600),
            .I(N__37594));
    InMux I__4332 (
            .O(N__37599),
            .I(N__37594));
    LocalMux I__4331 (
            .O(N__37594),
            .I(REG_mem_44_10));
    InMux I__4330 (
            .O(N__37591),
            .I(N__37585));
    InMux I__4329 (
            .O(N__37590),
            .I(N__37585));
    LocalMux I__4328 (
            .O(N__37585),
            .I(REG_mem_46_10));
    CascadeMux I__4327 (
            .O(N__37582),
            .I(N__37579));
    InMux I__4326 (
            .O(N__37579),
            .I(N__37576));
    LocalMux I__4325 (
            .O(N__37576),
            .I(N__37572));
    InMux I__4324 (
            .O(N__37575),
            .I(N__37569));
    Odrv12 I__4323 (
            .O(N__37572),
            .I(REG_mem_10_13));
    LocalMux I__4322 (
            .O(N__37569),
            .I(REG_mem_10_13));
    InMux I__4321 (
            .O(N__37564),
            .I(N__37561));
    LocalMux I__4320 (
            .O(N__37561),
            .I(N__37558));
    Glb2LocalMux I__4319 (
            .O(N__37558),
            .I(N__37555));
    GlobalMux I__4318 (
            .O(N__37555),
            .I(pll_clk_unbuf));
    IoInMux I__4317 (
            .O(N__37552),
            .I(N__37549));
    LocalMux I__4316 (
            .O(N__37549),
            .I(N__37546));
    Span4Mux_s3_h I__4315 (
            .O(N__37546),
            .I(N__37543));
    Span4Mux_v I__4314 (
            .O(N__37543),
            .I(N__37540));
    Span4Mux_v I__4313 (
            .O(N__37540),
            .I(N__37537));
    Span4Mux_h I__4312 (
            .O(N__37537),
            .I(N__37534));
    Odrv4 I__4311 (
            .O(N__37534),
            .I(GB_BUFFER_pll_clk_unbuf_THRU_CO));
    InMux I__4310 (
            .O(N__37531),
            .I(N__37528));
    LocalMux I__4309 (
            .O(N__37528),
            .I(N__37525));
    Span4Mux_v I__4308 (
            .O(N__37525),
            .I(N__37521));
    InMux I__4307 (
            .O(N__37524),
            .I(N__37518));
    Odrv4 I__4306 (
            .O(N__37521),
            .I(REG_mem_43_7));
    LocalMux I__4305 (
            .O(N__37518),
            .I(REG_mem_43_7));
    InMux I__4304 (
            .O(N__37513),
            .I(N__37509));
    InMux I__4303 (
            .O(N__37512),
            .I(N__37506));
    LocalMux I__4302 (
            .O(N__37509),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_12 ));
    LocalMux I__4301 (
            .O(N__37506),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_12 ));
    InMux I__4300 (
            .O(N__37501),
            .I(N__37497));
    InMux I__4299 (
            .O(N__37500),
            .I(N__37494));
    LocalMux I__4298 (
            .O(N__37497),
            .I(REG_mem_41_10));
    LocalMux I__4297 (
            .O(N__37494),
            .I(REG_mem_41_10));
    CascadeMux I__4296 (
            .O(N__37489),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13397_cascade_ ));
    InMux I__4295 (
            .O(N__37486),
            .I(N__37483));
    LocalMux I__4294 (
            .O(N__37483),
            .I(N__37480));
    Span4Mux_v I__4293 (
            .O(N__37480),
            .I(N__37477));
    Span4Mux_h I__4292 (
            .O(N__37477),
            .I(N__37474));
    Odrv4 I__4291 (
            .O(N__37474),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11630 ));
    InMux I__4290 (
            .O(N__37471),
            .I(N__37468));
    LocalMux I__4289 (
            .O(N__37468),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12487 ));
    InMux I__4288 (
            .O(N__37465),
            .I(N__37461));
    InMux I__4287 (
            .O(N__37464),
            .I(N__37458));
    LocalMux I__4286 (
            .O(N__37461),
            .I(REG_mem_42_12));
    LocalMux I__4285 (
            .O(N__37458),
            .I(REG_mem_42_12));
    InMux I__4284 (
            .O(N__37453),
            .I(N__37450));
    LocalMux I__4283 (
            .O(N__37450),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12488 ));
    InMux I__4282 (
            .O(N__37447),
            .I(N__37441));
    InMux I__4281 (
            .O(N__37446),
            .I(N__37441));
    LocalMux I__4280 (
            .O(N__37441),
            .I(REG_mem_43_12));
    CascadeMux I__4279 (
            .O(N__37438),
            .I(N__37435));
    InMux I__4278 (
            .O(N__37435),
            .I(N__37432));
    LocalMux I__4277 (
            .O(N__37432),
            .I(N__37428));
    InMux I__4276 (
            .O(N__37431),
            .I(N__37425));
    Odrv4 I__4275 (
            .O(N__37428),
            .I(REG_mem_31_12));
    LocalMux I__4274 (
            .O(N__37425),
            .I(REG_mem_31_12));
    CascadeMux I__4273 (
            .O(N__37420),
            .I(N__37417));
    InMux I__4272 (
            .O(N__37417),
            .I(N__37414));
    LocalMux I__4271 (
            .O(N__37414),
            .I(N__37410));
    InMux I__4270 (
            .O(N__37413),
            .I(N__37407));
    Odrv4 I__4269 (
            .O(N__37410),
            .I(REG_mem_44_12));
    LocalMux I__4268 (
            .O(N__37407),
            .I(REG_mem_44_12));
    InMux I__4267 (
            .O(N__37402),
            .I(N__37399));
    LocalMux I__4266 (
            .O(N__37399),
            .I(N__37396));
    Odrv4 I__4265 (
            .O(N__37396),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12493 ));
    InMux I__4264 (
            .O(N__37393),
            .I(N__37387));
    InMux I__4263 (
            .O(N__37392),
            .I(N__37387));
    LocalMux I__4262 (
            .O(N__37387),
            .I(REG_mem_45_12));
    InMux I__4261 (
            .O(N__37384),
            .I(N__37381));
    LocalMux I__4260 (
            .O(N__37381),
            .I(N__37378));
    Span4Mux_v I__4259 (
            .O(N__37378),
            .I(N__37375));
    Span4Mux_v I__4258 (
            .O(N__37375),
            .I(N__37371));
    InMux I__4257 (
            .O(N__37374),
            .I(N__37368));
    Odrv4 I__4256 (
            .O(N__37371),
            .I(REG_mem_9_10));
    LocalMux I__4255 (
            .O(N__37368),
            .I(REG_mem_9_10));
    InMux I__4254 (
            .O(N__37363),
            .I(N__37359));
    InMux I__4253 (
            .O(N__37362),
            .I(N__37356));
    LocalMux I__4252 (
            .O(N__37359),
            .I(REG_mem_42_11));
    LocalMux I__4251 (
            .O(N__37356),
            .I(REG_mem_42_11));
    CascadeMux I__4250 (
            .O(N__37351),
            .I(N__37347));
    InMux I__4249 (
            .O(N__37350),
            .I(N__37344));
    InMux I__4248 (
            .O(N__37347),
            .I(N__37341));
    LocalMux I__4247 (
            .O(N__37344),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_12 ));
    LocalMux I__4246 (
            .O(N__37341),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_12 ));
    InMux I__4245 (
            .O(N__37336),
            .I(N__37333));
    LocalMux I__4244 (
            .O(N__37333),
            .I(N__37329));
    InMux I__4243 (
            .O(N__37332),
            .I(N__37326));
    Odrv12 I__4242 (
            .O(N__37329),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_12 ));
    LocalMux I__4241 (
            .O(N__37326),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_12 ));
    CascadeMux I__4240 (
            .O(N__37321),
            .I(N__37317));
    InMux I__4239 (
            .O(N__37320),
            .I(N__37314));
    InMux I__4238 (
            .O(N__37317),
            .I(N__37311));
    LocalMux I__4237 (
            .O(N__37314),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_12 ));
    LocalMux I__4236 (
            .O(N__37311),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_12 ));
    CascadeMux I__4235 (
            .O(N__37306),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12494_cascade_ ));
    CascadeMux I__4234 (
            .O(N__37303),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14252_cascade_ ));
    CascadeMux I__4233 (
            .O(N__37300),
            .I(N__37297));
    InMux I__4232 (
            .O(N__37297),
            .I(N__37294));
    LocalMux I__4231 (
            .O(N__37294),
            .I(N__37291));
    Odrv12 I__4230 (
            .O(N__37291),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12481 ));
    InMux I__4229 (
            .O(N__37288),
            .I(N__37285));
    LocalMux I__4228 (
            .O(N__37285),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12476 ));
    CascadeMux I__4227 (
            .O(N__37282),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13292_cascade_ ));
    InMux I__4226 (
            .O(N__37279),
            .I(N__37276));
    LocalMux I__4225 (
            .O(N__37276),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12475 ));
    CascadeMux I__4224 (
            .O(N__37273),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13295_cascade_ ));
    InMux I__4223 (
            .O(N__37270),
            .I(N__37267));
    LocalMux I__4222 (
            .O(N__37267),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14255 ));
    InMux I__4221 (
            .O(N__37264),
            .I(N__37261));
    LocalMux I__4220 (
            .O(N__37261),
            .I(N__37258));
    Span4Mux_v I__4219 (
            .O(N__37258),
            .I(N__37255));
    Odrv4 I__4218 (
            .O(N__37255),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11643 ));
    InMux I__4217 (
            .O(N__37252),
            .I(N__37246));
    InMux I__4216 (
            .O(N__37251),
            .I(N__37246));
    LocalMux I__4215 (
            .O(N__37246),
            .I(REG_mem_11_3));
    CascadeMux I__4214 (
            .O(N__37243),
            .I(N__37240));
    InMux I__4213 (
            .O(N__37240),
            .I(N__37237));
    LocalMux I__4212 (
            .O(N__37237),
            .I(N__37233));
    InMux I__4211 (
            .O(N__37236),
            .I(N__37230));
    Odrv12 I__4210 (
            .O(N__37233),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_11 ));
    LocalMux I__4209 (
            .O(N__37230),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_11 ));
    InMux I__4208 (
            .O(N__37225),
            .I(N__37222));
    LocalMux I__4207 (
            .O(N__37222),
            .I(N__37219));
    Span4Mux_v I__4206 (
            .O(N__37219),
            .I(N__37215));
    InMux I__4205 (
            .O(N__37218),
            .I(N__37212));
    Odrv4 I__4204 (
            .O(N__37215),
            .I(REG_mem_10_14));
    LocalMux I__4203 (
            .O(N__37212),
            .I(REG_mem_10_14));
    CascadeMux I__4202 (
            .O(N__37207),
            .I(N__37203));
    InMux I__4201 (
            .O(N__37206),
            .I(N__37200));
    InMux I__4200 (
            .O(N__37203),
            .I(N__37197));
    LocalMux I__4199 (
            .O(N__37200),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_12 ));
    LocalMux I__4198 (
            .O(N__37197),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_12 ));
    InMux I__4197 (
            .O(N__37192),
            .I(N__37188));
    InMux I__4196 (
            .O(N__37191),
            .I(N__37185));
    LocalMux I__4195 (
            .O(N__37188),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_12 ));
    LocalMux I__4194 (
            .O(N__37185),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_12 ));
    InMux I__4193 (
            .O(N__37180),
            .I(N__37174));
    InMux I__4192 (
            .O(N__37179),
            .I(N__37174));
    LocalMux I__4191 (
            .O(N__37174),
            .I(REG_mem_42_7));
    InMux I__4190 (
            .O(N__37171),
            .I(N__37168));
    LocalMux I__4189 (
            .O(N__37168),
            .I(N__37164));
    InMux I__4188 (
            .O(N__37167),
            .I(N__37161));
    Odrv4 I__4187 (
            .O(N__37164),
            .I(REG_mem_44_9));
    LocalMux I__4186 (
            .O(N__37161),
            .I(REG_mem_44_9));
    CascadeMux I__4185 (
            .O(N__37156),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12800_cascade_ ));
    InMux I__4184 (
            .O(N__37153),
            .I(N__37150));
    LocalMux I__4183 (
            .O(N__37150),
            .I(N__37147));
    Span4Mux_h I__4182 (
            .O(N__37147),
            .I(N__37143));
    InMux I__4181 (
            .O(N__37146),
            .I(N__37140));
    Odrv4 I__4180 (
            .O(N__37143),
            .I(REG_mem_45_9));
    LocalMux I__4179 (
            .O(N__37140),
            .I(REG_mem_45_9));
    InMux I__4178 (
            .O(N__37135),
            .I(N__37132));
    LocalMux I__4177 (
            .O(N__37132),
            .I(N__37129));
    Span4Mux_v I__4176 (
            .O(N__37129),
            .I(N__37126));
    Odrv4 I__4175 (
            .O(N__37126),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12803 ));
    InMux I__4174 (
            .O(N__37123),
            .I(N__37120));
    LocalMux I__4173 (
            .O(N__37120),
            .I(N__37117));
    Span4Mux_v I__4172 (
            .O(N__37117),
            .I(N__37114));
    Span4Mux_v I__4171 (
            .O(N__37114),
            .I(N__37110));
    InMux I__4170 (
            .O(N__37113),
            .I(N__37107));
    Odrv4 I__4169 (
            .O(N__37110),
            .I(REG_mem_58_15));
    LocalMux I__4168 (
            .O(N__37107),
            .I(REG_mem_58_15));
    InMux I__4167 (
            .O(N__37102),
            .I(N__37098));
    InMux I__4166 (
            .O(N__37101),
            .I(N__37095));
    LocalMux I__4165 (
            .O(N__37098),
            .I(REG_mem_12_3));
    LocalMux I__4164 (
            .O(N__37095),
            .I(REG_mem_12_3));
    InMux I__4163 (
            .O(N__37090),
            .I(N__37087));
    LocalMux I__4162 (
            .O(N__37087),
            .I(N__37084));
    Span4Mux_v I__4161 (
            .O(N__37084),
            .I(N__37081));
    Odrv4 I__4160 (
            .O(N__37081),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11625 ));
    CascadeMux I__4159 (
            .O(N__37078),
            .I(N__37075));
    InMux I__4158 (
            .O(N__37075),
            .I(N__37071));
    InMux I__4157 (
            .O(N__37074),
            .I(N__37068));
    LocalMux I__4156 (
            .O(N__37071),
            .I(REG_mem_43_11));
    LocalMux I__4155 (
            .O(N__37068),
            .I(REG_mem_43_11));
    CascadeMux I__4154 (
            .O(N__37063),
            .I(N__37060));
    InMux I__4153 (
            .O(N__37060),
            .I(N__37057));
    LocalMux I__4152 (
            .O(N__37057),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13457 ));
    InMux I__4151 (
            .O(N__37054),
            .I(N__37051));
    LocalMux I__4150 (
            .O(N__37051),
            .I(N__37048));
    Span4Mux_v I__4149 (
            .O(N__37048),
            .I(N__37045));
    Odrv4 I__4148 (
            .O(N__37045),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11990 ));
    CascadeMux I__4147 (
            .O(N__37042),
            .I(N__37039));
    InMux I__4146 (
            .O(N__37039),
            .I(N__37033));
    InMux I__4145 (
            .O(N__37038),
            .I(N__37033));
    LocalMux I__4144 (
            .O(N__37033),
            .I(REG_mem_10_3));
    InMux I__4143 (
            .O(N__37030),
            .I(N__37024));
    InMux I__4142 (
            .O(N__37029),
            .I(N__37024));
    LocalMux I__4141 (
            .O(N__37024),
            .I(REG_mem_51_3));
    InMux I__4140 (
            .O(N__37021),
            .I(N__37017));
    InMux I__4139 (
            .O(N__37020),
            .I(N__37014));
    LocalMux I__4138 (
            .O(N__37017),
            .I(REG_mem_51_10));
    LocalMux I__4137 (
            .O(N__37014),
            .I(REG_mem_51_10));
    CascadeMux I__4136 (
            .O(N__37009),
            .I(N__37005));
    InMux I__4135 (
            .O(N__37008),
            .I(N__37002));
    InMux I__4134 (
            .O(N__37005),
            .I(N__36999));
    LocalMux I__4133 (
            .O(N__37002),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_3 ));
    LocalMux I__4132 (
            .O(N__36999),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_3 ));
    InMux I__4131 (
            .O(N__36994),
            .I(N__36991));
    LocalMux I__4130 (
            .O(N__36991),
            .I(N__36987));
    InMux I__4129 (
            .O(N__36990),
            .I(N__36984));
    Odrv12 I__4128 (
            .O(N__36987),
            .I(REG_mem_63_0));
    LocalMux I__4127 (
            .O(N__36984),
            .I(REG_mem_63_0));
    CascadeMux I__4126 (
            .O(N__36979),
            .I(N__36976));
    InMux I__4125 (
            .O(N__36976),
            .I(N__36973));
    LocalMux I__4124 (
            .O(N__36973),
            .I(N__36969));
    InMux I__4123 (
            .O(N__36972),
            .I(N__36966));
    Odrv4 I__4122 (
            .O(N__36969),
            .I(REG_mem_6_3));
    LocalMux I__4121 (
            .O(N__36966),
            .I(REG_mem_6_3));
    CascadeMux I__4120 (
            .O(N__36961),
            .I(N__36958));
    InMux I__4119 (
            .O(N__36958),
            .I(N__36955));
    LocalMux I__4118 (
            .O(N__36955),
            .I(N__36951));
    InMux I__4117 (
            .O(N__36954),
            .I(N__36948));
    Odrv12 I__4116 (
            .O(N__36951),
            .I(REG_mem_43_3));
    LocalMux I__4115 (
            .O(N__36948),
            .I(REG_mem_43_3));
    InMux I__4114 (
            .O(N__36943),
            .I(N__36937));
    InMux I__4113 (
            .O(N__36942),
            .I(N__36937));
    LocalMux I__4112 (
            .O(N__36937),
            .I(REG_mem_41_3));
    CascadeMux I__4111 (
            .O(N__36934),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13454_cascade_ ));
    InMux I__4110 (
            .O(N__36931),
            .I(N__36925));
    InMux I__4109 (
            .O(N__36930),
            .I(N__36925));
    LocalMux I__4108 (
            .O(N__36925),
            .I(REG_mem_42_3));
    CascadeMux I__4107 (
            .O(N__36922),
            .I(N__36919));
    InMux I__4106 (
            .O(N__36919),
            .I(N__36913));
    InMux I__4105 (
            .O(N__36918),
            .I(N__36913));
    LocalMux I__4104 (
            .O(N__36913),
            .I(REG_mem_11_14));
    InMux I__4103 (
            .O(N__36910),
            .I(N__36907));
    LocalMux I__4102 (
            .O(N__36907),
            .I(N__36903));
    InMux I__4101 (
            .O(N__36906),
            .I(N__36900));
    Odrv4 I__4100 (
            .O(N__36903),
            .I(REG_mem_5_14));
    LocalMux I__4099 (
            .O(N__36900),
            .I(REG_mem_5_14));
    InMux I__4098 (
            .O(N__36895),
            .I(N__36892));
    LocalMux I__4097 (
            .O(N__36892),
            .I(N__36888));
    InMux I__4096 (
            .O(N__36891),
            .I(N__36885));
    Odrv4 I__4095 (
            .O(N__36888),
            .I(REG_mem_6_14));
    LocalMux I__4094 (
            .O(N__36885),
            .I(REG_mem_6_14));
    InMux I__4093 (
            .O(N__36880),
            .I(N__36877));
    LocalMux I__4092 (
            .O(N__36877),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13022 ));
    InMux I__4091 (
            .O(N__36874),
            .I(N__36868));
    InMux I__4090 (
            .O(N__36873),
            .I(N__36868));
    LocalMux I__4089 (
            .O(N__36868),
            .I(REG_mem_49_3));
    CascadeMux I__4088 (
            .O(N__36865),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13244_cascade_ ));
    InMux I__4087 (
            .O(N__36862),
            .I(N__36859));
    LocalMux I__4086 (
            .O(N__36859),
            .I(N__36856));
    Span4Mux_v I__4085 (
            .O(N__36856),
            .I(N__36853));
    Odrv4 I__4084 (
            .O(N__36853),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13247 ));
    InMux I__4083 (
            .O(N__36850),
            .I(N__36846));
    InMux I__4082 (
            .O(N__36849),
            .I(N__36843));
    LocalMux I__4081 (
            .O(N__36846),
            .I(REG_mem_18_3));
    LocalMux I__4080 (
            .O(N__36843),
            .I(REG_mem_18_3));
    InMux I__4079 (
            .O(N__36838),
            .I(N__36834));
    InMux I__4078 (
            .O(N__36837),
            .I(N__36831));
    LocalMux I__4077 (
            .O(N__36834),
            .I(REG_mem_17_14));
    LocalMux I__4076 (
            .O(N__36831),
            .I(REG_mem_17_14));
    InMux I__4075 (
            .O(N__36826),
            .I(N__36823));
    LocalMux I__4074 (
            .O(N__36823),
            .I(N__36820));
    Odrv4 I__4073 (
            .O(N__36820),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12247 ));
    InMux I__4072 (
            .O(N__36817),
            .I(N__36814));
    LocalMux I__4071 (
            .O(N__36814),
            .I(N__36811));
    Odrv4 I__4070 (
            .O(N__36811),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13484 ));
    CascadeMux I__4069 (
            .O(N__36808),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11647_cascade_ ));
    InMux I__4068 (
            .O(N__36805),
            .I(N__36802));
    LocalMux I__4067 (
            .O(N__36802),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11648 ));
    InMux I__4066 (
            .O(N__36799),
            .I(N__36796));
    LocalMux I__4065 (
            .O(N__36796),
            .I(N__36793));
    Span4Mux_v I__4064 (
            .O(N__36793),
            .I(N__36790));
    Span4Mux_v I__4063 (
            .O(N__36790),
            .I(N__36787));
    Odrv4 I__4062 (
            .O(N__36787),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13487 ));
    InMux I__4061 (
            .O(N__36784),
            .I(N__36780));
    CascadeMux I__4060 (
            .O(N__36783),
            .I(N__36777));
    LocalMux I__4059 (
            .O(N__36780),
            .I(N__36774));
    InMux I__4058 (
            .O(N__36777),
            .I(N__36771));
    Odrv4 I__4057 (
            .O(N__36774),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_10 ));
    LocalMux I__4056 (
            .O(N__36771),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_10 ));
    InMux I__4055 (
            .O(N__36766),
            .I(N__36760));
    InMux I__4054 (
            .O(N__36765),
            .I(N__36760));
    LocalMux I__4053 (
            .O(N__36760),
            .I(REG_mem_16_3));
    InMux I__4052 (
            .O(N__36757),
            .I(N__36751));
    InMux I__4051 (
            .O(N__36756),
            .I(N__36751));
    LocalMux I__4050 (
            .O(N__36751),
            .I(REG_mem_17_3));
    InMux I__4049 (
            .O(N__36748),
            .I(N__36745));
    LocalMux I__4048 (
            .O(N__36745),
            .I(N__36742));
    Span4Mux_v I__4047 (
            .O(N__36742),
            .I(N__36739));
    Odrv4 I__4046 (
            .O(N__36739),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13814 ));
    CascadeMux I__4045 (
            .O(N__36736),
            .I(N__36733));
    InMux I__4044 (
            .O(N__36733),
            .I(N__36730));
    LocalMux I__4043 (
            .O(N__36730),
            .I(N__36727));
    Span12Mux_v I__4042 (
            .O(N__36727),
            .I(N__36723));
    InMux I__4041 (
            .O(N__36726),
            .I(N__36720));
    Odrv12 I__4040 (
            .O(N__36723),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_15 ));
    LocalMux I__4039 (
            .O(N__36720),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_15 ));
    InMux I__4038 (
            .O(N__36715),
            .I(N__36712));
    LocalMux I__4037 (
            .O(N__36712),
            .I(N__36709));
    Span4Mux_v I__4036 (
            .O(N__36709),
            .I(N__36705));
    CascadeMux I__4035 (
            .O(N__36708),
            .I(N__36702));
    Span4Mux_v I__4034 (
            .O(N__36705),
            .I(N__36699));
    InMux I__4033 (
            .O(N__36702),
            .I(N__36696));
    Odrv4 I__4032 (
            .O(N__36699),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_3 ));
    LocalMux I__4031 (
            .O(N__36696),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_3 ));
    CascadeMux I__4030 (
            .O(N__36691),
            .I(N__36688));
    InMux I__4029 (
            .O(N__36688),
            .I(N__36685));
    LocalMux I__4028 (
            .O(N__36685),
            .I(N__36682));
    Span4Mux_v I__4027 (
            .O(N__36682),
            .I(N__36679));
    Odrv4 I__4026 (
            .O(N__36679),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12190 ));
    InMux I__4025 (
            .O(N__36676),
            .I(N__36672));
    CascadeMux I__4024 (
            .O(N__36675),
            .I(N__36669));
    LocalMux I__4023 (
            .O(N__36672),
            .I(N__36666));
    InMux I__4022 (
            .O(N__36669),
            .I(N__36663));
    Odrv12 I__4021 (
            .O(N__36666),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_0 ));
    LocalMux I__4020 (
            .O(N__36663),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_0 ));
    CascadeMux I__4019 (
            .O(N__36658),
            .I(N__36654));
    InMux I__4018 (
            .O(N__36657),
            .I(N__36651));
    InMux I__4017 (
            .O(N__36654),
            .I(N__36648));
    LocalMux I__4016 (
            .O(N__36651),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_3 ));
    LocalMux I__4015 (
            .O(N__36648),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_3 ));
    InMux I__4014 (
            .O(N__36643),
            .I(N__36639));
    InMux I__4013 (
            .O(N__36642),
            .I(N__36636));
    LocalMux I__4012 (
            .O(N__36639),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_15 ));
    LocalMux I__4011 (
            .O(N__36636),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_15 ));
    InMux I__4010 (
            .O(N__36631),
            .I(N__36628));
    LocalMux I__4009 (
            .O(N__36628),
            .I(N__36625));
    Span4Mux_v I__4008 (
            .O(N__36625),
            .I(N__36622));
    Span4Mux_h I__4007 (
            .O(N__36622),
            .I(N__36618));
    InMux I__4006 (
            .O(N__36621),
            .I(N__36615));
    Odrv4 I__4005 (
            .O(N__36618),
            .I(REG_mem_23_3));
    LocalMux I__4004 (
            .O(N__36615),
            .I(REG_mem_23_3));
    CascadeMux I__4003 (
            .O(N__36610),
            .I(N__36607));
    InMux I__4002 (
            .O(N__36607),
            .I(N__36601));
    InMux I__4001 (
            .O(N__36606),
            .I(N__36601));
    LocalMux I__4000 (
            .O(N__36601),
            .I(REG_mem_17_15));
    CascadeMux I__3999 (
            .O(N__36598),
            .I(N__36594));
    InMux I__3998 (
            .O(N__36597),
            .I(N__36591));
    InMux I__3997 (
            .O(N__36594),
            .I(N__36588));
    LocalMux I__3996 (
            .O(N__36591),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_15 ));
    LocalMux I__3995 (
            .O(N__36588),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_15 ));
    CascadeMux I__3994 (
            .O(N__36583),
            .I(N__36580));
    InMux I__3993 (
            .O(N__36580),
            .I(N__36577));
    LocalMux I__3992 (
            .O(N__36577),
            .I(N__36574));
    Span4Mux_h I__3991 (
            .O(N__36574),
            .I(N__36570));
    CascadeMux I__3990 (
            .O(N__36573),
            .I(N__36567));
    Span4Mux_v I__3989 (
            .O(N__36570),
            .I(N__36564));
    InMux I__3988 (
            .O(N__36567),
            .I(N__36561));
    Odrv4 I__3987 (
            .O(N__36564),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_10 ));
    LocalMux I__3986 (
            .O(N__36561),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_10 ));
    InMux I__3985 (
            .O(N__36556),
            .I(N__36552));
    CascadeMux I__3984 (
            .O(N__36555),
            .I(N__36549));
    LocalMux I__3983 (
            .O(N__36552),
            .I(N__36546));
    InMux I__3982 (
            .O(N__36549),
            .I(N__36543));
    Odrv4 I__3981 (
            .O(N__36546),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_3 ));
    LocalMux I__3980 (
            .O(N__36543),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_3 ));
    CascadeMux I__3979 (
            .O(N__36538),
            .I(N__36534));
    InMux I__3978 (
            .O(N__36537),
            .I(N__36531));
    InMux I__3977 (
            .O(N__36534),
            .I(N__36528));
    LocalMux I__3976 (
            .O(N__36531),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_9 ));
    LocalMux I__3975 (
            .O(N__36528),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_9 ));
    InMux I__3974 (
            .O(N__36523),
            .I(N__36520));
    LocalMux I__3973 (
            .O(N__36520),
            .I(N__36517));
    Span4Mux_v I__3972 (
            .O(N__36517),
            .I(N__36514));
    Span4Mux_v I__3971 (
            .O(N__36514),
            .I(N__36511));
    Span4Mux_v I__3970 (
            .O(N__36511),
            .I(N__36508));
    Odrv4 I__3969 (
            .O(N__36508),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11530 ));
    InMux I__3968 (
            .O(N__36505),
            .I(N__36501));
    InMux I__3967 (
            .O(N__36504),
            .I(N__36498));
    LocalMux I__3966 (
            .O(N__36501),
            .I(N__36495));
    LocalMux I__3965 (
            .O(N__36498),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_12 ));
    Odrv4 I__3964 (
            .O(N__36495),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_12 ));
    InMux I__3963 (
            .O(N__36490),
            .I(N__36487));
    LocalMux I__3962 (
            .O(N__36487),
            .I(N__36483));
    CascadeMux I__3961 (
            .O(N__36486),
            .I(N__36480));
    Span4Mux_h I__3960 (
            .O(N__36483),
            .I(N__36477));
    InMux I__3959 (
            .O(N__36480),
            .I(N__36474));
    Odrv4 I__3958 (
            .O(N__36477),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_15 ));
    LocalMux I__3957 (
            .O(N__36474),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_15 ));
    CascadeMux I__3956 (
            .O(N__36469),
            .I(N__36465));
    InMux I__3955 (
            .O(N__36468),
            .I(N__36462));
    InMux I__3954 (
            .O(N__36465),
            .I(N__36459));
    LocalMux I__3953 (
            .O(N__36462),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_9 ));
    LocalMux I__3952 (
            .O(N__36459),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_9 ));
    CascadeMux I__3951 (
            .O(N__36454),
            .I(N__36450));
    InMux I__3950 (
            .O(N__36453),
            .I(N__36445));
    InMux I__3949 (
            .O(N__36450),
            .I(N__36445));
    LocalMux I__3948 (
            .O(N__36445),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_9 ));
    InMux I__3947 (
            .O(N__36442),
            .I(N__36439));
    LocalMux I__3946 (
            .O(N__36439),
            .I(N__36436));
    Span4Mux_v I__3945 (
            .O(N__36436),
            .I(N__36433));
    Odrv4 I__3944 (
            .O(N__36433),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12463 ));
    InMux I__3943 (
            .O(N__36430),
            .I(N__36426));
    InMux I__3942 (
            .O(N__36429),
            .I(N__36423));
    LocalMux I__3941 (
            .O(N__36426),
            .I(REG_mem_16_15));
    LocalMux I__3940 (
            .O(N__36423),
            .I(REG_mem_16_15));
    CascadeMux I__3939 (
            .O(N__36418),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12833_cascade_ ));
    InMux I__3938 (
            .O(N__36415),
            .I(N__36412));
    LocalMux I__3937 (
            .O(N__36412),
            .I(N__36409));
    Span4Mux_h I__3936 (
            .O(N__36409),
            .I(N__36406));
    Odrv4 I__3935 (
            .O(N__36406),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12070 ));
    CascadeMux I__3934 (
            .O(N__36403),
            .I(N__36399));
    InMux I__3933 (
            .O(N__36402),
            .I(N__36396));
    InMux I__3932 (
            .O(N__36399),
            .I(N__36393));
    LocalMux I__3931 (
            .O(N__36396),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_15 ));
    LocalMux I__3930 (
            .O(N__36393),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_15 ));
    CascadeMux I__3929 (
            .O(N__36388),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12788_cascade_ ));
    InMux I__3928 (
            .O(N__36385),
            .I(N__36382));
    LocalMux I__3927 (
            .O(N__36382),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12791 ));
    InMux I__3926 (
            .O(N__36379),
            .I(N__36376));
    LocalMux I__3925 (
            .O(N__36376),
            .I(N__36373));
    Odrv4 I__3924 (
            .O(N__36373),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12460 ));
    InMux I__3923 (
            .O(N__36370),
            .I(N__36364));
    InMux I__3922 (
            .O(N__36369),
            .I(N__36364));
    LocalMux I__3921 (
            .O(N__36364),
            .I(REG_mem_55_9));
    InMux I__3920 (
            .O(N__36361),
            .I(N__36355));
    InMux I__3919 (
            .O(N__36360),
            .I(N__36355));
    LocalMux I__3918 (
            .O(N__36355),
            .I(REG_mem_26_9));
    CascadeMux I__3917 (
            .O(N__36352),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13028_cascade_ ));
    CascadeMux I__3916 (
            .O(N__36349),
            .I(N__36345));
    InMux I__3915 (
            .O(N__36348),
            .I(N__36340));
    InMux I__3914 (
            .O(N__36345),
            .I(N__36340));
    LocalMux I__3913 (
            .O(N__36340),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_9 ));
    CascadeMux I__3912 (
            .O(N__36337),
            .I(N__36333));
    InMux I__3911 (
            .O(N__36336),
            .I(N__36328));
    InMux I__3910 (
            .O(N__36333),
            .I(N__36328));
    LocalMux I__3909 (
            .O(N__36328),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_9 ));
    InMux I__3908 (
            .O(N__36325),
            .I(N__36322));
    LocalMux I__3907 (
            .O(N__36322),
            .I(\usb3_if_inst.usb3_data_in_latched_10 ));
    InMux I__3906 (
            .O(N__36319),
            .I(N__36316));
    LocalMux I__3905 (
            .O(N__36316),
            .I(\usb3_if_inst.usb3_data_in_latched_11 ));
    InMux I__3904 (
            .O(N__36313),
            .I(N__36310));
    LocalMux I__3903 (
            .O(N__36310),
            .I(\usb3_if_inst.usb3_data_in_latched_12 ));
    InMux I__3902 (
            .O(N__36307),
            .I(N__36304));
    LocalMux I__3901 (
            .O(N__36304),
            .I(N__36301));
    Span4Mux_h I__3900 (
            .O(N__36301),
            .I(N__36298));
    Odrv4 I__3899 (
            .O(N__36298),
            .I(\usb3_if_inst.usb3_data_in_latched_13 ));
    CascadeMux I__3898 (
            .O(N__36295),
            .I(N__36291));
    InMux I__3897 (
            .O(N__36294),
            .I(N__36286));
    InMux I__3896 (
            .O(N__36291),
            .I(N__36286));
    LocalMux I__3895 (
            .O(N__36286),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_9 ));
    InMux I__3894 (
            .O(N__36283),
            .I(N__36280));
    LocalMux I__3893 (
            .O(N__36280),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12461 ));
    CascadeMux I__3892 (
            .O(N__36277),
            .I(N__36274));
    InMux I__3891 (
            .O(N__36274),
            .I(N__36271));
    LocalMux I__3890 (
            .O(N__36271),
            .I(N__36268));
    Odrv4 I__3889 (
            .O(N__36268),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13208 ));
    InMux I__3888 (
            .O(N__36265),
            .I(N__36262));
    LocalMux I__3887 (
            .O(N__36262),
            .I(N__36258));
    InMux I__3886 (
            .O(N__36261),
            .I(N__36255));
    Odrv4 I__3885 (
            .O(N__36258),
            .I(REG_mem_26_12));
    LocalMux I__3884 (
            .O(N__36255),
            .I(REG_mem_26_12));
    CascadeMux I__3883 (
            .O(N__36250),
            .I(N__36246));
    CascadeMux I__3882 (
            .O(N__36249),
            .I(N__36243));
    InMux I__3881 (
            .O(N__36246),
            .I(N__36238));
    InMux I__3880 (
            .O(N__36243),
            .I(N__36238));
    LocalMux I__3879 (
            .O(N__36238),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_12 ));
    CascadeMux I__3878 (
            .O(N__36235),
            .I(N__36231));
    InMux I__3877 (
            .O(N__36234),
            .I(N__36226));
    InMux I__3876 (
            .O(N__36231),
            .I(N__36226));
    LocalMux I__3875 (
            .O(N__36226),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_12 ));
    InMux I__3874 (
            .O(N__36223),
            .I(N__36217));
    InMux I__3873 (
            .O(N__36222),
            .I(N__36217));
    LocalMux I__3872 (
            .O(N__36217),
            .I(REG_mem_55_12));
    CascadeMux I__3871 (
            .O(N__36214),
            .I(N__36211));
    InMux I__3870 (
            .O(N__36211),
            .I(N__36208));
    LocalMux I__3869 (
            .O(N__36208),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12292 ));
    InMux I__3868 (
            .O(N__36205),
            .I(N__36202));
    LocalMux I__3867 (
            .O(N__36202),
            .I(N__36199));
    Span4Mux_v I__3866 (
            .O(N__36199),
            .I(N__36196));
    Odrv4 I__3865 (
            .O(N__36196),
            .I(FIFO_D10_c_10));
    InMux I__3864 (
            .O(N__36193),
            .I(N__36190));
    LocalMux I__3863 (
            .O(N__36190),
            .I(N__36186));
    CascadeMux I__3862 (
            .O(N__36189),
            .I(N__36183));
    Span4Mux_h I__3861 (
            .O(N__36186),
            .I(N__36180));
    InMux I__3860 (
            .O(N__36183),
            .I(N__36177));
    Odrv4 I__3859 (
            .O(N__36180),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_12 ));
    LocalMux I__3858 (
            .O(N__36177),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_12 ));
    CascadeMux I__3857 (
            .O(N__36172),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13100_cascade_ ));
    InMux I__3856 (
            .O(N__36169),
            .I(N__36166));
    LocalMux I__3855 (
            .O(N__36166),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12372 ));
    InMux I__3854 (
            .O(N__36163),
            .I(N__36160));
    LocalMux I__3853 (
            .O(N__36160),
            .I(N__36157));
    Odrv4 I__3852 (
            .O(N__36157),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12293 ));
    InMux I__3851 (
            .O(N__36154),
            .I(N__36151));
    LocalMux I__3850 (
            .O(N__36151),
            .I(N__36148));
    Odrv12 I__3849 (
            .O(N__36148),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12298 ));
    InMux I__3848 (
            .O(N__36145),
            .I(N__36142));
    LocalMux I__3847 (
            .O(N__36142),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13220 ));
    InMux I__3846 (
            .O(N__36139),
            .I(N__36136));
    LocalMux I__3845 (
            .O(N__36136),
            .I(N__36133));
    Odrv4 I__3844 (
            .O(N__36133),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14189 ));
    CascadeMux I__3843 (
            .O(N__36130),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11670_cascade_ ));
    InMux I__3842 (
            .O(N__36127),
            .I(N__36124));
    LocalMux I__3841 (
            .O(N__36124),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13223 ));
    CascadeMux I__3840 (
            .O(N__36121),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11576_cascade_ ));
    InMux I__3839 (
            .O(N__36118),
            .I(N__36115));
    LocalMux I__3838 (
            .O(N__36115),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13097 ));
    CascadeMux I__3837 (
            .O(N__36112),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11577_cascade_ ));
    InMux I__3836 (
            .O(N__36109),
            .I(N__36106));
    LocalMux I__3835 (
            .O(N__36106),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14054 ));
    InMux I__3834 (
            .O(N__36103),
            .I(N__36100));
    LocalMux I__3833 (
            .O(N__36100),
            .I(N__36097));
    Span4Mux_h I__3832 (
            .O(N__36097),
            .I(N__36094));
    Span4Mux_v I__3831 (
            .O(N__36094),
            .I(N__36090));
    CascadeMux I__3830 (
            .O(N__36093),
            .I(N__36087));
    Span4Mux_v I__3829 (
            .O(N__36090),
            .I(N__36084));
    InMux I__3828 (
            .O(N__36087),
            .I(N__36081));
    Odrv4 I__3827 (
            .O(N__36084),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_15 ));
    LocalMux I__3826 (
            .O(N__36081),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_15 ));
    InMux I__3825 (
            .O(N__36076),
            .I(N__36073));
    LocalMux I__3824 (
            .O(N__36073),
            .I(N__36070));
    Span4Mux_v I__3823 (
            .O(N__36070),
            .I(N__36067));
    Span4Mux_v I__3822 (
            .O(N__36067),
            .I(N__36063));
    InMux I__3821 (
            .O(N__36066),
            .I(N__36060));
    Odrv4 I__3820 (
            .O(N__36063),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_15 ));
    LocalMux I__3819 (
            .O(N__36060),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_15 ));
    CascadeMux I__3818 (
            .O(N__36055),
            .I(N__36051));
    InMux I__3817 (
            .O(N__36054),
            .I(N__36048));
    InMux I__3816 (
            .O(N__36051),
            .I(N__36045));
    LocalMux I__3815 (
            .O(N__36048),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_13 ));
    LocalMux I__3814 (
            .O(N__36045),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_13 ));
    InMux I__3813 (
            .O(N__36040),
            .I(N__36037));
    LocalMux I__3812 (
            .O(N__36037),
            .I(N__36033));
    InMux I__3811 (
            .O(N__36036),
            .I(N__36030));
    Odrv4 I__3810 (
            .O(N__36033),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_13 ));
    LocalMux I__3809 (
            .O(N__36030),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_13 ));
    InMux I__3808 (
            .O(N__36025),
            .I(N__36021));
    CascadeMux I__3807 (
            .O(N__36024),
            .I(N__36018));
    LocalMux I__3806 (
            .O(N__36021),
            .I(N__36015));
    InMux I__3805 (
            .O(N__36018),
            .I(N__36012));
    Odrv12 I__3804 (
            .O(N__36015),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_12 ));
    LocalMux I__3803 (
            .O(N__36012),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_12 ));
    CascadeMux I__3802 (
            .O(N__36007),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12878_cascade_ ));
    InMux I__3801 (
            .O(N__36004),
            .I(N__36000));
    CascadeMux I__3800 (
            .O(N__36003),
            .I(N__35997));
    LocalMux I__3799 (
            .O(N__36000),
            .I(N__35994));
    InMux I__3798 (
            .O(N__35997),
            .I(N__35991));
    Odrv4 I__3797 (
            .O(N__35994),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_12 ));
    LocalMux I__3796 (
            .O(N__35991),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_12 ));
    CascadeMux I__3795 (
            .O(N__35986),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12881_cascade_ ));
    CascadeMux I__3794 (
            .O(N__35983),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13094_cascade_ ));
    InMux I__3793 (
            .O(N__35980),
            .I(N__35976));
    CascadeMux I__3792 (
            .O(N__35979),
            .I(N__35973));
    LocalMux I__3791 (
            .O(N__35976),
            .I(N__35970));
    InMux I__3790 (
            .O(N__35973),
            .I(N__35967));
    Odrv4 I__3789 (
            .O(N__35970),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_12 ));
    LocalMux I__3788 (
            .O(N__35967),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_12 ));
    InMux I__3787 (
            .O(N__35962),
            .I(N__35959));
    LocalMux I__3786 (
            .O(N__35959),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12354 ));
    CascadeMux I__3785 (
            .O(N__35956),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14030_cascade_ ));
    InMux I__3784 (
            .O(N__35953),
            .I(N__35950));
    LocalMux I__3783 (
            .O(N__35950),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14024 ));
    InMux I__3782 (
            .O(N__35947),
            .I(N__35944));
    LocalMux I__3781 (
            .O(N__35944),
            .I(N__35941));
    Odrv4 I__3780 (
            .O(N__35941),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11559 ));
    InMux I__3779 (
            .O(N__35938),
            .I(N__35934));
    InMux I__3778 (
            .O(N__35937),
            .I(N__35931));
    LocalMux I__3777 (
            .O(N__35934),
            .I(REG_mem_5_12));
    LocalMux I__3776 (
            .O(N__35931),
            .I(REG_mem_5_12));
    CascadeMux I__3775 (
            .O(N__35926),
            .I(N__35923));
    InMux I__3774 (
            .O(N__35923),
            .I(N__35917));
    InMux I__3773 (
            .O(N__35922),
            .I(N__35917));
    LocalMux I__3772 (
            .O(N__35917),
            .I(REG_mem_26_13));
    InMux I__3771 (
            .O(N__35914),
            .I(N__35911));
    LocalMux I__3770 (
            .O(N__35911),
            .I(N__35908));
    Span4Mux_v I__3769 (
            .O(N__35908),
            .I(N__35904));
    InMux I__3768 (
            .O(N__35907),
            .I(N__35901));
    Odrv4 I__3767 (
            .O(N__35904),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_12 ));
    LocalMux I__3766 (
            .O(N__35901),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_12 ));
    InMux I__3765 (
            .O(N__35896),
            .I(N__35892));
    CascadeMux I__3764 (
            .O(N__35895),
            .I(N__35889));
    LocalMux I__3763 (
            .O(N__35892),
            .I(N__35886));
    InMux I__3762 (
            .O(N__35889),
            .I(N__35883));
    Odrv12 I__3761 (
            .O(N__35886),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_13 ));
    LocalMux I__3760 (
            .O(N__35883),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_13 ));
    InMux I__3759 (
            .O(N__35878),
            .I(N__35875));
    LocalMux I__3758 (
            .O(N__35875),
            .I(N__35871));
    InMux I__3757 (
            .O(N__35874),
            .I(N__35868));
    Odrv4 I__3756 (
            .O(N__35871),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_13 ));
    LocalMux I__3755 (
            .O(N__35868),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_13 ));
    CascadeMux I__3754 (
            .O(N__35863),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13184_cascade_ ));
    CascadeMux I__3753 (
            .O(N__35860),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12890_cascade_ ));
    InMux I__3752 (
            .O(N__35857),
            .I(N__35854));
    LocalMux I__3751 (
            .O(N__35854),
            .I(N__35851));
    Odrv4 I__3750 (
            .O(N__35851),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13187 ));
    CascadeMux I__3749 (
            .O(N__35848),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12893_cascade_ ));
    InMux I__3748 (
            .O(N__35845),
            .I(N__35842));
    LocalMux I__3747 (
            .O(N__35842),
            .I(N__35839));
    Odrv12 I__3746 (
            .O(N__35839),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12464 ));
    InMux I__3745 (
            .O(N__35836),
            .I(N__35832));
    InMux I__3744 (
            .O(N__35835),
            .I(N__35829));
    LocalMux I__3743 (
            .O(N__35832),
            .I(REG_mem_58_9));
    LocalMux I__3742 (
            .O(N__35829),
            .I(REG_mem_58_9));
    CascadeMux I__3741 (
            .O(N__35824),
            .I(N__35820));
    InMux I__3740 (
            .O(N__35823),
            .I(N__35815));
    InMux I__3739 (
            .O(N__35820),
            .I(N__35815));
    LocalMux I__3738 (
            .O(N__35815),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_9 ));
    InMux I__3737 (
            .O(N__35812),
            .I(N__35809));
    LocalMux I__3736 (
            .O(N__35809),
            .I(N__35806));
    Odrv4 I__3735 (
            .O(N__35806),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11675 ));
    InMux I__3734 (
            .O(N__35803),
            .I(N__35799));
    CascadeMux I__3733 (
            .O(N__35802),
            .I(N__35796));
    LocalMux I__3732 (
            .O(N__35799),
            .I(N__35793));
    InMux I__3731 (
            .O(N__35796),
            .I(N__35790));
    Odrv12 I__3730 (
            .O(N__35793),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_15 ));
    LocalMux I__3729 (
            .O(N__35790),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_15 ));
    InMux I__3728 (
            .O(N__35785),
            .I(N__35782));
    LocalMux I__3727 (
            .O(N__35782),
            .I(N__35778));
    CascadeMux I__3726 (
            .O(N__35781),
            .I(N__35775));
    Span4Mux_v I__3725 (
            .O(N__35778),
            .I(N__35772));
    InMux I__3724 (
            .O(N__35775),
            .I(N__35769));
    Odrv4 I__3723 (
            .O(N__35772),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_14 ));
    LocalMux I__3722 (
            .O(N__35769),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_14 ));
    InMux I__3721 (
            .O(N__35764),
            .I(N__35761));
    LocalMux I__3720 (
            .O(N__35761),
            .I(N__35758));
    Span4Mux_v I__3719 (
            .O(N__35758),
            .I(N__35754));
    InMux I__3718 (
            .O(N__35757),
            .I(N__35751));
    Odrv4 I__3717 (
            .O(N__35754),
            .I(REG_mem_12_7));
    LocalMux I__3716 (
            .O(N__35751),
            .I(REG_mem_12_7));
    InMux I__3715 (
            .O(N__35746),
            .I(N__35743));
    LocalMux I__3714 (
            .O(N__35743),
            .I(N__35739));
    InMux I__3713 (
            .O(N__35742),
            .I(N__35736));
    Odrv12 I__3712 (
            .O(N__35739),
            .I(REG_mem_8_10));
    LocalMux I__3711 (
            .O(N__35736),
            .I(REG_mem_8_10));
    CascadeMux I__3710 (
            .O(N__35731),
            .I(N__35728));
    InMux I__3709 (
            .O(N__35728),
            .I(N__35722));
    InMux I__3708 (
            .O(N__35727),
            .I(N__35722));
    LocalMux I__3707 (
            .O(N__35722),
            .I(REG_mem_15_14));
    CascadeMux I__3706 (
            .O(N__35719),
            .I(N__35716));
    InMux I__3705 (
            .O(N__35716),
            .I(N__35713));
    LocalMux I__3704 (
            .O(N__35713),
            .I(N__35710));
    Span4Mux_v I__3703 (
            .O(N__35710),
            .I(N__35707));
    Span4Mux_h I__3702 (
            .O(N__35707),
            .I(N__35703));
    CascadeMux I__3701 (
            .O(N__35706),
            .I(N__35700));
    Span4Mux_v I__3700 (
            .O(N__35703),
            .I(N__35697));
    InMux I__3699 (
            .O(N__35700),
            .I(N__35694));
    Odrv4 I__3698 (
            .O(N__35697),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_13 ));
    LocalMux I__3697 (
            .O(N__35694),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_13 ));
    InMux I__3696 (
            .O(N__35689),
            .I(N__35686));
    LocalMux I__3695 (
            .O(N__35686),
            .I(N__35683));
    Span4Mux_v I__3694 (
            .O(N__35683),
            .I(N__35680));
    Span4Mux_h I__3693 (
            .O(N__35680),
            .I(N__35677));
    Sp12to4 I__3692 (
            .O(N__35677),
            .I(N__35673));
    InMux I__3691 (
            .O(N__35676),
            .I(N__35670));
    Odrv12 I__3690 (
            .O(N__35673),
            .I(REG_mem_63_3));
    LocalMux I__3689 (
            .O(N__35670),
            .I(REG_mem_63_3));
    InMux I__3688 (
            .O(N__35665),
            .I(N__35662));
    LocalMux I__3687 (
            .O(N__35662),
            .I(N__35658));
    InMux I__3686 (
            .O(N__35661),
            .I(N__35655));
    Odrv12 I__3685 (
            .O(N__35658),
            .I(REG_mem_63_9));
    LocalMux I__3684 (
            .O(N__35655),
            .I(REG_mem_63_9));
    CascadeMux I__3683 (
            .O(N__35650),
            .I(N__35647));
    InMux I__3682 (
            .O(N__35647),
            .I(N__35644));
    LocalMux I__3681 (
            .O(N__35644),
            .I(N__35641));
    Odrv4 I__3680 (
            .O(N__35641),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13124 ));
    InMux I__3679 (
            .O(N__35638),
            .I(N__35634));
    CascadeMux I__3678 (
            .O(N__35637),
            .I(N__35631));
    LocalMux I__3677 (
            .O(N__35634),
            .I(N__35628));
    InMux I__3676 (
            .O(N__35631),
            .I(N__35625));
    Odrv12 I__3675 (
            .O(N__35628),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_9 ));
    LocalMux I__3674 (
            .O(N__35625),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_9 ));
    CascadeMux I__3673 (
            .O(N__35620),
            .I(N__35617));
    InMux I__3672 (
            .O(N__35617),
            .I(N__35613));
    InMux I__3671 (
            .O(N__35616),
            .I(N__35610));
    LocalMux I__3670 (
            .O(N__35613),
            .I(REG_mem_55_10));
    LocalMux I__3669 (
            .O(N__35610),
            .I(REG_mem_55_10));
    CascadeMux I__3668 (
            .O(N__35605),
            .I(N__35602));
    InMux I__3667 (
            .O(N__35602),
            .I(N__35596));
    InMux I__3666 (
            .O(N__35601),
            .I(N__35596));
    LocalMux I__3665 (
            .O(N__35596),
            .I(REG_mem_49_10));
    InMux I__3664 (
            .O(N__35593),
            .I(N__35590));
    LocalMux I__3663 (
            .O(N__35590),
            .I(N__35587));
    Odrv4 I__3662 (
            .O(N__35587),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11674 ));
    InMux I__3661 (
            .O(N__35584),
            .I(N__35578));
    InMux I__3660 (
            .O(N__35583),
            .I(N__35578));
    LocalMux I__3659 (
            .O(N__35578),
            .I(REG_mem_13_14));
    CascadeMux I__3658 (
            .O(N__35575),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13664_cascade_ ));
    InMux I__3657 (
            .O(N__35572),
            .I(N__35569));
    LocalMux I__3656 (
            .O(N__35569),
            .I(N__35566));
    Span4Mux_v I__3655 (
            .O(N__35566),
            .I(N__35563));
    Odrv4 I__3654 (
            .O(N__35563),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13667 ));
    InMux I__3653 (
            .O(N__35560),
            .I(N__35554));
    InMux I__3652 (
            .O(N__35559),
            .I(N__35554));
    LocalMux I__3651 (
            .O(N__35554),
            .I(REG_mem_12_14));
    InMux I__3650 (
            .O(N__35551),
            .I(N__35545));
    InMux I__3649 (
            .O(N__35550),
            .I(N__35545));
    LocalMux I__3648 (
            .O(N__35545),
            .I(REG_mem_14_14));
    CascadeMux I__3647 (
            .O(N__35542),
            .I(N__35539));
    InMux I__3646 (
            .O(N__35539),
            .I(N__35535));
    InMux I__3645 (
            .O(N__35538),
            .I(N__35532));
    LocalMux I__3644 (
            .O(N__35535),
            .I(REG_mem_42_9));
    LocalMux I__3643 (
            .O(N__35532),
            .I(REG_mem_42_9));
    InMux I__3642 (
            .O(N__35527),
            .I(N__35524));
    LocalMux I__3641 (
            .O(N__35524),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12854 ));
    InMux I__3640 (
            .O(N__35521),
            .I(N__35518));
    LocalMux I__3639 (
            .O(N__35518),
            .I(N__35515));
    Span4Mux_v I__3638 (
            .O(N__35515),
            .I(N__35512));
    Span4Mux_h I__3637 (
            .O(N__35512),
            .I(N__35509));
    Span4Mux_v I__3636 (
            .O(N__35509),
            .I(N__35506));
    Odrv4 I__3635 (
            .O(N__35506),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12959 ));
    InMux I__3634 (
            .O(N__35503),
            .I(N__35500));
    LocalMux I__3633 (
            .O(N__35500),
            .I(N__35497));
    Span4Mux_v I__3632 (
            .O(N__35497),
            .I(N__35494));
    Odrv4 I__3631 (
            .O(N__35494),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14300 ));
    InMux I__3630 (
            .O(N__35491),
            .I(N__35488));
    LocalMux I__3629 (
            .O(N__35488),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11501 ));
    CascadeMux I__3628 (
            .O(N__35485),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11500_cascade_ ));
    InMux I__3627 (
            .O(N__35482),
            .I(N__35479));
    LocalMux I__3626 (
            .O(N__35479),
            .I(N__35476));
    Span4Mux_v I__3625 (
            .O(N__35476),
            .I(N__35473));
    Odrv4 I__3624 (
            .O(N__35473),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12467 ));
    InMux I__3623 (
            .O(N__35470),
            .I(N__35467));
    LocalMux I__3622 (
            .O(N__35467),
            .I(N__35464));
    Span4Mux_v I__3621 (
            .O(N__35464),
            .I(N__35461));
    Odrv4 I__3620 (
            .O(N__35461),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13127 ));
    InMux I__3619 (
            .O(N__35458),
            .I(N__35455));
    LocalMux I__3618 (
            .O(N__35455),
            .I(N__35451));
    CascadeMux I__3617 (
            .O(N__35454),
            .I(N__35448));
    Span4Mux_h I__3616 (
            .O(N__35451),
            .I(N__35445));
    InMux I__3615 (
            .O(N__35448),
            .I(N__35442));
    Odrv4 I__3614 (
            .O(N__35445),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_10 ));
    LocalMux I__3613 (
            .O(N__35442),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_10 ));
    InMux I__3612 (
            .O(N__35437),
            .I(N__35434));
    LocalMux I__3611 (
            .O(N__35434),
            .I(N__35431));
    Span4Mux_h I__3610 (
            .O(N__35431),
            .I(N__35428));
    Odrv4 I__3609 (
            .O(N__35428),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12962 ));
    InMux I__3608 (
            .O(N__35425),
            .I(N__35421));
    InMux I__3607 (
            .O(N__35424),
            .I(N__35418));
    LocalMux I__3606 (
            .O(N__35421),
            .I(REG_mem_48_10));
    LocalMux I__3605 (
            .O(N__35418),
            .I(REG_mem_48_10));
    InMux I__3604 (
            .O(N__35413),
            .I(N__35410));
    LocalMux I__3603 (
            .O(N__35410),
            .I(N__35407));
    Span4Mux_h I__3602 (
            .O(N__35407),
            .I(N__35404));
    Odrv4 I__3601 (
            .O(N__35404),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13025 ));
    InMux I__3600 (
            .O(N__35401),
            .I(N__35398));
    LocalMux I__3599 (
            .O(N__35398),
            .I(N__35394));
    InMux I__3598 (
            .O(N__35397),
            .I(N__35391));
    Odrv4 I__3597 (
            .O(N__35394),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_9 ));
    LocalMux I__3596 (
            .O(N__35391),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_9 ));
    InMux I__3595 (
            .O(N__35386),
            .I(N__35383));
    LocalMux I__3594 (
            .O(N__35383),
            .I(N__35379));
    CascadeMux I__3593 (
            .O(N__35382),
            .I(N__35376));
    Span12Mux_s8_h I__3592 (
            .O(N__35379),
            .I(N__35373));
    InMux I__3591 (
            .O(N__35376),
            .I(N__35370));
    Odrv12 I__3590 (
            .O(N__35373),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_15 ));
    LocalMux I__3589 (
            .O(N__35370),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_15 ));
    CascadeMux I__3588 (
            .O(N__35365),
            .I(N__35362));
    InMux I__3587 (
            .O(N__35362),
            .I(N__35359));
    LocalMux I__3586 (
            .O(N__35359),
            .I(N__35355));
    CascadeMux I__3585 (
            .O(N__35358),
            .I(N__35352));
    Span4Mux_h I__3584 (
            .O(N__35355),
            .I(N__35349));
    InMux I__3583 (
            .O(N__35352),
            .I(N__35346));
    Odrv4 I__3582 (
            .O(N__35349),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_15 ));
    LocalMux I__3581 (
            .O(N__35346),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_15 ));
    CascadeMux I__3580 (
            .O(N__35341),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12857_cascade_ ));
    InMux I__3579 (
            .O(N__35338),
            .I(N__35335));
    LocalMux I__3578 (
            .O(N__35335),
            .I(N__35332));
    Odrv4 I__3577 (
            .O(N__35332),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12035 ));
    CascadeMux I__3576 (
            .O(N__35329),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14150_cascade_ ));
    InMux I__3575 (
            .O(N__35326),
            .I(N__35320));
    InMux I__3574 (
            .O(N__35325),
            .I(N__35320));
    LocalMux I__3573 (
            .O(N__35320),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_15 ));
    InMux I__3572 (
            .O(N__35317),
            .I(N__35313));
    CascadeMux I__3571 (
            .O(N__35316),
            .I(N__35310));
    LocalMux I__3570 (
            .O(N__35313),
            .I(N__35307));
    InMux I__3569 (
            .O(N__35310),
            .I(N__35304));
    Odrv4 I__3568 (
            .O(N__35307),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_15 ));
    LocalMux I__3567 (
            .O(N__35304),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_15 ));
    InMux I__3566 (
            .O(N__35299),
            .I(N__35296));
    LocalMux I__3565 (
            .O(N__35296),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12034 ));
    CascadeMux I__3564 (
            .O(N__35293),
            .I(N__35289));
    InMux I__3563 (
            .O(N__35292),
            .I(N__35284));
    InMux I__3562 (
            .O(N__35289),
            .I(N__35284));
    LocalMux I__3561 (
            .O(N__35284),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_15 ));
    InMux I__3560 (
            .O(N__35281),
            .I(N__35278));
    LocalMux I__3559 (
            .O(N__35278),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12043 ));
    InMux I__3558 (
            .O(N__35275),
            .I(N__35269));
    InMux I__3557 (
            .O(N__35274),
            .I(N__35269));
    LocalMux I__3556 (
            .O(N__35269),
            .I(REG_mem_50_9));
    InMux I__3555 (
            .O(N__35266),
            .I(N__35260));
    InMux I__3554 (
            .O(N__35265),
            .I(N__35260));
    LocalMux I__3553 (
            .O(N__35260),
            .I(REG_mem_51_9));
    InMux I__3552 (
            .O(N__35257),
            .I(N__35251));
    InMux I__3551 (
            .O(N__35256),
            .I(N__35251));
    LocalMux I__3550 (
            .O(N__35251),
            .I(REG_mem_55_15));
    InMux I__3549 (
            .O(N__35248),
            .I(N__35245));
    LocalMux I__3548 (
            .O(N__35245),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12031 ));
    CascadeMux I__3547 (
            .O(N__35242),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12032_cascade_ ));
    CascadeMux I__3546 (
            .O(N__35239),
            .I(N__35235));
    InMux I__3545 (
            .O(N__35238),
            .I(N__35230));
    InMux I__3544 (
            .O(N__35235),
            .I(N__35230));
    LocalMux I__3543 (
            .O(N__35230),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_15 ));
    CascadeMux I__3542 (
            .O(N__35227),
            .I(N__35223));
    InMux I__3541 (
            .O(N__35226),
            .I(N__35218));
    InMux I__3540 (
            .O(N__35223),
            .I(N__35218));
    LocalMux I__3539 (
            .O(N__35218),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_15 ));
    InMux I__3538 (
            .O(N__35215),
            .I(N__35212));
    LocalMux I__3537 (
            .O(N__35212),
            .I(N__35209));
    Span4Mux_h I__3536 (
            .O(N__35209),
            .I(N__35206));
    Span4Mux_v I__3535 (
            .O(N__35206),
            .I(N__35203));
    Odrv4 I__3534 (
            .O(N__35203),
            .I(FIFO_D11_c_11));
    InMux I__3533 (
            .O(N__35200),
            .I(N__35197));
    LocalMux I__3532 (
            .O(N__35197),
            .I(N__35194));
    Span12Mux_h I__3531 (
            .O(N__35194),
            .I(N__35191));
    Odrv12 I__3530 (
            .O(N__35191),
            .I(FIFO_D12_c_12));
    InMux I__3529 (
            .O(N__35188),
            .I(N__35185));
    LocalMux I__3528 (
            .O(N__35185),
            .I(N__35182));
    Odrv4 I__3527 (
            .O(N__35182),
            .I(\usb3_if_inst.usb3_data_in_latched_15 ));
    CascadeMux I__3526 (
            .O(N__35179),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13166_cascade_ ));
    CascadeMux I__3525 (
            .O(N__35176),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13169_cascade_ ));
    InMux I__3524 (
            .O(N__35173),
            .I(N__35170));
    LocalMux I__3523 (
            .O(N__35170),
            .I(N__35167));
    Odrv4 I__3522 (
            .O(N__35167),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12446 ));
    CascadeMux I__3521 (
            .O(N__35164),
            .I(N__35161));
    InMux I__3520 (
            .O(N__35161),
            .I(N__35158));
    LocalMux I__3519 (
            .O(N__35158),
            .I(N__35155));
    Span4Mux_v I__3518 (
            .O(N__35155),
            .I(N__35152));
    Odrv4 I__3517 (
            .O(N__35152),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12466 ));
    CascadeMux I__3516 (
            .O(N__35149),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14330_cascade_ ));
    InMux I__3515 (
            .O(N__35146),
            .I(N__35143));
    LocalMux I__3514 (
            .O(N__35143),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11516 ));
    CascadeMux I__3513 (
            .O(N__35140),
            .I(N__35136));
    InMux I__3512 (
            .O(N__35139),
            .I(N__35133));
    InMux I__3511 (
            .O(N__35136),
            .I(N__35130));
    LocalMux I__3510 (
            .O(N__35133),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_14 ));
    LocalMux I__3509 (
            .O(N__35130),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_14 ));
    CascadeMux I__3508 (
            .O(N__35125),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11531_cascade_ ));
    CascadeMux I__3507 (
            .O(N__35122),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11509_cascade_ ));
    InMux I__3506 (
            .O(N__35119),
            .I(N__35116));
    LocalMux I__3505 (
            .O(N__35116),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14186 ));
    InMux I__3504 (
            .O(N__35113),
            .I(N__35109));
    InMux I__3503 (
            .O(N__35112),
            .I(N__35106));
    LocalMux I__3502 (
            .O(N__35109),
            .I(REG_mem_58_12));
    LocalMux I__3501 (
            .O(N__35106),
            .I(REG_mem_58_12));
    InMux I__3500 (
            .O(N__35101),
            .I(N__35095));
    InMux I__3499 (
            .O(N__35100),
            .I(N__35095));
    LocalMux I__3498 (
            .O(N__35095),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_12 ));
    InMux I__3497 (
            .O(N__35092),
            .I(N__35089));
    LocalMux I__3496 (
            .O(N__35089),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11510 ));
    CascadeMux I__3495 (
            .O(N__35086),
            .I(N__35082));
    InMux I__3494 (
            .O(N__35085),
            .I(N__35077));
    InMux I__3493 (
            .O(N__35082),
            .I(N__35077));
    LocalMux I__3492 (
            .O(N__35077),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_12 ));
    InMux I__3491 (
            .O(N__35074),
            .I(N__35068));
    InMux I__3490 (
            .O(N__35073),
            .I(N__35068));
    LocalMux I__3489 (
            .O(N__35068),
            .I(REG_mem_58_13));
    CascadeMux I__3488 (
            .O(N__35065),
            .I(N__35061));
    InMux I__3487 (
            .O(N__35064),
            .I(N__35058));
    InMux I__3486 (
            .O(N__35061),
            .I(N__35055));
    LocalMux I__3485 (
            .O(N__35058),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_13 ));
    LocalMux I__3484 (
            .O(N__35055),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_13 ));
    CascadeMux I__3483 (
            .O(N__35050),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11830_cascade_ ));
    InMux I__3482 (
            .O(N__35047),
            .I(N__35043));
    CascadeMux I__3481 (
            .O(N__35046),
            .I(N__35040));
    LocalMux I__3480 (
            .O(N__35043),
            .I(N__35037));
    InMux I__3479 (
            .O(N__35040),
            .I(N__35034));
    Odrv4 I__3478 (
            .O(N__35037),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_10 ));
    LocalMux I__3477 (
            .O(N__35034),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_10 ));
    InMux I__3476 (
            .O(N__35029),
            .I(N__35026));
    LocalMux I__3475 (
            .O(N__35026),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13490 ));
    CascadeMux I__3474 (
            .O(N__35023),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11792_cascade_ ));
    InMux I__3473 (
            .O(N__35020),
            .I(N__35017));
    LocalMux I__3472 (
            .O(N__35017),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11791 ));
    InMux I__3471 (
            .O(N__35014),
            .I(N__35011));
    LocalMux I__3470 (
            .O(N__35011),
            .I(N__35008));
    Odrv4 I__3469 (
            .O(N__35008),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13493 ));
    InMux I__3468 (
            .O(N__35005),
            .I(N__34999));
    InMux I__3467 (
            .O(N__35004),
            .I(N__34999));
    LocalMux I__3466 (
            .O(N__34999),
            .I(REG_mem_36_3));
    InMux I__3465 (
            .O(N__34996),
            .I(N__34990));
    InMux I__3464 (
            .O(N__34995),
            .I(N__34990));
    LocalMux I__3463 (
            .O(N__34990),
            .I(REG_mem_37_3));
    InMux I__3462 (
            .O(N__34987),
            .I(N__34984));
    LocalMux I__3461 (
            .O(N__34984),
            .I(N__34981));
    Odrv4 I__3460 (
            .O(N__34981),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14003 ));
    CascadeMux I__3459 (
            .O(N__34978),
            .I(N__34975));
    InMux I__3458 (
            .O(N__34975),
            .I(N__34972));
    LocalMux I__3457 (
            .O(N__34972),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14099 ));
    CascadeMux I__3456 (
            .O(N__34969),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11975_cascade_ ));
    InMux I__3455 (
            .O(N__34966),
            .I(N__34963));
    LocalMux I__3454 (
            .O(N__34963),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11976 ));
    InMux I__3453 (
            .O(N__34960),
            .I(N__34957));
    LocalMux I__3452 (
            .O(N__34957),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11523 ));
    CascadeMux I__3451 (
            .O(N__34954),
            .I(N__34951));
    InMux I__3450 (
            .O(N__34951),
            .I(N__34948));
    LocalMux I__3449 (
            .O(N__34948),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12806 ));
    InMux I__3448 (
            .O(N__34945),
            .I(N__34942));
    LocalMux I__3447 (
            .O(N__34942),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12809 ));
    InMux I__3446 (
            .O(N__34939),
            .I(N__34936));
    LocalMux I__3445 (
            .O(N__34936),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13322 ));
    CascadeMux I__3444 (
            .O(N__34933),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13274_cascade_ ));
    CascadeMux I__3443 (
            .O(N__34930),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12339_cascade_ ));
    InMux I__3442 (
            .O(N__34927),
            .I(N__34924));
    LocalMux I__3441 (
            .O(N__34924),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12327 ));
    InMux I__3440 (
            .O(N__34921),
            .I(N__34915));
    InMux I__3439 (
            .O(N__34920),
            .I(N__34915));
    LocalMux I__3438 (
            .O(N__34915),
            .I(REG_mem_63_13));
    CascadeMux I__3437 (
            .O(N__34912),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13052_cascade_ ));
    CascadeMux I__3436 (
            .O(N__34909),
            .I(N__34905));
    InMux I__3435 (
            .O(N__34908),
            .I(N__34902));
    InMux I__3434 (
            .O(N__34905),
            .I(N__34899));
    LocalMux I__3433 (
            .O(N__34902),
            .I(N__34896));
    LocalMux I__3432 (
            .O(N__34899),
            .I(N__34893));
    Odrv12 I__3431 (
            .O(N__34896),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_3 ));
    Odrv4 I__3430 (
            .O(N__34893),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_3 ));
    InMux I__3429 (
            .O(N__34888),
            .I(N__34885));
    LocalMux I__3428 (
            .O(N__34885),
            .I(N__34882));
    Odrv12 I__3427 (
            .O(N__34882),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13055 ));
    CascadeMux I__3426 (
            .O(N__34879),
            .I(N__34875));
    InMux I__3425 (
            .O(N__34878),
            .I(N__34872));
    InMux I__3424 (
            .O(N__34875),
            .I(N__34869));
    LocalMux I__3423 (
            .O(N__34872),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_3 ));
    LocalMux I__3422 (
            .O(N__34869),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_3 ));
    CascadeMux I__3421 (
            .O(N__34864),
            .I(N__34861));
    InMux I__3420 (
            .O(N__34861),
            .I(N__34858));
    LocalMux I__3419 (
            .O(N__34858),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14336 ));
    InMux I__3418 (
            .O(N__34855),
            .I(N__34849));
    InMux I__3417 (
            .O(N__34854),
            .I(N__34849));
    LocalMux I__3416 (
            .O(N__34849),
            .I(REG_mem_26_3));
    CascadeMux I__3415 (
            .O(N__34846),
            .I(N__34842));
    InMux I__3414 (
            .O(N__34845),
            .I(N__34837));
    InMux I__3413 (
            .O(N__34842),
            .I(N__34837));
    LocalMux I__3412 (
            .O(N__34837),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_3 ));
    InMux I__3411 (
            .O(N__34834),
            .I(N__34831));
    LocalMux I__3410 (
            .O(N__34831),
            .I(N__34828));
    Odrv4 I__3409 (
            .O(N__34828),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12012 ));
    CascadeMux I__3408 (
            .O(N__34825),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11991_cascade_ ));
    CascadeMux I__3407 (
            .O(N__34822),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14312_cascade_ ));
    InMux I__3406 (
            .O(N__34819),
            .I(N__34815));
    InMux I__3405 (
            .O(N__34818),
            .I(N__34812));
    LocalMux I__3404 (
            .O(N__34815),
            .I(REG_mem_5_10));
    LocalMux I__3403 (
            .O(N__34812),
            .I(REG_mem_5_10));
    InMux I__3402 (
            .O(N__34807),
            .I(N__34801));
    InMux I__3401 (
            .O(N__34806),
            .I(N__34801));
    LocalMux I__3400 (
            .O(N__34801),
            .I(REG_mem_10_10));
    InMux I__3399 (
            .O(N__34798),
            .I(N__34792));
    InMux I__3398 (
            .O(N__34797),
            .I(N__34792));
    LocalMux I__3397 (
            .O(N__34792),
            .I(REG_mem_11_10));
    CascadeMux I__3396 (
            .O(N__34789),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14180_cascade_ ));
    InMux I__3395 (
            .O(N__34786),
            .I(N__34783));
    LocalMux I__3394 (
            .O(N__34783),
            .I(N__34780));
    Odrv12 I__3393 (
            .O(N__34780),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14183 ));
    CascadeMux I__3392 (
            .O(N__34777),
            .I(N__34773));
    CascadeMux I__3391 (
            .O(N__34776),
            .I(N__34770));
    InMux I__3390 (
            .O(N__34773),
            .I(N__34767));
    InMux I__3389 (
            .O(N__34770),
            .I(N__34764));
    LocalMux I__3388 (
            .O(N__34767),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_3 ));
    LocalMux I__3387 (
            .O(N__34764),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_3 ));
    InMux I__3386 (
            .O(N__34759),
            .I(N__34756));
    LocalMux I__3385 (
            .O(N__34756),
            .I(N__34752));
    CascadeMux I__3384 (
            .O(N__34755),
            .I(N__34749));
    Span4Mux_v I__3383 (
            .O(N__34752),
            .I(N__34746));
    InMux I__3382 (
            .O(N__34749),
            .I(N__34743));
    Odrv4 I__3381 (
            .O(N__34746),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_3 ));
    LocalMux I__3380 (
            .O(N__34743),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_3 ));
    CascadeMux I__3379 (
            .O(N__34738),
            .I(N__34734));
    CascadeMux I__3378 (
            .O(N__34737),
            .I(N__34731));
    InMux I__3377 (
            .O(N__34734),
            .I(N__34728));
    InMux I__3376 (
            .O(N__34731),
            .I(N__34725));
    LocalMux I__3375 (
            .O(N__34728),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_3 ));
    LocalMux I__3374 (
            .O(N__34725),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_3 ));
    InMux I__3373 (
            .O(N__34720),
            .I(N__34717));
    LocalMux I__3372 (
            .O(N__34717),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14096 ));
    CascadeMux I__3371 (
            .O(N__34714),
            .I(N__34711));
    InMux I__3370 (
            .O(N__34711),
            .I(N__34707));
    CascadeMux I__3369 (
            .O(N__34710),
            .I(N__34704));
    LocalMux I__3368 (
            .O(N__34707),
            .I(N__34701));
    InMux I__3367 (
            .O(N__34704),
            .I(N__34698));
    Odrv12 I__3366 (
            .O(N__34701),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_3 ));
    LocalMux I__3365 (
            .O(N__34698),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_3 ));
    InMux I__3364 (
            .O(N__34693),
            .I(N__34687));
    InMux I__3363 (
            .O(N__34692),
            .I(N__34687));
    LocalMux I__3362 (
            .O(N__34687),
            .I(REG_mem_31_3));
    CascadeMux I__3361 (
            .O(N__34684),
            .I(N__34680));
    InMux I__3360 (
            .O(N__34683),
            .I(N__34677));
    InMux I__3359 (
            .O(N__34680),
            .I(N__34674));
    LocalMux I__3358 (
            .O(N__34677),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_3 ));
    LocalMux I__3357 (
            .O(N__34674),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_3 ));
    CascadeMux I__3356 (
            .O(N__34669),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14000_cascade_ ));
    CascadeMux I__3355 (
            .O(N__34666),
            .I(N__34662));
    InMux I__3354 (
            .O(N__34665),
            .I(N__34657));
    InMux I__3353 (
            .O(N__34662),
            .I(N__34657));
    LocalMux I__3352 (
            .O(N__34657),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_3 ));
    InMux I__3351 (
            .O(N__34654),
            .I(N__34651));
    LocalMux I__3350 (
            .O(N__34651),
            .I(N__34647));
    CascadeMux I__3349 (
            .O(N__34650),
            .I(N__34644));
    Span4Mux_h I__3348 (
            .O(N__34647),
            .I(N__34641));
    InMux I__3347 (
            .O(N__34644),
            .I(N__34638));
    Odrv4 I__3346 (
            .O(N__34641),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_9 ));
    LocalMux I__3345 (
            .O(N__34638),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_9 ));
    CascadeMux I__3344 (
            .O(N__34633),
            .I(N__34630));
    InMux I__3343 (
            .O(N__34630),
            .I(N__34626));
    CascadeMux I__3342 (
            .O(N__34629),
            .I(N__34623));
    LocalMux I__3341 (
            .O(N__34626),
            .I(N__34620));
    InMux I__3340 (
            .O(N__34623),
            .I(N__34617));
    Odrv12 I__3339 (
            .O(N__34620),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_9 ));
    LocalMux I__3338 (
            .O(N__34617),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_9 ));
    CascadeMux I__3337 (
            .O(N__34612),
            .I(N__34609));
    InMux I__3336 (
            .O(N__34609),
            .I(N__34606));
    LocalMux I__3335 (
            .O(N__34606),
            .I(N__34603));
    Span4Mux_v I__3334 (
            .O(N__34603),
            .I(N__34599));
    InMux I__3333 (
            .O(N__34602),
            .I(N__34596));
    Odrv4 I__3332 (
            .O(N__34599),
            .I(REG_mem_63_14));
    LocalMux I__3331 (
            .O(N__34596),
            .I(REG_mem_63_14));
    InMux I__3330 (
            .O(N__34591),
            .I(N__34587));
    InMux I__3329 (
            .O(N__34590),
            .I(N__34584));
    LocalMux I__3328 (
            .O(N__34587),
            .I(REG_mem_6_10));
    LocalMux I__3327 (
            .O(N__34584),
            .I(REG_mem_6_10));
    InMux I__3326 (
            .O(N__34579),
            .I(N__34576));
    LocalMux I__3325 (
            .O(N__34576),
            .I(N__34573));
    Sp12to4 I__3324 (
            .O(N__34573),
            .I(N__34569));
    InMux I__3323 (
            .O(N__34572),
            .I(N__34566));
    Odrv12 I__3322 (
            .O(N__34569),
            .I(REG_mem_49_14));
    LocalMux I__3321 (
            .O(N__34566),
            .I(REG_mem_49_14));
    CascadeMux I__3320 (
            .O(N__34561),
            .I(N__34558));
    InMux I__3319 (
            .O(N__34558),
            .I(N__34555));
    LocalMux I__3318 (
            .O(N__34555),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12974 ));
    CascadeMux I__3317 (
            .O(N__34552),
            .I(N__34548));
    InMux I__3316 (
            .O(N__34551),
            .I(N__34545));
    InMux I__3315 (
            .O(N__34548),
            .I(N__34542));
    LocalMux I__3314 (
            .O(N__34545),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_14 ));
    LocalMux I__3313 (
            .O(N__34542),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_14 ));
    CascadeMux I__3312 (
            .O(N__34537),
            .I(N__34533));
    InMux I__3311 (
            .O(N__34536),
            .I(N__34528));
    InMux I__3310 (
            .O(N__34533),
            .I(N__34528));
    LocalMux I__3309 (
            .O(N__34528),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_14 ));
    CascadeMux I__3308 (
            .O(N__34525),
            .I(N__34522));
    InMux I__3307 (
            .O(N__34522),
            .I(N__34519));
    LocalMux I__3306 (
            .O(N__34519),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12271 ));
    CascadeMux I__3305 (
            .O(N__34516),
            .I(N__34512));
    InMux I__3304 (
            .O(N__34515),
            .I(N__34509));
    InMux I__3303 (
            .O(N__34512),
            .I(N__34506));
    LocalMux I__3302 (
            .O(N__34509),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_14 ));
    LocalMux I__3301 (
            .O(N__34506),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_14 ));
    InMux I__3300 (
            .O(N__34501),
            .I(N__34498));
    LocalMux I__3299 (
            .O(N__34498),
            .I(N__34495));
    Odrv4 I__3298 (
            .O(N__34495),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12191 ));
    InMux I__3297 (
            .O(N__34492),
            .I(N__34488));
    InMux I__3296 (
            .O(N__34491),
            .I(N__34485));
    LocalMux I__3295 (
            .O(N__34488),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_10 ));
    LocalMux I__3294 (
            .O(N__34485),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_10 ));
    InMux I__3293 (
            .O(N__34480),
            .I(N__34476));
    InMux I__3292 (
            .O(N__34479),
            .I(N__34473));
    LocalMux I__3291 (
            .O(N__34476),
            .I(N__34470));
    LocalMux I__3290 (
            .O(N__34473),
            .I(N__34467));
    Odrv4 I__3289 (
            .O(N__34470),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_3 ));
    Odrv4 I__3288 (
            .O(N__34467),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_3 ));
    InMux I__3287 (
            .O(N__34462),
            .I(N__34456));
    InMux I__3286 (
            .O(N__34461),
            .I(N__34456));
    LocalMux I__3285 (
            .O(N__34456),
            .I(REG_mem_44_14));
    InMux I__3284 (
            .O(N__34453),
            .I(N__34450));
    LocalMux I__3283 (
            .O(N__34450),
            .I(N__34446));
    InMux I__3282 (
            .O(N__34449),
            .I(N__34443));
    Odrv4 I__3281 (
            .O(N__34446),
            .I(REG_mem_31_14));
    LocalMux I__3280 (
            .O(N__34443),
            .I(REG_mem_31_14));
    InMux I__3279 (
            .O(N__34438),
            .I(N__34435));
    LocalMux I__3278 (
            .O(N__34435),
            .I(N__34432));
    Odrv4 I__3277 (
            .O(N__34432),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12272 ));
    CascadeMux I__3276 (
            .O(N__34429),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13190_cascade_ ));
    InMux I__3275 (
            .O(N__34426),
            .I(N__34423));
    LocalMux I__3274 (
            .O(N__34423),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12248 ));
    InMux I__3273 (
            .O(N__34420),
            .I(N__34417));
    LocalMux I__3272 (
            .O(N__34417),
            .I(N__34414));
    Odrv4 I__3271 (
            .O(N__34414),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13193 ));
    InMux I__3270 (
            .O(N__34411),
            .I(N__34405));
    InMux I__3269 (
            .O(N__34410),
            .I(N__34405));
    LocalMux I__3268 (
            .O(N__34405),
            .I(REG_mem_18_14));
    InMux I__3267 (
            .O(N__34402),
            .I(N__34396));
    InMux I__3266 (
            .O(N__34401),
            .I(N__34396));
    LocalMux I__3265 (
            .O(N__34396),
            .I(REG_mem_19_14));
    CascadeMux I__3264 (
            .O(N__34393),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13160_cascade_ ));
    InMux I__3263 (
            .O(N__34390),
            .I(N__34387));
    LocalMux I__3262 (
            .O(N__34387),
            .I(N__34384));
    Span4Mux_v I__3261 (
            .O(N__34384),
            .I(N__34381));
    Span4Mux_v I__3260 (
            .O(N__34381),
            .I(N__34378));
    Odrv4 I__3259 (
            .O(N__34378),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12185 ));
    InMux I__3258 (
            .O(N__34375),
            .I(N__34372));
    LocalMux I__3257 (
            .O(N__34372),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13163 ));
    InMux I__3256 (
            .O(N__34369),
            .I(N__34365));
    InMux I__3255 (
            .O(N__34368),
            .I(N__34362));
    LocalMux I__3254 (
            .O(N__34365),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_9 ));
    LocalMux I__3253 (
            .O(N__34362),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_9 ));
    InMux I__3252 (
            .O(N__34357),
            .I(N__34354));
    LocalMux I__3251 (
            .O(N__34354),
            .I(N__34351));
    Span4Mux_v I__3250 (
            .O(N__34351),
            .I(N__34348));
    Odrv4 I__3249 (
            .O(N__34348),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13475 ));
    InMux I__3248 (
            .O(N__34345),
            .I(N__34342));
    LocalMux I__3247 (
            .O(N__34342),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13331 ));
    InMux I__3246 (
            .O(N__34339),
            .I(N__34336));
    LocalMux I__3245 (
            .O(N__34336),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11534 ));
    CascadeMux I__3244 (
            .O(N__34333),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13106_cascade_ ));
    InMux I__3243 (
            .O(N__34330),
            .I(N__34327));
    LocalMux I__3242 (
            .O(N__34327),
            .I(N__34324));
    Odrv4 I__3241 (
            .O(N__34324),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13109 ));
    InMux I__3240 (
            .O(N__34321),
            .I(N__34315));
    InMux I__3239 (
            .O(N__34320),
            .I(N__34315));
    LocalMux I__3238 (
            .O(N__34315),
            .I(REG_mem_46_14));
    CascadeMux I__3237 (
            .O(N__34312),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13046_cascade_ ));
    InMux I__3236 (
            .O(N__34309),
            .I(N__34306));
    LocalMux I__3235 (
            .O(N__34306),
            .I(N__34303));
    Odrv4 I__3234 (
            .O(N__34303),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13049 ));
    CascadeMux I__3233 (
            .O(N__34300),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12980_cascade_ ));
    InMux I__3232 (
            .O(N__34297),
            .I(N__34291));
    InMux I__3231 (
            .O(N__34296),
            .I(N__34291));
    LocalMux I__3230 (
            .O(N__34291),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_9 ));
    InMux I__3229 (
            .O(N__34288),
            .I(N__34284));
    InMux I__3228 (
            .O(N__34287),
            .I(N__34281));
    LocalMux I__3227 (
            .O(N__34284),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_9 ));
    LocalMux I__3226 (
            .O(N__34281),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_9 ));
    InMux I__3225 (
            .O(N__34276),
            .I(N__34273));
    LocalMux I__3224 (
            .O(N__34273),
            .I(N__34269));
    CascadeMux I__3223 (
            .O(N__34272),
            .I(N__34266));
    Span12Mux_s6_h I__3222 (
            .O(N__34269),
            .I(N__34263));
    InMux I__3221 (
            .O(N__34266),
            .I(N__34260));
    Odrv12 I__3220 (
            .O(N__34263),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_10 ));
    LocalMux I__3219 (
            .O(N__34260),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_10 ));
    CascadeMux I__3218 (
            .O(N__34255),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13817_cascade_ ));
    InMux I__3217 (
            .O(N__34252),
            .I(N__34249));
    LocalMux I__3216 (
            .O(N__34249),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13226 ));
    CascadeMux I__3215 (
            .O(N__34246),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11513_cascade_ ));
    InMux I__3214 (
            .O(N__34243),
            .I(N__34240));
    LocalMux I__3213 (
            .O(N__34240),
            .I(N__34237));
    Span12Mux_v I__3212 (
            .O(N__34237),
            .I(N__34234));
    Odrv12 I__3211 (
            .O(N__34234),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11525 ));
    CascadeMux I__3210 (
            .O(N__34231),
            .I(N__34227));
    InMux I__3209 (
            .O(N__34230),
            .I(N__34222));
    InMux I__3208 (
            .O(N__34227),
            .I(N__34222));
    LocalMux I__3207 (
            .O(N__34222),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_10 ));
    CascadeMux I__3206 (
            .O(N__34219),
            .I(N__34215));
    InMux I__3205 (
            .O(N__34218),
            .I(N__34212));
    InMux I__3204 (
            .O(N__34215),
            .I(N__34209));
    LocalMux I__3203 (
            .O(N__34212),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_10 ));
    LocalMux I__3202 (
            .O(N__34209),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_10 ));
    InMux I__3201 (
            .O(N__34204),
            .I(N__34201));
    LocalMux I__3200 (
            .O(N__34201),
            .I(N__34198));
    Span12Mux_h I__3199 (
            .O(N__34198),
            .I(N__34195));
    Odrv12 I__3198 (
            .O(N__34195),
            .I(FIFO_D13_c_13));
    InMux I__3197 (
            .O(N__34192),
            .I(N__34189));
    LocalMux I__3196 (
            .O(N__34189),
            .I(N__34186));
    Span4Mux_v I__3195 (
            .O(N__34186),
            .I(N__34183));
    IoSpan4Mux I__3194 (
            .O(N__34183),
            .I(N__34180));
    Odrv4 I__3193 (
            .O(N__34180),
            .I(FIFO_D14_c_14));
    InMux I__3192 (
            .O(N__34177),
            .I(N__34174));
    LocalMux I__3191 (
            .O(N__34174),
            .I(N__34171));
    Span4Mux_h I__3190 (
            .O(N__34171),
            .I(N__34168));
    Span4Mux_v I__3189 (
            .O(N__34168),
            .I(N__34165));
    Odrv4 I__3188 (
            .O(N__34165),
            .I(FIFO_D15_c_15));
    InMux I__3187 (
            .O(N__34162),
            .I(N__34159));
    LocalMux I__3186 (
            .O(N__34159),
            .I(\usb3_if_inst.usb3_data_in_latched_14 ));
    InMux I__3185 (
            .O(N__34156),
            .I(N__34150));
    InMux I__3184 (
            .O(N__34155),
            .I(N__34150));
    LocalMux I__3183 (
            .O(N__34150),
            .I(REG_mem_31_9));
    InMux I__3182 (
            .O(N__34147),
            .I(N__34144));
    LocalMux I__3181 (
            .O(N__34144),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11578 ));
    CascadeMux I__3180 (
            .O(N__34141),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11579_cascade_ ));
    InMux I__3179 (
            .O(N__34138),
            .I(N__34135));
    LocalMux I__3178 (
            .O(N__34135),
            .I(N__34132));
    Odrv4 I__3177 (
            .O(N__34132),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13271 ));
    InMux I__3176 (
            .O(N__34129),
            .I(N__34123));
    InMux I__3175 (
            .O(N__34128),
            .I(N__34123));
    LocalMux I__3174 (
            .O(N__34123),
            .I(REG_mem_36_10));
    InMux I__3173 (
            .O(N__34120),
            .I(N__34114));
    InMux I__3172 (
            .O(N__34119),
            .I(N__34114));
    LocalMux I__3171 (
            .O(N__34114),
            .I(REG_mem_37_10));
    CascadeMux I__3170 (
            .O(N__34111),
            .I(N__34107));
    CascadeMux I__3169 (
            .O(N__34110),
            .I(N__34104));
    InMux I__3168 (
            .O(N__34107),
            .I(N__34099));
    InMux I__3167 (
            .O(N__34104),
            .I(N__34099));
    LocalMux I__3166 (
            .O(N__34099),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_10 ));
    InMux I__3165 (
            .O(N__34096),
            .I(N__34090));
    InMux I__3164 (
            .O(N__34095),
            .I(N__34090));
    LocalMux I__3163 (
            .O(N__34090),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_14 ));
    InMux I__3162 (
            .O(N__34087),
            .I(N__34083));
    CascadeMux I__3161 (
            .O(N__34086),
            .I(N__34080));
    LocalMux I__3160 (
            .O(N__34083),
            .I(N__34077));
    InMux I__3159 (
            .O(N__34080),
            .I(N__34074));
    Odrv12 I__3158 (
            .O(N__34077),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_14 ));
    LocalMux I__3157 (
            .O(N__34074),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_14 ));
    InMux I__3156 (
            .O(N__34069),
            .I(N__34066));
    LocalMux I__3155 (
            .O(N__34066),
            .I(N__34063));
    Odrv4 I__3154 (
            .O(N__34063),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11584 ));
    InMux I__3153 (
            .O(N__34060),
            .I(N__34057));
    LocalMux I__3152 (
            .O(N__34057),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13268 ));
    CascadeMux I__3151 (
            .O(N__34054),
            .I(N__34050));
    InMux I__3150 (
            .O(N__34053),
            .I(N__34045));
    InMux I__3149 (
            .O(N__34050),
            .I(N__34045));
    LocalMux I__3148 (
            .O(N__34045),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_3 ));
    CascadeMux I__3147 (
            .O(N__34042),
            .I(N__34038));
    InMux I__3146 (
            .O(N__34041),
            .I(N__34033));
    InMux I__3145 (
            .O(N__34038),
            .I(N__34033));
    LocalMux I__3144 (
            .O(N__34033),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_3 ));
    CascadeMux I__3143 (
            .O(N__34030),
            .I(N__34026));
    CascadeMux I__3142 (
            .O(N__34029),
            .I(N__34023));
    InMux I__3141 (
            .O(N__34026),
            .I(N__34018));
    InMux I__3140 (
            .O(N__34023),
            .I(N__34018));
    LocalMux I__3139 (
            .O(N__34018),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_3 ));
    InMux I__3138 (
            .O(N__34015),
            .I(N__34011));
    CascadeMux I__3137 (
            .O(N__34014),
            .I(N__34008));
    LocalMux I__3136 (
            .O(N__34011),
            .I(N__34005));
    InMux I__3135 (
            .O(N__34008),
            .I(N__34002));
    Odrv4 I__3134 (
            .O(N__34005),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_10 ));
    LocalMux I__3133 (
            .O(N__34002),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_10 ));
    InMux I__3132 (
            .O(N__33997),
            .I(N__33994));
    LocalMux I__3131 (
            .O(N__33994),
            .I(N__33991));
    Odrv4 I__3130 (
            .O(N__33991),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11549 ));
    InMux I__3129 (
            .O(N__33988),
            .I(N__33984));
    CascadeMux I__3128 (
            .O(N__33987),
            .I(N__33981));
    LocalMux I__3127 (
            .O(N__33984),
            .I(N__33978));
    InMux I__3126 (
            .O(N__33981),
            .I(N__33975));
    Odrv4 I__3125 (
            .O(N__33978),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_3 ));
    LocalMux I__3124 (
            .O(N__33975),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_3 ));
    InMux I__3123 (
            .O(N__33970),
            .I(N__33966));
    CascadeMux I__3122 (
            .O(N__33969),
            .I(N__33963));
    LocalMux I__3121 (
            .O(N__33966),
            .I(N__33960));
    InMux I__3120 (
            .O(N__33963),
            .I(N__33957));
    Odrv4 I__3119 (
            .O(N__33960),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_3 ));
    LocalMux I__3118 (
            .O(N__33957),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_3 ));
    CascadeMux I__3117 (
            .O(N__33952),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12998_cascade_ ));
    CascadeMux I__3116 (
            .O(N__33949),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13001_cascade_ ));
    CascadeMux I__3115 (
            .O(N__33946),
            .I(N__33942));
    CascadeMux I__3114 (
            .O(N__33945),
            .I(N__33939));
    InMux I__3113 (
            .O(N__33942),
            .I(N__33934));
    InMux I__3112 (
            .O(N__33939),
            .I(N__33934));
    LocalMux I__3111 (
            .O(N__33934),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_3 ));
    CascadeMux I__3110 (
            .O(N__33931),
            .I(N__33928));
    InMux I__3109 (
            .O(N__33928),
            .I(N__33925));
    LocalMux I__3108 (
            .O(N__33925),
            .I(N__33922));
    Span4Mux_v I__3107 (
            .O(N__33922),
            .I(N__33918));
    InMux I__3106 (
            .O(N__33921),
            .I(N__33915));
    Odrv4 I__3105 (
            .O(N__33918),
            .I(REG_mem_26_14));
    LocalMux I__3104 (
            .O(N__33915),
            .I(REG_mem_26_14));
    InMux I__3103 (
            .O(N__33910),
            .I(N__33907));
    LocalMux I__3102 (
            .O(N__33907),
            .I(N__33904));
    Span4Mux_v I__3101 (
            .O(N__33904),
            .I(N__33901));
    Odrv4 I__3100 (
            .O(N__33901),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12355 ));
    InMux I__3099 (
            .O(N__33898),
            .I(N__33895));
    LocalMux I__3098 (
            .O(N__33895),
            .I(N__33892));
    Span4Mux_v I__3097 (
            .O(N__33892),
            .I(N__33889));
    Odrv4 I__3096 (
            .O(N__33889),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13196 ));
    CascadeMux I__3095 (
            .O(N__33886),
            .I(N__33882));
    InMux I__3094 (
            .O(N__33885),
            .I(N__33877));
    InMux I__3093 (
            .O(N__33882),
            .I(N__33877));
    LocalMux I__3092 (
            .O(N__33877),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_3 ));
    CascadeMux I__3091 (
            .O(N__33874),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14264_cascade_ ));
    CascadeMux I__3090 (
            .O(N__33871),
            .I(N__33867));
    CascadeMux I__3089 (
            .O(N__33870),
            .I(N__33864));
    InMux I__3088 (
            .O(N__33867),
            .I(N__33859));
    InMux I__3087 (
            .O(N__33864),
            .I(N__33859));
    LocalMux I__3086 (
            .O(N__33859),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_10 ));
    InMux I__3085 (
            .O(N__33856),
            .I(N__33853));
    LocalMux I__3084 (
            .O(N__33853),
            .I(N__33850));
    Odrv4 I__3083 (
            .O(N__33850),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12965 ));
    InMux I__3082 (
            .O(N__33847),
            .I(N__33844));
    LocalMux I__3081 (
            .O(N__33844),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11635 ));
    InMux I__3080 (
            .O(N__33841),
            .I(N__33838));
    LocalMux I__3079 (
            .O(N__33838),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11548 ));
    InMux I__3078 (
            .O(N__33835),
            .I(N__33832));
    LocalMux I__3077 (
            .O(N__33832),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13262 ));
    InMux I__3076 (
            .O(N__33829),
            .I(N__33826));
    LocalMux I__3075 (
            .O(N__33826),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11546 ));
    InMux I__3074 (
            .O(N__33823),
            .I(N__33817));
    InMux I__3073 (
            .O(N__33822),
            .I(N__33817));
    LocalMux I__3072 (
            .O(N__33817),
            .I(REG_mem_18_10));
    InMux I__3071 (
            .O(N__33814),
            .I(N__33808));
    InMux I__3070 (
            .O(N__33813),
            .I(N__33808));
    LocalMux I__3069 (
            .O(N__33808),
            .I(REG_mem_19_10));
    InMux I__3068 (
            .O(N__33805),
            .I(N__33802));
    LocalMux I__3067 (
            .O(N__33802),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14228 ));
    InMux I__3066 (
            .O(N__33799),
            .I(N__33796));
    LocalMux I__3065 (
            .O(N__33796),
            .I(N__33793));
    Span4Mux_h I__3064 (
            .O(N__33793),
            .I(N__33790));
    Odrv4 I__3063 (
            .O(N__33790),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11528 ));
    InMux I__3062 (
            .O(N__33787),
            .I(N__33784));
    LocalMux I__3061 (
            .O(N__33784),
            .I(N__33781));
    Span4Mux_v I__3060 (
            .O(N__33781),
            .I(N__33777));
    InMux I__3059 (
            .O(N__33780),
            .I(N__33774));
    Odrv4 I__3058 (
            .O(N__33777),
            .I(REG_mem_58_14));
    LocalMux I__3057 (
            .O(N__33774),
            .I(REG_mem_58_14));
    InMux I__3056 (
            .O(N__33769),
            .I(N__33763));
    InMux I__3055 (
            .O(N__33768),
            .I(N__33763));
    LocalMux I__3054 (
            .O(N__33763),
            .I(REG_mem_37_14));
    CascadeMux I__3053 (
            .O(N__33760),
            .I(N__33756));
    InMux I__3052 (
            .O(N__33759),
            .I(N__33751));
    InMux I__3051 (
            .O(N__33756),
            .I(N__33751));
    LocalMux I__3050 (
            .O(N__33751),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_14 ));
    InMux I__3049 (
            .O(N__33748),
            .I(N__33742));
    InMux I__3048 (
            .O(N__33747),
            .I(N__33742));
    LocalMux I__3047 (
            .O(N__33742),
            .I(REG_mem_31_10));
    CascadeMux I__3046 (
            .O(N__33739),
            .I(N__33735));
    CascadeMux I__3045 (
            .O(N__33738),
            .I(N__33732));
    InMux I__3044 (
            .O(N__33735),
            .I(N__33729));
    InMux I__3043 (
            .O(N__33732),
            .I(N__33726));
    LocalMux I__3042 (
            .O(N__33729),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_10 ));
    LocalMux I__3041 (
            .O(N__33726),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_10 ));
    CascadeMux I__3040 (
            .O(N__33721),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13898_cascade_ ));
    CascadeMux I__3039 (
            .O(N__33718),
            .I(N__33714));
    InMux I__3038 (
            .O(N__33717),
            .I(N__33711));
    InMux I__3037 (
            .O(N__33714),
            .I(N__33708));
    LocalMux I__3036 (
            .O(N__33711),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_10 ));
    LocalMux I__3035 (
            .O(N__33708),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_10 ));
    InMux I__3034 (
            .O(N__33703),
            .I(N__33700));
    LocalMux I__3033 (
            .O(N__33700),
            .I(N__33697));
    Odrv4 I__3032 (
            .O(N__33697),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13901 ));
    CascadeMux I__3031 (
            .O(N__33694),
            .I(N__33690));
    InMux I__3030 (
            .O(N__33693),
            .I(N__33685));
    InMux I__3029 (
            .O(N__33690),
            .I(N__33685));
    LocalMux I__3028 (
            .O(N__33685),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_10 ));
    InMux I__3027 (
            .O(N__33682),
            .I(N__33679));
    LocalMux I__3026 (
            .O(N__33679),
            .I(N__33676));
    Odrv4 I__3025 (
            .O(N__33676),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11527 ));
    InMux I__3024 (
            .O(N__33673),
            .I(N__33669));
    InMux I__3023 (
            .O(N__33672),
            .I(N__33666));
    LocalMux I__3022 (
            .O(N__33669),
            .I(REG_mem_16_10));
    LocalMux I__3021 (
            .O(N__33666),
            .I(REG_mem_16_10));
    InMux I__3020 (
            .O(N__33661),
            .I(N__33657));
    InMux I__3019 (
            .O(N__33660),
            .I(N__33654));
    LocalMux I__3018 (
            .O(N__33657),
            .I(REG_mem_55_14));
    LocalMux I__3017 (
            .O(N__33654),
            .I(REG_mem_55_14));
    CascadeMux I__3016 (
            .O(N__33649),
            .I(N__33645));
    InMux I__3015 (
            .O(N__33648),
            .I(N__33640));
    InMux I__3014 (
            .O(N__33645),
            .I(N__33640));
    LocalMux I__3013 (
            .O(N__33640),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_14 ));
    InMux I__3012 (
            .O(N__33637),
            .I(N__33631));
    InMux I__3011 (
            .O(N__33636),
            .I(N__33631));
    LocalMux I__3010 (
            .O(N__33631),
            .I(REG_mem_48_14));
    InMux I__3009 (
            .O(N__33628),
            .I(N__33625));
    LocalMux I__3008 (
            .O(N__33625),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12332 ));
    InMux I__3007 (
            .O(N__33622),
            .I(N__33619));
    LocalMux I__3006 (
            .O(N__33619),
            .I(N__33615));
    CascadeMux I__3005 (
            .O(N__33618),
            .I(N__33612));
    Span4Mux_h I__3004 (
            .O(N__33615),
            .I(N__33609));
    InMux I__3003 (
            .O(N__33612),
            .I(N__33606));
    Odrv4 I__3002 (
            .O(N__33609),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_14 ));
    LocalMux I__3001 (
            .O(N__33606),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_14 ));
    CascadeMux I__3000 (
            .O(N__33601),
            .I(N__33598));
    InMux I__2999 (
            .O(N__33598),
            .I(N__33595));
    LocalMux I__2998 (
            .O(N__33595),
            .I(N__33592));
    Odrv4 I__2997 (
            .O(N__33592),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12331 ));
    CascadeMux I__2996 (
            .O(N__33589),
            .I(N__33586));
    InMux I__2995 (
            .O(N__33586),
            .I(N__33582));
    CascadeMux I__2994 (
            .O(N__33585),
            .I(N__33579));
    LocalMux I__2993 (
            .O(N__33582),
            .I(N__33576));
    InMux I__2992 (
            .O(N__33579),
            .I(N__33573));
    Odrv4 I__2991 (
            .O(N__33576),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_10 ));
    LocalMux I__2990 (
            .O(N__33573),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_10 ));
    InMux I__2989 (
            .O(N__33568),
            .I(N__33564));
    InMux I__2988 (
            .O(N__33567),
            .I(N__33561));
    LocalMux I__2987 (
            .O(N__33564),
            .I(REG_mem_36_14));
    LocalMux I__2986 (
            .O(N__33561),
            .I(REG_mem_36_14));
    CascadeMux I__2985 (
            .O(N__33556),
            .I(N__33552));
    InMux I__2984 (
            .O(N__33555),
            .I(N__33547));
    InMux I__2983 (
            .O(N__33552),
            .I(N__33547));
    LocalMux I__2982 (
            .O(N__33547),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_14 ));
    CascadeMux I__2981 (
            .O(N__33544),
            .I(N__33540));
    InMux I__2980 (
            .O(N__33543),
            .I(N__33535));
    InMux I__2979 (
            .O(N__33540),
            .I(N__33535));
    LocalMux I__2978 (
            .O(N__33535),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_14 ));
    CascadeMux I__2977 (
            .O(N__33532),
            .I(N__33528));
    CascadeMux I__2976 (
            .O(N__33531),
            .I(N__33525));
    InMux I__2975 (
            .O(N__33528),
            .I(N__33522));
    InMux I__2974 (
            .O(N__33525),
            .I(N__33519));
    LocalMux I__2973 (
            .O(N__33522),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_14 ));
    LocalMux I__2972 (
            .O(N__33519),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_14 ));
    CascadeMux I__2971 (
            .O(N__33514),
            .I(N__33510));
    InMux I__2970 (
            .O(N__33513),
            .I(N__33507));
    InMux I__2969 (
            .O(N__33510),
            .I(N__33504));
    LocalMux I__2968 (
            .O(N__33507),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_14 ));
    LocalMux I__2967 (
            .O(N__33504),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_14 ));
    CascadeMux I__2966 (
            .O(N__33499),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12977_cascade_ ));
    InMux I__2965 (
            .O(N__33496),
            .I(N__33493));
    LocalMux I__2964 (
            .O(N__33493),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11572 ));
    CascadeMux I__2963 (
            .O(N__33490),
            .I(N__33487));
    InMux I__2962 (
            .O(N__33487),
            .I(N__33484));
    LocalMux I__2961 (
            .O(N__33484),
            .I(N__33480));
    InMux I__2960 (
            .O(N__33483),
            .I(N__33477));
    Odrv12 I__2959 (
            .O(N__33480),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_14 ));
    LocalMux I__2958 (
            .O(N__33477),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_14 ));
    CascadeMux I__2957 (
            .O(N__33472),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12866_cascade_ ));
    InMux I__2956 (
            .O(N__33469),
            .I(N__33466));
    LocalMux I__2955 (
            .O(N__33466),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12869 ));
    InMux I__2954 (
            .O(N__33463),
            .I(N__33460));
    LocalMux I__2953 (
            .O(N__33460),
            .I(N__33456));
    CascadeMux I__2952 (
            .O(N__33459),
            .I(N__33453));
    Span4Mux_v I__2951 (
            .O(N__33456),
            .I(N__33450));
    InMux I__2950 (
            .O(N__33453),
            .I(N__33447));
    Odrv4 I__2949 (
            .O(N__33450),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_10 ));
    LocalMux I__2948 (
            .O(N__33447),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_10 ));
    CascadeMux I__2947 (
            .O(N__33442),
            .I(N__33439));
    InMux I__2946 (
            .O(N__33439),
            .I(N__33435));
    CascadeMux I__2945 (
            .O(N__33438),
            .I(N__33432));
    LocalMux I__2944 (
            .O(N__33435),
            .I(N__33429));
    InMux I__2943 (
            .O(N__33432),
            .I(N__33426));
    Odrv4 I__2942 (
            .O(N__33429),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_14 ));
    LocalMux I__2941 (
            .O(N__33426),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_14 ));
    InMux I__2940 (
            .O(N__33421),
            .I(N__33417));
    InMux I__2939 (
            .O(N__33420),
            .I(N__33414));
    LocalMux I__2938 (
            .O(N__33417),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_14 ));
    LocalMux I__2937 (
            .O(N__33414),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_14 ));
    InMux I__2936 (
            .O(N__33409),
            .I(N__33406));
    LocalMux I__2935 (
            .O(N__33406),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14270 ));
    CascadeMux I__2934 (
            .O(N__33403),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13328_cascade_ ));
    CascadeMux I__2933 (
            .O(N__33400),
            .I(N__33396));
    InMux I__2932 (
            .O(N__33399),
            .I(N__33391));
    InMux I__2931 (
            .O(N__33396),
            .I(N__33391));
    LocalMux I__2930 (
            .O(N__33391),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_14 ));
    InMux I__2929 (
            .O(N__33388),
            .I(N__33385));
    LocalMux I__2928 (
            .O(N__33385),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12776 ));
    CascadeMux I__2927 (
            .O(N__33382),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14384_cascade_ ));
    CascadeMux I__2926 (
            .O(N__33379),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14387_cascade_ ));
    InMux I__2925 (
            .O(N__33376),
            .I(N__33373));
    LocalMux I__2924 (
            .O(N__33373),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12779 ));
    CascadeMux I__2923 (
            .O(N__33370),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12071_cascade_ ));
    CascadeMux I__2922 (
            .O(N__33367),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13688_cascade_ ));
    CascadeMux I__2921 (
            .O(N__33364),
            .I(N__33361));
    InMux I__2920 (
            .O(N__33361),
            .I(N__33355));
    InMux I__2919 (
            .O(N__33360),
            .I(N__33355));
    LocalMux I__2918 (
            .O(N__33355),
            .I(REG_mem_23_14));
    CascadeMux I__2917 (
            .O(N__33352),
            .I(N__33348));
    InMux I__2916 (
            .O(N__33351),
            .I(N__33343));
    InMux I__2915 (
            .O(N__33348),
            .I(N__33343));
    LocalMux I__2914 (
            .O(N__33343),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_14 ));
    InMux I__2913 (
            .O(N__33340),
            .I(N__33337));
    LocalMux I__2912 (
            .O(N__33337),
            .I(N__33333));
    InMux I__2911 (
            .O(N__33336),
            .I(N__33330));
    Odrv12 I__2910 (
            .O(N__33333),
            .I(REG_mem_58_10));
    LocalMux I__2909 (
            .O(N__33330),
            .I(REG_mem_58_10));
    CascadeMux I__2908 (
            .O(N__33325),
            .I(N__33321));
    InMux I__2907 (
            .O(N__33324),
            .I(N__33316));
    InMux I__2906 (
            .O(N__33321),
            .I(N__33316));
    LocalMux I__2905 (
            .O(N__33316),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_10 ));
    InMux I__2904 (
            .O(N__33313),
            .I(N__33310));
    LocalMux I__2903 (
            .O(N__33310),
            .I(N__33307));
    Odrv12 I__2902 (
            .O(N__33307),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11524 ));
    CascadeMux I__2901 (
            .O(N__33304),
            .I(N__33301));
    InMux I__2900 (
            .O(N__33301),
            .I(N__33295));
    InMux I__2899 (
            .O(N__33300),
            .I(N__33295));
    LocalMux I__2898 (
            .O(N__33295),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_10 ));
    InMux I__2897 (
            .O(N__33292),
            .I(N__33286));
    InMux I__2896 (
            .O(N__33291),
            .I(N__33286));
    LocalMux I__2895 (
            .O(N__33286),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_10 ));
    CascadeMux I__2894 (
            .O(N__33283),
            .I(N__33279));
    InMux I__2893 (
            .O(N__33282),
            .I(N__33274));
    InMux I__2892 (
            .O(N__33279),
            .I(N__33274));
    LocalMux I__2891 (
            .O(N__33274),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_10 ));
    CascadeMux I__2890 (
            .O(N__33271),
            .I(N__33267));
    InMux I__2889 (
            .O(N__33270),
            .I(N__33264));
    InMux I__2888 (
            .O(N__33267),
            .I(N__33261));
    LocalMux I__2887 (
            .O(N__33264),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_10 ));
    LocalMux I__2886 (
            .O(N__33261),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_10 ));
    CascadeMux I__2885 (
            .O(N__33256),
            .I(N__33252));
    CascadeMux I__2884 (
            .O(N__33255),
            .I(N__33249));
    InMux I__2883 (
            .O(N__33252),
            .I(N__33244));
    InMux I__2882 (
            .O(N__33249),
            .I(N__33244));
    LocalMux I__2881 (
            .O(N__33244),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_10 ));
    CascadeMux I__2880 (
            .O(N__33241),
            .I(N__33237));
    InMux I__2879 (
            .O(N__33240),
            .I(N__33232));
    InMux I__2878 (
            .O(N__33237),
            .I(N__33232));
    LocalMux I__2877 (
            .O(N__33232),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_10 ));
    InMux I__2876 (
            .O(N__33229),
            .I(N__33226));
    LocalMux I__2875 (
            .O(N__33226),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14048 ));
    CascadeMux I__2874 (
            .O(N__33223),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14036_cascade_ ));
    CascadeMux I__2873 (
            .O(N__33220),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12129_cascade_ ));
    InMux I__2872 (
            .O(N__33217),
            .I(N__33214));
    LocalMux I__2871 (
            .O(N__33214),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12126 ));
    InMux I__2870 (
            .O(N__33211),
            .I(N__33205));
    InMux I__2869 (
            .O(N__33210),
            .I(N__33205));
    LocalMux I__2868 (
            .O(N__33205),
            .I(REG_mem_13_7));
    InMux I__2867 (
            .O(N__33202),
            .I(N__33196));
    InMux I__2866 (
            .O(N__33201),
            .I(N__33196));
    LocalMux I__2865 (
            .O(N__33196),
            .I(REG_mem_26_10));
    InMux I__2864 (
            .O(N__33193),
            .I(N__33190));
    LocalMux I__2863 (
            .O(N__33190),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11545 ));
    CascadeMux I__2862 (
            .O(N__33187),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13265_cascade_ ));
    InMux I__2861 (
            .O(N__33184),
            .I(N__33181));
    LocalMux I__2860 (
            .O(N__33181),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11621 ));
    CascadeMux I__2859 (
            .O(N__33178),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13298_cascade_ ));
    InMux I__2858 (
            .O(N__33175),
            .I(N__33172));
    LocalMux I__2857 (
            .O(N__33172),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13259 ));
    InMux I__2856 (
            .O(N__33169),
            .I(N__33166));
    LocalMux I__2855 (
            .O(N__33166),
            .I(N__33163));
    Odrv4 I__2854 (
            .O(N__33163),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14006 ));
    CascadeMux I__2853 (
            .O(N__33160),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14009_cascade_ ));
    InMux I__2852 (
            .O(N__33157),
            .I(N__33154));
    LocalMux I__2851 (
            .O(N__33154),
            .I(N__33151));
    Odrv4 I__2850 (
            .O(N__33151),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11627 ));
    InMux I__2849 (
            .O(N__33148),
            .I(N__33145));
    LocalMux I__2848 (
            .O(N__33145),
            .I(N__33142));
    Odrv12 I__2847 (
            .O(N__33142),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12914 ));
    InMux I__2846 (
            .O(N__33139),
            .I(N__33136));
    LocalMux I__2845 (
            .O(N__33136),
            .I(N__33133));
    Span4Mux_v I__2844 (
            .O(N__33133),
            .I(N__33130));
    Odrv4 I__2843 (
            .O(N__33130),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12917 ));
    CascadeMux I__2842 (
            .O(N__33127),
            .I(N__33123));
    InMux I__2841 (
            .O(N__33126),
            .I(N__33118));
    InMux I__2840 (
            .O(N__33123),
            .I(N__33118));
    LocalMux I__2839 (
            .O(N__33118),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_10 ));
    CascadeMux I__2838 (
            .O(N__33115),
            .I(N__33111));
    CascadeMux I__2837 (
            .O(N__33114),
            .I(N__33108));
    InMux I__2836 (
            .O(N__33111),
            .I(N__33103));
    InMux I__2835 (
            .O(N__33108),
            .I(N__33103));
    LocalMux I__2834 (
            .O(N__33103),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_10 ));
    CascadeMux I__2833 (
            .O(N__33100),
            .I(N__33097));
    InMux I__2832 (
            .O(N__33097),
            .I(N__33094));
    LocalMux I__2831 (
            .O(N__33094),
            .I(N__33091));
    Odrv4 I__2830 (
            .O(N__33091),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13256 ));
    CascadeMux I__2829 (
            .O(N__33088),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12842_cascade_ ));
    CascadeMux I__2828 (
            .O(N__33085),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12845_cascade_ ));
    CascadeMux I__2827 (
            .O(N__33082),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11636_cascade_ ));
    CascadeMux I__2826 (
            .O(N__33079),
            .I(N__33075));
    InMux I__2825 (
            .O(N__33078),
            .I(N__33072));
    InMux I__2824 (
            .O(N__33075),
            .I(N__33069));
    LocalMux I__2823 (
            .O(N__33072),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_10 ));
    LocalMux I__2822 (
            .O(N__33069),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_10 ));
    CascadeMux I__2821 (
            .O(N__33064),
            .I(N__33060));
    CascadeMux I__2820 (
            .O(N__33063),
            .I(N__33057));
    InMux I__2819 (
            .O(N__33060),
            .I(N__33054));
    InMux I__2818 (
            .O(N__33057),
            .I(N__33051));
    LocalMux I__2817 (
            .O(N__33054),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_14 ));
    LocalMux I__2816 (
            .O(N__33051),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_14 ));
    CascadeMux I__2815 (
            .O(N__33046),
            .I(N__33042));
    InMux I__2814 (
            .O(N__33045),
            .I(N__33037));
    InMux I__2813 (
            .O(N__33042),
            .I(N__33037));
    LocalMux I__2812 (
            .O(N__33037),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_9 ));
    CascadeMux I__2811 (
            .O(N__33034),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12956_cascade_ ));
    CascadeMux I__2810 (
            .O(N__33031),
            .I(N__33027));
    InMux I__2809 (
            .O(N__33030),
            .I(N__33022));
    InMux I__2808 (
            .O(N__33027),
            .I(N__33022));
    LocalMux I__2807 (
            .O(N__33022),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_9 ));
    CascadeMux I__2806 (
            .O(N__33019),
            .I(N__33015));
    CascadeMux I__2805 (
            .O(N__33018),
            .I(N__33012));
    InMux I__2804 (
            .O(N__33015),
            .I(N__33007));
    InMux I__2803 (
            .O(N__33012),
            .I(N__33007));
    LocalMux I__2802 (
            .O(N__33007),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_9 ));
    InMux I__2801 (
            .O(N__33004),
            .I(N__33001));
    LocalMux I__2800 (
            .O(N__33001),
            .I(N__32998));
    Odrv4 I__2799 (
            .O(N__32998),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13199 ));
    InMux I__2798 (
            .O(N__32995),
            .I(N__32992));
    LocalMux I__2797 (
            .O(N__32992),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12839 ));
    CascadeMux I__2796 (
            .O(N__32989),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11573_cascade_ ));
    InMux I__2795 (
            .O(N__32986),
            .I(N__32983));
    LocalMux I__2794 (
            .O(N__32983),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11543 ));
    CascadeMux I__2793 (
            .O(N__32980),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13628_cascade_ ));
    CascadeMux I__2792 (
            .O(N__32977),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13472_cascade_ ));
    CascadeMux I__2791 (
            .O(N__32974),
            .I(N__32970));
    InMux I__2790 (
            .O(N__32973),
            .I(N__32965));
    InMux I__2789 (
            .O(N__32970),
            .I(N__32965));
    LocalMux I__2788 (
            .O(N__32965),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_14 ));
    CascadeMux I__2787 (
            .O(N__32962),
            .I(N__32958));
    InMux I__2786 (
            .O(N__32961),
            .I(N__32953));
    InMux I__2785 (
            .O(N__32958),
            .I(N__32953));
    LocalMux I__2784 (
            .O(N__32953),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_14 ));
    CascadeMux I__2783 (
            .O(N__32950),
            .I(N__32946));
    InMux I__2782 (
            .O(N__32949),
            .I(N__32941));
    InMux I__2781 (
            .O(N__32946),
            .I(N__32941));
    LocalMux I__2780 (
            .O(N__32941),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_14 ));
    CascadeMux I__2779 (
            .O(N__32938),
            .I(N__32934));
    InMux I__2778 (
            .O(N__32937),
            .I(N__32931));
    InMux I__2777 (
            .O(N__32934),
            .I(N__32928));
    LocalMux I__2776 (
            .O(N__32931),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_14 ));
    LocalMux I__2775 (
            .O(N__32928),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_14 ));
    InMux I__2774 (
            .O(N__32923),
            .I(N__32920));
    LocalMux I__2773 (
            .O(N__32920),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12836 ));
    CascadeMux I__2772 (
            .O(N__32917),
            .I(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14273_cascade_ ));
    IoInMux I__2771 (
            .O(N__32914),
            .I(N__32911));
    LocalMux I__2770 (
            .O(N__32911),
            .I(N__32908));
    Span4Mux_s0_v I__2769 (
            .O(N__32908),
            .I(N__32905));
    Span4Mux_v I__2768 (
            .O(N__32905),
            .I(N__32902));
    Sp12to4 I__2767 (
            .O(N__32902),
            .I(N__32899));
    Span12Mux_h I__2766 (
            .O(N__32899),
            .I(N__32896));
    Span12Mux_v I__2765 (
            .O(N__32896),
            .I(N__32893));
    Odrv12 I__2764 (
            .O(N__32893),
            .I(ICE_SYSCLK_c));
    INV \INVbluejay_data_inst.bluejay_data_out_i14C  (
            .O(\INVbluejay_data_inst.bluejay_data_out_i14C_net ),
            .I(N__97391));
    INV \INVusb3_if_inst.dc32_fifo_data_in_i9C  (
            .O(\INVusb3_if_inst.dc32_fifo_data_in_i9C_net ),
            .I(N__93452));
    INV \INVbluejay_data_inst.bluejay_data_out_i9C  (
            .O(\INVbluejay_data_inst.bluejay_data_out_i9C_net ),
            .I(N__97427));
    INV \INVusb3_if_inst.state_FSM_i3C  (
            .O(\INVusb3_if_inst.state_FSM_i3C_net ),
            .I(N__93404));
    INV \INVusb3_if_inst.dc32_fifo_data_in_i2C  (
            .O(\INVusb3_if_inst.dc32_fifo_data_in_i2C_net ),
            .I(N__93447));
    INV \INVbluejay_data_inst.bluejay_data_out_i16C  (
            .O(\INVbluejay_data_inst.bluejay_data_out_i16C_net ),
            .I(N__97367));
    INV \INVusb3_if_inst.state_FSM_i2C  (
            .O(\INVusb3_if_inst.state_FSM_i2C_net ),
            .I(N__93377));
    INV \INVusb3_if_inst.num_lines_clocked_out_i8C  (
            .O(\INVusb3_if_inst.num_lines_clocked_out_i8C_net ),
            .I(N__93388));
    INV \INVusb3_if_inst.num_lines_clocked_out_i0C  (
            .O(\INVusb3_if_inst.num_lines_clocked_out_i0C_net ),
            .I(N__93375));
    INV \INVusb3_if_inst.state_timeout_counter_i0_i3C  (
            .O(\INVusb3_if_inst.state_timeout_counter_i0_i3C_net ),
            .I(N__93362));
    INV \INVusb3_if_inst.state_timeout_counter_i0_i1C  (
            .O(\INVusb3_if_inst.state_timeout_counter_i0_i1C_net ),
            .I(N__93346));
    INV \INVusb3_if_inst.FT_RD_internal_75C  (
            .O(\INVusb3_if_inst.FT_RD_internal_75C_net ),
            .I(N__93315));
    INV \INVusb3_if_inst.state_timeout_counter_i0_i2C  (
            .O(\INVusb3_if_inst.state_timeout_counter_i0_i2C_net ),
            .I(N__93288));
    INV \INVusb3_if_inst.state_FSM_i5C  (
            .O(\INVusb3_if_inst.state_FSM_i5C_net ),
            .I(N__93322));
    INV \INVusb3_if_inst.dc32_fifo_data_in_i16C  (
            .O(\INVusb3_if_inst.dc32_fifo_data_in_i16C_net ),
            .I(N__93320));
    INV \INVusb3_if_inst.dc32_fifo_data_in_i15C  (
            .O(\INVusb3_if_inst.dc32_fifo_data_in_i15C_net ),
            .I(N__93277));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\usb3_if_inst.n10667 ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_23_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_13_0_));
    defparam IN_MUX_bfv_23_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_14_0_ (
            .carryinitin(\timing_controller_inst.n10595 ),
            .carryinitout(bfn_23_14_0_));
    defparam IN_MUX_bfv_23_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_15_0_ (
            .carryinitin(\timing_controller_inst.n10603 ),
            .carryinitout(bfn_23_15_0_));
    defparam IN_MUX_bfv_23_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_16_0_ (
            .carryinitin(\timing_controller_inst.n10611 ),
            .carryinitout(bfn_23_16_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(\spi0.n10701 ),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_24_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_11_0_));
    defparam IN_MUX_bfv_24_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_12_0_ (
            .carryinitin(\pc_tx.n10719 ),
            .carryinitout(bfn_24_12_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(\pc_rx.n10710 ),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_23_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_5_0_));
    defparam IN_MUX_bfv_23_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_6_0_ (
            .carryinitin(n10677),
            .carryinitout(bfn_23_6_0_));
    defparam IN_MUX_bfv_23_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_7_0_ (
            .carryinitin(n10685),
            .carryinitout(bfn_23_7_0_));
    defparam IN_MUX_bfv_23_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_8_0_ (
            .carryinitin(n10693),
            .carryinitout(bfn_23_8_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(\bluejay_data_inst.n10650 ),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(\bluejay_data_inst.n10583_THRU_CRY_4_THRU_CO ),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(\bluejay_data_inst.n10584_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_16_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_14_0_ (
            .carryinitin(\bluejay_data_inst.n10585_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_16_14_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(\bluejay_data_inst.n10586_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_16_15_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB clk_gb (
            .USERSIGNALTOGLOBALBUFFER(N__37552),
            .GLOBALBUFFEROUTPUT(SLM_CLK_c));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12836_bdd_4_lut_LC_1_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12836_bdd_4_lut_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12836_bdd_4_lut_LC_1_7_0 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12836_bdd_4_lut_LC_1_7_0  (
            .in0(N__92563),
            .in1(N__32923),
            .in2(N__33064),
            .in3(N__32937),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12839 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9894_3_lut_LC_1_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9894_3_lut_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9894_3_lut_LC_1_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9894_3_lut_LC_1_7_1  (
            .in0(N__85816),
            .in1(N__34330),
            .in2(_gnd_net_),
            .in3(N__34309),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11181_LC_1_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11181_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11181_LC_1_7_2 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11181_LC_1_7_2  (
            .in0(N__92565),
            .in1(N__88811),
            .in2(N__33442),
            .in3(N__33787),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12836 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14270_bdd_4_lut_LC_1_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14270_bdd_4_lut_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14270_bdd_4_lut_LC_1_7_3 .LUT_INIT=16'b1011101010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14270_bdd_4_lut_LC_1_7_3  (
            .in0(N__33409),
            .in1(N__92564),
            .in2(N__33532),
            .in3(N__33513),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14273_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9924_3_lut_LC_1_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9924_3_lut_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9924_3_lut_LC_1_7_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9924_3_lut_LC_1_7_4  (
            .in0(_gnd_net_),
            .in1(N__85817),
            .in2(N__32917),
            .in3(N__32995),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11573_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11884_LC_1_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11884_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11884_LC_1_7_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11884_LC_1_7_5  (
            .in0(N__33496),
            .in1(N__81467),
            .in2(N__32989),
            .in3(N__90341),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13628_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13628_bdd_4_lut_LC_1_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13628_bdd_4_lut_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13628_bdd_4_lut_LC_1_7_6 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13628_bdd_4_lut_LC_1_7_6  (
            .in0(N__81466),
            .in1(N__32986),
            .in2(N__32980),
            .in3(N__33004),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13631 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11530_LC_1_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11530_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11530_LC_1_8_0 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11530_LC_1_8_0  (
            .in0(N__33682),
            .in1(N__33799),
            .in2(N__85568),
            .in3(N__92562),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13256 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11729_LC_1_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11729_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11729_LC_1_8_1 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11729_LC_1_8_1  (
            .in0(N__32949),
            .in1(N__92599),
            .in2(N__33931),
            .in3(N__88241),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13472_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13472_bdd_4_lut_LC_1_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13472_bdd_4_lut_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13472_bdd_4_lut_LC_1_8_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13472_bdd_4_lut_LC_1_8_2  (
            .in0(N__32961),
            .in1(N__92561),
            .in2(N__32977),
            .in3(N__32973),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13475 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2480_2481_LC_1_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2480_2481_LC_1_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2480_2481_LC_1_8_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2480_2481_LC_1_8_3  (
            .in0(N__41767),
            .in1(N__95369),
            .in2(N__32974),
            .in3(N__96942),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93223),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2384_2385_LC_1_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2384_2385_LC_1_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2384_2385_LC_1_8_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2384_2385_LC_1_8_4  (
            .in0(N__95367),
            .in1(N__41766),
            .in2(N__32962),
            .in3(N__96008),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93223),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2672_2673_LC_1_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2672_2673_LC_1_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2672_2673_LC_1_8_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2672_2673_LC_1_8_5  (
            .in0(N__41768),
            .in1(N__95370),
            .in2(N__32950),
            .in3(N__79742),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93223),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5456_5457_LC_1_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5456_5457_LC_1_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5456_5457_LC_1_8_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5456_5457_LC_1_8_6  (
            .in0(N__95368),
            .in1(N__41769),
            .in2(N__32938),
            .in3(N__96009),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93223),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5552_5553_LC_1_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5552_5553_LC_1_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5552_5553_LC_1_8_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5552_5553_LC_1_8_7  (
            .in0(N__41770),
            .in1(N__95371),
            .in2(N__33063),
            .in3(N__96943),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93223),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3233_3234_LC_1_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3233_3234_LC_1_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3233_3234_LC_1_9_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3233_3234_LC_1_9_0  (
            .in0(N__95379),
            .in1(N__56548),
            .in2(N__33046),
            .in3(N__80313),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11281_LC_1_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11281_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11281_LC_1_9_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11281_LC_1_9_1  (
            .in0(N__92211),
            .in1(N__88032),
            .in2(N__33019),
            .in3(N__34654),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12956_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12956_bdd_4_lut_LC_1_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12956_bdd_4_lut_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12956_bdd_4_lut_LC_1_9_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12956_bdd_4_lut_LC_1_9_2  (
            .in0(N__33045),
            .in1(N__92210),
            .in2(N__33034),
            .in3(N__33030),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12959 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3137_3138_LC_1_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3137_3138_LC_1_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3137_3138_LC_1_9_3 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3137_3138_LC_1_9_3  (
            .in0(N__56546),
            .in1(N__95380),
            .in2(N__33031),
            .in3(N__82950),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2948_2949_LC_1_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2948_2949_LC_1_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2948_2949_LC_1_9_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2948_2949_LC_1_9_4  (
            .in0(N__95378),
            .in1(N__48812),
            .in2(N__33738),
            .in3(N__77936),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3425_3426_LC_1_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3425_3426_LC_1_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3425_3426_LC_1_9_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3425_3426_LC_1_9_5  (
            .in0(N__56547),
            .in1(N__95381),
            .in2(N__33018),
            .in3(N__83298),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13196_bdd_4_lut_LC_1_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13196_bdd_4_lut_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13196_bdd_4_lut_LC_1_9_6 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13196_bdd_4_lut_LC_1_9_6  (
            .in0(N__33628),
            .in1(N__85625),
            .in2(N__33601),
            .in3(N__33898),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5060_5061_LC_1_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5060_5061_LC_1_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5060_5061_LC_1_9_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5060_5061_LC_1_9_7  (
            .in0(N__48813),
            .in1(N__95382),
            .in2(N__33585),
            .in3(N__77443),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93220),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13256_bdd_4_lut_LC_1_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13256_bdd_4_lut_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13256_bdd_4_lut_LC_1_10_0 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13256_bdd_4_lut_LC_1_10_0  (
            .in0(N__85624),
            .in1(N__33313),
            .in2(N__33100),
            .in3(N__34243),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11246_LC_1_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11246_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11246_LC_1_10_1 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11246_LC_1_10_1  (
            .in0(N__88240),
            .in1(N__92318),
            .in2(N__36583),
            .in3(N__33340),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12914 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11186_LC_1_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11186_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11186_LC_1_10_2 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11186_LC_1_10_2  (
            .in0(N__92317),
            .in1(N__33463),
            .in2(N__45394),
            .in3(N__88239),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12842_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12842_bdd_4_lut_LC_1_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12842_bdd_4_lut_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12842_bdd_4_lut_LC_1_10_3 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12842_bdd_4_lut_LC_1_10_3  (
            .in0(N__33078),
            .in1(N__92316),
            .in2(N__33088),
            .in3(N__34276),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12845_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9987_3_lut_LC_1_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9987_3_lut_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9987_3_lut_LC_1_10_4 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9987_3_lut_LC_1_10_4  (
            .in0(N__85623),
            .in1(N__33139),
            .in2(N__33085),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11636_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12358_LC_1_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12358_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12358_LC_1_10_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12358_LC_1_10_5  (
            .in0(N__33847),
            .in1(N__81472),
            .in2(N__33082),
            .in3(N__90340),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9896_3_lut_LC_1_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9896_3_lut_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9896_3_lut_LC_1_10_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9896_3_lut_LC_1_10_6  (
            .in0(N__38512),
            .in1(N__88238),
            .in2(_gnd_net_),
            .in3(N__33673),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5828_5829_LC_1_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5828_5829_LC_1_11_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5828_5829_LC_1_11_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5828_5829_LC_1_11_0  (
            .in0(N__48866),
            .in1(N__94221),
            .in2(N__33079),
            .in3(N__70715),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93221),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2564_2565_LC_1_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2564_2565_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2564_2565_LC_1_11_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2564_2565_LC_1_11_1  (
            .in0(N__33201),
            .in1(N__48865),
            .in2(_gnd_net_),
            .in3(N__70317),
            .lcout(REG_mem_26_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93221),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9972_3_lut_LC_1_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9972_3_lut_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9972_3_lut_LC_1_11_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9972_3_lut_LC_1_11_2  (
            .in0(N__34786),
            .in1(_gnd_net_),
            .in2(N__85621),
            .in3(N__38362),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11621 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12153_LC_1_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12153_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12153_LC_1_11_3 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12153_LC_1_11_3  (
            .in0(N__33202),
            .in1(N__92129),
            .in2(N__88618),
            .in3(N__33270),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14006 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13262_bdd_4_lut_LC_1_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13262_bdd_4_lut_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13262_bdd_4_lut_LC_1_11_4 .LUT_INIT=16'b1111101000001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13262_bdd_4_lut_LC_1_11_4  (
            .in0(N__33829),
            .in1(N__33193),
            .in2(N__85622),
            .in3(N__33835),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13265_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11625_LC_1_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11625_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11625_LC_1_11_5 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11625_LC_1_11_5  (
            .in0(N__90339),
            .in1(N__33157),
            .in2(N__33187),
            .in3(N__81471),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13298_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13298_bdd_4_lut_LC_1_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13298_bdd_4_lut_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13298_bdd_4_lut_LC_1_11_6 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13298_bdd_4_lut_LC_1_11_6  (
            .in0(N__81470),
            .in1(N__33184),
            .in2(N__33178),
            .in3(N__33175),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14006_bdd_4_lut_LC_1_12_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14006_bdd_4_lut_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14006_bdd_4_lut_LC_1_12_0 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14006_bdd_4_lut_LC_1_12_0  (
            .in0(N__92115),
            .in1(N__33169),
            .in2(N__33115),
            .in3(N__33126),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14009_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9978_3_lut_LC_1_12_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9978_3_lut_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9978_3_lut_LC_1_12_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9978_3_lut_LC_1_12_1  (
            .in0(N__85344),
            .in1(_gnd_net_),
            .in2(N__33160),
            .in3(N__33703),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12914_bdd_4_lut_LC_1_12_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12914_bdd_4_lut_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12914_bdd_4_lut_LC_1_12_2 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12914_bdd_4_lut_LC_1_12_2  (
            .in0(N__92114),
            .in1(N__33148),
            .in2(N__33256),
            .in3(N__33240),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12917 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2468_2469_LC_1_12_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2468_2469_LC_1_12_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2468_2469_LC_1_12_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2468_2469_LC_1_12_3  (
            .in0(N__48869),
            .in1(N__95387),
            .in2(N__33127),
            .in3(N__97045),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93224),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2372_2373_LC_1_12_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2372_2373_LC_1_12_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2372_2373_LC_1_12_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2372_2373_LC_1_12_4  (
            .in0(N__95385),
            .in1(N__48868),
            .in2(N__33114),
            .in3(N__96004),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93224),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2660_2661_LC_1_12_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2660_2661_LC_1_12_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2660_2661_LC_1_12_5 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2660_2661_LC_1_12_5  (
            .in0(N__48870),
            .in1(N__79744),
            .in2(N__33271),
            .in3(N__95389),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93224),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5444_5445_LC_1_12_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5444_5445_LC_1_12_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5444_5445_LC_1_12_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5444_5445_LC_1_12_6  (
            .in0(N__95386),
            .in1(N__48871),
            .in2(N__33255),
            .in3(N__96005),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93224),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5540_5541_LC_1_12_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5540_5541_LC_1_12_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5540_5541_LC_1_12_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5540_5541_LC_1_12_7  (
            .in0(N__48872),
            .in1(N__95388),
            .in2(N__33241),
            .in3(N__97046),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93224),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14048_bdd_4_lut_LC_1_13_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14048_bdd_4_lut_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14048_bdd_4_lut_LC_1_13_0 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14048_bdd_4_lut_LC_1_13_0  (
            .in0(N__92140),
            .in1(N__33229),
            .in2(N__48478),
            .in3(N__38581),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12193_LC_1_13_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12193_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12193_LC_1_13_1 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12193_LC_1_13_1  (
            .in0(N__87903),
            .in1(N__92142),
            .in2(N__38890),
            .in3(N__38707),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14048 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12178_LC_1_13_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12178_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12178_LC_1_13_2 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12178_LC_1_13_2  (
            .in0(N__92141),
            .in1(N__87902),
            .in2(N__38761),
            .in3(N__45790),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14036_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14036_bdd_4_lut_LC_1_13_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14036_bdd_4_lut_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14036_bdd_4_lut_LC_1_13_3 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14036_bdd_4_lut_LC_1_13_3  (
            .in0(N__33211),
            .in1(N__35764),
            .in2(N__33223),
            .in3(N__92139),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12129_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11819_LC_1_13_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11819_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11819_LC_1_13_4 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11819_LC_1_13_4  (
            .in0(N__90084),
            .in1(N__85343),
            .in2(N__33220),
            .in3(N__33217),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1307_1308_LC_1_13_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1307_1308_LC_1_13_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1307_1308_LC_1_13_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1307_1308_LC_1_13_5  (
            .in0(N__33210),
            .in1(N__63471),
            .in2(_gnd_net_),
            .in3(N__70141),
            .lcout(REG_mem_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93227),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5636_5637_LC_1_13_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5636_5637_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5636_5637_LC_1_13_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5636_5637_LC_1_13_7  (
            .in0(N__48867),
            .in1(N__33336),
            .in2(_gnd_net_),
            .in3(N__79994),
            .lcout(REG_mem_58_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93227),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i164_165_LC_1_14_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i164_165_LC_1_14_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i164_165_LC_1_14_0 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i164_165_LC_1_14_0  (
            .in0(N__95396),
            .in1(N__48853),
            .in2(N__33325),
            .in3(N__80320),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3236_3237_LC_1_14_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3236_3237_LC_1_14_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3236_3237_LC_1_14_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3236_3237_LC_1_14_1  (
            .in0(N__80321),
            .in1(N__33291),
            .in2(N__48893),
            .in3(N__95400),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9875_3_lut_LC_1_14_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9875_3_lut_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9875_3_lut_LC_1_14_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9875_3_lut_LC_1_14_2  (
            .in0(N__33324),
            .in1(_gnd_net_),
            .in2(N__33304),
            .in3(N__87716),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11524 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i68_69_LC_1_14_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i68_69_LC_1_14_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i68_69_LC_1_14_3 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i68_69_LC_1_14_3  (
            .in0(N__82953),
            .in1(N__33300),
            .in2(N__48894),
            .in3(N__95401),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3140_3141_LC_1_14_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3140_3141_LC_1_14_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3140_3141_LC_1_14_4 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3140_3141_LC_1_14_4  (
            .in0(N__95398),
            .in1(N__48855),
            .in2(N__33283),
            .in3(N__82952),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3242_3243_LC_1_14_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3242_3243_LC_1_14_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3242_3243_LC_1_14_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3242_3243_LC_1_14_5  (
            .in0(N__80322),
            .in1(N__95399),
            .in2(N__46537),
            .in3(N__37332),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2180_2181_LC_1_14_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2180_2181_LC_1_14_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2180_2181_LC_1_14_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2180_2181_LC_1_14_6  (
            .in0(N__95397),
            .in1(N__48854),
            .in2(N__34014),
            .in3(N__76331),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93233),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9929_3_lut_LC_1_14_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9929_3_lut_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9929_3_lut_LC_1_14_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9929_3_lut_LC_1_14_7  (
            .in0(N__87717),
            .in1(N__33292),
            .in2(_gnd_net_),
            .in3(N__33282),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11578 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12776_bdd_4_lut_LC_2_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12776_bdd_4_lut_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12776_bdd_4_lut_LC_2_5_0 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12776_bdd_4_lut_LC_2_5_0  (
            .in0(N__36103),
            .in1(N__92660),
            .in2(N__35365),
            .in3(N__33388),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12779 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11134_LC_2_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11134_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11134_LC_2_5_1 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11134_LC_2_5_1  (
            .in0(N__92662),
            .in1(N__35317),
            .in2(N__88879),
            .in3(N__62032),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12776 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12468_LC_2_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12468_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12468_LC_2_5_2 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12468_LC_2_5_2  (
            .in0(N__54166),
            .in1(N__92663),
            .in2(N__36736),
            .in3(N__88808),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14384_bdd_4_lut_LC_2_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14384_bdd_4_lut_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14384_bdd_4_lut_LC_2_5_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14384_bdd_4_lut_LC_2_5_3  (
            .in0(N__92661),
            .in1(N__36490),
            .in2(N__33382),
            .in3(N__35386),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14387_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10422_3_lut_LC_2_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10422_3_lut_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10422_3_lut_LC_2_5_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10422_3_lut_LC_2_5_4  (
            .in0(N__85567),
            .in1(_gnd_net_),
            .in2(N__33379),
            .in3(N__33376),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12071_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11899_LC_2_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11899_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11899_LC_2_5_5 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11899_LC_2_5_5  (
            .in0(N__81480),
            .in1(N__36415),
            .in2(N__33370),
            .in3(N__90300),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13688_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13688_bdd_4_lut_LC_2_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13688_bdd_4_lut_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13688_bdd_4_lut_LC_2_5_6 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13688_bdd_4_lut_LC_2_5_6  (
            .in0(N__44698),
            .in1(N__81479),
            .in2(N__33367),
            .in3(N__37849),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13691 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10623_3_lut_LC_2_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10623_3_lut_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10623_3_lut_LC_2_6_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10623_3_lut_LC_2_6_0  (
            .in0(N__33351),
            .in1(_gnd_net_),
            .in2(N__33364),
            .in3(N__88331),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12272 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2288_2289_LC_2_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2288_2289_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2288_2289_LC_2_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2288_2289_LC_2_6_1  (
            .in0(N__41613),
            .in1(N__33360),
            .in2(_gnd_net_),
            .in3(N__75065),
            .lcout(REG_mem_23_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2192_2193_LC_2_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2192_2193_LC_2_6_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2192_2193_LC_2_6_2 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2192_2193_LC_2_6_2  (
            .in0(N__41685),
            .in1(N__95689),
            .in2(N__33352),
            .in3(N__76350),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5264_5265_LC_2_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5264_5265_LC_2_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5264_5265_LC_2_6_3 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5264_5265_LC_2_6_3  (
            .in0(N__76351),
            .in1(N__33483),
            .in2(N__95759),
            .in3(N__41687),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6020_6021_LC_2_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6020_6021_LC_2_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6020_6021_LC_2_6_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6020_6021_LC_2_6_4  (
            .in0(N__48846),
            .in1(N__95691),
            .in2(N__33459),
            .in3(N__77892),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3248_3249_LC_2_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3248_3249_LC_2_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3248_3249_LC_2_6_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3248_3249_LC_2_6_5  (
            .in0(N__95688),
            .in1(N__41686),
            .in2(N__33618),
            .in3(N__80323),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5744_5745_LC_2_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5744_5745_LC_2_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5744_5745_LC_2_6_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5744_5745_LC_2_6_6  (
            .in0(N__41688),
            .in1(N__95690),
            .in2(N__33438),
            .in3(N__79750),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6032_6033_LC_2_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6032_6033_LC_2_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6032_6033_LC_2_6_7 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6032_6033_LC_2_6_7  (
            .in0(N__77891),
            .in1(N__33420),
            .in2(N__95760),
            .in3(N__41689),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93239),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12383_LC_2_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12383_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12383_LC_2_7_0 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12383_LC_2_7_0  (
            .in0(N__88810),
            .in1(N__92560),
            .in2(N__34612),
            .in3(N__33421),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11590_LC_2_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11590_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11590_LC_2_7_1 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11590_LC_2_7_1  (
            .in0(N__33543),
            .in1(N__34453),
            .in2(N__92659),
            .in3(N__88809),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13328_bdd_4_lut_LC_2_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13328_bdd_4_lut_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13328_bdd_4_lut_LC_2_7_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13328_bdd_4_lut_LC_2_7_2  (
            .in0(N__33555),
            .in1(N__92556),
            .in2(N__33403),
            .in3(N__33399),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2864_2865_LC_2_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2864_2865_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2864_2865_LC_2_7_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2864_2865_LC_2_7_3  (
            .in0(N__95698),
            .in1(N__41647),
            .in2(N__33400),
            .in3(N__70986),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2768_2769_LC_2_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2768_2769_LC_2_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2768_2769_LC_2_7_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2768_2769_LC_2_7_4  (
            .in0(N__41646),
            .in1(N__95701),
            .in2(N__33556),
            .in3(N__70706),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2960_2961_LC_2_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2960_2961_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2960_2961_LC_2_7_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2960_2961_LC_2_7_5  (
            .in0(N__95699),
            .in1(N__41648),
            .in2(N__33544),
            .in3(N__77893),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5840_5841_LC_2_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5840_5841_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5840_5841_LC_2_7_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5840_5841_LC_2_7_6  (
            .in0(N__41649),
            .in1(N__95702),
            .in2(N__33531),
            .in3(N__70707),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5936_5937_LC_2_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5936_5937_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5936_5937_LC_2_7_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5936_5937_LC_2_7_7  (
            .in0(N__95700),
            .in1(N__41650),
            .in2(N__33514),
            .in3(N__70987),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93234),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12974_bdd_4_lut_LC_2_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12974_bdd_4_lut_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12974_bdd_4_lut_LC_2_8_0 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12974_bdd_4_lut_LC_2_8_0  (
            .in0(N__34579),
            .in1(N__92425),
            .in2(N__34561),
            .in3(N__33637),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12977_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9923_3_lut_LC_2_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9923_3_lut_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9923_3_lut_LC_2_8_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9923_3_lut_LC_2_8_1  (
            .in0(_gnd_net_),
            .in1(N__85440),
            .in2(N__33499),
            .in3(N__33469),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11206_LC_2_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11206_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11206_LC_2_8_2 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11206_LC_2_8_2  (
            .in0(N__33661),
            .in1(N__92426),
            .in2(N__33490),
            .in3(N__88617),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12866_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12866_bdd_4_lut_LC_2_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12866_bdd_4_lut_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12866_bdd_4_lut_LC_2_8_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12866_bdd_4_lut_LC_2_8_3  (
            .in0(N__92424),
            .in1(N__33648),
            .in2(N__33472),
            .in3(N__34515),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12869 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2096_2097_LC_2_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2096_2097_LC_2_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2096_2097_LC_2_8_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2096_2097_LC_2_8_4  (
            .in0(N__41721),
            .in1(N__95374),
            .in2(N__34552),
            .in3(N__77013),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93228),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5360_5361_LC_2_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5360_5361_LC_2_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5360_5361_LC_2_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5360_5361_LC_2_8_5  (
            .in0(N__33660),
            .in1(N__41720),
            .in2(_gnd_net_),
            .in3(N__77230),
            .lcout(REG_mem_55_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93228),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5168_5169_LC_2_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5168_5169_LC_2_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5168_5169_LC_2_8_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5168_5169_LC_2_8_6  (
            .in0(N__41722),
            .in1(N__95375),
            .in2(N__33649),
            .in3(N__77014),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93228),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4688_4689_LC_2_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4688_4689_LC_2_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4688_4689_LC_2_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4688_4689_LC_2_8_7  (
            .in0(N__33636),
            .in1(N__41719),
            .in2(_gnd_net_),
            .in3(N__75566),
            .lcout(REG_mem_48_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93228),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2756_2757_LC_2_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2756_2757_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2756_2757_LC_2_9_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2756_2757_LC_2_9_0  (
            .in0(N__48811),
            .in1(N__95377),
            .in2(N__33718),
            .in3(N__70713),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93225),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10706_3_lut_LC_2_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10706_3_lut_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10706_3_lut_LC_2_9_1 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10706_3_lut_LC_2_9_1  (
            .in0(N__33769),
            .in1(N__33568),
            .in2(N__88774),
            .in3(_gnd_net_),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10683_3_lut_LC_2_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10683_3_lut_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10683_3_lut_LC_2_9_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10683_3_lut_LC_2_9_2  (
            .in0(N__34087),
            .in1(N__88613),
            .in2(_gnd_net_),
            .in3(N__33759),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10682_3_lut_LC_2_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10682_3_lut_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10682_3_lut_LC_2_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10682_3_lut_LC_2_9_3  (
            .in0(N__88612),
            .in1(N__33622),
            .in2(_gnd_net_),
            .in3(N__35785),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12962_bdd_4_lut_LC_2_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12962_bdd_4_lut_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12962_bdd_4_lut_LC_2_9_4 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12962_bdd_4_lut_LC_2_9_4  (
            .in0(N__35458),
            .in1(N__92321),
            .in2(N__33589),
            .in3(N__35437),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12965 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3536_3537_LC_2_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3536_3537_LC_2_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3536_3537_LC_2_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3536_3537_LC_2_9_5  (
            .in0(N__33567),
            .in1(N__41723),
            .in2(_gnd_net_),
            .in3(N__54094),
            .lcout(REG_mem_36_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93225),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3632_3633_LC_2_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3632_3633_LC_2_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3632_3633_LC_2_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3632_3633_LC_2_9_6  (
            .in0(N__41724),
            .in1(N__33768),
            .in2(_gnd_net_),
            .in3(N__63727),
            .lcout(REG_mem_37_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93225),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3344_3345_LC_2_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3344_3345_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3344_3345_LC_2_9_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3344_3345_LC_2_9_7  (
            .in0(N__95376),
            .in1(N__41725),
            .in2(N__33760),
            .in3(N__80599),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93225),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3044_3045_LC_2_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3044_3045_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3044_3045_LC_2_10_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3044_3045_LC_2_10_0  (
            .in0(N__33747),
            .in1(N__72515),
            .in2(_gnd_net_),
            .in3(N__48878),
            .lcout(REG_mem_31_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93219),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12063_LC_2_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12063_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12063_LC_2_10_1 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12063_LC_2_10_1  (
            .in0(N__88610),
            .in1(N__33748),
            .in2(N__33739),
            .in3(N__92408),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13898_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13898_bdd_4_lut_LC_2_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13898_bdd_4_lut_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13898_bdd_4_lut_LC_2_10_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13898_bdd_4_lut_LC_2_10_2  (
            .in0(N__92407),
            .in1(N__33693),
            .in2(N__33721),
            .in3(N__33717),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13901 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2852_2853_LC_2_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2852_2853_LC_2_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2852_2853_LC_2_10_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2852_2853_LC_2_10_3  (
            .in0(N__48880),
            .in1(N__95373),
            .in2(N__33694),
            .in3(N__70897),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93219),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9878_3_lut_LC_2_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9878_3_lut_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9878_3_lut_LC_2_10_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9878_3_lut_LC_2_10_4  (
            .in0(N__34819),
            .in1(N__88608),
            .in2(_gnd_net_),
            .in3(N__38314),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11527 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9899_3_lut_LC_2_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9899_3_lut_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9899_3_lut_LC_2_10_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9899_3_lut_LC_2_10_5  (
            .in0(N__88609),
            .in1(_gnd_net_),
            .in2(N__33871),
            .in3(N__34492),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11548 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1604_1605_LC_2_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1604_1605_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1604_1605_LC_2_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1604_1605_LC_2_10_6  (
            .in0(N__33672),
            .in1(N__48877),
            .in2(_gnd_net_),
            .in3(N__65686),
            .lcout(REG_mem_16_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93219),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2084_2085_LC_2_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2084_2085_LC_2_10_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2084_2085_LC_2_10_7 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2084_2085_LC_2_10_7  (
            .in0(N__48879),
            .in1(N__95372),
            .in2(N__33870),
            .in3(N__76975),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93219),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9986_3_lut_LC_2_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9986_3_lut_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9986_3_lut_LC_2_11_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9986_3_lut_LC_2_11_0  (
            .in0(N__35413),
            .in1(N__85480),
            .in2(_gnd_net_),
            .in3(N__33856),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11535_LC_2_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11535_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11535_LC_2_11_1 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11535_LC_2_11_1  (
            .in0(N__85481),
            .in1(N__33841),
            .in2(N__92654),
            .in3(N__33997),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9897_3_lut_LC_2_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9897_3_lut_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9897_3_lut_LC_2_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9897_3_lut_LC_2_11_2  (
            .in0(N__88374),
            .in1(N__33814),
            .in2(_gnd_net_),
            .in3(N__33823),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11546 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1796_1797_LC_2_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1796_1797_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1796_1797_LC_2_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1796_1797_LC_2_11_3  (
            .in0(N__33822),
            .in1(N__48881),
            .in2(_gnd_net_),
            .in3(N__67509),
            .lcout(REG_mem_18_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93226),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1892_1893_LC_2_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1892_1893_LC_2_11_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1892_1893_LC_2_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1892_1893_LC_2_11_4  (
            .in0(N__48882),
            .in1(N__33813),
            .in2(_gnd_net_),
            .in3(N__72115),
            .lcout(REG_mem_19_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93226),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14228_bdd_4_lut_LC_2_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14228_bdd_4_lut_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14228_bdd_4_lut_LC_2_11_5 .LUT_INIT=16'b1010110110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14228_bdd_4_lut_LC_2_11_5  (
            .in0(N__33805),
            .in1(N__37486),
            .in2(N__81399),
            .in3(N__34138),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9879_3_lut_LC_2_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9879_3_lut_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9879_3_lut_LC_2_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9879_3_lut_LC_2_11_6  (
            .in0(N__88373),
            .in1(N__43423),
            .in2(_gnd_net_),
            .in3(N__34591),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11528 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5648_5649_LC_2_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5648_5649_LC_2_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5648_5649_LC_2_11_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5648_5649_LC_2_11_7  (
            .in0(N__33780),
            .in1(N__79935),
            .in2(_gnd_net_),
            .in3(N__41726),
            .lcout(REG_mem_58_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93226),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11325_LC_2_12_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11325_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11325_LC_2_12_0 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11325_LC_2_12_0  (
            .in0(N__91871),
            .in1(N__88031),
            .in2(N__33946),
            .in3(N__35689),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12998_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12998_bdd_4_lut_LC_2_12_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12998_bdd_4_lut_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12998_bdd_4_lut_LC_2_12_1 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12998_bdd_4_lut_LC_2_12_1  (
            .in0(N__34480),
            .in1(N__91870),
            .in2(N__33952),
            .in3(N__38629),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13001_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12438_LC_2_12_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12438_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12438_LC_2_12_2 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12438_LC_2_12_2  (
            .in0(N__85329),
            .in1(N__34888),
            .in2(N__33949),
            .in3(N__90221),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2639_2640_LC_2_12_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2639_2640_LC_2_12_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2639_2640_LC_2_12_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2639_2640_LC_2_12_3  (
            .in0(N__61343),
            .in1(N__95384),
            .in2(N__34737),
            .in3(N__79745),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93229),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5999_6000_LC_2_12_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5999_6000_LC_2_12_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5999_6000_LC_2_12_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5999_6000_LC_2_12_4  (
            .in0(N__95383),
            .in1(N__61344),
            .in2(N__33945),
            .in3(N__77943),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93229),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2576_2577_LC_2_12_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2576_2577_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2576_2577_LC_2_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2576_2577_LC_2_12_5  (
            .in0(N__33921),
            .in1(N__41765),
            .in2(_gnd_net_),
            .in3(N__70383),
            .lcout(REG_mem_26_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93229),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11490_LC_2_12_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11490_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11490_LC_2_12_6 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11490_LC_2_12_6  (
            .in0(N__91872),
            .in1(N__41905),
            .in2(N__85437),
            .in3(N__33910),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13196 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i143_144_LC_2_13_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i143_144_LC_2_13_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i143_144_LC_2_13_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i143_144_LC_2_13_0  (
            .in0(N__61107),
            .in1(N__95393),
            .in2(N__33886),
            .in3(N__80300),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12368_LC_2_13_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12368_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12368_LC_2_13_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12368_LC_2_13_1  (
            .in0(N__91995),
            .in1(N__87726),
            .in2(N__34030),
            .in3(N__34041),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14264_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14264_bdd_4_lut_LC_2_13_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14264_bdd_4_lut_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14264_bdd_4_lut_LC_2_13_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14264_bdd_4_lut_LC_2_13_2  (
            .in0(N__33885),
            .in1(N__91994),
            .in2(N__33874),
            .in3(N__34053),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11523 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i47_48_LC_2_13_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i47_48_LC_2_13_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i47_48_LC_2_13_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i47_48_LC_2_13_3  (
            .in0(N__95392),
            .in1(N__61112),
            .in2(N__34054),
            .in3(N__82940),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i239_240_LC_2_13_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i239_240_LC_2_13_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i239_240_LC_2_13_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i239_240_LC_2_13_4  (
            .in0(N__61108),
            .in1(N__95394),
            .in2(N__34042),
            .in3(N__80600),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i335_336_LC_2_13_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i335_336_LC_2_13_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i335_336_LC_2_13_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i335_336_LC_2_13_5  (
            .in0(N__95391),
            .in1(N__61111),
            .in2(N__34029),
            .in3(N__83389),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3215_3216_LC_2_13_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3215_3216_LC_2_13_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3215_3216_LC_2_13_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3215_3216_LC_2_13_6  (
            .in0(N__61109),
            .in1(N__95395),
            .in2(N__33969),
            .in3(N__80301),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3119_3120_LC_2_13_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3119_3120_LC_2_13_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3119_3120_LC_2_13_7 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3119_3120_LC_2_13_7  (
            .in0(N__95390),
            .in1(N__61110),
            .in2(N__33987),
            .in3(N__82939),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93235),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9935_3_lut_LC_2_14_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9935_3_lut_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9935_3_lut_LC_2_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9935_3_lut_LC_2_14_0  (
            .in0(N__34129),
            .in1(N__88043),
            .in2(_gnd_net_),
            .in3(N__34120),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11584 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9900_3_lut_LC_2_14_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9900_3_lut_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9900_3_lut_LC_2_14_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9900_3_lut_LC_2_14_1  (
            .in0(N__88041),
            .in1(N__34015),
            .in2(_gnd_net_),
            .in3(N__38911),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11549 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10142_3_lut_LC_2_14_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10142_3_lut_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10142_3_lut_LC_2_14_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10142_3_lut_LC_2_14_2  (
            .in0(N__33988),
            .in1(N__88040),
            .in2(_gnd_net_),
            .in3(N__33970),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9930_3_lut_LC_2_14_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9930_3_lut_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9930_3_lut_LC_2_14_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9930_3_lut_LC_2_14_3  (
            .in0(N__88042),
            .in1(_gnd_net_),
            .in2(N__34111),
            .in3(N__34218),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11579_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13268_bdd_4_lut_LC_2_14_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13268_bdd_4_lut_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13268_bdd_4_lut_LC_2_14_4 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13268_bdd_4_lut_LC_2_14_4  (
            .in0(N__85325),
            .in1(N__34147),
            .in2(N__34141),
            .in3(N__34060),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3524_3525_LC_2_14_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3524_3525_LC_2_14_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3524_3525_LC_2_14_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3524_3525_LC_2_14_5  (
            .in0(N__54098),
            .in1(N__34128),
            .in2(_gnd_net_),
            .in3(N__48850),
            .lcout(REG_mem_36_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93240),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3620_3621_LC_2_14_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3620_3621_LC_2_14_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3620_3621_LC_2_14_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3620_3621_LC_2_14_6  (
            .in0(N__48851),
            .in1(N__34119),
            .in2(_gnd_net_),
            .in3(N__63733),
            .lcout(REG_mem_37_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93240),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3332_3333_LC_2_14_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3332_3333_LC_2_14_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3332_3333_LC_2_14_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3332_3333_LC_2_14_7  (
            .in0(N__80576),
            .in1(N__48852),
            .in2(N__34110),
            .in3(N__95407),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93240),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10536_3_lut_LC_2_15_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10536_3_lut_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10536_3_lut_LC_2_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10536_3_lut_LC_2_15_0  (
            .in0(N__87594),
            .in1(N__34096),
            .in2(_gnd_net_),
            .in3(N__35139),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12185 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5642_5643_LC_2_15_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5642_5643_LC_2_15_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5642_5643_LC_2_15_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5642_5643_LC_2_15_1  (
            .in0(N__35112),
            .in1(N__46580),
            .in2(_gnd_net_),
            .in3(N__79968),
            .lcout(REG_mem_58_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93247),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i368_369_LC_2_15_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i368_369_LC_2_15_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i368_369_LC_2_15_2 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i368_369_LC_2_15_2  (
            .in0(N__83386),
            .in1(N__41783),
            .in2(N__95634),
            .in3(N__34095),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93247),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3440_3441_LC_2_15_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3440_3441_LC_2_15_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3440_3441_LC_2_15_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3440_3441_LC_2_15_3  (
            .in0(N__41782),
            .in1(N__95403),
            .in2(N__34086),
            .in3(N__83388),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93247),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11555_LC_2_15_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11555_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11555_LC_2_15_4 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11555_LC_2_15_4  (
            .in0(N__91992),
            .in1(N__34069),
            .in2(N__50677),
            .in3(N__85231),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9876_3_lut_LC_2_15_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9876_3_lut_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9876_3_lut_LC_2_15_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9876_3_lut_LC_2_15_5  (
            .in0(N__35047),
            .in1(N__34230),
            .in2(_gnd_net_),
            .in3(N__87595),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11525 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i356_357_LC_2_15_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i356_357_LC_2_15_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i356_357_LC_2_15_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i356_357_LC_2_15_6  (
            .in0(N__83385),
            .in1(N__48898),
            .in2(N__34231),
            .in3(N__95408),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93247),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3428_3429_LC_2_15_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3428_3429_LC_2_15_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3428_3429_LC_2_15_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3428_3429_LC_2_15_7  (
            .in0(N__48897),
            .in1(N__95402),
            .in2(N__34219),
            .in3(N__83387),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93247),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.usb3_data_in_latched__i14_LC_3_1_3 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i14_LC_3_1_3 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i14_LC_3_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i14_LC_3_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34204),
            .lcout(\usb3_if_inst.usb3_data_in_latched_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93303),
            .ce(),
            .sr(N__73756));
    defparam \usb3_if_inst.usb3_data_in_latched__i15_LC_3_2_0 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i15_LC_3_2_0 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i15_LC_3_2_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i15_LC_3_2_0  (
            .in0(N__34192),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\usb3_if_inst.usb3_data_in_latched_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93289),
            .ce(),
            .sr(N__73755));
    defparam \usb3_if_inst.usb3_data_in_latched__i16_LC_3_2_5 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i16_LC_3_2_5 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i16_LC_3_2_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i16_LC_3_2_5  (
            .in0(N__34177),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\usb3_if_inst.usb3_data_in_latched_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93289),
            .ce(),
            .sr(N__73755));
    defparam \usb3_if_inst.dc32_fifo_data_in_i15_LC_3_3_1 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i15_LC_3_3_1 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i15_LC_3_3_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i15_LC_3_3_1  (
            .in0(_gnd_net_),
            .in1(N__34162),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(dc32_fifo_data_in_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.dc32_fifo_data_in_i15C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3041_3042_LC_3_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3041_3042_LC_3_5_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3041_3042_LC_3_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3041_3042_LC_3_5_0  (
            .in0(N__34155),
            .in1(N__56457),
            .in2(_gnd_net_),
            .in3(N__72565),
            .lcout(REG_mem_31_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11301_LC_3_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11301_LC_3_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11301_LC_3_5_1 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11301_LC_3_5_1  (
            .in0(N__90976),
            .in1(N__34156),
            .in2(N__34633),
            .in3(N__88589),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12980_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12980_bdd_4_lut_LC_3_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12980_bdd_4_lut_LC_3_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12980_bdd_4_lut_LC_3_5_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12980_bdd_4_lut_LC_3_5_2  (
            .in0(N__34297),
            .in1(N__90975),
            .in2(N__34300),
            .in3(N__34288),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12983 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2849_2850_LC_3_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2849_2850_LC_3_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2849_2850_LC_3_5_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2849_2850_LC_3_5_3  (
            .in0(N__95442),
            .in1(N__34296),
            .in2(N__56549),
            .in3(N__70988),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2753_2754_LC_3_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2753_2754_LC_3_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2753_2754_LC_3_5_4 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2753_2754_LC_3_5_4  (
            .in0(N__34287),
            .in1(N__95444),
            .in2(N__70728),
            .in3(N__56458),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5924_5925_LC_3_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5924_5925_LC_3_5_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5924_5925_LC_3_5_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5924_5925_LC_3_5_5  (
            .in0(N__95443),
            .in1(N__48725),
            .in2(N__34272),
            .in3(N__70989),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5825_5826_LC_3_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5825_5826_LC_3_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5825_5826_LC_3_5_6 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5825_5826_LC_3_5_6  (
            .in0(N__34368),
            .in1(N__95445),
            .in2(N__70729),
            .in3(N__56459),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93255),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11520_LC_3_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11520_LC_3_5_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11520_LC_3_5_7 .LUT_INIT=16'b1100101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11520_LC_3_5_7  (
            .in0(N__34420),
            .in1(N__34339),
            .in2(N__90350),
            .in3(N__81469),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13814_bdd_4_lut_LC_3_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13814_bdd_4_lut_LC_3_6_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13814_bdd_4_lut_LC_3_6_0 .LUT_INIT=16'b1011101010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13814_bdd_4_lut_LC_3_6_0  (
            .in0(N__36748),
            .in1(N__90973),
            .in2(N__41827),
            .in3(N__41326),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13817_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9864_3_lut_LC_3_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9864_3_lut_LC_3_6_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9864_3_lut_LC_3_6_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9864_3_lut_LC_3_6_1  (
            .in0(N__35572),
            .in1(_gnd_net_),
            .in2(N__34255),
            .in3(N__85563),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11513_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13226_bdd_4_lut_LC_3_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13226_bdd_4_lut_LC_3_6_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13226_bdd_4_lut_LC_3_6_2 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13226_bdd_4_lut_LC_3_6_2  (
            .in0(N__81468),
            .in1(N__34252),
            .in2(N__34246),
            .in3(N__34375),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11450_LC_3_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11450_LC_3_6_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11450_LC_3_6_3 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11450_LC_3_6_3  (
            .in0(N__90974),
            .in1(N__85566),
            .in2(N__36691),
            .in3(N__34501),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13160_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13160_bdd_4_lut_LC_3_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13160_bdd_4_lut_LC_3_6_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13160_bdd_4_lut_LC_3_6_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13160_bdd_4_lut_LC_3_6_4  (
            .in0(N__85565),
            .in1(N__41008),
            .in2(N__34393),
            .in3(N__34390),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10817_3_lut_LC_3_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10817_3_lut_LC_3_6_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10817_3_lut_LC_3_6_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10817_3_lut_LC_3_6_5  (
            .in0(N__34369),
            .in1(N__88804),
            .in2(_gnd_net_),
            .in3(N__35401),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12466 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9885_3_lut_LC_3_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9885_3_lut_LC_3_6_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9885_3_lut_LC_3_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9885_3_lut_LC_3_6_6  (
            .in0(N__85564),
            .in1(N__34357),
            .in2(_gnd_net_),
            .in3(N__34345),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2447_2448_LC_3_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2447_2448_LC_3_7_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2447_2448_LC_3_7_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2447_2448_LC_3_7_0  (
            .in0(N__61373),
            .in1(N__95528),
            .in2(N__34755),
            .in3(N__97036),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93241),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4496_4497_LC_3_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4496_4497_LC_3_7_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4496_4497_LC_3_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4496_4497_LC_3_7_1  (
            .in0(N__34320),
            .in1(N__41529),
            .in2(_gnd_net_),
            .in3(N__89124),
            .lcout(REG_mem_46_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93241),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11405_LC_3_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11405_LC_3_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11405_LC_3_7_2 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11405_LC_3_7_2  (
            .in0(N__92658),
            .in1(N__41845),
            .in2(N__88803),
            .in3(N__41440),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13106_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13106_bdd_4_lut_LC_3_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13106_bdd_4_lut_LC_3_7_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13106_bdd_4_lut_LC_3_7_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13106_bdd_4_lut_LC_3_7_3  (
            .in0(N__39793),
            .in1(N__92656),
            .in2(N__34333),
            .in3(N__38068),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11355_LC_3_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11355_LC_3_7_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11355_LC_3_7_4 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11355_LC_3_7_4  (
            .in0(N__92657),
            .in1(N__34321),
            .in2(N__88802),
            .in3(N__40231),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13046_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13046_bdd_4_lut_LC_3_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13046_bdd_4_lut_LC_3_7_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13046_bdd_4_lut_LC_3_7_5 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13046_bdd_4_lut_LC_3_7_5  (
            .in0(N__34462),
            .in1(N__92655),
            .in2(N__34312),
            .in3(N__38260),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13049 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4304_4305_LC_3_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4304_4305_LC_3_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4304_4305_LC_3_7_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4304_4305_LC_3_7_6  (
            .in0(N__41528),
            .in1(N__34461),
            .in2(_gnd_net_),
            .in3(N__71763),
            .lcout(REG_mem_44_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93241),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3056_3057_LC_3_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3056_3057_LC_3_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3056_3057_LC_3_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3056_3057_LC_3_7_7  (
            .in0(N__34449),
            .in1(N__41527),
            .in2(_gnd_net_),
            .in3(N__72564),
            .lcout(REG_mem_31_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93241),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10599_3_lut_LC_3_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10599_3_lut_LC_3_8_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10599_3_lut_LC_3_8_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10599_3_lut_LC_3_8_0  (
            .in0(N__88611),
            .in1(N__34402),
            .in2(_gnd_net_),
            .in3(N__34411),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11475_LC_3_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11475_LC_3_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11475_LC_3_8_1 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11475_LC_3_8_1  (
            .in0(N__92555),
            .in1(N__85439),
            .in2(N__34525),
            .in3(N__34438),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13190_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13190_bdd_4_lut_LC_3_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13190_bdd_4_lut_LC_3_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13190_bdd_4_lut_LC_3_8_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13190_bdd_4_lut_LC_3_8_2  (
            .in0(N__85438),
            .in1(N__36826),
            .in2(N__34429),
            .in3(N__34426),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13193 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1808_1809_LC_3_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1808_1809_LC_3_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1808_1809_LC_3_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1808_1809_LC_3_8_3  (
            .in0(N__34410),
            .in1(N__41558),
            .in2(_gnd_net_),
            .in3(N__67499),
            .lcout(REG_mem_18_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1904_1905_LC_3_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1904_1905_LC_3_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1904_1905_LC_3_8_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1904_1905_LC_3_8_4  (
            .in0(N__41559),
            .in1(N__34401),
            .in2(_gnd_net_),
            .in3(N__72113),
            .lcout(REG_mem_19_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5711_5712_LC_3_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5711_5712_LC_3_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5711_5712_LC_3_8_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5711_5712_LC_3_8_5  (
            .in0(N__95740),
            .in1(N__61398),
            .in2(N__34710),
            .in3(N__79741),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5423_5424_LC_3_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5423_5424_LC_3_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5423_5424_LC_3_8_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5423_5424_LC_3_8_6  (
            .in0(N__61397),
            .in1(N__95741),
            .in2(N__34909),
            .in3(N__95955),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4784_4785_LC_3_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4784_4785_LC_3_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4784_4785_LC_3_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4784_4785_LC_3_8_7  (
            .in0(N__34572),
            .in1(N__41560),
            .in2(_gnd_net_),
            .in3(N__62984),
            .lcout(REG_mem_49_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93236),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11296_LC_3_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11296_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11296_LC_3_9_0 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11296_LC_3_9_0  (
            .in0(N__92545),
            .in1(N__88607),
            .in2(N__40000),
            .in3(N__38530),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12974 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2000_2001_LC_3_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2000_2001_LC_3_9_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2000_2001_LC_3_9_1 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2000_2001_LC_3_9_1  (
            .in0(N__41667),
            .in1(N__95424),
            .in2(N__34537),
            .in3(N__77441),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10622_3_lut_LC_3_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10622_3_lut_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10622_3_lut_LC_3_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10622_3_lut_LC_3_9_2  (
            .in0(N__34551),
            .in1(N__34536),
            .in2(_gnd_net_),
            .in3(N__88606),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5072_5073_LC_3_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5072_5073_LC_3_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5072_5073_LC_3_9_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5072_5073_LC_3_9_3  (
            .in0(N__41668),
            .in1(N__95425),
            .in2(N__34516),
            .in3(N__77442),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10542_3_lut_LC_3_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10542_3_lut_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10542_3_lut_LC_3_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10542_3_lut_LC_3_9_4  (
            .in0(N__36895),
            .in1(N__88605),
            .in2(_gnd_net_),
            .in3(N__39697),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12191 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1988_1989_LC_3_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1988_1989_LC_3_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1988_1989_LC_3_9_5 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1988_1989_LC_3_9_5  (
            .in0(N__48810),
            .in1(N__34491),
            .in2(N__77479),
            .in3(N__95427),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2735_2736_LC_3_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2735_2736_LC_3_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2735_2736_LC_3_9_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2735_2736_LC_3_9_6  (
            .in0(N__95423),
            .in1(N__61399),
            .in2(N__34684),
            .in3(N__70676),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5807_5808_LC_3_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5807_5808_LC_3_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5807_5808_LC_3_9_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5807_5808_LC_3_9_7  (
            .in0(N__70675),
            .in1(N__34479),
            .in2(N__61405),
            .in3(N__95426),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93230),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3023_3024_LC_3_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3023_3024_LC_3_10_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3023_3024_LC_3_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3023_3024_LC_3_10_0  (
            .in0(N__34692),
            .in1(N__61263),
            .in2(_gnd_net_),
            .in3(N__72514),
            .lcout(REG_mem_31_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93222),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12148_LC_3_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12148_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12148_LC_3_10_1 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12148_LC_3_10_1  (
            .in0(N__92401),
            .in1(N__88604),
            .in2(N__34777),
            .in3(N__34693),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14000_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14000_bdd_4_lut_LC_3_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14000_bdd_4_lut_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14000_bdd_4_lut_LC_3_10_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14000_bdd_4_lut_LC_3_10_2  (
            .in0(N__34683),
            .in1(N__92400),
            .in2(N__34669),
            .in3(N__34665),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14003 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2831_2832_LC_3_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2831_2832_LC_3_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2831_2832_LC_3_10_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2831_2832_LC_3_10_3  (
            .in0(N__61262),
            .in1(N__95422),
            .in2(N__34666),
            .in3(N__70896),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93222),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3329_3330_LC_3_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3329_3330_LC_3_10_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3329_3330_LC_3_10_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3329_3330_LC_3_10_4  (
            .in0(N__95420),
            .in1(N__56605),
            .in2(N__34650),
            .in3(N__80598),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93222),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i161_162_LC_3_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i161_162_LC_3_10_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i161_162_LC_3_10_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i161_162_LC_3_10_5  (
            .in0(N__56603),
            .in1(N__95421),
            .in2(N__40125),
            .in3(N__80167),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93222),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2945_2946_LC_3_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2945_2946_LC_3_10_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2945_2946_LC_3_10_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2945_2946_LC_3_10_6  (
            .in0(N__95419),
            .in1(N__56604),
            .in2(N__34629),
            .in3(N__77840),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93222),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6128_6129_LC_3_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6128_6129_LC_3_10_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6128_6129_LC_3_10_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6128_6129_LC_3_10_7  (
            .in0(N__41561),
            .in1(N__67672),
            .in2(_gnd_net_),
            .in3(N__34602),
            .lcout(REG_mem_63_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93222),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i644_645_LC_3_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i644_645_LC_3_11_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i644_645_LC_3_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i644_645_LC_3_11_0  (
            .in0(N__48876),
            .in1(N__34590),
            .in2(_gnd_net_),
            .in3(N__66430),
            .lcout(REG_mem_6_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1028_1029_LC_3_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1028_1029_LC_3_11_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1028_1029_LC_3_11_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1028_1029_LC_3_11_1  (
            .in0(N__34806),
            .in1(N__48873),
            .in2(_gnd_net_),
            .in3(N__66973),
            .lcout(REG_mem_10_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1124_1125_LC_3_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1124_1125_LC_3_11_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1124_1125_LC_3_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1124_1125_LC_3_11_2  (
            .in0(N__48874),
            .in1(N__34797),
            .in2(_gnd_net_),
            .in3(N__66829),
            .lcout(REG_mem_11_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i548_549_LC_3_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i548_549_LC_3_11_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i548_549_LC_3_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i548_549_LC_3_11_3  (
            .in0(N__34818),
            .in1(N__48875),
            .in2(_gnd_net_),
            .in3(N__67888),
            .lcout(REG_mem_5_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12303_LC_3_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12303_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12303_LC_3_11_4 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12303_LC_3_11_4  (
            .in0(N__92541),
            .in1(N__34807),
            .in2(N__88372),
            .in3(N__34798),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14180_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14180_bdd_4_lut_LC_3_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14180_bdd_4_lut_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14180_bdd_4_lut_LC_3_11_5 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14180_bdd_4_lut_LC_3_11_5  (
            .in0(N__35746),
            .in1(N__92540),
            .in2(N__34789),
            .in3(N__37384),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2927_2928_LC_3_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2927_2928_LC_3_11_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2927_2928_LC_3_11_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2927_2928_LC_3_11_6  (
            .in0(N__61251),
            .in1(N__94974),
            .in2(N__34776),
            .in3(N__77904),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5723_5724_LC_3_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5723_5724_LC_3_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5723_5724_LC_3_11_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5723_5724_LC_3_11_7  (
            .in0(N__94973),
            .in1(N__63382),
            .in2(N__38670),
            .in3(N__79786),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93231),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14096_bdd_4_lut_LC_3_12_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14096_bdd_4_lut_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14096_bdd_4_lut_LC_3_12_0 .LUT_INIT=16'b1100101111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14096_bdd_4_lut_LC_3_12_0  (
            .in0(N__34759),
            .in1(N__34720),
            .in2(N__92209),
            .in3(N__34878),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14099 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12228_LC_3_12_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12228_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12228_LC_3_12_1 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12228_LC_3_12_1  (
            .in0(N__88030),
            .in1(N__91869),
            .in2(N__34738),
            .in3(N__34855),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14096 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11365_LC_3_12_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11365_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11365_LC_3_12_2 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11365_LC_3_12_2  (
            .in0(N__91868),
            .in1(N__88029),
            .in2(N__34714),
            .in3(N__45730),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13052_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13052_bdd_4_lut_LC_3_12_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13052_bdd_4_lut_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13052_bdd_4_lut_LC_3_12_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13052_bdd_4_lut_LC_3_12_3  (
            .in0(N__34845),
            .in1(N__91864),
            .in2(N__34912),
            .in3(N__34908),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13055 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2351_2352_LC_3_12_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2351_2352_LC_3_12_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2351_2352_LC_3_12_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2351_2352_LC_3_12_4  (
            .in0(N__95642),
            .in1(N__61345),
            .in2(N__34879),
            .in3(N__96010),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93237),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14336_bdd_4_lut_LC_3_12_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14336_bdd_4_lut_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14336_bdd_4_lut_LC_3_12_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14336_bdd_4_lut_LC_3_12_5  (
            .in0(N__90134),
            .in1(N__36862),
            .in2(N__34864),
            .in3(N__35470),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2543_2544_LC_3_12_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2543_2544_LC_3_12_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2543_2544_LC_3_12_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2543_2544_LC_3_12_6  (
            .in0(N__34854),
            .in1(_gnd_net_),
            .in2(N__61332),
            .in3(N__70378),
            .lcout(REG_mem_26_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93237),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5519_5520_LC_3_12_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5519_5520_LC_3_12_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5519_5520_LC_3_12_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5519_5520_LC_3_12_7  (
            .in0(N__97047),
            .in1(N__95643),
            .in2(N__34846),
            .in3(N__61264),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93237),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10342_3_lut_LC_3_13_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10342_3_lut_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10342_3_lut_LC_3_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10342_3_lut_LC_3_13_0  (
            .in0(N__90142),
            .in1(N__35014),
            .in2(_gnd_net_),
            .in3(N__37054),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11991_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12408_LC_3_13_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12408_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12408_LC_3_13_1 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12408_LC_3_13_1  (
            .in0(N__81016),
            .in1(N__34834),
            .in2(N__34825),
            .in3(N__81416),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14312_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i4_LC_3_13_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i4_LC_3_13_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i4_LC_3_13_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i4_LC_3_13_2  (
            .in0(N__34966),
            .in1(N__81015),
            .in2(N__34822),
            .in3(N__34945),
            .lcout(REG_out_raw_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97342),
            .ce(N__80880),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11231_LC_3_13_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11231_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11231_LC_3_13_3 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11231_LC_3_13_3  (
            .in0(N__37090),
            .in1(N__38719),
            .in2(N__90229),
            .in3(N__85324),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10326_3_lut_LC_3_13_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10326_3_lut_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10326_3_lut_LC_3_13_4 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10326_3_lut_LC_3_13_4  (
            .in0(N__85323),
            .in1(N__34987),
            .in2(N__34978),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11975_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10327_3_lut_LC_3_13_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10327_3_lut_LC_3_13_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10327_3_lut_LC_3_13_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10327_3_lut_LC_3_13_5  (
            .in0(N__36799),
            .in1(_gnd_net_),
            .in2(N__34969),
            .in3(N__90141),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11976 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12806_bdd_4_lut_LC_3_13_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12806_bdd_4_lut_LC_3_13_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12806_bdd_4_lut_LC_3_13_6 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12806_bdd_4_lut_LC_3_13_6  (
            .in0(N__90143),
            .in1(N__34960),
            .in2(N__34954),
            .in3(N__35947),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12809 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13322_bdd_4_lut_LC_3_14_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13322_bdd_4_lut_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13322_bdd_4_lut_LC_3_14_0 .LUT_INIT=16'b1011101010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13322_bdd_4_lut_LC_3_14_0  (
            .in0(N__34939),
            .in1(N__91745),
            .in2(N__38029),
            .in3(N__35878),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11585_LC_3_14_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11585_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11585_LC_3_14_1 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11585_LC_3_14_1  (
            .in0(N__91747),
            .in1(N__36040),
            .in2(N__88332),
            .in3(N__35074),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11545_LC_3_14_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11545_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11545_LC_3_14_2 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11545_LC_3_14_2  (
            .in0(N__34921),
            .in1(N__91746),
            .in2(N__35719),
            .in3(N__88036),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13274_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13274_bdd_4_lut_LC_3_14_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13274_bdd_4_lut_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13274_bdd_4_lut_LC_3_14_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13274_bdd_4_lut_LC_3_14_3  (
            .in0(N__91744),
            .in1(N__35064),
            .in2(N__34933),
            .in3(N__39925),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12339_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11266_LC_3_14_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11266_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11266_LC_3_14_4 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11266_LC_3_14_4  (
            .in0(N__85322),
            .in1(N__90018),
            .in2(N__34930),
            .in3(N__34927),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6125_6126_LC_3_14_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6125_6126_LC_3_14_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6125_6126_LC_3_14_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6125_6126_LC_3_14_5  (
            .in0(N__46858),
            .in1(N__34920),
            .in2(_gnd_net_),
            .in3(N__67716),
            .lcout(REG_mem_63_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93248),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5645_5646_LC_3_14_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5645_5646_LC_3_14_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5645_5646_LC_3_14_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5645_5646_LC_3_14_6  (
            .in0(N__35073),
            .in1(N__46860),
            .in2(_gnd_net_),
            .in3(N__79989),
            .lcout(REG_mem_58_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93248),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5933_5934_LC_3_14_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5933_5934_LC_3_14_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5933_5934_LC_3_14_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5933_5934_LC_3_14_7  (
            .in0(N__46859),
            .in1(N__95644),
            .in2(N__35065),
            .in3(N__70974),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93248),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10181_3_lut_LC_3_15_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10181_3_lut_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10181_3_lut_LC_3_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10181_3_lut_LC_3_15_0  (
            .in0(N__87736),
            .in1(N__34996),
            .in2(_gnd_net_),
            .in3(N__35005),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11830_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11749_LC_3_15_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11749_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11749_LC_3_15_1 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11749_LC_3_15_1  (
            .in0(N__85230),
            .in1(N__91991),
            .in2(N__35050),
            .in3(N__42364),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i260_261_LC_3_15_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i260_261_LC_3_15_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i260_261_LC_3_15_2 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i260_261_LC_3_15_2  (
            .in0(N__48896),
            .in1(N__95632),
            .in2(N__35046),
            .in3(N__80601),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93256),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10143_3_lut_LC_3_15_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10143_3_lut_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10143_3_lut_LC_3_15_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10143_3_lut_LC_3_15_3  (
            .in0(N__38833),
            .in1(N__87735),
            .in2(_gnd_net_),
            .in3(N__36715),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11792_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13490_bdd_4_lut_LC_3_15_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13490_bdd_4_lut_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13490_bdd_4_lut_LC_3_15_4 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13490_bdd_4_lut_LC_3_15_4  (
            .in0(N__35029),
            .in1(N__85229),
            .in2(N__35023),
            .in3(N__35020),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3503_3504_LC_3_15_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3503_3504_LC_3_15_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3503_3504_LC_3_15_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3503_3504_LC_3_15_5  (
            .in0(N__35004),
            .in1(N__61250),
            .in2(_gnd_net_),
            .in3(N__54109),
            .lcout(REG_mem_36_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93256),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3599_3600_LC_3_15_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3599_3600_LC_3_15_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3599_3600_LC_3_15_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3599_3600_LC_3_15_6  (
            .in0(N__61249),
            .in1(N__34995),
            .in2(_gnd_net_),
            .in3(N__63729),
            .lcout(REG_mem_37_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93256),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i272_273_LC_3_15_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i272_273_LC_3_15_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i272_273_LC_3_15_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i272_273_LC_3_15_7  (
            .in0(N__95631),
            .in1(N__80594),
            .in2(N__35140),
            .in3(N__41671),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93256),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9882_3_lut_LC_3_16_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9882_3_lut_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9882_3_lut_LC_3_16_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9882_3_lut_LC_3_16_0  (
            .in0(N__38800),
            .in1(N__38782),
            .in2(_gnd_net_),
            .in3(N__87446),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11531_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12353_LC_3_16_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12353_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12353_LC_3_16_1 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12353_LC_3_16_1  (
            .in0(N__91786),
            .in1(N__36523),
            .in2(N__35125),
            .in3(N__85202),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9860_3_lut_LC_3_16_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9860_3_lut_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9860_3_lut_LC_3_16_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9860_3_lut_LC_3_16_2  (
            .in0(N__35914),
            .in1(N__87444),
            .in2(_gnd_net_),
            .in3(N__35085),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11509_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14186_bdd_4_lut_LC_3_16_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14186_bdd_4_lut_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14186_bdd_4_lut_LC_3_16_3 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14186_bdd_4_lut_LC_3_16_3  (
            .in0(N__35092),
            .in1(N__85201),
            .in2(N__35122),
            .in3(N__35119),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14189 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5738_5739_LC_3_16_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5738_5739_LC_3_16_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5738_5739_LC_3_16_4 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5738_5739_LC_3_16_4  (
            .in0(N__79793),
            .in1(N__35100),
            .in2(N__95771),
            .in3(N__46554),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93266),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2666_2667_LC_3_16_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2666_2667_LC_3_16_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2666_2667_LC_3_16_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2666_2667_LC_3_16_5  (
            .in0(N__46552),
            .in1(N__95735),
            .in2(N__36189),
            .in3(N__79794),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93266),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9861_3_lut_LC_3_16_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9861_3_lut_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9861_3_lut_LC_3_16_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9861_3_lut_LC_3_16_6  (
            .in0(N__35113),
            .in1(N__35101),
            .in2(_gnd_net_),
            .in3(N__87445),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11510 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5450_5451_LC_3_16_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5450_5451_LC_3_16_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5450_5451_LC_3_16_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5450_5451_LC_3_16_7  (
            .in0(N__46553),
            .in1(N__95736),
            .in2(N__35086),
            .in3(N__96013),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93266),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.usb3_data_in_latched__i12_LC_5_1_1 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i12_LC_5_1_1 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i12_LC_5_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i12_LC_5_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35215),
            .lcout(\usb3_if_inst.usb3_data_in_latched_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93334),
            .ce(),
            .sr(N__73747));
    defparam \usb3_if_inst.usb3_data_in_latched__i13_LC_5_1_3 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i13_LC_5_1_3 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i13_LC_5_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i13_LC_5_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35200),
            .lcout(\usb3_if_inst.usb3_data_in_latched_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93334),
            .ce(),
            .sr(N__73747));
    defparam \usb3_if_inst.dc32_fifo_data_in_i16_LC_5_2_7 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i16_LC_5_2_7 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i16_LC_5_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i16_LC_5_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35188),
            .lcout(dc32_fifo_data_in_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.dc32_fifo_data_in_i16C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11470_LC_5_3_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11470_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11470_LC_5_3_0 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11470_LC_5_3_0  (
            .in0(N__85812),
            .in1(N__36283),
            .in2(N__92665),
            .in3(N__36379),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13166_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13166_bdd_4_lut_LC_5_3_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13166_bdd_4_lut_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13166_bdd_4_lut_LC_5_3_1 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13166_bdd_4_lut_LC_5_3_1  (
            .in0(N__39472),
            .in1(N__85810),
            .in2(N__35179),
            .in3(N__35173),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13169_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_LC_5_3_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_LC_5_3_2 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_LC_5_3_2  (
            .in0(N__90347),
            .in1(N__35146),
            .in2(N__35176),
            .in3(N__81478),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10797_3_lut_LC_5_3_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10797_3_lut_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10797_3_lut_LC_5_3_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10797_3_lut_LC_5_3_3  (
            .in0(N__88337),
            .in1(N__35266),
            .in2(_gnd_net_),
            .in3(N__35275),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12446 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_LC_5_3_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_LC_5_3_4 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_LC_5_3_4  (
            .in0(N__92593),
            .in1(N__85813),
            .in2(N__35164),
            .in3(N__35482),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14330_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14330_bdd_4_lut_LC_5_3_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14330_bdd_4_lut_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14330_bdd_4_lut_LC_5_3_5 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14330_bdd_4_lut_LC_5_3_5  (
            .in0(N__35845),
            .in1(N__85811),
            .in2(N__35149),
            .in3(N__36442),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4865_4866_LC_5_3_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4865_4866_LC_5_3_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4865_4866_LC_5_3_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4865_4866_LC_5_3_6  (
            .in0(N__35274),
            .in1(N__56330),
            .in2(_gnd_net_),
            .in3(N__73054),
            .lcout(REG_mem_50_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93305),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4961_4962_LC_5_3_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4961_4962_LC_5_3_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4961_4962_LC_5_3_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4961_4962_LC_5_3_7  (
            .in0(N__56329),
            .in1(N__35265),
            .in2(_gnd_net_),
            .in3(N__72263),
            .lcout(REG_mem_51_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93305),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5363_5364_LC_5_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5363_5364_LC_5_4_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5363_5364_LC_5_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5363_5364_LC_5_4_0  (
            .in0(N__62273),
            .in1(N__35256),
            .in2(_gnd_net_),
            .in3(N__77247),
            .lcout(REG_mem_55_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10382_3_lut_LC_5_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10382_3_lut_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10382_3_lut_LC_5_4_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10382_3_lut_LC_5_4_1  (
            .in0(N__35238),
            .in1(N__88234),
            .in2(_gnd_net_),
            .in3(N__36597),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12031 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10383_3_lut_LC_5_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10383_3_lut_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10383_3_lut_LC_5_4_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10383_3_lut_LC_5_4_2  (
            .in0(N__35226),
            .in1(_gnd_net_),
            .in2(N__88535),
            .in3(N__35257),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12032_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11879_LC_5_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11879_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11879_LC_5_4_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11879_LC_5_4_3  (
            .in0(N__35248),
            .in1(N__85456),
            .in2(N__35242),
            .in3(N__92589),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1619_1620_LC_5_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1619_1620_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1619_1620_LC_5_4_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1619_1620_LC_5_4_4  (
            .in0(N__36429),
            .in1(_gnd_net_),
            .in2(N__62360),
            .in3(N__65685),
            .lcout(REG_mem_16_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5171_5172_LC_5_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5171_5172_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5171_5172_LC_5_4_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5171_5172_LC_5_4_5  (
            .in0(N__95538),
            .in1(N__62269),
            .in2(N__35239),
            .in3(N__77038),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5267_5268_LC_5_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5267_5268_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5267_5268_LC_5_4_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5267_5268_LC_5_4_6  (
            .in0(N__62268),
            .in1(N__95539),
            .in2(N__35227),
            .in3(N__76336),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4646_4647_LC_5_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4646_4647_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4646_4647_LC_5_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4646_4647_LC_5_4_7  (
            .in0(N__39342),
            .in1(N__71295),
            .in2(_gnd_net_),
            .in3(N__75576),
            .lcout(REG_mem_48_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93290),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10386_3_lut_LC_5_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10386_3_lut_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10386_3_lut_LC_5_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10386_3_lut_LC_5_5_0  (
            .in0(N__37123),
            .in1(N__35326),
            .in2(_gnd_net_),
            .in3(N__88233),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12035 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12273_LC_5_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12273_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12273_LC_5_5_1 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12273_LC_5_5_1  (
            .in0(N__35281),
            .in1(N__85815),
            .in2(N__92596),
            .in3(N__37693),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14150_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14150_bdd_4_lut_LC_5_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14150_bdd_4_lut_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14150_bdd_4_lut_LC_5_5_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14150_bdd_4_lut_LC_5_5_2  (
            .in0(N__85814),
            .in1(N__35338),
            .in2(N__35329),
            .in3(N__35299),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12083 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i449_450_LC_5_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i449_450_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i449_450_LC_5_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i449_450_LC_5_5_3  (
            .in0(N__37872),
            .in1(N__56353),
            .in2(_gnd_net_),
            .in3(N__72710),
            .lcout(REG_mem_4_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93278),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5747_5748_LC_5_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5747_5748_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5747_5748_LC_5_5_4 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5747_5748_LC_5_5_4  (
            .in0(N__79739),
            .in1(N__35325),
            .in2(N__95703),
            .in3(N__62357),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93278),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2675_2676_LC_5_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2675_2676_LC_5_5_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2675_2676_LC_5_5_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2675_2676_LC_5_5_5  (
            .in0(N__62355),
            .in1(N__95540),
            .in2(N__35316),
            .in3(N__79740),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93278),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10385_3_lut_LC_5_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10385_3_lut_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10385_3_lut_LC_5_5_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10385_3_lut_LC_5_5_6  (
            .in0(N__36076),
            .in1(N__88232),
            .in2(_gnd_net_),
            .in3(N__35292),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12034 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5459_5460_LC_5_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5459_5460_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5459_5460_LC_5_5_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5459_5460_LC_5_5_7  (
            .in0(N__62356),
            .in1(N__95541),
            .in2(N__35293),
            .in3(N__96006),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93278),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10394_3_lut_LC_5_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10394_3_lut_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10394_3_lut_LC_5_6_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10394_3_lut_LC_5_6_0  (
            .in0(N__35803),
            .in1(_gnd_net_),
            .in2(N__88534),
            .in3(N__36643),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12043 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5921_5922_LC_5_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5921_5922_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5921_5922_LC_5_6_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5921_5922_LC_5_6_1  (
            .in0(N__95531),
            .in1(N__35397),
            .in2(N__56568),
            .in3(N__70950),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5030_5031_LC_5_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5030_5031_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5030_5031_LC_5_6_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5030_5031_LC_5_6_2  (
            .in0(N__71456),
            .in1(N__95533),
            .in2(N__39423),
            .in3(N__77467),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2771_2772_LC_5_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2771_2772_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2771_2772_LC_5_6_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2771_2772_LC_5_6_3  (
            .in0(N__95530),
            .in1(N__62218),
            .in2(N__35382),
            .in3(N__70663),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4097_4098_LC_5_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4097_4098_LC_5_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4097_4098_LC_5_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4097_4098_LC_5_6_4  (
            .in0(N__35538),
            .in1(N__56490),
            .in2(_gnd_net_),
            .in3(N__68085),
            .lcout(REG_mem_42_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10025_3_lut_LC_5_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10025_3_lut_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10025_3_lut_LC_5_6_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10025_3_lut_LC_5_6_5  (
            .in0(N__39588),
            .in1(N__88228),
            .in2(_gnd_net_),
            .in3(N__36657),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11674 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2195_2196_LC_5_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2195_2196_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2195_2196_LC_5_6_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2195_2196_LC_5_6_6  (
            .in0(N__62216),
            .in1(N__95532),
            .in2(N__36403),
            .in3(N__76325),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2387_2388_LC_5_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2387_2388_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2387_2388_LC_5_6_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2387_2388_LC_5_6_7  (
            .in0(N__95529),
            .in1(N__62217),
            .in2(N__35358),
            .in3(N__96007),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93267),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12854_bdd_4_lut_LC_5_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12854_bdd_4_lut_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12854_bdd_4_lut_LC_5_7_0 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12854_bdd_4_lut_LC_5_7_0  (
            .in0(N__92594),
            .in1(N__39673),
            .in2(N__45289),
            .in3(N__35527),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12857_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9852_3_lut_LC_5_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9852_3_lut_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9852_3_lut_LC_5_7_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9852_3_lut_LC_5_7_1  (
            .in0(N__85723),
            .in1(_gnd_net_),
            .in2(N__35341),
            .in3(N__37135),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11201_LC_5_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11201_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11201_LC_5_7_2 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11201_LC_5_7_2  (
            .in0(N__92595),
            .in1(N__43465),
            .in2(N__35542),
            .in3(N__87425),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12854 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4676_4677_LC_5_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4676_4677_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4676_4677_LC_5_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4676_4677_LC_5_7_3  (
            .in0(N__35424),
            .in1(N__48708),
            .in2(_gnd_net_),
            .in3(N__75558),
            .lcout(REG_mem_48_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93257),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9851_3_lut_LC_5_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9851_3_lut_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9851_3_lut_LC_5_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9851_3_lut_LC_5_7_4  (
            .in0(N__37765),
            .in1(N__35521),
            .in2(_gnd_net_),
            .in3(N__85722),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11500_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14300_bdd_4_lut_LC_5_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14300_bdd_4_lut_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14300_bdd_4_lut_LC_5_7_5 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14300_bdd_4_lut_LC_5_7_5  (
            .in0(N__35503),
            .in1(N__35491),
            .in2(N__35485),
            .in3(N__81442),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10818_3_lut_LC_5_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10818_3_lut_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10818_3_lut_LC_5_7_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10818_3_lut_LC_5_7_6  (
            .in0(N__35638),
            .in1(N__87424),
            .in2(_gnd_net_),
            .in3(N__35665),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13124_bdd_4_lut_LC_5_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13124_bdd_4_lut_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13124_bdd_4_lut_LC_5_8_0 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13124_bdd_4_lut_LC_5_8_0  (
            .in0(N__36556),
            .in1(N__92414),
            .in2(N__35650),
            .in3(N__38212),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5156_5157_LC_5_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5156_5157_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5156_5157_LC_5_8_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5156_5157_LC_5_8_1  (
            .in0(N__48751),
            .in1(N__95409),
            .in2(N__35454),
            .in3(N__76911),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93249),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11291_LC_5_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11291_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11291_LC_5_8_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11291_LC_5_8_2  (
            .in0(N__36784),
            .in1(N__92415),
            .in2(N__35620),
            .in3(N__87886),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12962 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13022_bdd_4_lut_LC_5_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13022_bdd_4_lut_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13022_bdd_4_lut_LC_5_8_3 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13022_bdd_4_lut_LC_5_8_3  (
            .in0(N__92413),
            .in1(N__36880),
            .in2(N__35605),
            .in3(N__35425),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13025 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1712_1713_LC_5_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1712_1713_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1712_1713_LC_5_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1712_1713_LC_5_8_4  (
            .in0(N__36837),
            .in1(N__41751),
            .in2(_gnd_net_),
            .in3(N__66573),
            .lcout(REG_mem_17_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93249),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5348_5349_LC_5_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5348_5349_LC_5_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5348_5349_LC_5_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5348_5349_LC_5_8_5  (
            .in0(N__35616),
            .in1(N__48711),
            .in2(_gnd_net_),
            .in3(N__77236),
            .lcout(REG_mem_55_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93249),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4772_4773_LC_5_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4772_4773_LC_5_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4772_4773_LC_5_8_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4772_4773_LC_5_8_6  (
            .in0(N__48710),
            .in1(N__62983),
            .in2(_gnd_net_),
            .in3(N__35601),
            .lcout(REG_mem_49_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93249),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11720_LC_5_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11720_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11720_LC_5_8_7 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11720_LC_5_8_7  (
            .in0(N__85348),
            .in1(N__35593),
            .in2(N__92597),
            .in3(N__35812),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1328_1329_LC_5_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1328_1329_LC_5_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1328_1329_LC_5_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1328_1329_LC_5_9_0  (
            .in0(N__41745),
            .in1(N__35583),
            .in2(_gnd_net_),
            .in3(N__70138),
            .lcout(REG_mem_13_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93242),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11894_LC_5_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11894_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11894_LC_5_9_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11894_LC_5_9_1  (
            .in0(N__35551),
            .in1(N__92320),
            .in2(N__35731),
            .in3(N__87715),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13664_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13664_bdd_4_lut_LC_5_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13664_bdd_4_lut_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13664_bdd_4_lut_LC_5_9_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13664_bdd_4_lut_LC_5_9_2  (
            .in0(N__92319),
            .in1(N__35584),
            .in2(N__35575),
            .in3(N__35560),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1232_1233_LC_5_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1232_1233_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1232_1233_LC_5_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1232_1233_LC_5_9_3  (
            .in0(N__35559),
            .in1(N__41744),
            .in2(_gnd_net_),
            .in3(N__59601),
            .lcout(REG_mem_12_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93242),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1424_1425_LC_5_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1424_1425_LC_5_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1424_1425_LC_5_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1424_1425_LC_5_9_4  (
            .in0(N__41746),
            .in1(N__35550),
            .in2(_gnd_net_),
            .in3(N__74765),
            .lcout(REG_mem_14_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93242),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1520_1521_LC_5_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1520_1521_LC_5_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1520_1521_LC_5_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1520_1521_LC_5_9_5  (
            .in0(N__35727),
            .in1(N__41747),
            .in2(_gnd_net_),
            .in3(N__64007),
            .lcout(REG_mem_15_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93242),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4385_4386_LC_5_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4385_4386_LC_5_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4385_4386_LC_5_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4385_4386_LC_5_9_6  (
            .in0(N__37146),
            .in1(N__56565),
            .in2(_gnd_net_),
            .in3(N__71865),
            .lcout(REG_mem_45_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93242),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6029_6030_LC_5_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6029_6030_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6029_6030_LC_5_9_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6029_6030_LC_5_9_7  (
            .in0(N__46899),
            .in1(N__94876),
            .in2(N__35706),
            .in3(N__77841),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93242),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10368_3_lut_LC_5_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10368_3_lut_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10368_3_lut_LC_5_10_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10368_3_lut_LC_5_10_0  (
            .in0(N__87713),
            .in1(N__39874),
            .in2(_gnd_net_),
            .in3(N__36994),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12017 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2858_2859_LC_5_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2858_2859_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2858_2859_LC_5_10_1 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2858_2859_LC_5_10_1  (
            .in0(N__46406),
            .in1(N__94831),
            .in2(N__36024),
            .in3(N__70860),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1199_1200_LC_5_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1199_1200_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1199_1200_LC_5_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1199_1200_LC_5_10_2  (
            .in0(N__61286),
            .in1(N__37101),
            .in2(_gnd_net_),
            .in3(N__59632),
            .lcout(REG_mem_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6095_6096_LC_5_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6095_6096_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6095_6096_LC_5_10_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6095_6096_LC_5_10_3  (
            .in0(N__35676),
            .in1(N__61287),
            .in2(_gnd_net_),
            .in3(N__67670),
            .lcout(REG_mem_63_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6113_6114_LC_5_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6113_6114_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6113_6114_LC_5_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6113_6114_LC_5_10_4  (
            .in0(N__67671),
            .in1(N__35661),
            .in2(_gnd_net_),
            .in3(N__56567),
            .lcout(REG_mem_63_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11430_LC_5_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11430_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11430_LC_5_10_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11430_LC_5_10_5  (
            .in0(N__37008),
            .in1(N__92010),
            .in2(N__42013),
            .in3(N__87714),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6017_6018_LC_5_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6017_6018_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6017_6018_LC_5_10_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6017_6018_LC_5_10_6  (
            .in0(N__94830),
            .in1(N__56566),
            .in2(N__35637),
            .in3(N__77833),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1508_1509_LC_5_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1508_1509_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1508_1509_LC_5_10_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1508_1509_LC_5_10_7  (
            .in0(N__38388),
            .in1(N__48744),
            .in2(_gnd_net_),
            .in3(N__64008),
            .lcout(REG_mem_15_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93232),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10815_3_lut_LC_5_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10815_3_lut_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10815_3_lut_LC_5_11_0 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10815_3_lut_LC_5_11_0  (
            .in0(N__35823),
            .in1(N__35836),
            .in2(N__88371),
            .in3(_gnd_net_),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12464 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5633_5634_LC_5_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5633_5634_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5633_5634_LC_5_11_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5633_5634_LC_5_11_1  (
            .in0(N__56512),
            .in1(N__35835),
            .in2(_gnd_net_),
            .in3(N__79970),
            .lcout(REG_mem_58_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93243),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5729_5730_LC_5_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5729_5730_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5729_5730_LC_5_11_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5729_5730_LC_5_11_2  (
            .in0(N__94970),
            .in1(N__56513),
            .in2(N__35824),
            .in3(N__79743),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93243),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10026_3_lut_LC_5_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10026_3_lut_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10026_3_lut_LC_5_11_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10026_3_lut_LC_5_11_3  (
            .in0(N__36631),
            .in1(N__88097),
            .in2(_gnd_net_),
            .in3(N__40192),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11675 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5939_5940_LC_5_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5939_5940_LC_5_11_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5939_5940_LC_5_11_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5939_5940_LC_5_11_4  (
            .in0(N__94971),
            .in1(N__62400),
            .in2(N__35802),
            .in3(N__70928),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93243),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3152_3153_LC_5_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3152_3153_LC_5_11_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3152_3153_LC_5_11_5 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3152_3153_LC_5_11_5  (
            .in0(N__41801),
            .in1(N__94972),
            .in2(N__35781),
            .in3(N__82909),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93243),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1211_1212_LC_5_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1211_1212_LC_5_11_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1211_1212_LC_5_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1211_1212_LC_5_11_6  (
            .in0(N__35757),
            .in1(N__63398),
            .in2(_gnd_net_),
            .in3(N__59633),
            .lcout(REG_mem_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93243),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i836_837_LC_5_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i836_837_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i836_837_LC_5_11_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i836_837_LC_5_11_7  (
            .in0(N__35742),
            .in1(N__48755),
            .in2(_gnd_net_),
            .in3(N__67322),
            .lcout(REG_mem_8_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93243),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11480_LC_5_12_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11480_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11480_LC_5_12_0 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11480_LC_5_12_0  (
            .in0(N__92006),
            .in1(N__87581),
            .in2(N__37078),
            .in3(N__37363),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13184_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13184_bdd_4_lut_LC_5_12_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13184_bdd_4_lut_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13184_bdd_4_lut_LC_5_12_1 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13184_bdd_4_lut_LC_5_12_1  (
            .in0(N__42172),
            .in1(N__92004),
            .in2(N__35863),
            .in3(N__40042),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11226_LC_5_12_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11226_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11226_LC_5_12_2 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11226_LC_5_12_2  (
            .in0(N__92005),
            .in1(N__87580),
            .in2(N__45688),
            .in3(N__45544),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12890_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12890_bdd_4_lut_LC_5_12_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12890_bdd_4_lut_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12890_bdd_4_lut_LC_5_12_3 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12890_bdd_4_lut_LC_5_12_3  (
            .in0(N__39976),
            .in1(N__92003),
            .in2(N__35860),
            .in3(N__45241),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12893_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12448_LC_5_12_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12448_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12448_LC_5_12_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12448_LC_5_12_4  (
            .in0(N__35857),
            .in1(N__90101),
            .in2(N__35848),
            .in3(N__85241),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12168_LC_5_12_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12168_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12168_LC_5_12_5 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12168_LC_5_12_5  (
            .in0(N__87582),
            .in1(N__92007),
            .in2(N__36979),
            .in3(N__41425),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14024 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10649_3_lut_LC_5_12_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10649_3_lut_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10649_3_lut_LC_5_12_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10649_3_lut_LC_5_12_6  (
            .in0(N__35938),
            .in1(N__87579),
            .in2(_gnd_net_),
            .in3(N__40279),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4298_4299_LC_5_13_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4298_4299_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4298_4299_LC_5_13_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4298_4299_LC_5_13_0  (
            .in0(N__37413),
            .in1(N__46483),
            .in2(_gnd_net_),
            .in3(N__71755),
            .lcout(REG_mem_44_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2090_2091_LC_5_13_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2090_2091_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2090_2091_LC_5_13_1 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2090_2091_LC_5_13_1  (
            .in0(N__95347),
            .in1(N__46407),
            .in2(N__35979),
            .in3(N__77041),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12173_LC_5_13_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12173_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12173_LC_5_13_2 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12173_LC_5_13_2  (
            .in0(N__36054),
            .in1(N__91993),
            .in2(N__35926),
            .in3(N__87578),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14030_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14030_bdd_4_lut_LC_5_13_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14030_bdd_4_lut_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14030_bdd_4_lut_LC_5_13_3 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14030_bdd_4_lut_LC_5_13_3  (
            .in0(N__38332),
            .in1(N__91775),
            .in2(N__35956),
            .in3(N__35896),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14024_bdd_4_lut_LC_5_13_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14024_bdd_4_lut_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14024_bdd_4_lut_LC_5_13_4 .LUT_INIT=16'b1111101000001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14024_bdd_4_lut_LC_5_13_4  (
            .in0(N__38476),
            .in1(N__38560),
            .in2(N__92131),
            .in3(N__35953),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i554_555_LC_5_13_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i554_555_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i554_555_LC_5_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i554_555_LC_5_13_5  (
            .in0(N__46482),
            .in1(N__35937),
            .in2(_gnd_net_),
            .in3(N__67887),
            .lcout(REG_mem_5_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2573_2574_LC_5_13_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2573_2574_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2573_2574_LC_5_13_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2573_2574_LC_5_13_6  (
            .in0(N__35922),
            .in1(N__46994),
            .in2(_gnd_net_),
            .in3(N__70373),
            .lcout(REG_mem_26_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2762_2763_LC_5_13_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2762_2763_LC_5_13_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2762_2763_LC_5_13_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2762_2763_LC_5_13_7  (
            .in0(N__95348),
            .in1(N__46408),
            .in2(N__36003),
            .in3(N__70716),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93258),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10644_3_lut_LC_5_14_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10644_3_lut_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10644_3_lut_LC_5_14_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10644_3_lut_LC_5_14_0  (
            .in0(N__87431),
            .in1(N__37206),
            .in2(_gnd_net_),
            .in3(N__37192),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5546_5547_LC_5_14_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5546_5547_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5546_5547_LC_5_14_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5546_5547_LC_5_14_1  (
            .in0(N__97037),
            .in1(N__35907),
            .in2(N__95410),
            .in3(N__46409),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2477_2478_LC_5_14_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2477_2478_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2477_2478_LC_5_14_2 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2477_2478_LC_5_14_2  (
            .in0(N__46984),
            .in1(N__94978),
            .in2(N__35895),
            .in3(N__97040),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5549_5550_LC_5_14_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5549_5550_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5549_5550_LC_5_14_3 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5549_5550_LC_5_14_3  (
            .in0(N__97038),
            .in1(N__35874),
            .in2(N__95411),
            .in3(N__46986),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2483_2484_LC_5_14_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2483_2484_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2483_2484_LC_5_14_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2483_2484_LC_5_14_4  (
            .in0(N__62329),
            .in1(N__94979),
            .in2(N__36093),
            .in3(N__97041),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5555_5556_LC_5_14_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5555_5556_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5555_5556_LC_5_14_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5555_5556_LC_5_14_5  (
            .in0(N__97039),
            .in1(N__36066),
            .in2(N__95412),
            .in3(N__62330),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2669_2670_LC_5_14_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2669_2670_LC_5_14_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2669_2670_LC_5_14_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2669_2670_LC_5_14_6  (
            .in0(N__46985),
            .in1(N__94980),
            .in2(N__36055),
            .in3(N__79797),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5741_5742_LC_5_14_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5741_5742_LC_5_14_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5741_5742_LC_5_14_7 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5741_5742_LC_5_14_7  (
            .in0(N__79796),
            .in1(N__36036),
            .in2(N__95413),
            .in3(N__46987),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93268),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11216_LC_5_15_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11216_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11216_LC_5_15_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11216_LC_5_15_0  (
            .in0(N__39049),
            .in1(N__91590),
            .in2(N__37438),
            .in3(N__87301),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12878_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12878_bdd_4_lut_LC_5_15_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12878_bdd_4_lut_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12878_bdd_4_lut_LC_5_15_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12878_bdd_4_lut_LC_5_15_1  (
            .in0(N__91587),
            .in1(N__36025),
            .in2(N__36007),
            .in3(N__36004),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12881_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11420_LC_5_15_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11420_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11420_LC_5_15_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11420_LC_5_15_2  (
            .in0(N__36169),
            .in1(N__90035),
            .in2(N__35986),
            .in3(N__85110),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13094_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13094_bdd_4_lut_LC_5_15_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13094_bdd_4_lut_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13094_bdd_4_lut_LC_5_15_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13094_bdd_4_lut_LC_5_15_3  (
            .in0(N__90034),
            .in1(N__35962),
            .in2(N__35983),
            .in3(N__40321),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13097 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13208_bdd_4_lut_LC_5_15_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13208_bdd_4_lut_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13208_bdd_4_lut_LC_5_15_4 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13208_bdd_4_lut_LC_5_15_4  (
            .in0(N__38440),
            .in1(N__91589),
            .in2(N__36277),
            .in3(N__35980),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11400_LC_5_15_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11400_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11400_LC_5_15_5 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11400_LC_5_15_5  (
            .in0(N__87302),
            .in1(N__36193),
            .in2(N__91990),
            .in3(N__36265),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13100_bdd_4_lut_LC_5_15_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13100_bdd_4_lut_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13100_bdd_4_lut_LC_5_15_6 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13100_bdd_4_lut_LC_5_15_6  (
            .in0(N__37513),
            .in1(N__91588),
            .in2(N__36172),
            .in3(N__38194),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13220_bdd_4_lut_LC_5_16_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13220_bdd_4_lut_LC_5_16_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13220_bdd_4_lut_LC_5_16_0 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13220_bdd_4_lut_LC_5_16_0  (
            .in0(N__85227),
            .in1(N__36145),
            .in2(N__36214),
            .in3(N__36163),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11510_LC_5_16_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11510_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11510_LC_5_16_1 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11510_LC_5_16_1  (
            .in0(N__36154),
            .in1(N__85228),
            .in2(N__92130),
            .in3(N__44293),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13220 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10021_3_lut_LC_5_16_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10021_3_lut_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10021_3_lut_LC_5_16_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10021_3_lut_LC_5_16_2  (
            .in0(N__36139),
            .in1(N__90065),
            .in2(_gnd_net_),
            .in3(N__39106),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11670_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12403_LC_5_16_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12403_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12403_LC_5_16_3 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12403_LC_5_16_3  (
            .in0(N__80993),
            .in1(N__37264),
            .in2(N__36130),
            .in3(N__81348),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14054 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9927_3_lut_LC_5_16_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9927_3_lut_LC_5_16_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9927_3_lut_LC_5_16_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9927_3_lut_LC_5_16_4  (
            .in0(N__85226),
            .in1(N__44137),
            .in2(_gnd_net_),
            .in3(N__45658),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11576_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9928_3_lut_LC_5_16_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9928_3_lut_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9928_3_lut_LC_5_16_5 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9928_3_lut_LC_5_16_5  (
            .in0(N__90066),
            .in1(N__36127),
            .in2(N__36121),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11577_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i13_LC_5_16_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i13_LC_5_16_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i13_LC_5_16_6 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i13_LC_5_16_6  (
            .in0(N__36118),
            .in1(N__80992),
            .in2(N__36112),
            .in3(N__36109),
            .lcout(REG_out_raw_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97343),
            .ce(N__80867),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11505_LC_5_17_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11505_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11505_LC_5_17_0 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11505_LC_5_17_0  (
            .in0(N__87430),
            .in1(N__91784),
            .in2(N__36250),
            .in3(N__38851),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2570_2571_LC_5_17_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2570_2571_LC_5_17_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2570_2571_LC_5_17_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2570_2571_LC_5_17_1  (
            .in0(N__36261),
            .in1(N__46539),
            .in2(_gnd_net_),
            .in3(N__70374),
            .lcout(REG_mem_26_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93304),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2186_2187_LC_5_17_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2186_2187_LC_5_17_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2186_2187_LC_5_17_2 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2186_2187_LC_5_17_2  (
            .in0(N__46538),
            .in1(N__95633),
            .in2(N__36249),
            .in3(N__76323),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93304),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5258_5259_LC_5_17_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5258_5259_LC_5_17_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5258_5259_LC_5_17_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5258_5259_LC_5_17_3  (
            .in0(N__76324),
            .in1(N__46541),
            .in2(N__36235),
            .in3(N__95630),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93304),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5354_5355_LC_5_17_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5354_5355_LC_5_17_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5354_5355_LC_5_17_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5354_5355_LC_5_17_5  (
            .in0(N__36222),
            .in1(N__46540),
            .in2(_gnd_net_),
            .in3(N__77248),
            .lcout(REG_mem_55_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93304),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10869_3_lut_LC_5_17_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10869_3_lut_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10869_3_lut_LC_5_17_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10869_3_lut_LC_5_17_6  (
            .in0(N__87429),
            .in1(N__36234),
            .in2(_gnd_net_),
            .in3(N__36223),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10643_3_lut_LC_5_17_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10643_3_lut_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10643_3_lut_LC_5_17_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10643_3_lut_LC_5_17_7  (
            .in0(N__40093),
            .in1(N__87428),
            .in2(_gnd_net_),
            .in3(N__40633),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.usb3_data_in_latched__i11_LC_6_1_4 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i11_LC_6_1_4 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i11_LC_6_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i11_LC_6_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36205),
            .lcout(\usb3_if_inst.usb3_data_in_latched_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93335),
            .ce(),
            .sr(N__73754));
    defparam \usb3_if_inst.state_FSM_i5_LC_6_2_0 .C_ON=1'b0;
    defparam \usb3_if_inst.state_FSM_i5_LC_6_2_0 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.state_FSM_i5_LC_6_2_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \usb3_if_inst.state_FSM_i5_LC_6_2_0  (
            .in0(N__73708),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57261),
            .lcout(\usb3_if_inst.n551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_FSM_i5C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.dc32_fifo_data_in_i1_LC_6_2_1 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i1_LC_6_2_1 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i1_LC_6_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i1_LC_6_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44887),
            .lcout(dc32_fifo_data_in_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_FSM_i5C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.dc32_fifo_data_in_i10_LC_6_2_2 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i10_LC_6_2_2 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i10_LC_6_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i10_LC_6_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37711),
            .lcout(dc32_fifo_data_in_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_FSM_i5C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.dc32_fifo_data_in_i11_LC_6_2_3 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i11_LC_6_2_3 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i11_LC_6_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i11_LC_6_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36325),
            .lcout(dc32_fifo_data_in_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_FSM_i5C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.dc32_fifo_data_in_i12_LC_6_2_4 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i12_LC_6_2_4 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i12_LC_6_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i12_LC_6_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36319),
            .lcout(dc32_fifo_data_in_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_FSM_i5C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.dc32_fifo_data_in_i13_LC_6_2_5 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i13_LC_6_2_5 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i13_LC_6_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i13_LC_6_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36313),
            .lcout(dc32_fifo_data_in_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_FSM_i5C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.dc32_fifo_data_in_i14_LC_6_2_6 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i14_LC_6_2_6 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i14_LC_6_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i14_LC_6_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36307),
            .lcout(dc32_fifo_data_in_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_FSM_i5C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4115_4116_LC_6_3_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4115_4116_LC_6_3_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4115_4116_LC_6_3_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4115_4116_LC_6_3_0  (
            .in0(N__37827),
            .in1(N__62244),
            .in2(_gnd_net_),
            .in3(N__68087),
            .lcout(REG_mem_42_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4211_4212_LC_6_3_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4211_4212_LC_6_3_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4211_4212_LC_6_3_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4211_4212_LC_6_3_1  (
            .in0(N__62243),
            .in1(N__37815),
            .in2(_gnd_net_),
            .in3(N__68299),
            .lcout(REG_mem_43_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5249_5250_LC_6_3_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5249_5250_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5249_5250_LC_6_3_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5249_5250_LC_6_3_2  (
            .in0(N__76307),
            .in1(N__56332),
            .in2(N__36295),
            .in3(N__95720),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10812_3_lut_LC_6_3_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10812_3_lut_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10812_3_lut_LC_6_3_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10812_3_lut_LC_6_3_3  (
            .in0(N__88336),
            .in1(N__36294),
            .in2(_gnd_net_),
            .in3(N__36370),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12461 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5345_5346_LC_6_3_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5345_5346_LC_6_3_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5345_5346_LC_6_3_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5345_5346_LC_6_3_4  (
            .in0(N__36369),
            .in1(N__56331),
            .in2(_gnd_net_),
            .in3(N__77231),
            .lcout(REG_mem_55_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i176_177_LC_6_3_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i176_177_LC_6_3_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i176_177_LC_6_3_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i176_177_LC_6_3_5  (
            .in0(N__41612),
            .in1(N__95718),
            .in2(N__41025),
            .in3(N__80319),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2054_2055_LC_6_3_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2054_2055_LC_6_3_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2054_2055_LC_6_3_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2054_2055_LC_6_3_6  (
            .in0(N__95717),
            .in1(N__71330),
            .in2(N__37666),
            .in3(N__76976),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5237_5238_LC_6_3_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5237_5238_LC_6_3_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5237_5238_LC_6_3_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5237_5238_LC_6_3_7  (
            .in0(N__62852),
            .in1(N__95719),
            .in2(N__47973),
            .in3(N__76306),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93307),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2561_2562_LC_6_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2561_2562_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2561_2562_LC_6_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2561_2562_LC_6_4_0  (
            .in0(N__36360),
            .in1(N__56352),
            .in2(_gnd_net_),
            .in3(N__70384),
            .lcout(REG_mem_26_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11345_LC_6_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11345_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11345_LC_6_4_1 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11345_LC_6_4_1  (
            .in0(N__88054),
            .in1(N__36361),
            .in2(N__92668),
            .in3(N__36468),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13028_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13028_bdd_4_lut_LC_6_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13028_bdd_4_lut_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13028_bdd_4_lut_LC_6_4_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13028_bdd_4_lut_LC_6_4_2  (
            .in0(N__36336),
            .in1(N__92605),
            .in2(N__36352),
            .in3(N__36348),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13031 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2465_2466_LC_6_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2465_2466_LC_6_4_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2465_2466_LC_6_4_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2465_2466_LC_6_4_3  (
            .in0(N__95534),
            .in1(N__56518),
            .in2(N__36349),
            .in3(N__97034),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2369_2370_LC_6_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2369_2370_LC_6_4_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2369_2370_LC_6_4_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2369_2370_LC_6_4_4  (
            .in0(N__56516),
            .in1(N__95536),
            .in2(N__36337),
            .in3(N__95998),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2657_2658_LC_6_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2657_2658_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2657_2658_LC_6_4_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2657_2658_LC_6_4_5  (
            .in0(N__95535),
            .in1(N__56519),
            .in2(N__36469),
            .in3(N__79746),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5441_5442_LC_6_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5441_5442_LC_6_4_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5441_5442_LC_6_4_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5441_5442_LC_6_4_6  (
            .in0(N__56517),
            .in1(N__95537),
            .in2(N__36454),
            .in3(N__95999),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93292),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10814_3_lut_LC_6_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10814_3_lut_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10814_3_lut_LC_6_4_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10814_3_lut_LC_6_4_7  (
            .in0(N__88053),
            .in1(N__38143),
            .in2(_gnd_net_),
            .in3(N__36453),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12463 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12830_bdd_4_lut_LC_6_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12830_bdd_4_lut_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12830_bdd_4_lut_LC_6_5_0 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12830_bdd_4_lut_LC_6_5_0  (
            .in0(N__37936),
            .in1(N__92420),
            .in2(N__36610),
            .in3(N__36430),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12833_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10421_3_lut_LC_6_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10421_3_lut_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10421_3_lut_LC_6_5_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10421_3_lut_LC_6_5_1  (
            .in0(N__36385),
            .in1(_gnd_net_),
            .in2(N__36418),
            .in3(N__85515),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12070 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11148_LC_6_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11148_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11148_LC_6_5_2 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11148_LC_6_5_2  (
            .in0(N__92567),
            .in1(N__36402),
            .in2(N__41401),
            .in3(N__88051),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12788_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12788_bdd_4_lut_LC_6_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12788_bdd_4_lut_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12788_bdd_4_lut_LC_6_5_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12788_bdd_4_lut_LC_6_5_3  (
            .in0(N__92419),
            .in1(N__41944),
            .in2(N__36388),
            .in3(N__39757),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10811_3_lut_LC_6_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10811_3_lut_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10811_3_lut_LC_6_5_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10811_3_lut_LC_6_5_4  (
            .in0(N__38233),
            .in1(N__88050),
            .in2(_gnd_net_),
            .in3(N__36537),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12460 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11166_LC_6_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11166_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11166_LC_6_5_5 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11166_LC_6_5_5  (
            .in0(N__88052),
            .in1(N__37891),
            .in2(N__92598),
            .in3(N__53689),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12812 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1715_1716_LC_6_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1715_1716_LC_6_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1715_1716_LC_6_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1715_1716_LC_6_5_6  (
            .in0(N__36606),
            .in1(N__62359),
            .in2(_gnd_net_),
            .in3(N__66582),
            .lcout(REG_mem_17_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93280),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5075_5076_LC_6_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5075_5076_LC_6_5_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5075_5076_LC_6_5_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5075_5076_LC_6_5_7  (
            .in0(N__62358),
            .in1(N__95342),
            .in2(N__36598),
            .in3(N__77465),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93280),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5732_5733_LC_6_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5732_5733_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5732_5733_LC_6_6_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5732_5733_LC_6_6_0  (
            .in0(N__95336),
            .in1(N__48692),
            .in2(N__36573),
            .in3(N__79702),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5894_5895_LC_6_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5894_5895_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5894_5895_LC_6_6_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5894_5895_LC_6_6_1  (
            .in0(N__71329),
            .in1(N__95338),
            .in2(N__36675),
            .in3(N__70949),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5135_5136_LC_6_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5135_5136_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5135_5136_LC_6_6_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5135_5136_LC_6_6_2  (
            .in0(N__61404),
            .in1(N__95334),
            .in2(N__36555),
            .in3(N__76917),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4175_4176_LC_6_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4175_4176_LC_6_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4175_4176_LC_6_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4175_4176_LC_6_6_3  (
            .in0(N__36954),
            .in1(N__61403),
            .in2(_gnd_net_),
            .in3(N__68288),
            .lcout(REG_mem_43_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5153_5154_LC_6_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5153_5154_LC_6_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5153_5154_LC_6_6_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5153_5154_LC_6_6_4  (
            .in0(N__95335),
            .in1(N__56520),
            .in2(N__36538),
            .in3(N__76918),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9881_3_lut_LC_6_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9881_3_lut_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9881_3_lut_LC_6_6_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9881_3_lut_LC_6_6_5  (
            .in0(N__39568),
            .in1(N__88044),
            .in2(_gnd_net_),
            .in3(N__36504),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5834_5835_LC_6_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5834_5835_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5834_5835_LC_6_6_6 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5834_5835_LC_6_6_6  (
            .in0(N__46308),
            .in1(N__70705),
            .in2(N__95626),
            .in3(N__36505),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2867_2868_LC_6_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2867_2868_LC_6_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2867_2868_LC_6_6_7 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2867_2868_LC_6_6_7  (
            .in0(N__62407),
            .in1(N__95337),
            .in2(N__36486),
            .in3(N__70948),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93270),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2963_2964_LC_6_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2963_2964_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2963_2964_LC_6_7_0 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2963_2964_LC_6_7_0  (
            .in0(N__95218),
            .in1(N__36726),
            .in2(N__62429),
            .in3(N__77832),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3407_3408_LC_6_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3407_3408_LC_6_7_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3407_3408_LC_6_7_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3407_3408_LC_6_7_1  (
            .in0(N__61333),
            .in1(N__95220),
            .in2(N__36708),
            .in3(N__83344),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10541_3_lut_LC_6_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10541_3_lut_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10541_3_lut_LC_6_7_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10541_3_lut_LC_6_7_2  (
            .in0(N__36910),
            .in1(N__87422),
            .in2(_gnd_net_),
            .in3(N__38293),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9999_3_lut_LC_6_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9999_3_lut_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9999_3_lut_LC_6_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9999_3_lut_LC_6_7_3  (
            .in0(N__87423),
            .in1(N__43021),
            .in2(_gnd_net_),
            .in3(N__36850),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11648 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10367_3_lut_LC_6_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10367_3_lut_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10367_3_lut_LC_6_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10367_3_lut_LC_6_7_4  (
            .in0(N__36676),
            .in1(N__87421),
            .in2(_gnd_net_),
            .in3(N__41989),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2063_2064_LC_6_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2063_2064_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2063_2064_LC_6_7_5 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2063_2064_LC_6_7_5  (
            .in0(N__76915),
            .in1(N__61340),
            .in2(N__36658),
            .in3(N__95222),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3143_3144_LC_6_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3143_3144_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3143_3144_LC_6_7_6 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3143_3144_LC_6_7_6  (
            .in0(N__95219),
            .in1(N__37236),
            .in2(N__47296),
            .in3(N__82908),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5843_5844_LC_6_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5843_5844_LC_6_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5843_5844_LC_6_7_7 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5843_5844_LC_6_7_7  (
            .in0(N__36642),
            .in1(N__95221),
            .in2(N__70717),
            .in3(N__62411),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93260),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2255_2256_LC_6_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2255_2256_LC_6_8_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2255_2256_LC_6_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2255_2256_LC_6_8_0  (
            .in0(N__36621),
            .in1(N__61349),
            .in2(_gnd_net_),
            .in3(N__75049),
            .lcout(REG_mem_23_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1775_1776_LC_6_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1775_1776_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1775_1776_LC_6_8_1 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1775_1776_LC_6_8_1  (
            .in0(N__61347),
            .in1(N__36849),
            .in2(N__67512),
            .in3(_gnd_net_),
            .lcout(REG_mem_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10598_3_lut_LC_6_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10598_3_lut_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10598_3_lut_LC_6_8_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10598_3_lut_LC_6_8_2  (
            .in0(N__38169),
            .in1(N__87755),
            .in2(_gnd_net_),
            .in3(N__36838),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9998_3_lut_LC_6_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9998_3_lut_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9998_3_lut_LC_6_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9998_3_lut_LC_6_8_3  (
            .in0(N__87756),
            .in1(N__36757),
            .in2(_gnd_net_),
            .in3(N__36766),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11647_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13484_bdd_4_lut_LC_6_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13484_bdd_4_lut_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13484_bdd_4_lut_LC_6_8_4 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13484_bdd_4_lut_LC_6_8_4  (
            .in0(N__85280),
            .in1(N__36817),
            .in2(N__36808),
            .in3(N__36805),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5252_5253_LC_6_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5252_5253_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5252_5253_LC_6_8_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5252_5253_LC_6_8_5  (
            .in0(N__48693),
            .in1(N__94875),
            .in2(N__36783),
            .in3(N__76283),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1583_1584_LC_6_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1583_1584_LC_6_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1583_1584_LC_6_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1583_1584_LC_6_8_6  (
            .in0(N__36765),
            .in1(N__61348),
            .in2(_gnd_net_),
            .in3(N__65640),
            .lcout(REG_mem_16_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1679_1680_LC_6_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1679_1680_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1679_1680_LC_6_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1679_1680_LC_6_8_7  (
            .in0(N__61346),
            .in1(N__36756),
            .in2(_gnd_net_),
            .in3(N__66530),
            .lcout(REG_mem_17_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93251),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11993_LC_6_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11993_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11993_LC_6_9_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11993_LC_6_9_0  (
            .in0(N__37225),
            .in1(N__92135),
            .in2(N__36922),
            .in3(N__87754),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13814 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2651_2652_LC_6_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2651_2652_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2651_2652_LC_6_9_1 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2651_2652_LC_6_9_1  (
            .in0(N__79637),
            .in1(N__63311),
            .in2(N__37920),
            .in3(N__94877),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93245),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1136_1137_LC_6_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1136_1137_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1136_1137_LC_6_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1136_1137_LC_6_9_2  (
            .in0(N__36918),
            .in1(N__41748),
            .in2(_gnd_net_),
            .in3(N__66802),
            .lcout(REG_mem_11_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93245),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i560_561_LC_6_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i560_561_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i560_561_LC_6_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i560_561_LC_6_9_3  (
            .in0(N__41749),
            .in1(N__36906),
            .in2(_gnd_net_),
            .in3(N__67854),
            .lcout(REG_mem_5_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93245),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i656_657_LC_6_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i656_657_LC_6_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i656_657_LC_6_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i656_657_LC_6_9_4  (
            .in0(N__36891),
            .in1(N__41750),
            .in2(_gnd_net_),
            .in3(N__66416),
            .lcout(REG_mem_6_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93245),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11335_LC_6_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11335_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11335_LC_6_9_5 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11335_LC_6_9_5  (
            .in0(N__87753),
            .in1(N__38245),
            .in2(N__92409),
            .in3(N__37021),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13022 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4289_4290_LC_6_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4289_4290_LC_6_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4289_4290_LC_6_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4289_4290_LC_6_9_6  (
            .in0(N__37167),
            .in1(N__56415),
            .in2(_gnd_net_),
            .in3(N__71699),
            .lcout(REG_mem_44_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93245),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1316_1317_LC_6_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1316_1317_LC_6_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1316_1317_LC_6_9_7 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1316_1317_LC_6_9_7  (
            .in0(N__38376),
            .in1(N__48709),
            .in2(N__70137),
            .in3(_gnd_net_),
            .lcout(REG_mem_13_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93245),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4751_4752_LC_6_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4751_4752_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4751_4752_LC_6_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4751_4752_LC_6_10_0  (
            .in0(N__36873),
            .in1(N__61387),
            .in2(_gnd_net_),
            .in3(N__63001),
            .lcout(REG_mem_49_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11540_LC_6_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11540_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11540_LC_6_10_1 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11540_LC_6_10_1  (
            .in0(N__92009),
            .in1(N__88125),
            .in2(N__38458),
            .in3(N__37030),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13244_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13244_bdd_4_lut_LC_6_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13244_bdd_4_lut_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13244_bdd_4_lut_LC_6_10_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13244_bdd_4_lut_LC_6_10_2  (
            .in0(N__36874),
            .in1(N__92008),
            .in2(N__36865),
            .in3(N__38272),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4943_4944_LC_6_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4943_4944_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4943_4944_LC_6_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4943_4944_LC_6_10_3  (
            .in0(N__61384),
            .in1(N__72245),
            .in2(_gnd_net_),
            .in3(N__37029),
            .lcout(REG_mem_51_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4964_4965_LC_6_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4964_4965_LC_6_10_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4964_4965_LC_6_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4964_4965_LC_6_10_4  (
            .in0(N__72246),
            .in1(N__37020),
            .in2(_gnd_net_),
            .in3(N__48648),
            .lcout(REG_mem_51_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5231_5232_LC_6_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5231_5232_LC_6_10_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5231_5232_LC_6_10_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5231_5232_LC_6_10_5  (
            .in0(N__61386),
            .in1(N__94874),
            .in2(N__37009),
            .in3(N__76211),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6086_6087_LC_6_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6086_6087_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6086_6087_LC_6_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6086_6087_LC_6_10_6  (
            .in0(N__36990),
            .in1(N__71331),
            .in2(_gnd_net_),
            .in3(N__67669),
            .lcout(REG_mem_63_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i623_624_LC_6_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i623_624_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i623_624_LC_6_10_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i623_624_LC_6_10_7  (
            .in0(N__61385),
            .in1(N__36972),
            .in2(_gnd_net_),
            .in3(N__66425),
            .lcout(REG_mem_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93238),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3983_3984_LC_6_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3983_3984_LC_6_11_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3983_3984_LC_6_11_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3983_3984_LC_6_11_0  (
            .in0(N__36942),
            .in1(N__61389),
            .in2(_gnd_net_),
            .in3(N__66022),
            .lcout(REG_mem_41_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93246),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11695_LC_6_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11695_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11695_LC_6_11_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11695_LC_6_11_1  (
            .in0(N__92288),
            .in1(N__88096),
            .in2(N__36961),
            .in3(N__36931),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13454_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13454_bdd_4_lut_LC_6_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13454_bdd_4_lut_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13454_bdd_4_lut_LC_6_11_2 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13454_bdd_4_lut_LC_6_11_2  (
            .in0(N__36943),
            .in1(N__38542),
            .in2(N__36934),
            .in3(N__92285),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13457 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4079_4080_LC_6_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4079_4080_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4079_4080_LC_6_11_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4079_4080_LC_6_11_3  (
            .in0(N__61388),
            .in1(N__36930),
            .in2(_gnd_net_),
            .in3(N__68045),
            .lcout(REG_mem_42_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93246),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11157_LC_6_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11157_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11157_LC_6_11_4 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11157_LC_6_11_4  (
            .in0(N__88095),
            .in1(N__92287),
            .in2(N__43753),
            .in3(N__40069),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12800_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12800_bdd_4_lut_LC_6_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12800_bdd_4_lut_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12800_bdd_4_lut_LC_6_11_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12800_bdd_4_lut_LC_6_11_5  (
            .in0(N__92284),
            .in1(N__37171),
            .in2(N__37156),
            .in3(N__37153),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5651_5652_LC_6_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5651_5652_LC_6_11_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5651_5652_LC_6_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5651_5652_LC_6_11_6  (
            .in0(N__37113),
            .in1(N__62425),
            .in2(_gnd_net_),
            .in3(N__79969),
            .lcout(REG_mem_58_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93246),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14306_bdd_4_lut_LC_6_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14306_bdd_4_lut_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14306_bdd_4_lut_LC_6_11_7 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14306_bdd_4_lut_LC_6_11_7  (
            .in0(N__92286),
            .in1(N__45619),
            .in2(N__45445),
            .in3(N__37102),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11625 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11395_LC_6_12_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11395_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11395_LC_6_12_0 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11395_LC_6_12_0  (
            .in0(N__37252),
            .in1(N__91479),
            .in2(N__37042),
            .in3(N__87576),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13088 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4199_4200_LC_6_12_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4199_4200_LC_6_12_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4199_4200_LC_6_12_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4199_4200_LC_6_12_1  (
            .in0(N__37074),
            .in1(N__47155),
            .in2(_gnd_net_),
            .in3(N__68265),
            .lcout(REG_mem_43_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93252),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10341_3_lut_LC_6_12_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10341_3_lut_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10341_3_lut_LC_6_12_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10341_3_lut_LC_6_12_2  (
            .in0(N__85170),
            .in1(_gnd_net_),
            .in2(N__37063),
            .in3(N__38686),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11990 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11859_LC_6_12_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11859_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11859_LC_6_12_3 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11859_LC_6_12_3  (
            .in0(N__87577),
            .in1(N__38497),
            .in2(N__91863),
            .in3(N__38416),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13652 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1007_1008_LC_6_12_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1007_1008_LC_6_12_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1007_1008_LC_6_12_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1007_1008_LC_6_12_4  (
            .in0(N__37038),
            .in1(N__61396),
            .in2(_gnd_net_),
            .in3(N__66971),
            .lcout(REG_mem_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93252),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1103_1104_LC_6_12_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1103_1104_LC_6_12_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1103_1104_LC_6_12_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1103_1104_LC_6_12_5  (
            .in0(N__61395),
            .in1(N__37251),
            .in2(_gnd_net_),
            .in3(N__66817),
            .lcout(REG_mem_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93252),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13754_bdd_4_lut_LC_6_12_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13754_bdd_4_lut_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13754_bdd_4_lut_LC_6_12_6 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13754_bdd_4_lut_LC_6_12_6  (
            .in0(N__40210),
            .in1(N__91478),
            .in2(N__37243),
            .in3(N__45502),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13757 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1040_1041_LC_6_12_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1040_1041_LC_6_12_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1040_1041_LC_6_12_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1040_1041_LC_6_12_7  (
            .in0(N__66972),
            .in1(N__37218),
            .in2(_gnd_net_),
            .in3(N__41669),
            .lcout(REG_mem_10_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93252),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10832_3_lut_LC_6_13_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10832_3_lut_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10832_3_lut_LC_6_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10832_3_lut_LC_6_13_0  (
            .in0(N__87432),
            .in1(N__40159),
            .in2(_gnd_net_),
            .in3(N__40351),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12481 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i266_267_LC_6_13_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i266_267_LC_6_13_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i266_267_LC_6_13_1 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i266_267_LC_6_13_1  (
            .in0(N__46394),
            .in1(N__95345),
            .in2(N__37207),
            .in3(N__80554),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i362_363_LC_6_13_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i362_363_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i362_363_LC_6_13_2 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i362_363_LC_6_13_2  (
            .in0(N__95344),
            .in1(N__37191),
            .in2(N__46472),
            .in3(N__83374),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3338_3339_LC_6_13_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3338_3339_LC_6_13_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3338_3339_LC_6_13_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3338_3339_LC_6_13_3  (
            .in0(N__46395),
            .in1(N__95346),
            .in2(N__37351),
            .in3(N__80555),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12003_LC_6_13_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12003_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12003_LC_6_13_4 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12003_LC_6_13_4  (
            .in0(N__91602),
            .in1(N__37531),
            .in2(N__87712),
            .in3(N__37180),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13826 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4091_4092_LC_6_13_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4091_4092_LC_6_13_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4091_4092_LC_6_13_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4091_4092_LC_6_13_5  (
            .in0(N__37179),
            .in1(N__63230),
            .in2(_gnd_net_),
            .in3(N__68049),
            .lcout(REG_mem_42_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3146_3147_LC_6_13_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3146_3147_LC_6_13_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3146_3147_LC_6_13_6 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3146_3147_LC_6_13_6  (
            .in0(N__95343),
            .in1(N__82910),
            .in2(N__37321),
            .in3(N__46396),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4103_4104_LC_6_13_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4103_4104_LC_6_13_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4103_4104_LC_6_13_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4103_4104_LC_6_13_7  (
            .in0(N__37362),
            .in1(N__47156),
            .in2(_gnd_net_),
            .in3(N__68050),
            .lcout(REG_mem_42_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93261),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10827_3_lut_LC_6_14_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10827_3_lut_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10827_3_lut_LC_6_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10827_3_lut_LC_6_14_0  (
            .in0(N__37350),
            .in1(N__87529),
            .in2(_gnd_net_),
            .in3(N__38955),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10826_3_lut_LC_6_14_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10826_3_lut_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10826_3_lut_LC_6_14_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10826_3_lut_LC_6_14_1  (
            .in0(N__87528),
            .in1(N__37336),
            .in2(_gnd_net_),
            .in3(N__37320),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12475 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10845_3_lut_LC_6_14_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10845_3_lut_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10845_3_lut_LC_6_14_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10845_3_lut_LC_6_14_2  (
            .in0(N__45766),
            .in1(N__87530),
            .in2(_gnd_net_),
            .in3(N__38812),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12494_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12373_LC_6_14_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12373_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12373_LC_6_14_3 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12373_LC_6_14_3  (
            .in0(N__91330),
            .in1(N__37402),
            .in2(N__37306),
            .in3(N__85169),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14252_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14252_bdd_4_lut_LC_6_14_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14252_bdd_4_lut_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14252_bdd_4_lut_LC_6_14_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14252_bdd_4_lut_LC_6_14_4  (
            .in0(N__85167),
            .in1(N__37453),
            .in2(N__37303),
            .in3(N__37471),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11570_LC_6_14_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11570_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11570_LC_6_14_5 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11570_LC_6_14_5  (
            .in0(N__91329),
            .in1(N__85168),
            .in2(N__37300),
            .in3(N__40288),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13292_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13292_bdd_4_lut_LC_6_14_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13292_bdd_4_lut_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13292_bdd_4_lut_LC_6_14_6 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13292_bdd_4_lut_LC_6_14_6  (
            .in0(N__85166),
            .in1(N__37288),
            .in2(N__37282),
            .in3(N__37279),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13295_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9994_3_lut_LC_6_14_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9994_3_lut_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9994_3_lut_LC_6_14_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9994_3_lut_LC_6_14_7  (
            .in0(N__90054),
            .in1(_gnd_net_),
            .in2(N__37273),
            .in3(N__37270),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10838_3_lut_LC_6_15_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10838_3_lut_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10838_3_lut_LC_6_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10838_3_lut_LC_6_15_0  (
            .in0(N__87298),
            .in1(N__42448),
            .in2(_gnd_net_),
            .in3(N__42304),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1037_1038_LC_6_15_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1037_1038_LC_6_15_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1037_1038_LC_6_15_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1037_1038_LC_6_15_1  (
            .in0(N__37575),
            .in1(N__46989),
            .in2(_gnd_net_),
            .in3(N__66974),
            .lcout(REG_mem_10_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4106_4107_LC_6_15_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4106_4107_LC_6_15_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4106_4107_LC_6_15_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4106_4107_LC_6_15_2  (
            .in0(N__46384),
            .in1(N__37464),
            .in2(_gnd_net_),
            .in3(N__68075),
            .lcout(REG_mem_42_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10839_3_lut_LC_6_15_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10839_3_lut_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10839_3_lut_LC_6_15_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10839_3_lut_LC_6_15_3  (
            .in0(N__37447),
            .in1(N__37465),
            .in2(_gnd_net_),
            .in3(N__87299),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12488 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4202_4203_LC_6_15_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4202_4203_LC_6_15_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4202_4203_LC_6_15_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4202_4203_LC_6_15_4  (
            .in0(N__46385),
            .in1(N__37446),
            .in2(_gnd_net_),
            .in3(N__68292),
            .lcout(REG_mem_43_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3050_3051_LC_6_15_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3050_3051_LC_6_15_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3050_3051_LC_6_15_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3050_3051_LC_6_15_5  (
            .in0(N__37431),
            .in1(N__46386),
            .in2(_gnd_net_),
            .in3(N__72551),
            .lcout(REG_mem_31_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10844_3_lut_LC_6_15_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10844_3_lut_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10844_3_lut_LC_6_15_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10844_3_lut_LC_6_15_6  (
            .in0(N__87300),
            .in1(_gnd_net_),
            .in2(N__37420),
            .in3(N__37393),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4394_4395_LC_6_15_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4394_4395_LC_6_15_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4394_4395_LC_6_15_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4394_4395_LC_6_15_7  (
            .in0(N__37392),
            .in1(N__46387),
            .in2(_gnd_net_),
            .in3(N__71904),
            .lcout(REG_mem_45_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93281),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i932_933_LC_6_16_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i932_933_LC_6_16_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i932_933_LC_6_16_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i932_933_LC_6_16_0  (
            .in0(N__48764),
            .in1(N__37374),
            .in2(_gnd_net_),
            .in3(N__67197),
            .lcout(REG_mem_9_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4187_4188_LC_6_16_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4187_4188_LC_6_16_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4187_4188_LC_6_16_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4187_4188_LC_6_16_1  (
            .in0(N__37524),
            .in1(N__63312),
            .in2(_gnd_net_),
            .in3(N__68293),
            .lcout(REG_mem_43_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2474_2475_LC_6_16_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2474_2475_LC_6_16_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2474_2475_LC_6_16_2 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2474_2475_LC_6_16_2  (
            .in0(N__46397),
            .in1(N__37512),
            .in2(N__97060),
            .in3(N__95628),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5447_5448_LC_6_16_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5447_5448_LC_6_16_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5447_5448_LC_6_16_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5447_5448_LC_6_16_3  (
            .in0(N__95627),
            .in1(N__47157),
            .in2(N__47697),
            .in3(N__96003),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5165_5166_LC_6_16_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5165_5166_LC_6_16_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5165_5166_LC_6_16_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5165_5166_LC_6_16_4  (
            .in0(N__46988),
            .in1(N__95629),
            .in2(N__40548),
            .in3(N__77047),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4004_4005_LC_6_16_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4004_4005_LC_6_16_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4004_4005_LC_6_16_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4004_4005_LC_6_16_5  (
            .in0(N__37500),
            .in1(N__48761),
            .in2(_gnd_net_),
            .in3(N__66027),
            .lcout(REG_mem_41_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4100_4101_LC_6_16_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4100_4101_LC_6_16_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4100_4101_LC_6_16_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4100_4101_LC_6_16_6  (
            .in0(N__48762),
            .in1(N__37641),
            .in2(_gnd_net_),
            .in3(N__68076),
            .lcout(REG_mem_42_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4196_4197_LC_6_16_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4196_4197_LC_6_16_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4196_4197_LC_6_16_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4196_4197_LC_6_16_7  (
            .in0(N__37626),
            .in1(N__48763),
            .in2(_gnd_net_),
            .in3(N__68294),
            .lcout(REG_mem_43_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93293),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13394_bdd_4_lut_LC_6_17_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13394_bdd_4_lut_LC_6_17_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13394_bdd_4_lut_LC_6_17_0 .LUT_INIT=16'b1011101010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13394_bdd_4_lut_LC_6_17_0  (
            .in0(N__37615),
            .in1(N__91766),
            .in2(N__40525),
            .in3(N__37501),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13397_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9981_3_lut_LC_6_17_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9981_3_lut_LC_6_17_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9981_3_lut_LC_6_17_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9981_3_lut_LC_6_17_1  (
            .in0(N__85051),
            .in1(_gnd_net_),
            .in2(N__37489),
            .in3(N__37648),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11630 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11435_LC_6_17_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11435_LC_6_17_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11435_LC_6_17_2 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11435_LC_6_17_2  (
            .in0(N__37591),
            .in1(N__91767),
            .in2(N__87467),
            .in3(N__48502),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13142_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13142_bdd_4_lut_LC_6_17_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13142_bdd_4_lut_LC_6_17_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13142_bdd_4_lut_LC_6_17_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13142_bdd_4_lut_LC_6_17_3  (
            .in0(N__91765),
            .in1(N__37609),
            .in2(N__37651),
            .in3(N__37600),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11645_LC_6_17_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11645_LC_6_17_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11645_LC_6_17_4 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11645_LC_6_17_4  (
            .in0(N__37642),
            .in1(N__91768),
            .in2(N__87468),
            .in3(N__37630),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4388_4389_LC_6_17_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4388_4389_LC_6_17_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4388_4389_LC_6_17_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4388_4389_LC_6_17_5  (
            .in0(N__48766),
            .in1(N__37608),
            .in2(_gnd_net_),
            .in3(N__71908),
            .lcout(REG_mem_45_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93306),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4292_4293_LC_6_17_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4292_4293_LC_6_17_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4292_4293_LC_6_17_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4292_4293_LC_6_17_6  (
            .in0(N__37599),
            .in1(N__48765),
            .in2(_gnd_net_),
            .in3(N__71764),
            .lcout(REG_mem_44_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93306),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4484_4485_LC_6_17_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4484_4485_LC_6_17_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4484_4485_LC_6_17_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4484_4485_LC_6_17_7  (
            .in0(N__48767),
            .in1(N__37590),
            .in2(_gnd_net_),
            .in3(N__89115),
            .lcout(REG_mem_46_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93306),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12293_LC_6_18_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12293_LC_6_18_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12293_LC_6_18_1 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12293_LC_6_18_1  (
            .in0(N__91785),
            .in1(N__42427),
            .in2(N__37582),
            .in3(N__87223),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14174 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i4_1_lut_LC_6_19_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i4_1_lut_LC_6_19_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i4_1_lut_LC_6_19_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i4_1_lut_LC_6_19_0  (
            .in0(N__89964),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_pll_clk_unbuf_THRU_LUT4_0_LC_6_19_7.C_ON=1'b0;
    defparam GB_BUFFER_pll_clk_unbuf_THRU_LUT4_0_LC_6_19_7.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_pll_clk_unbuf_THRU_LUT4_0_LC_6_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_pll_clk_unbuf_THRU_LUT4_0_LC_6_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37564),
            .lcout(GB_BUFFER_pll_clk_unbuf_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.usb3_data_in_latched__i10_LC_7_1_2 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i10_LC_7_1_2 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i10_LC_7_1_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i10_LC_7_1_2  (
            .in0(N__37723),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\usb3_if_inst.usb3_data_in_latched_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93350),
            .ce(),
            .sr(N__73746));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10371_3_lut_LC_7_2_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10371_3_lut_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10371_3_lut_LC_7_2_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10371_3_lut_LC_7_2_0  (
            .in0(N__39331),
            .in1(N__43441),
            .in2(_gnd_net_),
            .in3(N__88334),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12020 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3878_3879_LC_7_2_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3878_3879_LC_7_2_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3878_3879_LC_7_2_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3878_3879_LC_7_2_1  (
            .in0(N__65888),
            .in1(N__71358),
            .in2(_gnd_net_),
            .in3(N__39636),
            .lcout(REG_mem_40_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93336),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6131_6132_LC_7_2_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6131_6132_LC_7_2_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6131_6132_LC_7_2_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6131_6132_LC_7_2_2  (
            .in0(N__62198),
            .in1(N__37701),
            .in2(_gnd_net_),
            .in3(N__67717),
            .lcout(REG_mem_63_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93336),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10395_3_lut_LC_7_2_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10395_3_lut_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10395_3_lut_LC_7_2_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10395_3_lut_LC_7_2_3  (
            .in0(N__88335),
            .in1(_gnd_net_),
            .in2(N__37705),
            .in3(N__37680),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12044 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6035_6036_LC_7_2_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6035_6036_LC_7_2_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6035_6036_LC_7_2_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6035_6036_LC_7_2_4  (
            .in0(N__94600),
            .in1(N__62255),
            .in2(N__37681),
            .in3(N__77850),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93336),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i179_180_LC_7_2_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i179_180_LC_7_2_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i179_180_LC_7_2_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i179_180_LC_7_2_5  (
            .in0(N__62254),
            .in1(N__94601),
            .in2(N__44733),
            .in3(N__80297),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93336),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11236_LC_7_2_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11236_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11236_LC_7_2_6 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11236_LC_7_2_6  (
            .in0(N__85633),
            .in1(N__92587),
            .in2(N__41146),
            .in3(N__37861),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12860_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12860_bdd_4_lut_LC_7_2_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12860_bdd_4_lut_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12860_bdd_4_lut_LC_7_2_7 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12860_bdd_4_lut_LC_7_2_7  (
            .in0(N__40108),
            .in1(N__42973),
            .in2(N__37669),
            .in3(N__85632),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12863 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13502_bdd_4_lut_LC_7_3_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13502_bdd_4_lut_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13502_bdd_4_lut_LC_7_3_0 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13502_bdd_4_lut_LC_7_3_0  (
            .in0(N__91230),
            .in1(N__39505),
            .in2(N__39550),
            .in3(N__37665),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10350_3_lut_LC_7_3_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10350_3_lut_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10350_3_lut_LC_7_3_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10350_3_lut_LC_7_3_1  (
            .in0(N__37828),
            .in1(N__88674),
            .in2(_gnd_net_),
            .in3(N__37816),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11999 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11650_LC_7_3_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11650_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11650_LC_7_3_2 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11650_LC_7_3_2  (
            .in0(N__88675),
            .in1(N__43276),
            .in2(N__91661),
            .in3(N__69991),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13400_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13400_bdd_4_lut_LC_7_3_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13400_bdd_4_lut_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13400_bdd_4_lut_LC_7_3_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13400_bdd_4_lut_LC_7_3_3  (
            .in0(N__37987),
            .in1(N__91229),
            .in2(N__37804),
            .in3(N__39835),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13403_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10419_3_lut_LC_7_3_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10419_3_lut_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10419_3_lut_LC_7_3_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10419_3_lut_LC_7_3_4  (
            .in0(N__85809),
            .in1(_gnd_net_),
            .in2(N__37801),
            .in3(N__39385),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12068_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12013_LC_7_3_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12013_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12013_LC_7_3_5 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12013_LC_7_3_5  (
            .in0(N__81482),
            .in1(N__90231),
            .in2(N__37798),
            .in3(N__39433),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12268_LC_7_3_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12268_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12268_LC_7_3_6 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12268_LC_7_3_6  (
            .in0(N__91234),
            .in1(N__85824),
            .in2(N__37795),
            .in3(N__37777),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12932_bdd_4_lut_LC_7_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12932_bdd_4_lut_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12932_bdd_4_lut_LC_7_4_0 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12932_bdd_4_lut_LC_7_4_0  (
            .in0(N__39286),
            .in1(N__92666),
            .in2(N__37735),
            .in3(N__39394),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12935 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9846_3_lut_LC_7_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9846_3_lut_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9846_3_lut_LC_7_4_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9846_3_lut_LC_7_4_1  (
            .in0(N__37753),
            .in1(N__85391),
            .in2(_gnd_net_),
            .in3(N__37741),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11495 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3617_3618_LC_7_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3617_3618_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3617_3618_LC_7_4_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3617_3618_LC_7_4_2  (
            .in0(N__37731),
            .in1(N__56515),
            .in2(_gnd_net_),
            .in3(N__63728),
            .lcout(REG_mem_37_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93308),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13232_bdd_4_lut_LC_7_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13232_bdd_4_lut_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13232_bdd_4_lut_LC_7_4_3 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13232_bdd_4_lut_LC_7_4_3  (
            .in0(N__92667),
            .in1(N__43483),
            .in2(N__39373),
            .in3(N__43159),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13235_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9843_3_lut_LC_7_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9843_3_lut_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9843_3_lut_LC_7_4_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9843_3_lut_LC_7_4_4  (
            .in0(N__85390),
            .in1(_gnd_net_),
            .in2(N__37894),
            .in3(N__45358),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11492 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3809_3810_LC_7_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3809_3810_LC_7_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3809_3810_LC_7_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3809_3810_LC_7_4_5  (
            .in0(N__56514),
            .in1(N__39405),
            .in2(_gnd_net_),
            .in3(N__61881),
            .lcout(REG_mem_39_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93308),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4550_4551_LC_7_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4550_4551_LC_7_4_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4550_4551_LC_7_4_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4550_4551_LC_7_4_6  (
            .in0(N__37890),
            .in1(N__71325),
            .in2(_gnd_net_),
            .in3(N__66269),
            .lcout(REG_mem_47_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93308),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10694_3_lut_LC_7_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10694_3_lut_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10694_3_lut_LC_7_4_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10694_3_lut_LC_7_4_7  (
            .in0(N__37879),
            .in1(N__88045),
            .in2(_gnd_net_),
            .in3(N__45430),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12920_bdd_4_lut_LC_7_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12920_bdd_4_lut_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12920_bdd_4_lut_LC_7_5_0 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12920_bdd_4_lut_LC_7_5_0  (
            .in0(N__43375),
            .in1(N__92647),
            .in2(N__38050),
            .in3(N__39478),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12923_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10410_3_lut_LC_7_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10410_3_lut_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10410_3_lut_LC_7_5_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10410_3_lut_LC_7_5_1  (
            .in0(N__85389),
            .in1(_gnd_net_),
            .in2(N__37852),
            .in3(N__37834),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12059 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11241_LC_7_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11241_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11241_LC_7_5_2 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11241_LC_7_5_2  (
            .in0(N__38098),
            .in1(N__92649),
            .in2(N__88333),
            .in3(N__48919),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12896_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12896_bdd_4_lut_LC_7_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12896_bdd_4_lut_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12896_bdd_4_lut_LC_7_5_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12896_bdd_4_lut_LC_7_5_3  (
            .in0(N__37960),
            .in1(N__92566),
            .in2(N__37837),
            .in3(N__39739),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12899 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12812_bdd_4_lut_LC_7_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12812_bdd_4_lut_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12812_bdd_4_lut_LC_7_5_4 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12812_bdd_4_lut_LC_7_5_4  (
            .in0(N__37948),
            .in1(N__92646),
            .in2(N__39604),
            .in3(N__37966),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12815 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1331_1332_LC_7_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1331_1332_LC_7_5_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1331_1332_LC_7_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1331_1332_LC_7_5_5  (
            .in0(N__37959),
            .in1(N__62315),
            .in2(_gnd_net_),
            .in3(N__70133),
            .lcout(REG_mem_13_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93294),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4262_4263_LC_7_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4262_4263_LC_7_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4262_4263_LC_7_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4262_4263_LC_7_5_6  (
            .in0(N__37947),
            .in1(N__71405),
            .in2(_gnd_net_),
            .in3(N__71737),
            .lcout(REG_mem_44_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93294),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11176_LC_7_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11176_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11176_LC_7_5_7 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11176_LC_7_5_7  (
            .in0(N__92648),
            .in1(N__88046),
            .in2(N__43318),
            .in3(N__51847),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12830 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12078_LC_7_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12078_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12078_LC_7_6_0 .LUT_INIT=16'b1011110010110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12078_LC_7_6_0  (
            .in0(N__38122),
            .in1(N__92388),
            .in2(N__88669),
            .in3(N__41311),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13916_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13916_bdd_4_lut_LC_7_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13916_bdd_4_lut_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13916_bdd_4_lut_LC_7_6_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13916_bdd_4_lut_LC_7_6_1  (
            .in0(N__92386),
            .in1(N__41293),
            .in2(N__37930),
            .in3(N__38001),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12168_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11794_LC_7_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11794_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11794_LC_7_6_2 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11794_LC_7_6_2  (
            .in0(N__90222),
            .in1(N__85388),
            .in2(N__37927),
            .in3(N__37900),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13478 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12083_LC_7_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12083_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12083_LC_7_6_3 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12083_LC_7_6_3  (
            .in0(N__92389),
            .in1(N__88442),
            .in2(N__38113),
            .in3(N__37924),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13922_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13922_bdd_4_lut_LC_7_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13922_bdd_4_lut_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13922_bdd_4_lut_LC_7_6_4 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13922_bdd_4_lut_LC_7_6_4  (
            .in0(N__38086),
            .in1(N__43357),
            .in2(N__37903),
            .in3(N__92387),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3035_3036_LC_7_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3035_3036_LC_7_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3035_3036_LC_7_6_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3035_3036_LC_7_6_5  (
            .in0(N__63436),
            .in1(N__38121),
            .in2(_gnd_net_),
            .in3(N__72540),
            .lcout(REG_mem_31_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93282),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2555_2556_LC_7_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2555_2556_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2555_2556_LC_7_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2555_2556_LC_7_6_6  (
            .in0(N__38109),
            .in1(N__63437),
            .in2(_gnd_net_),
            .in3(N__70379),
            .lcout(REG_mem_26_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93282),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1427_1428_LC_7_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1427_1428_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1427_1428_LC_7_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1427_1428_LC_7_6_7  (
            .in0(N__38097),
            .in1(N__62316),
            .in2(_gnd_net_),
            .in3(N__74761),
            .lcout(REG_mem_14_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93282),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2363_2364_LC_7_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2363_2364_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2363_2364_LC_7_7_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2363_2364_LC_7_7_0  (
            .in0(N__63485),
            .in1(N__95049),
            .in2(N__38085),
            .in3(N__95892),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3920_3921_LC_7_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3920_3921_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3920_3921_LC_7_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3920_3921_LC_7_7_1  (
            .in0(N__38061),
            .in1(N__41791),
            .in2(_gnd_net_),
            .in3(N__65804),
            .lcout(REG_mem_40_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i851_852_LC_7_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i851_852_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i851_852_LC_7_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i851_852_LC_7_7_2  (
            .in0(N__38046),
            .in1(N__62384),
            .in2(_gnd_net_),
            .in3(N__67236),
            .lcout(REG_mem_8_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3728_3729_LC_7_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3728_3729_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3728_3729_LC_7_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3728_3729_LC_7_7_3  (
            .in0(N__41916),
            .in1(N__41790),
            .in2(_gnd_net_),
            .in3(N__59279),
            .lcout(REG_mem_38_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5453_5454_LC_7_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5453_5454_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5453_5454_LC_7_7_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5453_5454_LC_7_7_4  (
            .in0(N__46731),
            .in1(N__95051),
            .in2(N__38019),
            .in3(N__95893),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2843_2844_LC_7_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2843_2844_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2843_2844_LC_7_7_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2843_2844_LC_7_7_5  (
            .in0(N__95048),
            .in1(N__63486),
            .in2(N__38002),
            .in3(N__70938),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2438_2439_LC_7_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2438_2439_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2438_2439_LC_7_7_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2438_2439_LC_7_7_6  (
            .in0(N__71404),
            .in1(N__95050),
            .in2(N__37983),
            .in3(N__96988),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4400_4401_LC_7_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4400_4401_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4400_4401_LC_7_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4400_4401_LC_7_7_7  (
            .in0(N__38256),
            .in1(N__41792),
            .in2(_gnd_net_),
            .in3(N__71888),
            .lcout(REG_mem_45_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93271),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4868_4869_LC_7_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4868_4869_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4868_4869_LC_7_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4868_4869_LC_7_8_0  (
            .in0(N__38244),
            .in1(N__48731),
            .in2(_gnd_net_),
            .in3(N__73018),
            .lcout(REG_mem_50_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93262),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5057_5058_LC_7_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5057_5058_LC_7_8_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5057_5058_LC_7_8_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5057_5058_LC_7_8_1  (
            .in0(N__77387),
            .in1(N__38223),
            .in2(N__95456),
            .in3(N__56624),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93262),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5039_5040_LC_7_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5039_5040_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5039_5040_LC_7_8_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5039_5040_LC_7_8_2  (
            .in0(N__61372),
            .in1(N__95080),
            .in2(N__38211),
            .in3(N__77389),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93262),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2378_2379_LC_7_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2378_2379_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2378_2379_LC_7_8_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2378_2379_LC_7_8_3  (
            .in0(N__95078),
            .in1(N__46347),
            .in2(N__38187),
            .in3(N__95891),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93262),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1616_1617_LC_7_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1616_1617_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1616_1617_LC_7_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1616_1617_LC_7_8_4  (
            .in0(N__38170),
            .in1(N__41793),
            .in2(_gnd_net_),
            .in3(N__65605),
            .lcout(REG_mem_16_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93262),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5066_5067_LC_7_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5066_5067_LC_7_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5066_5067_LC_7_8_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5066_5067_LC_7_8_5  (
            .in0(N__77388),
            .in1(N__38151),
            .in2(N__95457),
            .in3(N__46348),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93262),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10868_3_lut_LC_7_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10868_3_lut_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10868_3_lut_LC_7_8_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10868_3_lut_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(N__87752),
            .in2(N__38155),
            .in3(N__39771),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5537_5538_LC_7_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5537_5538_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5537_5538_LC_7_8_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5537_5538_LC_7_8_7  (
            .in0(N__95079),
            .in1(N__38133),
            .in2(N__56626),
            .in3(N__96934),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93262),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6011_6012_LC_7_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6011_6012_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6011_6012_LC_7_9_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6011_6012_LC_7_9_0  (
            .in0(N__38406),
            .in1(N__95053),
            .in2(N__63538),
            .in3(N__77951),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93253),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12283_LC_7_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12283_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12283_LC_7_9_1 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12283_LC_7_9_1  (
            .in0(N__38341),
            .in1(N__92521),
            .in2(N__88408),
            .in3(N__38395),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14162_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14162_bdd_4_lut_LC_7_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14162_bdd_4_lut_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14162_bdd_4_lut_LC_7_9_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14162_bdd_4_lut_LC_7_9_2  (
            .in0(N__92520),
            .in1(N__38377),
            .in2(N__38365),
            .in3(N__38350),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1220_1221_LC_7_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1220_1221_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1220_1221_LC_7_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1220_1221_LC_7_9_3  (
            .in0(N__38349),
            .in1(N__48732),
            .in2(_gnd_net_),
            .in3(N__59565),
            .lcout(REG_mem_12_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93253),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1412_1413_LC_7_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1412_1413_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1412_1413_LC_7_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1412_1413_LC_7_9_4  (
            .in0(N__48733),
            .in1(N__38340),
            .in2(_gnd_net_),
            .in3(N__74749),
            .lcout(REG_mem_14_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93253),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2381_2382_LC_7_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2381_2382_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2381_2382_LC_7_9_5 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2381_2382_LC_7_9_5  (
            .in0(N__95052),
            .in1(N__38325),
            .in2(N__95990),
            .in3(N__46732),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93253),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i452_453_LC_7_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i452_453_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i452_453_LC_7_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i452_453_LC_7_9_6  (
            .in0(N__48734),
            .in1(N__38304),
            .in2(_gnd_net_),
            .in3(N__72668),
            .lcout(REG_mem_4_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93253),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i464_465_LC_7_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i464_465_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i464_465_LC_7_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i464_465_LC_7_9_7  (
            .in0(N__72667),
            .in1(N__38289),
            .in2(_gnd_net_),
            .in3(N__41785),
            .lcout(REG_mem_4_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93253),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4655_4656_LC_7_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4655_4656_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4655_4656_LC_7_10_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4655_4656_LC_7_10_0  (
            .in0(N__75513),
            .in1(_gnd_net_),
            .in2(N__61341),
            .in3(N__38271),
            .lcout(REG_mem_48_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3887_3888_LC_7_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3887_3888_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3887_3888_LC_7_10_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3887_3888_LC_7_10_1  (
            .in0(N__38541),
            .in1(N__61281),
            .in2(_gnd_net_),
            .in3(N__65860),
            .lcout(REG_mem_40_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4976_4977_LC_7_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4976_4977_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4976_4977_LC_7_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4976_4977_LC_7_10_2  (
            .in0(N__38523),
            .in1(N__41786),
            .in2(_gnd_net_),
            .in3(N__72244),
            .lcout(REG_mem_51_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1700_1701_LC_7_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1700_1701_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1700_1701_LC_7_10_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1700_1701_LC_7_10_3  (
            .in0(N__38508),
            .in1(N__48842),
            .in2(_gnd_net_),
            .in3(N__66579),
            .lcout(REG_mem_17_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6107_6108_LC_7_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6107_6108_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6107_6108_LC_7_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6107_6108_LC_7_10_4  (
            .in0(N__38493),
            .in1(N__63537),
            .in2(_gnd_net_),
            .in3(N__67668),
            .lcout(REG_mem_63_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i527_528_LC_7_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i527_528_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i527_528_LC_7_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i527_528_LC_7_10_5  (
            .in0(N__38469),
            .in1(N__61282),
            .in2(_gnd_net_),
            .in3(N__67875),
            .lcout(REG_mem_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4847_4848_LC_7_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4847_4848_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4847_4848_LC_7_10_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4847_4848_LC_7_10_6  (
            .in0(N__61280),
            .in1(N__38451),
            .in2(_gnd_net_),
            .in3(N__73017),
            .lcout(REG_mem_50_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1994_1995_LC_7_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1994_1995_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1994_1995_LC_7_10_7 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1994_1995_LC_7_10_7  (
            .in0(N__77391),
            .in1(N__95054),
            .in2(N__38433),
            .in3(N__46451),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93244),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13700_bdd_4_lut_LC_7_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13700_bdd_4_lut_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13700_bdd_4_lut_LC_7_11_0 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13700_bdd_4_lut_LC_7_11_0  (
            .in0(N__39943),
            .in1(N__92282),
            .in2(N__38653),
            .in3(N__45091),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3899_3900_LC_7_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3899_3900_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3899_3900_LC_7_11_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3899_3900_LC_7_11_1  (
            .in0(N__39000),
            .in1(N__63532),
            .in2(_gnd_net_),
            .in3(N__65880),
            .lcout(REG_mem_40_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93254),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11904_LC_7_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11904_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11904_LC_7_11_2 .LUT_INIT=16'b1011110010110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11904_LC_7_11_2  (
            .in0(N__38671),
            .in1(N__92283),
            .in2(N__88069),
            .in3(N__38605),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13652_bdd_4_lut_LC_7_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13652_bdd_4_lut_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13652_bdd_4_lut_LC_7_11_3 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13652_bdd_4_lut_LC_7_11_3  (
            .in0(N__92281),
            .in1(N__38644),
            .in2(N__38596),
            .in3(N__39957),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12237_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11620_LC_7_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11620_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11620_LC_7_11_4 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11620_LC_7_11_4  (
            .in0(N__90022),
            .in1(N__85352),
            .in2(N__38638),
            .in3(N__38635),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5903_5904_LC_7_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5903_5904_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5903_5904_LC_7_11_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5903_5904_LC_7_11_5  (
            .in0(N__61268),
            .in1(N__94456),
            .in2(N__38622),
            .in3(N__70812),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93254),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5627_5628_LC_7_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5627_5628_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5627_5628_LC_7_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5627_5628_LC_7_11_6  (
            .in0(N__63531),
            .in1(N__38604),
            .in2(_gnd_net_),
            .in3(N__79936),
            .lcout(REG_mem_58_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93254),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5915_5916_LC_7_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5915_5916_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5915_5916_LC_7_11_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5915_5916_LC_7_11_7  (
            .in0(N__63533),
            .in1(N__94457),
            .in2(N__38595),
            .in3(N__70813),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93254),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i827_828_LC_7_12_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i827_828_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i827_828_LC_7_12_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i827_828_LC_7_12_0  (
            .in0(N__38571),
            .in1(N__63493),
            .in2(_gnd_net_),
            .in3(N__67301),
            .lcout(REG_mem_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i911_912_LC_7_12_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i911_912_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i911_912_LC_7_12_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i911_912_LC_7_12_1  (
            .in0(N__61304),
            .in1(N__38736),
            .in2(_gnd_net_),
            .in3(N__67194),
            .lcout(REG_mem_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i431_432_LC_7_12_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i431_432_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i431_432_LC_7_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i431_432_LC_7_12_2  (
            .in0(N__38553),
            .in1(N__61305),
            .in2(_gnd_net_),
            .in3(N__72716),
            .lcout(REG_mem_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2957_2958_LC_7_12_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2957_2958_LC_7_12_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2957_2958_LC_7_12_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2957_2958_LC_7_12_3  (
            .in0(N__95452),
            .in1(N__39021),
            .in2(N__47031),
            .in3(N__77950),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1499_1500_LC_7_12_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1499_1500_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1499_1500_LC_7_12_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1499_1500_LC_7_12_4  (
            .in0(N__38748),
            .in1(N__63491),
            .in2(_gnd_net_),
            .in3(N__64011),
            .lcout(REG_mem_15_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13088_bdd_4_lut_LC_7_12_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13088_bdd_4_lut_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13088_bdd_4_lut_LC_7_12_5 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13088_bdd_4_lut_LC_7_12_5  (
            .in0(N__91477),
            .in1(N__38737),
            .in2(N__38728),
            .in3(N__40054),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3995_3996_LC_7_12_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3995_3996_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3995_3996_LC_7_12_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3995_3996_LC_7_12_6  (
            .in0(N__38973),
            .in1(N__63492),
            .in2(_gnd_net_),
            .in3(N__66021),
            .lcout(REG_mem_41_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2861_2862_LC_7_12_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2861_2862_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2861_2862_LC_7_12_7 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2861_2862_LC_7_12_7  (
            .in0(N__46990),
            .in1(N__39084),
            .in2(N__95650),
            .in3(N__70882),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93263),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1115_1116_LC_7_13_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1115_1116_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1115_1116_LC_7_13_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1115_1116_LC_7_13_0  (
            .in0(N__38700),
            .in1(_gnd_net_),
            .in2(N__63536),
            .in3(N__66818),
            .lcout(REG_mem_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11595_LC_7_13_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11595_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11595_LC_7_13_1 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11595_LC_7_13_1  (
            .in0(N__38920),
            .in1(N__91601),
            .in2(N__87751),
            .in3(N__42481),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13334_bdd_4_lut_LC_7_13_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13334_bdd_4_lut_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13334_bdd_4_lut_LC_7_13_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13334_bdd_4_lut_LC_7_13_2  (
            .in0(N__91600),
            .in1(N__38680),
            .in2(N__38689),
            .in3(N__40171),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4367_4368_LC_7_13_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4367_4368_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4367_4368_LC_7_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4367_4368_LC_7_13_3  (
            .in0(N__38679),
            .in1(N__61056),
            .in2(_gnd_net_),
            .in3(N__71892),
            .lcout(REG_mem_45_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4463_4464_LC_7_13_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4463_4464_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4463_4464_LC_7_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4463_4464_LC_7_13_4  (
            .in0(N__61055),
            .in1(N__38919),
            .in2(_gnd_net_),
            .in3(N__89072),
            .lcout(REG_mem_46_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2276_2277_LC_7_13_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2276_2277_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2276_2277_LC_7_13_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2276_2277_LC_7_13_5  (
            .in0(N__38901),
            .in1(N__48759),
            .in2(_gnd_net_),
            .in3(N__75039),
            .lcout(REG_mem_23_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1019_1020_LC_7_13_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1019_1020_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1019_1020_LC_7_13_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1019_1020_LC_7_13_6  (
            .in0(N__38883),
            .in1(_gnd_net_),
            .in2(N__63535),
            .in3(N__66959),
            .lcout(REG_mem_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93272),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14354_bdd_4_lut_LC_7_13_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14354_bdd_4_lut_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14354_bdd_4_lut_LC_7_13_7 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14354_bdd_4_lut_LC_7_13_7  (
            .in0(N__90055),
            .in1(N__38872),
            .in2(N__38860),
            .in3(N__40420),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12486 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2282_2283_LC_7_14_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2282_2283_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2282_2283_LC_7_14_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2282_2283_LC_7_14_0  (
            .in0(N__75040),
            .in1(N__38844),
            .in2(_gnd_net_),
            .in3(N__46497),
            .lcout(REG_mem_23_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3311_3312_LC_7_14_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3311_3312_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3311_3312_LC_7_14_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3311_3312_LC_7_14_1  (
            .in0(N__61342),
            .in1(N__95449),
            .in2(N__38829),
            .in3(N__80556),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4586_4587_LC_7_14_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4586_4587_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4586_4587_LC_7_14_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4586_4587_LC_7_14_2  (
            .in0(N__38811),
            .in1(N__46492),
            .in2(_gnd_net_),
            .in3(N__66267),
            .lcout(REG_mem_47_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6122_6123_LC_7_14_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6122_6123_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6122_6123_LC_7_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6122_6123_LC_7_14_3  (
            .in0(N__46491),
            .in1(N__38793),
            .in2(_gnd_net_),
            .in3(N__67707),
            .lcout(REG_mem_63_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2375_2376_LC_7_14_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2375_2376_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2375_2376_LC_7_14_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2375_2376_LC_7_14_4  (
            .in0(N__95447),
            .in1(N__47213),
            .in2(N__44787),
            .in3(N__95989),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6026_6027_LC_7_14_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6026_6027_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6026_6027_LC_7_14_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6026_6027_LC_7_14_5  (
            .in0(N__77889),
            .in1(N__38778),
            .in2(N__46548),
            .in3(N__95450),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2954_2955_LC_7_14_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2954_2955_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2954_2955_LC_7_14_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2954_2955_LC_7_14_6  (
            .in0(N__95448),
            .in1(N__46493),
            .in2(N__39045),
            .in3(N__77890),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93283),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12113_LC_7_14_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12113_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12113_LC_7_14_7 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12113_LC_7_14_7  (
            .in0(N__87734),
            .in1(N__91328),
            .in2(N__39028),
            .in3(N__45709),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13958 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11998_LC_7_15_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11998_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11998_LC_7_15_0 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11998_LC_7_15_0  (
            .in0(N__90712),
            .in1(N__87297),
            .in2(N__39154),
            .in3(N__43795),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13820_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13820_bdd_4_lut_LC_7_15_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13820_bdd_4_lut_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13820_bdd_4_lut_LC_7_15_1 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13820_bdd_4_lut_LC_7_15_1  (
            .in0(N__38941),
            .in1(N__90710),
            .in2(N__39010),
            .in3(N__38929),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11710_LC_7_15_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11710_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11710_LC_7_15_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11710_LC_7_15_2  (
            .in0(N__38962),
            .in1(N__90053),
            .in2(N__39007),
            .in3(N__85102),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13466 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13826_bdd_4_lut_LC_7_15_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13826_bdd_4_lut_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13826_bdd_4_lut_LC_7_15_3 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13826_bdd_4_lut_LC_7_15_3  (
            .in0(N__39004),
            .in1(N__90711),
            .in2(N__38989),
            .in3(N__38977),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12195 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3434_3435_LC_7_15_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3434_3435_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3434_3435_LC_7_15_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3434_3435_LC_7_15_4  (
            .in0(N__95451),
            .in1(N__46487),
            .in2(N__38956),
            .in3(N__83375),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93295),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4379_4380_LC_7_15_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4379_4380_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4379_4380_LC_7_15_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4379_4380_LC_7_15_5  (
            .in0(N__63472),
            .in1(N__38940),
            .in2(_gnd_net_),
            .in3(N__71903),
            .lcout(REG_mem_45_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93295),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4283_4284_LC_7_15_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4283_4284_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4283_4284_LC_7_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4283_4284_LC_7_15_6  (
            .in0(N__38928),
            .in1(N__63473),
            .in2(_gnd_net_),
            .in3(N__71742),
            .lcout(REG_mem_44_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93295),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4475_4476_LC_7_15_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4475_4476_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4475_4476_LC_7_15_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4475_4476_LC_7_15_7  (
            .in0(N__89074),
            .in1(_gnd_net_),
            .in2(N__63530),
            .in3(N__39150),
            .lcout(REG_mem_46_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93295),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10857_3_lut_LC_7_16_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10857_3_lut_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10857_3_lut_LC_7_16_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10857_3_lut_LC_7_16_0  (
            .in0(N__46609),
            .in1(N__42394),
            .in2(_gnd_net_),
            .in3(N__87178),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11600_LC_7_16_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11600_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11600_LC_7_16_1 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11600_LC_7_16_1  (
            .in0(N__91368),
            .in1(N__39142),
            .in2(N__85165),
            .in3(N__39127),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13310_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13310_bdd_4_lut_LC_7_16_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13310_bdd_4_lut_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13310_bdd_4_lut_LC_7_16_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13310_bdd_4_lut_LC_7_16_2  (
            .in0(N__39115),
            .in1(N__85052),
            .in2(N__39109),
            .in3(N__39073),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2285_2286_LC_7_16_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2285_2286_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2285_2286_LC_7_16_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2285_2286_LC_7_16_3  (
            .in0(N__40701),
            .in1(N__46962),
            .in2(_gnd_net_),
            .in3(N__75041),
            .lcout(REG_mem_23_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93309),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13958_bdd_4_lut_LC_7_16_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13958_bdd_4_lut_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13958_bdd_4_lut_LC_7_16_4 .LUT_INIT=16'b1011101010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13958_bdd_4_lut_LC_7_16_4  (
            .in0(N__39097),
            .in1(N__91367),
            .in2(N__39901),
            .in3(N__39088),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10856_3_lut_LC_7_16_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10856_3_lut_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10856_3_lut_LC_7_16_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10856_3_lut_LC_7_16_5  (
            .in0(N__87177),
            .in1(N__39058),
            .in2(_gnd_net_),
            .in3(N__39067),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4682_4683_LC_7_16_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4682_4683_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4682_4683_LC_7_16_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4682_4683_LC_7_16_6  (
            .in0(N__39066),
            .in1(N__46509),
            .in2(_gnd_net_),
            .in3(N__75578),
            .lcout(REG_mem_48_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93309),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4778_4779_LC_7_16_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4778_4779_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4778_4779_LC_7_16_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4778_4779_LC_7_16_7  (
            .in0(N__46508),
            .in1(N__39057),
            .in2(_gnd_net_),
            .in3(N__63007),
            .lcout(REG_mem_49_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93309),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12902_bdd_4_lut_LC_7_17_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12902_bdd_4_lut_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12902_bdd_4_lut_LC_7_17_0 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12902_bdd_4_lut_LC_7_17_0  (
            .in0(N__44629),
            .in1(N__89943),
            .in2(N__39193),
            .in3(N__40531),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13034_bdd_4_lut_LC_7_17_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13034_bdd_4_lut_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13034_bdd_4_lut_LC_7_17_1 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13034_bdd_4_lut_LC_7_17_1  (
            .in0(N__89945),
            .in1(N__39220),
            .in2(N__42142),
            .in3(N__40462),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12387 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12968_bdd_4_lut_LC_7_17_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12968_bdd_4_lut_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12968_bdd_4_lut_LC_7_17_2 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12968_bdd_4_lut_LC_7_17_2  (
            .in0(N__40393),
            .in1(N__89944),
            .in2(N__45961),
            .in3(N__42868),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12405_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_11360_LC_7_17_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_11360_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_11360_LC_7_17_3 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_11360_LC_7_17_3  (
            .in0(N__39178),
            .in1(N__80953),
            .in2(N__39172),
            .in3(N__81245),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12794 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13076_bdd_4_lut_LC_7_17_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13076_bdd_4_lut_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13076_bdd_4_lut_LC_7_17_4 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13076_bdd_4_lut_LC_7_17_4  (
            .in0(N__40654),
            .in1(N__89946),
            .in2(N__44476),
            .in3(N__42673),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12375_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i14_LC_7_17_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i14_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i14_LC_7_17_5 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i14_LC_7_17_5  (
            .in0(N__39169),
            .in1(N__80952),
            .in2(N__39163),
            .in3(N__39160),
            .lcout(REG_out_raw_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97344),
            .ce(N__80872),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3_4_lut_LC_7_18_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3_4_lut_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3_4_lut_LC_7_18_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3_4_lut_LC_7_18_0  (
            .in0(N__50448),
            .in1(N__39303),
            .in2(N__50580),
            .in3(N__39204),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9760_4_lut_LC_7_18_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9760_4_lut_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9760_4_lut_LC_7_18_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9760_4_lut_LC_7_18_1  (
            .in0(N__80949),
            .in1(N__50449),
            .in2(N__50581),
            .in3(N__89880),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_i4_3_lut_LC_7_18_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_i4_3_lut_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_i4_3_lut_LC_7_18_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_i4_3_lut_LC_7_18_2  (
            .in0(N__89882),
            .in1(N__52574),
            .in2(_gnd_net_),
            .in3(N__39205),
            .lcout(rd_addr_nxt_c_6_N_465_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_i6_3_lut_LC_7_18_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_i6_3_lut_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_i6_3_lut_LC_7_18_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_i6_3_lut_LC_7_18_3  (
            .in0(N__80950),
            .in1(_gnd_net_),
            .in2(N__52579),
            .in3(N__39304),
            .lcout(rd_addr_nxt_c_6_N_465_5),
            .ltout(rd_addr_nxt_c_6_N_465_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i5_LC_7_18_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i5_LC_7_18_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i5_LC_7_18_4 .LUT_INIT=16'b0011000000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i5_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(N__73372),
            .in2(N__39247),
            .in3(_gnd_net_),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97345),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i3_1_lut_LC_7_18_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i3_1_lut_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i3_1_lut_LC_7_18_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i3_1_lut_LC_7_18_5  (
            .in0(N__85050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n6_adj_1150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i6_1_lut_LC_7_18_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i6_1_lut_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i6_1_lut_LC_7_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i6_1_lut_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80951),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11375_LC_7_18_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11375_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11375_LC_7_18_7 .LUT_INIT=16'b1011110010110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11375_LC_7_18_7  (
            .in0(N__39244),
            .in1(N__89881),
            .in2(N__85164),
            .in3(N__39235),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13034 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_2_lut_LC_7_19_0 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_2_lut_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_2_lut_LC_7_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_2_lut_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__87015),
            .in2(_gnd_net_),
            .in3(N__39214),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_0 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10637 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_3_lut_LC_7_19_1 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_3_lut_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_3_lut_LC_7_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_3_lut_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__91989),
            .in3(N__39211),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_1 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10637 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10638 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_4_lut_LC_7_19_2 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_4_lut_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_4_lut_LC_7_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_4_lut_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__84967),
            .in2(_gnd_net_),
            .in3(N__39208),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_2 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10638 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10639 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_5_lut_LC_7_19_3 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_5_lut_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_5_lut_LC_7_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_5_lut_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__89850),
            .in2(_gnd_net_),
            .in3(N__39196),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_3 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10639 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10640 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_6_lut_LC_7_19_4 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_6_lut_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_6_lut_LC_7_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_6_lut_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__81195),
            .in2(_gnd_net_),
            .in3(N__39307),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_4 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10640 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10641 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_7_lut_LC_7_19_5 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_7_lut_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_7_lut_LC_7_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_7_lut_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__80954),
            .in2(_gnd_net_),
            .in3(N__39292),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_5 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10641 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10642 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_8_lut_LC_7_19_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_8_lut_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_8_lut_LC_7_19_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_151_8_lut_LC_7_19_6  (
            .in0(N__44392),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39289),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_p1_w_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i467_468_LC_8_1_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i467_468_LC_8_1_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i467_468_LC_8_1_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i467_468_LC_8_1_0  (
            .in0(N__44673),
            .in1(N__62351),
            .in2(_gnd_net_),
            .in3(N__72701),
            .lcout(REG_mem_4_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93367),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10073_3_lut_LC_8_1_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10073_3_lut_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10073_3_lut_LC_8_1_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10073_3_lut_LC_8_1_1  (
            .in0(N__88004),
            .in1(N__39270),
            .in2(_gnd_net_),
            .in3(N__52132),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3521_3522_LC_8_1_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3521_3522_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3521_3522_LC_8_1_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3521_3522_LC_8_1_2  (
            .in0(N__56488),
            .in1(N__39282),
            .in2(_gnd_net_),
            .in3(N__54065),
            .lcout(REG_mem_36_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93367),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i353_354_LC_8_1_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i353_354_LC_8_1_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i353_354_LC_8_1_3 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i353_354_LC_8_1_3  (
            .in0(N__42984),
            .in1(N__56489),
            .in2(N__83384),
            .in3(N__94181),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93367),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5129_5130_LC_8_1_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5129_5130_LC_8_1_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5129_5130_LC_8_1_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5129_5130_LC_8_1_4  (
            .in0(N__94179),
            .in1(N__96815),
            .in2(N__39271),
            .in3(N__77037),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93367),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5225_5226_LC_8_1_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5225_5226_LC_8_1_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5225_5226_LC_8_1_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5225_5226_LC_8_1_5  (
            .in0(N__96816),
            .in1(N__94180),
            .in2(N__39259),
            .in3(N__76335),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93367),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10074_3_lut_LC_8_1_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10074_3_lut_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10074_3_lut_LC_8_1_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10074_3_lut_LC_8_1_6  (
            .in0(N__41236),
            .in1(N__39258),
            .in2(_gnd_net_),
            .in3(N__88005),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11723_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11715_LC_8_1_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11715_LC_8_1_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11715_LC_8_1_7 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11715_LC_8_1_7  (
            .in0(N__39358),
            .in1(N__85825),
            .in2(N__39352),
            .in3(N__92677),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10322_3_lut_LC_8_2_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10322_3_lut_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10322_3_lut_LC_8_2_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10322_3_lut_LC_8_2_0  (
            .in0(N__39349),
            .in1(_gnd_net_),
            .in2(N__40975),
            .in3(N__88002),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11971 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3923_3924_LC_8_2_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3923_3924_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3923_3924_LC_8_2_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3923_3924_LC_8_2_1  (
            .in0(N__40896),
            .in1(N__62253),
            .in2(_gnd_net_),
            .in3(N__65887),
            .lcout(REG_mem_40_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93352),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4883_4884_LC_8_2_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4883_4884_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4883_4884_LC_8_2_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4883_4884_LC_8_2_2  (
            .in0(N__62252),
            .in1(N__39330),
            .in2(_gnd_net_),
            .in3(N__73052),
            .lcout(REG_mem_50_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93352),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2150_2151_LC_8_2_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2150_2151_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2150_2151_LC_8_2_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2150_2151_LC_8_2_3  (
            .in0(N__94176),
            .in1(N__71357),
            .in2(N__39522),
            .in3(N__76312),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93352),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i137_138_LC_8_2_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i137_138_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i137_138_LC_8_2_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i137_138_LC_8_2_4  (
            .in0(N__96777),
            .in1(N__94178),
            .in2(N__40819),
            .in3(N__80293),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93352),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2177_2178_LC_8_2_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2177_2178_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2177_2178_LC_8_2_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2177_2178_LC_8_2_5  (
            .in0(N__94177),
            .in1(N__56409),
            .in2(N__41262),
            .in3(N__76313),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93352),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4307_4308_LC_8_2_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4307_4308_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4307_4308_LC_8_2_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4307_4308_LC_8_2_6  (
            .in0(N__62251),
            .in1(N__39318),
            .in2(_gnd_net_),
            .in3(N__71738),
            .lcout(REG_mem_44_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93352),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10364_3_lut_LC_8_2_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10364_3_lut_LC_8_2_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10364_3_lut_LC_8_2_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10364_3_lut_LC_8_2_7  (
            .in0(N__88003),
            .in1(N__39319),
            .in2(_gnd_net_),
            .in3(N__45163),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12013 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10358_3_lut_LC_8_3_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10358_3_lut_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10358_3_lut_LC_8_3_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10358_3_lut_LC_8_3_0  (
            .in0(N__87664),
            .in1(N__39811),
            .in2(_gnd_net_),
            .in3(N__41275),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12007 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11500_LC_8_3_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11500_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11500_LC_8_3_1 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11500_LC_8_3_1  (
            .in0(N__39460),
            .in1(N__81441),
            .in2(N__43210),
            .in3(N__90230),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13172_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13172_bdd_4_lut_LC_8_3_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13172_bdd_4_lut_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13172_bdd_4_lut_LC_8_3_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13172_bdd_4_lut_LC_8_3_2  (
            .in0(N__81440),
            .in1(N__39454),
            .in2(N__39448),
            .in3(N__39445),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10418_3_lut_LC_8_3_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10418_3_lut_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10418_3_lut_LC_8_3_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10418_3_lut_LC_8_3_3  (
            .in0(N__85808),
            .in1(N__39439),
            .in2(_gnd_net_),
            .in3(N__39529),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12067 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10334_3_lut_LC_8_3_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10334_3_lut_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10334_3_lut_LC_8_3_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10334_3_lut_LC_8_3_4  (
            .in0(N__87663),
            .in1(N__48079),
            .in2(_gnd_net_),
            .in3(N__39427),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11983 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11261_LC_8_3_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11261_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11261_LC_8_3_5 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11261_LC_8_3_5  (
            .in0(N__45310),
            .in1(N__92385),
            .in2(N__88812),
            .in3(N__39406),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12932 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13148_bdd_4_lut_LC_8_3_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13148_bdd_4_lut_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13148_bdd_4_lut_LC_8_3_6 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13148_bdd_4_lut_LC_8_3_6  (
            .in0(N__92384),
            .in1(N__39379),
            .in2(N__40024),
            .in3(N__42073),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11460_LC_8_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11460_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11460_LC_8_4_0 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11460_LC_8_4_0  (
            .in0(N__92651),
            .in1(N__87676),
            .in2(N__39718),
            .in3(N__43336),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i833_834_LC_8_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i833_834_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i833_834_LC_8_4_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i833_834_LC_8_4_1  (
            .in0(N__39369),
            .in1(N__56476),
            .in2(_gnd_net_),
            .in3(N__67311),
            .lcout(REG_mem_8_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93323),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11804_LC_8_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11804_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11804_LC_8_4_2 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11804_LC_8_4_2  (
            .in0(N__92653),
            .in1(N__87678),
            .in2(N__43150),
            .in3(N__43192),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13586_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13586_bdd_4_lut_LC_8_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13586_bdd_4_lut_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13586_bdd_4_lut_LC_8_4_3 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13586_bdd_4_lut_LC_8_4_3  (
            .in0(N__41887),
            .in1(N__92650),
            .in2(N__39532),
            .in3(N__39487),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11734_LC_8_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11734_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11734_LC_8_4_4 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11734_LC_8_4_4  (
            .in0(N__92652),
            .in1(N__87677),
            .in2(N__39499),
            .in3(N__39523),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13502 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2246_2247_LC_8_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2246_2247_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2246_2247_LC_8_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2246_2247_LC_8_4_5  (
            .in0(N__71523),
            .in1(N__39495),
            .in2(_gnd_net_),
            .in3(N__75051),
            .lcout(REG_mem_23_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93323),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1670_1671_LC_8_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1670_1671_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1670_1671_LC_8_4_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1670_1671_LC_8_4_6  (
            .in0(N__39486),
            .in1(N__71524),
            .in2(_gnd_net_),
            .in3(N__66578),
            .lcout(REG_mem_17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93323),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i425_426_LC_8_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i425_426_LC_8_4_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i425_426_LC_8_4_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i425_426_LC_8_4_7  (
            .in0(N__72709),
            .in1(N__48117),
            .in2(_gnd_net_),
            .in3(N__96807),
            .lcout(REG_mem_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93323),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11251_LC_8_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11251_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11251_LC_8_5_0 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11251_LC_8_5_0  (
            .in0(N__87647),
            .in1(N__45109),
            .in2(N__92588),
            .in3(N__43549),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12920 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10796_3_lut_LC_8_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10796_3_lut_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10796_3_lut_LC_8_5_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10796_3_lut_LC_8_5_1  (
            .in0(N__39658),
            .in1(N__87646),
            .in2(_gnd_net_),
            .in3(N__43258),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10445_3_lut_LC_8_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10445_3_lut_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10445_3_lut_LC_8_5_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10445_3_lut_LC_8_5_2  (
            .in0(N__85662),
            .in1(N__41209),
            .in2(_gnd_net_),
            .in3(N__53746),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12094 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12938_bdd_4_lut_LC_8_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12938_bdd_4_lut_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12938_bdd_4_lut_LC_8_5_3 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12938_bdd_4_lut_LC_8_5_3  (
            .in0(N__41218),
            .in1(N__92380),
            .in2(N__41353),
            .in3(N__39643),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12941_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10446_3_lut_LC_8_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10446_3_lut_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10446_3_lut_LC_8_5_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10446_3_lut_LC_8_5_4  (
            .in0(N__85663),
            .in1(_gnd_net_),
            .in2(N__39625),
            .in3(N__39622),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12095_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14078_bdd_4_lut_LC_8_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14078_bdd_4_lut_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14078_bdd_4_lut_LC_8_5_5 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14078_bdd_4_lut_LC_8_5_5  (
            .in0(N__81433),
            .in1(N__48016),
            .in2(N__39613),
            .in3(N__39610),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4358_4359_LC_8_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4358_4359_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4358_4359_LC_8_5_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4358_4359_LC_8_5_6  (
            .in0(_gnd_net_),
            .in1(N__39600),
            .in2(N__71568),
            .in3(N__71886),
            .lcout(REG_mem_45_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93310),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5240_5241_LC_8_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5240_5241_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5240_5241_LC_8_6_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5240_5241_LC_8_6_0  (
            .in0(N__94168),
            .in1(N__96391),
            .in2(N__75117),
            .in3(N__76255),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93296),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1967_1968_LC_8_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1967_1968_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1967_1968_LC_8_6_1 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1967_1968_LC_8_6_1  (
            .in0(N__61295),
            .in1(N__94171),
            .in2(N__39589),
            .in3(N__77439),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93296),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5930_5931_LC_8_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5930_5931_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5930_5931_LC_8_6_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5930_5931_LC_8_6_2  (
            .in0(N__94169),
            .in1(N__46579),
            .in2(N__39567),
            .in3(N__70937),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93296),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1973_1974_LC_8_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1973_1974_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1973_1974_LC_8_6_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1973_1974_LC_8_6_3  (
            .in0(N__62791),
            .in1(N__94172),
            .in2(N__55899),
            .in3(N__77440),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93296),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4277_4278_LC_8_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4277_4278_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4277_4278_LC_8_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4277_4278_LC_8_6_4  (
            .in0(N__51546),
            .in1(N__62792),
            .in2(_gnd_net_),
            .in3(N__71703),
            .lcout(REG_mem_44_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93296),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1958_1959_LC_8_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1958_1959_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1958_1959_LC_8_6_5 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1958_1959_LC_8_6_5  (
            .in0(N__39543),
            .in1(N__94170),
            .in2(N__77466),
            .in3(N__71528),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93296),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2003_2004_LC_8_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2003_2004_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2003_2004_LC_8_6_6 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2003_2004_LC_8_6_6  (
            .in0(N__77438),
            .in1(N__39750),
            .in2(N__94602),
            .in3(N__62317),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93296),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10655_3_lut_LC_8_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10655_3_lut_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10655_3_lut_LC_8_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10655_3_lut_LC_8_6_7  (
            .in0(N__39856),
            .in1(N__48223),
            .in2(_gnd_net_),
            .in3(N__87356),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1235_1236_LC_8_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1235_1236_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1235_1236_LC_8_7_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1235_1236_LC_8_7_0  (
            .in0(N__39729),
            .in1(_gnd_net_),
            .in2(N__62430),
            .in3(N__59600),
            .lcout(REG_mem_12_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2918_2919_LC_8_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2918_2919_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2918_2919_LC_8_7_1 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2918_2919_LC_8_7_1  (
            .in0(N__71561),
            .in1(N__95224),
            .in2(N__39714),
            .in3(N__77744),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i752_753_LC_8_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i752_753_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i752_753_LC_8_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i752_753_LC_8_7_2  (
            .in0(N__39684),
            .in1(N__41784),
            .in2(_gnd_net_),
            .in3(N__89649),
            .lcout(REG_mem_7_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3905_3906_LC_8_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3905_3906_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3905_3906_LC_8_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3905_3906_LC_8_7_3  (
            .in0(N__56555),
            .in1(N__39669),
            .in2(_gnd_net_),
            .in3(N__65803),
            .lcout(REG_mem_40_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4673_4674_LC_8_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4673_4674_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4673_4674_LC_8_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4673_4674_LC_8_7_4  (
            .in0(N__39654),
            .in1(N__56556),
            .in2(_gnd_net_),
            .in3(N__75473),
            .lcout(REG_mem_48_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3509_3510_LC_8_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3509_3510_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3509_3510_LC_8_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3509_3510_LC_8_7_5  (
            .in0(N__48090),
            .in1(N__62688),
            .in2(_gnd_net_),
            .in3(N__54041),
            .lcout(REG_mem_36_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1601_1602_LC_8_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1601_1602_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1601_1602_LC_8_7_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1601_1602_LC_8_7_6  (
            .in0(N__43287),
            .in1(N__65604),
            .in2(_gnd_net_),
            .in3(N__56557),
            .lcout(REG_mem_16_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2342_2343_LC_8_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2342_2343_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2342_2343_LC_8_7_7 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2342_2343_LC_8_7_7  (
            .in0(N__71560),
            .in1(N__95223),
            .in2(N__39831),
            .in3(N__95890),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93284),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i101_2_lut_3_lut_4_lut_LC_8_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i101_2_lut_3_lut_4_lut_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i101_2_lut_3_lut_4_lut_LC_8_8_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i101_2_lut_3_lut_4_lut_LC_8_8_0  (
            .in0(N__49539),
            .in1(N__49846),
            .in2(N__94595),
            .in3(N__42111),
            .lcout(n17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i102_2_lut_3_lut_4_lut_LC_8_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i102_2_lut_3_lut_4_lut_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i102_2_lut_3_lut_4_lut_LC_8_8_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i102_2_lut_3_lut_4_lut_LC_8_8_1  (
            .in0(N__42112),
            .in1(N__94142),
            .in2(N__49859),
            .in3(N__49541),
            .lcout(n49),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i85_2_lut_3_lut_4_lut_LC_8_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i85_2_lut_3_lut_4_lut_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i85_2_lut_3_lut_4_lut_LC_8_8_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i85_2_lut_3_lut_4_lut_LC_8_8_2  (
            .in0(N__49540),
            .in1(N__49850),
            .in2(N__94596),
            .in3(N__42113),
            .lcout(n25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i86_2_lut_3_lut_4_lut_LC_8_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i86_2_lut_3_lut_4_lut_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i86_2_lut_3_lut_4_lut_LC_8_8_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i86_2_lut_3_lut_4_lut_LC_8_8_3  (
            .in0(N__42114),
            .in1(N__94141),
            .in2(N__49858),
            .in3(N__49537),
            .lcout(n57),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i53_2_lut_3_lut_LC_8_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i53_2_lut_3_lut_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i53_2_lut_3_lut_LC_8_8_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i53_2_lut_3_lut_LC_8_8_4  (
            .in0(N__49538),
            .in1(N__49845),
            .in2(_gnd_net_),
            .in3(N__42110),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53 ),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n53_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5414_5415_LC_8_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5414_5415_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5414_5415_LC_8_8_5 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5414_5415_LC_8_8_5  (
            .in0(N__39804),
            .in1(N__71559),
            .in2(N__39814),
            .in3(N__94150),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93273),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4016_4017_LC_8_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4016_4017_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4016_4017_LC_8_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4016_4017_LC_8_8_6  (
            .in0(N__39783),
            .in1(N__41802),
            .in2(_gnd_net_),
            .in3(N__66003),
            .lcout(REG_mem_41_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93273),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5162_5163_LC_8_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5162_5163_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5162_5163_LC_8_8_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5162_5163_LC_8_8_7  (
            .in0(N__46452),
            .in1(N__94149),
            .in2(N__39772),
            .in3(N__76841),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93273),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i77_2_lut_3_lut_4_lut_LC_8_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i77_2_lut_3_lut_4_lut_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i77_2_lut_3_lut_4_lut_LC_8_9_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i77_2_lut_3_lut_4_lut_LC_8_9_0  (
            .in0(N__49547),
            .in1(N__49878),
            .in2(N__94599),
            .in3(N__41965),
            .lcout(n29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i78_2_lut_3_lut_4_lut_LC_8_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i78_2_lut_3_lut_4_lut_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i78_2_lut_3_lut_4_lut_LC_8_9_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i78_2_lut_3_lut_4_lut_LC_8_9_1  (
            .in0(N__41966),
            .in1(N__49549),
            .in2(N__49885),
            .in3(N__94160),
            .lcout(n61),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i93_2_lut_3_lut_4_lut_LC_8_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i93_2_lut_3_lut_4_lut_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i93_2_lut_3_lut_4_lut_LC_8_9_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i93_2_lut_3_lut_4_lut_LC_8_9_2  (
            .in0(N__49546),
            .in1(N__49877),
            .in2(N__94598),
            .in3(N__41967),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5837_5838_LC_8_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5837_5838_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5837_5838_LC_8_9_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5837_5838_LC_8_9_3  (
            .in0(N__46773),
            .in1(N__94162),
            .in2(N__39918),
            .in3(N__70570),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93264),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i45_2_lut_3_lut_LC_8_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i45_2_lut_3_lut_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i45_2_lut_3_lut_LC_8_9_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i45_2_lut_3_lut_LC_8_9_4  (
            .in0(N__49548),
            .in1(N__49882),
            .in2(_gnd_net_),
            .in3(N__41964),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2765_2766_LC_8_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2765_2766_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2765_2766_LC_8_9_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2765_2766_LC_8_9_5  (
            .in0(N__46772),
            .in1(N__94161),
            .in2(N__39894),
            .in3(N__70569),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93264),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i94_2_lut_3_lut_4_lut_LC_8_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i94_2_lut_3_lut_4_lut_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i94_2_lut_3_lut_4_lut_LC_8_9_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i94_2_lut_3_lut_4_lut_LC_8_9_6  (
            .in0(N__49545),
            .in1(N__49876),
            .in2(N__94597),
            .in3(N__41968),
            .lcout(n53),
            .ltout(n53_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1196_1197_LC_8_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1196_1197_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1196_1197_LC_8_9_7 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1196_1197_LC_8_9_7  (
            .in0(N__76003),
            .in1(N__59478),
            .in2(N__39877),
            .in3(_gnd_net_),
            .lcout(REG_mem_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93264),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5990_5991_LC_8_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5990_5991_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5990_5991_LC_8_10_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5990_5991_LC_8_10_0  (
            .in0(N__39867),
            .in1(N__71558),
            .in2(N__77968),
            .in3(N__95076),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5045_5046_LC_8_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5045_5046_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5045_5046_LC_8_10_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5045_5046_LC_8_10_1  (
            .in0(N__95075),
            .in1(N__62690),
            .in2(N__39852),
            .in3(N__77390),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1205_1206_LC_8_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1205_1206_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1205_1206_LC_8_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1205_1206_LC_8_10_2  (
            .in0(N__58671),
            .in1(N__62689),
            .in2(_gnd_net_),
            .in3(N__59564),
            .lcout(REG_mem_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i63_2_lut_3_lut_4_lut_LC_8_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i63_2_lut_3_lut_4_lut_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i63_2_lut_3_lut_4_lut_LC_8_10_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i63_2_lut_3_lut_4_lut_LC_8_10_3  (
            .in0(N__50026),
            .in1(N__49857),
            .in2(N__49594),
            .in3(N__43723),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n63 ),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n63_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2822_2823_LC_8_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2822_2823_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2822_2823_LC_8_10_4 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2822_2823_LC_8_10_4  (
            .in0(N__40017),
            .in1(N__71557),
            .in2(N__40027),
            .in3(N__95077),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4880_4881_LC_8_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4880_4881_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4880_4881_LC_8_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4880_4881_LC_8_10_5  (
            .in0(N__39987),
            .in1(N__41797),
            .in2(_gnd_net_),
            .in3(N__72981),
            .lcout(REG_mem_50_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i49_2_lut_3_lut_4_lut_LC_8_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i49_2_lut_3_lut_4_lut_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i49_2_lut_3_lut_4_lut_LC_8_10_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i49_2_lut_3_lut_4_lut_LC_8_10_6  (
            .in0(N__49856),
            .in1(N__50027),
            .in2(N__49595),
            .in3(N__43654),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4295_4296_LC_8_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4295_4296_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4295_4296_LC_8_10_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4295_4296_LC_8_10_7  (
            .in0(N__39969),
            .in1(N__47338),
            .in2(_gnd_net_),
            .in3(N__71657),
            .lcout(REG_mem_44_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93250),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5222_5223_LC_8_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5222_5223_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5222_5223_LC_8_11_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5222_5223_LC_8_11_0  (
            .in0(N__71498),
            .in1(N__93931),
            .in2(N__41379),
            .in3(N__76134),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5819_5820_LC_8_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5819_5820_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5819_5820_LC_8_11_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5819_5820_LC_8_11_1  (
            .in0(N__93929),
            .in1(N__63504),
            .in2(N__39958),
            .in3(N__70585),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i65_66_LC_8_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i65_66_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i65_66_LC_8_11_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i65_66_LC_8_11_2  (
            .in0(N__56599),
            .in1(N__93932),
            .in2(N__40144),
            .in3(N__82885),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5435_5436_LC_8_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5435_5436_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5435_5436_LC_8_11_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5435_5436_LC_8_11_3  (
            .in0(N__93928),
            .in1(N__63503),
            .in2(N__39942),
            .in3(N__95937),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10691_3_lut_LC_8_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10691_3_lut_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10691_3_lut_LC_8_11_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10691_3_lut_LC_8_11_4  (
            .in0(N__40143),
            .in1(N__87793),
            .in2(_gnd_net_),
            .in3(N__40132),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i74_75_LC_8_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i74_75_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i74_75_LC_8_11_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i74_75_LC_8_11_5  (
            .in0(N__93930),
            .in1(N__46456),
            .in2(N__40086),
            .in3(N__82886),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4481_4482_LC_8_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4481_4482_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4481_4482_LC_8_11_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4481_4482_LC_8_11_6  (
            .in0(N__89039),
            .in1(_gnd_net_),
            .in2(N__56620),
            .in3(N__40065),
            .lcout(REG_mem_46_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4466_4467_LC_8_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4466_4467_LC_8_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4466_4467_LC_8_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4466_4467_LC_8_11_7  (
            .in0(N__76695),
            .in1(N__57060),
            .in2(_gnd_net_),
            .in3(N__89038),
            .lcout(REG_mem_46_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93265),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i815_816_LC_8_12_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i815_816_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i815_816_LC_8_12_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i815_816_LC_8_12_0  (
            .in0(N__40053),
            .in1(N__61288),
            .in2(_gnd_net_),
            .in3(N__67266),
            .lcout(REG_mem_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3494_3495_LC_8_12_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3494_3495_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3494_3495_LC_8_12_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3494_3495_LC_8_12_1  (
            .in0(N__53757),
            .in1(N__71556),
            .in2(_gnd_net_),
            .in3(N__54064),
            .lcout(REG_mem_36_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3527_3528_LC_8_12_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3527_3528_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3527_3528_LC_8_12_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3527_3528_LC_8_12_2  (
            .in0(N__54063),
            .in1(N__40242),
            .in2(_gnd_net_),
            .in3(N__47314),
            .lcout(REG_mem_36_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3623_3624_LC_8_12_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3623_3624_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3623_3624_LC_8_12_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3623_3624_LC_8_12_3  (
            .in0(N__47311),
            .in1(N__40257),
            .in2(_gnd_net_),
            .in3(N__63712),
            .lcout(REG_mem_37_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3911_3912_LC_8_12_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3911_3912_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3911_3912_LC_8_12_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3911_3912_LC_8_12_4  (
            .in0(N__40038),
            .in1(N__47312),
            .in2(_gnd_net_),
            .in3(N__65879),
            .lcout(REG_mem_40_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4592_4593_LC_8_12_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4592_4593_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4592_4593_LC_8_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4592_4593_LC_8_12_5  (
            .in0(N__40221),
            .in1(N__41670),
            .in2(_gnd_net_),
            .in3(N__66255),
            .lcout(REG_mem_47_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3239_3240_LC_8_12_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3239_3240_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3239_3240_LC_8_12_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3239_3240_LC_8_12_6  (
            .in0(N__94233),
            .in1(N__47313),
            .in2(N__40209),
            .in3(N__80215),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2159_2160_LC_8_12_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2159_2160_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2159_2160_LC_8_12_7 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2159_2160_LC_8_12_7  (
            .in0(N__76195),
            .in1(N__61289),
            .in2(N__40188),
            .in3(N__94234),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93274),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4271_4272_LC_8_13_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4271_4272_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4271_4272_LC_8_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4271_4272_LC_8_13_0  (
            .in0(N__71710),
            .in1(N__40170),
            .in2(_gnd_net_),
            .in3(N__61290),
            .lcout(REG_mem_44_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3722_3723_LC_8_13_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3722_3723_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3722_3723_LC_8_13_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3722_3723_LC_8_13_1  (
            .in0(N__59282),
            .in1(N__40299),
            .in2(_gnd_net_),
            .in3(N__46455),
            .lcout(REG_mem_38_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i80_81_LC_8_13_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i80_81_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i80_81_LC_8_13_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i80_81_LC_8_13_2  (
            .in0(N__95446),
            .in1(N__41803),
            .in2(N__41046),
            .in3(N__82887),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3716_3717_LC_8_13_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3716_3717_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3716_3717_LC_8_13_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3716_3717_LC_8_13_3  (
            .in0(N__59281),
            .in1(_gnd_net_),
            .in2(N__50694),
            .in3(N__48760),
            .lcout(REG_mem_38_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3917_3918_LC_8_13_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3917_3918_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3917_3918_LC_8_13_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3917_3918_LC_8_13_4  (
            .in0(N__40410),
            .in1(N__46774),
            .in2(_gnd_net_),
            .in3(N__65896),
            .lcout(REG_mem_40_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3530_3531_LC_8_13_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3530_3531_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3530_3531_LC_8_13_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3530_3531_LC_8_13_5  (
            .in0(N__54072),
            .in1(N__40155),
            .in2(_gnd_net_),
            .in3(N__46454),
            .lcout(REG_mem_36_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3626_3627_LC_8_13_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3626_3627_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3626_3627_LC_8_13_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3626_3627_LC_8_13_6  (
            .in0(N__46453),
            .in1(_gnd_net_),
            .in2(N__40350),
            .in3(N__63713),
            .lcout(REG_mem_37_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1607_1608_LC_8_13_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1607_1608_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1607_1608_LC_8_13_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1607_1608_LC_8_13_7  (
            .in0(N__40764),
            .in1(N__47337),
            .in2(_gnd_net_),
            .in3(N__65664),
            .lcout(REG_mem_16_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93285),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1706_1707_LC_8_14_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1706_1707_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1706_1707_LC_8_14_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1706_1707_LC_8_14_0  (
            .in0(N__46462),
            .in1(N__40332),
            .in2(_gnd_net_),
            .in3(N__66587),
            .lcout(REG_mem_17_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93297),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11655_LC_8_14_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11655_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11655_LC_8_14_1 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11655_LC_8_14_1  (
            .in0(N__87427),
            .in1(N__91327),
            .in2(N__42466),
            .in3(N__44563),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13406_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13406_bdd_4_lut_LC_8_14_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13406_bdd_4_lut_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13406_bdd_4_lut_LC_8_14_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13406_bdd_4_lut_LC_8_14_2  (
            .in0(N__91325),
            .in1(N__40333),
            .in2(N__40324),
            .in3(N__40309),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1610_1611_LC_8_14_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1610_1611_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1610_1611_LC_8_14_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1610_1611_LC_8_14_3  (
            .in0(N__40308),
            .in1(N__46464),
            .in2(_gnd_net_),
            .in3(N__65665),
            .lcout(REG_mem_16_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93297),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10833_3_lut_LC_8_14_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10833_3_lut_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10833_3_lut_LC_8_14_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10833_3_lut_LC_8_14_4  (
            .in0(N__42052),
            .in1(N__40300),
            .in2(_gnd_net_),
            .in3(N__87426),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i845_846_LC_8_14_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i845_846_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i845_846_LC_8_14_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i845_846_LC_8_14_5  (
            .in0(N__40431),
            .in1(N__46775),
            .in2(_gnd_net_),
            .in3(N__67278),
            .lcout(REG_mem_8_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93297),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i458_459_LC_8_14_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i458_459_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i458_459_LC_8_14_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i458_459_LC_8_14_6  (
            .in0(N__46463),
            .in1(N__40272),
            .in2(_gnd_net_),
            .in3(N__72700),
            .lcout(REG_mem_4_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93297),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13424_bdd_4_lut_LC_8_14_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13424_bdd_4_lut_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13424_bdd_4_lut_LC_8_14_7 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13424_bdd_4_lut_LC_8_14_7  (
            .in0(N__40261),
            .in1(N__91326),
            .in2(N__44440),
            .in3(N__40246),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13427 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11983_LC_8_15_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11983_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11983_LC_8_15_0 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11983_LC_8_15_0  (
            .in0(N__87472),
            .in1(N__45583),
            .in2(N__42325),
            .in3(N__90709),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13802_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13802_bdd_4_lut_LC_8_15_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13802_bdd_4_lut_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13802_bdd_4_lut_LC_8_15_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13802_bdd_4_lut_LC_8_15_1  (
            .in0(N__90707),
            .in1(N__40414),
            .in2(N__40399),
            .in3(N__44326),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11316_LC_8_15_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11316_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11316_LC_8_15_2 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11316_LC_8_15_2  (
            .in0(N__89953),
            .in1(N__40384),
            .in2(N__40396),
            .in3(N__85101),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12968 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13712_bdd_4_lut_LC_8_15_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13712_bdd_4_lut_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13712_bdd_4_lut_LC_8_15_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13712_bdd_4_lut_LC_8_15_3  (
            .in0(N__90706),
            .in1(N__46627),
            .in2(N__40378),
            .in3(N__40369),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11909_LC_8_15_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11909_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11909_LC_8_15_4 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11909_LC_8_15_4  (
            .in0(N__40360),
            .in1(N__90708),
            .in2(N__87733),
            .in3(N__45808),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i743_744_LC_8_15_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i743_744_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i743_744_LC_8_15_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i743_744_LC_8_15_5  (
            .in0(N__40578),
            .in1(N__47310),
            .in2(_gnd_net_),
            .in3(N__89671),
            .lcout(REG_mem_7_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93311),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4301_4302_LC_8_15_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4301_4302_LC_8_15_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4301_4302_LC_8_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4301_4302_LC_8_15_6  (
            .in0(N__40368),
            .in1(N__46855),
            .in2(_gnd_net_),
            .in3(N__71711),
            .lcout(REG_mem_44_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93311),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4493_4494_LC_8_15_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4493_4494_LC_8_15_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4493_4494_LC_8_15_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4493_4494_LC_8_15_7  (
            .in0(N__46854),
            .in1(N__40359),
            .in2(_gnd_net_),
            .in3(N__89073),
            .lcout(REG_mem_46_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93311),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5357_5358_LC_8_16_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5357_5358_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5357_5358_LC_8_16_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5357_5358_LC_8_16_0  (
            .in0(N__40560),
            .in1(N__46856),
            .in2(_gnd_net_),
            .in3(N__77240),
            .lcout(REG_mem_55_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93324),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11739_LC_8_16_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11739_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11739_LC_8_16_1 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11739_LC_8_16_1  (
            .in0(N__91366),
            .in1(N__40561),
            .in2(N__40489),
            .in3(N__87176),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13508_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13508_bdd_4_lut_LC_8_16_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13508_bdd_4_lut_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13508_bdd_4_lut_LC_8_16_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13508_bdd_4_lut_LC_8_16_2  (
            .in0(N__40500),
            .in1(N__91364),
            .in2(N__40552),
            .in3(N__40549),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3908_3909_LC_8_16_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3908_3909_LC_8_16_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3908_3909_LC_8_16_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3908_3909_LC_8_16_3  (
            .in0(N__40518),
            .in1(N__48892),
            .in2(_gnd_net_),
            .in3(N__65897),
            .lcout(REG_mem_40_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93324),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5069_5070_LC_8_16_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5069_5070_LC_8_16_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5069_5070_LC_8_16_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5069_5070_LC_8_16_4  (
            .in0(N__47014),
            .in1(N__94237),
            .in2(N__40501),
            .in3(N__77456),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93324),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5261_5262_LC_8_16_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5261_5262_LC_8_16_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5261_5262_LC_8_16_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5261_5262_LC_8_16_5  (
            .in0(N__94235),
            .in1(N__47015),
            .in2(N__40488),
            .in3(N__76268),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93324),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1997_1998_LC_8_16_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1997_1998_LC_8_16_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1997_1998_LC_8_16_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1997_1998_LC_8_16_6  (
            .in0(N__47013),
            .in1(N__94236),
            .in2(N__40474),
            .in3(N__77455),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93324),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14066_bdd_4_lut_LC_8_16_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14066_bdd_4_lut_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14066_bdd_4_lut_LC_8_16_7 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14066_bdd_4_lut_LC_8_16_7  (
            .in0(N__91365),
            .in1(N__40690),
            .in2(N__42349),
            .in3(N__40473),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12258_LC_8_17_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12258_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12258_LC_8_17_0 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12258_LC_8_17_0  (
            .in0(N__40597),
            .in1(N__91569),
            .in2(N__87296),
            .in3(N__45604),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14174_bdd_4_lut_LC_8_17_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14174_bdd_4_lut_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14174_bdd_4_lut_LC_8_17_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14174_bdd_4_lut_LC_8_17_1  (
            .in0(N__91568),
            .in1(N__42409),
            .in2(N__40450),
            .in3(N__40435),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12075_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11380_LC_8_17_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11380_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11380_LC_8_17_2 .LUT_INIT=16'b1011100011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11380_LC_8_17_2  (
            .in0(N__40639),
            .in1(N__85006),
            .in2(N__40657),
            .in3(N__89942),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13076 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14126_bdd_4_lut_LC_8_17_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14126_bdd_4_lut_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14126_bdd_4_lut_LC_8_17_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14126_bdd_4_lut_LC_8_17_3  (
            .in0(N__91567),
            .in1(N__40615),
            .in2(N__40648),
            .in3(N__40606),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i170_171_LC_8_17_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i170_171_LC_8_17_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i170_171_LC_8_17_4 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i170_171_LC_8_17_4  (
            .in0(N__94238),
            .in1(N__40626),
            .in2(N__46587),
            .in3(N__80298),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93337),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1325_1326_LC_8_17_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1325_1326_LC_8_17_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1325_1326_LC_8_17_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1325_1326_LC_8_17_5  (
            .in0(N__46963),
            .in1(N__40614),
            .in2(_gnd_net_),
            .in3(N__70139),
            .lcout(REG_mem_13_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93337),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1229_1230_LC_8_17_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1229_1230_LC_8_17_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1229_1230_LC_8_17_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1229_1230_LC_8_17_6  (
            .in0(N__40605),
            .in1(N__46965),
            .in2(_gnd_net_),
            .in3(N__59651),
            .lcout(REG_mem_12_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93337),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1421_1422_LC_8_17_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1421_1422_LC_8_17_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1421_1422_LC_8_17_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1421_1422_LC_8_17_7  (
            .in0(N__46964),
            .in1(N__40596),
            .in2(_gnd_net_),
            .in3(N__74762),
            .lcout(REG_mem_14_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93337),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11221_LC_8_18_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11221_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11221_LC_8_18_0 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11221_LC_8_18_0  (
            .in0(N__91572),
            .in1(N__86919),
            .in2(N__47062),
            .in3(N__40588),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12884_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12884_bdd_4_lut_LC_8_18_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12884_bdd_4_lut_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12884_bdd_4_lut_LC_8_18_1 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12884_bdd_4_lut_LC_8_18_1  (
            .in0(N__46009),
            .in1(N__91570),
            .in2(N__40567),
            .in3(N__42244),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12887_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13154_bdd_4_lut_LC_8_18_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13154_bdd_4_lut_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13154_bdd_4_lut_LC_8_18_2 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13154_bdd_4_lut_LC_8_18_2  (
            .in0(N__44605),
            .in1(N__89876),
            .in2(N__40564),
            .in3(N__40714),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13157 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4685_4686_LC_8_18_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4685_4686_LC_8_18_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4685_4686_LC_8_18_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4685_4686_LC_8_18_3  (
            .in0(N__44640),
            .in1(N__46857),
            .in2(_gnd_net_),
            .in3(N__75584),
            .lcout(REG_mem_48_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93351),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12950_bdd_4_lut_LC_8_18_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12950_bdd_4_lut_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12950_bdd_4_lut_LC_8_18_4 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12950_bdd_4_lut_LC_8_18_4  (
            .in0(N__91571),
            .in1(N__40663),
            .in2(N__42199),
            .in3(N__42739),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12953 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3245_3246_LC_8_18_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3245_3246_LC_8_18_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3245_3246_LC_8_18_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3245_3246_LC_8_18_5  (
            .in0(N__46935),
            .in1(N__94244),
            .in2(N__42888),
            .in3(N__80302),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93351),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12203_LC_8_18_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12203_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12203_LC_8_18_6 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12203_LC_8_18_6  (
            .in0(N__91573),
            .in1(N__42694),
            .in2(N__40708),
            .in3(N__86920),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14066 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1799_1800_LC_8_19_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1799_1800_LC_8_19_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1799_1800_LC_8_19_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1799_1800_LC_8_19_1  (
            .in0(N__40782),
            .in1(N__47391),
            .in2(_gnd_net_),
            .in3(N__67504),
            .lcout(REG_mem_18_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5255_5256_LC_8_19_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5255_5256_LC_8_19_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5255_5256_LC_8_19_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5255_5256_LC_8_19_2  (
            .in0(N__76334),
            .in1(N__42903),
            .in2(N__47443),
            .in3(N__94243),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2183_2184_LC_8_19_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2183_2184_LC_8_19_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2183_2184_LC_8_19_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2183_2184_LC_8_19_3  (
            .in0(N__94239),
            .in1(N__47392),
            .in2(N__40804),
            .in3(N__76333),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i263_264_LC_8_19_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i263_264_LC_8_19_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i263_264_LC_8_19_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i263_264_LC_8_19_4  (
            .in0(N__47390),
            .in1(N__94242),
            .in2(N__40680),
            .in3(N__80608),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11276_LC_8_19_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11276_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11276_LC_8_19_5 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11276_LC_8_19_5  (
            .in0(N__42586),
            .in1(N__91574),
            .in2(N__40681),
            .in3(N__86861),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12950 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1991_1992_LC_8_19_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1991_1992_LC_8_19_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1991_1992_LC_8_19_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1991_1992_LC_8_19_6  (
            .in0(N__47389),
            .in1(N__94241),
            .in2(N__40738),
            .in3(N__77457),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5063_5064_LC_8_19_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5063_5064_LC_8_19_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5063_5064_LC_8_19_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5063_5064_LC_8_19_7  (
            .in0(N__94240),
            .in1(N__47393),
            .in2(N__44850),
            .in3(N__77458),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93366),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11685_LC_8_20_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11685_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11685_LC_8_20_0 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11685_LC_8_20_0  (
            .in0(N__91987),
            .in1(N__86921),
            .in2(N__42613),
            .in3(N__40803),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12483_LC_8_20_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12483_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12483_LC_8_20_1 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12483_LC_8_20_1  (
            .in0(N__89826),
            .in1(N__42622),
            .in2(N__85005),
            .in3(N__44746),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14366_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14366_bdd_4_lut_LC_8_20_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14366_bdd_4_lut_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14366_bdd_4_lut_LC_8_20_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14366_bdd_4_lut_LC_8_20_2  (
            .in0(N__40723),
            .in1(N__89825),
            .in2(N__40789),
            .in3(N__40753),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12463_LC_8_20_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12463_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12463_LC_8_20_3 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12463_LC_8_20_3  (
            .in0(N__86922),
            .in1(N__91988),
            .in2(N__40786),
            .in3(N__44503),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14378_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14378_bdd_4_lut_LC_8_20_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14378_bdd_4_lut_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14378_bdd_4_lut_LC_8_20_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14378_bdd_4_lut_LC_8_20_4  (
            .in0(N__91986),
            .in1(N__42286),
            .in2(N__40771),
            .in3(N__40768),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12471 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13436_bdd_4_lut_LC_8_20_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13436_bdd_4_lut_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13436_bdd_4_lut_LC_8_20_5 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13436_bdd_4_lut_LC_8_20_5  (
            .in0(N__44596),
            .in1(N__91985),
            .in2(N__40747),
            .in3(N__40737),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13439 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i3_LC_8_20_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i3_LC_8_20_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i3_LC_8_20_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i3_LC_8_20_6  (
            .in0(N__42717),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73482),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97356),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10049_3_lut_LC_9_1_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10049_3_lut_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10049_3_lut_LC_9_1_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10049_3_lut_LC_9_1_0  (
            .in0(N__40872),
            .in1(N__40884),
            .in2(_gnd_net_),
            .in3(N__88000),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3113_3114_LC_9_1_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3113_3114_LC_9_1_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3113_3114_LC_9_1_1 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3113_3114_LC_9_1_1  (
            .in0(N__96812),
            .in1(N__95546),
            .in2(N__40885),
            .in3(N__82869),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3209_3210_LC_9_1_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3209_3210_LC_9_1_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3209_3210_LC_9_1_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3209_3210_LC_9_1_2  (
            .in0(N__95545),
            .in1(N__96813),
            .in2(N__40873),
            .in3(N__80287),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i41_42_LC_9_1_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i41_42_LC_9_1_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i41_42_LC_9_1_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i41_42_LC_9_1_3  (
            .in0(N__96814),
            .in1(N__95549),
            .in2(N__40834),
            .in3(N__82871),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i83_84_LC_9_1_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i83_84_LC_9_1_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i83_84_LC_9_1_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i83_84_LC_9_1_4  (
            .in0(N__82872),
            .in1(N__44712),
            .in2(N__95704),
            .in3(N__62350),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3155_3156_LC_9_1_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3155_3156_LC_9_1_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3155_3156_LC_9_1_5 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3155_3156_LC_9_1_5  (
            .in0(N__62349),
            .in1(N__95547),
            .in2(N__40861),
            .in3(N__82870),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10337_3_lut_LC_9_1_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10337_3_lut_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10337_3_lut_LC_9_1_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10337_3_lut_LC_9_1_6  (
            .in0(N__40860),
            .in1(N__40845),
            .in2(_gnd_net_),
            .in3(N__88001),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11986 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3251_3252_LC_9_1_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3251_3252_LC_9_1_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3251_3252_LC_9_1_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3251_3252_LC_9_1_7  (
            .in0(N__80288),
            .in1(N__95548),
            .in2(N__40846),
            .in3(N__62352),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93380),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10004_3_lut_LC_9_2_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10004_3_lut_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10004_3_lut_LC_9_2_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10004_3_lut_LC_9_2_0  (
            .in0(N__40833),
            .in1(N__87661),
            .in2(_gnd_net_),
            .in3(N__40818),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11874_LC_9_2_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11874_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11874_LC_9_2_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11874_LC_9_2_1  (
            .in0(N__85806),
            .in1(N__92584),
            .in2(N__54145),
            .in3(N__43387),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13670_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13670_bdd_4_lut_LC_9_2_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13670_bdd_4_lut_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13670_bdd_4_lut_LC_9_2_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13670_bdd_4_lut_LC_9_2_2  (
            .in0(N__40957),
            .in1(N__85804),
            .in2(N__40951),
            .in3(N__42940),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13673 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12298_LC_9_2_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12298_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12298_LC_9_2_3 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12298_LC_9_2_3  (
            .in0(N__85807),
            .in1(N__40948),
            .in2(N__45187),
            .in3(N__92585),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14156 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13676_bdd_4_lut_LC_9_2_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13676_bdd_4_lut_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13676_bdd_4_lut_LC_9_2_4 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13676_bdd_4_lut_LC_9_2_4  (
            .in0(N__40942),
            .in1(N__85805),
            .in2(N__40930),
            .in3(N__45037),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13679_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12333_LC_9_2_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12333_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12333_LC_9_2_5 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12333_LC_9_2_5  (
            .in0(N__90386),
            .in1(N__81439),
            .in2(N__40912),
            .in3(N__40909),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10349_3_lut_LC_9_2_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10349_3_lut_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10349_3_lut_LC_9_2_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10349_3_lut_LC_9_2_6  (
            .in0(N__42034),
            .in1(N__40897),
            .in2(_gnd_net_),
            .in3(N__87662),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11998 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10082_3_lut_LC_9_3_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10082_3_lut_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10082_3_lut_LC_9_3_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10082_3_lut_LC_9_3_0  (
            .in0(N__41200),
            .in1(N__87648),
            .in2(_gnd_net_),
            .in3(N__53089),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11731 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10083_3_lut_LC_9_3_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10083_3_lut_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10083_3_lut_LC_9_3_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10083_3_lut_LC_9_3_1  (
            .in0(N__87649),
            .in1(N__40993),
            .in2(_gnd_net_),
            .in3(N__43039),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11732 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1121_1122_LC_9_3_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1121_1122_LC_9_3_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1121_1122_LC_9_3_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1121_1122_LC_9_3_2  (
            .in0(N__43170),
            .in1(N__56474),
            .in2(_gnd_net_),
            .in3(N__66816),
            .lcout(REG_mem_11_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93354),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i737_738_LC_9_3_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i737_738_LC_9_3_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i737_738_LC_9_3_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i737_738_LC_9_3_3  (
            .in0(N__56473),
            .in1(N__41154),
            .in2(_gnd_net_),
            .in3(N__89663),
            .lcout(REG_mem_7_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93354),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10695_3_lut_LC_9_3_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10695_3_lut_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10695_3_lut_LC_9_3_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10695_3_lut_LC_9_3_4  (
            .in0(N__41155),
            .in1(N__87650),
            .in2(_gnd_net_),
            .in3(N__56212),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13706_bdd_4_lut_LC_9_3_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13706_bdd_4_lut_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13706_bdd_4_lut_LC_9_3_5 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13706_bdd_4_lut_LC_9_3_5  (
            .in0(N__41062),
            .in1(N__81437),
            .in2(N__41131),
            .in3(N__45046),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13709 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14156_bdd_4_lut_LC_9_3_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14156_bdd_4_lut_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14156_bdd_4_lut_LC_9_3_6 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14156_bdd_4_lut_LC_9_3_6  (
            .in0(N__85748),
            .in1(N__41116),
            .in2(N__41110),
            .in3(N__41101),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12080_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14114_bdd_4_lut_LC_9_3_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14114_bdd_4_lut_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14114_bdd_4_lut_LC_9_3_7 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14114_bdd_4_lut_LC_9_3_7  (
            .in0(N__41092),
            .in1(N__81438),
            .in2(N__41086),
            .in3(N__41083),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13562_bdd_4_lut_LC_9_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13562_bdd_4_lut_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13562_bdd_4_lut_LC_9_4_0 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13562_bdd_4_lut_LC_9_4_0  (
            .in0(N__85661),
            .in1(N__48385),
            .in2(N__41077),
            .in3(N__41068),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13565 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10535_3_lut_LC_9_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10535_3_lut_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10535_3_lut_LC_9_4_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10535_3_lut_LC_9_4_1  (
            .in0(N__41056),
            .in1(N__87395),
            .in2(_gnd_net_),
            .in3(N__41029),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12184 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2273_2274_LC_9_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2273_2274_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2273_2274_LC_9_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2273_2274_LC_9_4_2  (
            .in0(N__56475),
            .in1(N__41244),
            .in2(_gnd_net_),
            .in3(N__75050),
            .lcout(REG_mem_23_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i326_327_LC_9_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i326_327_LC_9_4_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i326_327_LC_9_4_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i326_327_LC_9_4_3  (
            .in0(N__95290),
            .in1(N__71526),
            .in2(N__40992),
            .in3(N__83311),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4742_4743_LC_9_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4742_4743_LC_9_4_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4742_4743_LC_9_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4742_4743_LC_9_4_4  (
            .in0(N__71525),
            .in1(N__40968),
            .in2(_gnd_net_),
            .in3(N__63006),
            .lcout(REG_mem_49_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5510_5511_LC_9_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5510_5511_LC_9_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5510_5511_LC_9_4_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5510_5511_LC_9_4_5  (
            .in0(N__97059),
            .in1(N__41274),
            .in2(N__95616),
            .in3(N__71527),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10734_3_lut_LC_9_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10734_3_lut_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10734_3_lut_LC_9_4_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10734_3_lut_LC_9_4_6  (
            .in0(N__87396),
            .in1(N__41263),
            .in2(_gnd_net_),
            .in3(N__41245),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12383 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5321_5322_LC_9_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5321_5322_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5321_5322_LC_9_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5321_5322_LC_9_4_7  (
            .in0(N__41229),
            .in1(N__96782),
            .in2(_gnd_net_),
            .in3(N__77209),
            .lcout(REG_mem_55_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93338),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11271_LC_9_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11271_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11271_LC_9_5_0 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11271_LC_9_5_0  (
            .in0(N__41338),
            .in1(N__87393),
            .in2(N__41863),
            .in3(N__92373),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12938 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11410_LC_9_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11410_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11410_LC_9_5_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11410_LC_9_5_1  (
            .in0(N__87394),
            .in1(N__41169),
            .in2(N__92586),
            .in3(N__41181),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13112_bdd_4_lut_LC_9_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13112_bdd_4_lut_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13112_bdd_4_lut_LC_9_5_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13112_bdd_4_lut_LC_9_5_2  (
            .in0(N__42088),
            .in1(N__92372),
            .in2(N__41212),
            .in3(N__59335),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i38_39_LC_9_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i38_39_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i38_39_LC_9_5_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i38_39_LC_9_5_3  (
            .in0(N__71521),
            .in1(N__95289),
            .in2(N__41199),
            .in3(N__82904),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3302_3303_LC_9_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3302_3303_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3302_3303_LC_9_5_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3302_3303_LC_9_5_4  (
            .in0(N__95286),
            .in1(N__71522),
            .in2(N__41182),
            .in3(N__80603),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3398_3399_LC_9_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3398_3399_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3398_3399_LC_9_5_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3398_3399_LC_9_5_5  (
            .in0(N__71520),
            .in1(N__95288),
            .in2(N__41170),
            .in3(N__83313),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2291_2292_LC_9_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2291_2292_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2291_2292_LC_9_5_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2291_2292_LC_9_5_6  (
            .in0(N__62332),
            .in1(N__41394),
            .in2(_gnd_net_),
            .in3(N__75020),
            .lcout(REG_mem_23_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i329_330_LC_9_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i329_330_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i329_330_LC_9_5_7 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i329_330_LC_9_5_7  (
            .in0(N__96811),
            .in1(N__95287),
            .in2(N__51441),
            .in3(N__83312),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93325),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10335_3_lut_LC_9_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10335_3_lut_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10335_3_lut_LC_9_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10335_3_lut_LC_9_6_0  (
            .in0(N__87392),
            .in1(N__41362),
            .in2(_gnd_net_),
            .in3(N__41383),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11984 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5318_5319_LC_9_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5318_5319_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5318_5319_LC_9_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5318_5319_LC_9_6_1  (
            .in0(N__41361),
            .in1(N__71519),
            .in2(_gnd_net_),
            .in3(N__77202),
            .lcout(REG_mem_55_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3974_3975_LC_9_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3974_3975_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3974_3975_LC_9_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3974_3975_LC_9_6_2  (
            .in0(N__71517),
            .in1(N__41349),
            .in2(_gnd_net_),
            .in3(N__66008),
            .lcout(REG_mem_41_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4070_4071_LC_9_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4070_4071_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4070_4071_LC_9_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4070_4071_LC_9_6_3  (
            .in0(N__41337),
            .in1(N__71518),
            .in2(_gnd_net_),
            .in3(N__68071),
            .lcout(REG_mem_42_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i944_945_LC_9_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i944_945_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i944_945_LC_9_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i944_945_LC_9_6_4  (
            .in0(N__41322),
            .in1(N__41771),
            .in2(_gnd_net_),
            .in3(N__67154),
            .lcout(REG_mem_9_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2939_2940_LC_9_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2939_2940_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2939_2940_LC_9_6_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2939_2940_LC_9_6_5  (
            .in0(N__95284),
            .in1(N__63439),
            .in2(N__41310),
            .in3(N__77783),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2747_2748_LC_9_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2747_2748_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2747_2748_LC_9_6_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2747_2748_LC_9_6_6  (
            .in0(N__63438),
            .in1(N__95285),
            .in2(N__41292),
            .in3(N__70661),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2099_2100_LC_9_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2099_2100_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2099_2100_LC_9_6_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2099_2100_LC_9_6_7  (
            .in0(N__95283),
            .in1(N__62415),
            .in2(N__41940),
            .in3(N__76916),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93312),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10707_3_lut_LC_9_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10707_3_lut_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10707_3_lut_LC_9_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10707_3_lut_LC_9_7_0  (
            .in0(N__41872),
            .in1(N__41923),
            .in2(_gnd_net_),
            .in3(N__87355),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1574_1575_LC_9_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1574_1575_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1574_1575_LC_9_7_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1574_1575_LC_9_7_1  (
            .in0(N__41883),
            .in1(_gnd_net_),
            .in2(N__71586),
            .in3(N__65618),
            .lcout(REG_mem_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3824_3825_LC_9_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3824_3825_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3824_3825_LC_9_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3824_3825_LC_9_7_2  (
            .in0(N__41871),
            .in1(N__41772),
            .in2(_gnd_net_),
            .in3(N__61829),
            .lcout(REG_mem_39_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4166_4167_LC_9_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4166_4167_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4166_4167_LC_9_7_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4166_4167_LC_9_7_3  (
            .in0(N__41856),
            .in1(_gnd_net_),
            .in2(N__71587),
            .in3(N__68245),
            .lcout(REG_mem_43_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4208_4209_LC_9_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4208_4209_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4208_4209_LC_9_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4208_4209_LC_9_7_4  (
            .in0(N__68246),
            .in1(N__41838),
            .in2(_gnd_net_),
            .in3(N__41774),
            .lcout(REG_mem_43_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i848_849_LC_9_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i848_849_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i848_849_LC_9_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i848_849_LC_9_7_5  (
            .in0(N__67235),
            .in1(N__41814),
            .in2(_gnd_net_),
            .in3(N__41775),
            .lcout(REG_mem_8_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4112_4113_LC_9_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4112_4113_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4112_4113_LC_9_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4112_4113_LC_9_7_6  (
            .in0(N__41436),
            .in1(N__41773),
            .in2(_gnd_net_),
            .in3(N__68038),
            .lcout(REG_mem_42_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i719_720_LC_9_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i719_720_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i719_720_LC_9_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i719_720_LC_9_7_7  (
            .in0(N__41412),
            .in1(N__61246),
            .in2(_gnd_net_),
            .in3(N__89609),
            .lcout(REG_mem_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93298),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i13_2_lut_3_lut_4_lut_LC_9_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i13_2_lut_3_lut_4_lut_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i13_2_lut_3_lut_4_lut_LC_9_8_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i13_2_lut_3_lut_4_lut_LC_9_8_0  (
            .in0(N__50161),
            .in1(N__49034),
            .in2(N__50053),
            .in3(N__49120),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6433_2_lut_3_lut_4_lut_LC_9_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6433_2_lut_3_lut_4_lut_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6433_2_lut_3_lut_4_lut_LC_9_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6433_2_lut_3_lut_4_lut_LC_9_8_1  (
            .in0(N__49121),
            .in1(N__50029),
            .in2(N__49036),
            .in3(N__50162),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i1_3_lut_LC_9_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i1_3_lut_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i1_3_lut_LC_9_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i1_3_lut_LC_9_8_2  (
            .in0(N__48949),
            .in1(N__49035),
            .in2(_gnd_net_),
            .in3(N__49123),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_nxt_c_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i0_LC_9_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i0_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i0_LC_9_8_3 .LUT_INIT=16'b0001111010110100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i0_LC_9_8_3  (
            .in0(N__49124),
            .in1(N__50091),
            .in2(N__41995),
            .in3(N__50163),
            .lcout(wr_grey_sync_r_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93286),
            .ce(),
            .sr(N__73483));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i1_LC_9_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i1_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i1_LC_9_8_4 .LUT_INIT=16'b0110011000111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i1_LC_9_8_4  (
            .in0(N__50164),
            .in1(N__49068),
            .in2(N__50095),
            .in3(N__49125),
            .lcout(wr_grey_sync_r_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93286),
            .ce(),
            .sr(N__73483));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i3_3_lut_LC_9_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i3_3_lut_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i3_3_lut_LC_9_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i3_3_lut_LC_9_8_5  (
            .in0(N__49122),
            .in1(N__49912),
            .in2(_gnd_net_),
            .in3(N__50033),
            .lcout(wr_addr_nxt_c_2),
            .ltout(wr_addr_nxt_c_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i2_LC_9_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i2_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i2_LC_9_8_6 .LUT_INIT=16'b0101101000111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i2_LC_9_8_6  (
            .in0(N__49883),
            .in1(N__49632),
            .in2(N__41992),
            .in3(N__49126),
            .lcout(wr_grey_sync_r_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93286),
            .ce(),
            .sr(N__73483));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i3_LC_9_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i3_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i3_LC_9_8_7 .LUT_INIT=16'b0010011111011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i3_LC_9_8_7  (
            .in0(N__49127),
            .in1(N__49884),
            .in2(N__49636),
            .in3(N__49054),
            .lcout(wr_grey_sync_r_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93286),
            .ce(),
            .sr(N__73483));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5798_5799_LC_9_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5798_5799_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5798_5799_LC_9_9_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5798_5799_LC_9_9_0  (
            .in0(N__94593),
            .in1(N__41979),
            .in2(N__70633),
            .in3(N__71543),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i61_2_lut_3_lut_LC_9_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i61_2_lut_3_lut_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i61_2_lut_3_lut_LC_9_9_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i61_2_lut_3_lut_LC_9_9_1  (
            .in0(N__49544),
            .in1(N__41963),
            .in2(_gnd_net_),
            .in3(N__49805),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n61_adj_1154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6437_2_lut_3_lut_LC_9_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6437_2_lut_3_lut_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6437_2_lut_3_lut_LC_9_9_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6437_2_lut_3_lut_LC_9_9_2  (
            .in0(N__49806),
            .in1(N__42115),
            .in2(_gnd_net_),
            .in3(N__49543),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616 ),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7616_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3110_3111_LC_9_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3110_3111_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3110_3111_LC_9_9_3 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3110_3111_LC_9_9_3  (
            .in0(N__71541),
            .in1(N__42084),
            .in2(N__42091),
            .in3(N__94594),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2726_2727_LC_9_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2726_2727_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2726_2727_LC_9_9_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2726_2727_LC_9_9_4  (
            .in0(N__94592),
            .in1(N__71542),
            .in2(N__42069),
            .in3(N__70565),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3818_3819_LC_9_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3818_3819_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3818_3819_LC_9_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3818_3819_LC_9_9_5  (
            .in0(N__42045),
            .in1(N__46380),
            .in2(_gnd_net_),
            .in3(N__61880),
            .lcout(REG_mem_39_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i59_2_lut_3_lut_4_lut_LC_9_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i59_2_lut_3_lut_4_lut_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i59_2_lut_3_lut_4_lut_LC_9_9_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i59_2_lut_3_lut_4_lut_LC_9_9_6  (
            .in0(N__49804),
            .in1(N__49542),
            .in2(N__43591),
            .in3(N__50024),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4019_4020_LC_9_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4019_4020_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4019_4020_LC_9_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4019_4020_LC_9_9_7  (
            .in0(N__42027),
            .in1(N__62331),
            .in2(_gnd_net_),
            .in3(N__65979),
            .lcout(REG_mem_41_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93275),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i115_2_lut_3_lut_LC_9_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i115_2_lut_3_lut_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i115_2_lut_3_lut_LC_9_10_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i115_2_lut_3_lut_LC_9_10_0  (
            .in0(N__49512),
            .in1(N__94669),
            .in2(_gnd_net_),
            .in3(N__43609),
            .lcout(n10),
            .ltout(n10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5327_5328_LC_9_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5327_5328_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5327_5328_LC_9_10_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5327_5328_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__42006),
            .in2(N__42016),
            .in3(N__61220),
            .lcout(REG_mem_55_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93259),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i65_2_lut_3_lut_4_lut_LC_9_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i65_2_lut_3_lut_4_lut_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i65_2_lut_3_lut_4_lut_LC_9_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i65_2_lut_3_lut_4_lut_LC_9_10_2  (
            .in0(N__49510),
            .in1(N__49831),
            .in2(N__50055),
            .in3(N__43650),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1127_1128_LC_9_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1127_1128_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1127_1128_LC_9_10_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1127_1128_LC_9_10_3  (
            .in0(N__42510),
            .in1(N__47315),
            .in2(_gnd_net_),
            .in3(N__66717),
            .lcout(REG_mem_11_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93259),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3500_3501_LC_9_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3500_3501_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3500_3501_LC_9_10_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3500_3501_LC_9_10_4  (
            .in0(N__61512),
            .in1(_gnd_net_),
            .in2(N__75999),
            .in3(N__54029),
            .lcout(REG_mem_36_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93259),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i71_72_LC_9_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i71_72_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i71_72_LC_9_10_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i71_72_LC_9_10_5  (
            .in0(N__94670),
            .in1(N__47317),
            .in2(N__42189),
            .in3(N__82756),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93259),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i116_2_lut_3_lut_LC_9_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i116_2_lut_3_lut_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i116_2_lut_3_lut_LC_9_10_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i116_2_lut_3_lut_LC_9_10_6  (
            .in0(N__49511),
            .in1(N__94668),
            .in2(_gnd_net_),
            .in3(N__43610),
            .lcout(n42),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4007_4008_LC_9_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4007_4008_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4007_4008_LC_9_10_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4007_4008_LC_9_10_7  (
            .in0(N__42165),
            .in1(N__47316),
            .in2(_gnd_net_),
            .in3(N__65993),
            .lcout(REG_mem_41_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93259),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1709_1710_LC_9_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1709_1710_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1709_1710_LC_9_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1709_1710_LC_9_11_0  (
            .in0(N__46973),
            .in1(N__42153),
            .in2(_gnd_net_),
            .in3(N__66566),
            .lcout(REG_mem_17_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12233_LC_9_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12233_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12233_LC_9_11_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12233_LC_9_11_1  (
            .in0(N__42265),
            .in1(N__91948),
            .in2(N__42256),
            .in3(N__87914),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14102_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14102_bdd_4_lut_LC_9_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14102_bdd_4_lut_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14102_bdd_4_lut_LC_9_11_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14102_bdd_4_lut_LC_9_11_2  (
            .in0(N__91947),
            .in1(N__42154),
            .in2(N__42145),
            .in3(N__42124),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1613_1614_LC_9_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1613_1614_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1613_1614_LC_9_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1613_1614_LC_9_11_3  (
            .in0(N__42123),
            .in1(N__46975),
            .in2(_gnd_net_),
            .in3(N__65669),
            .lcout(REG_mem_16_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1805_1806_LC_9_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1805_1806_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1805_1806_LC_9_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1805_1806_LC_9_11_4  (
            .in0(N__46974),
            .in1(N__42264),
            .in2(_gnd_net_),
            .in3(N__67421),
            .lcout(REG_mem_18_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1901_1902_LC_9_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1901_1902_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1901_1902_LC_9_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1901_1902_LC_9_11_5  (
            .in0(N__42252),
            .in1(N__46976),
            .in2(_gnd_net_),
            .in3(N__72019),
            .lcout(REG_mem_19_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i455_456_LC_9_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i455_456_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i455_456_LC_9_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i455_456_LC_9_11_6  (
            .in0(N__42234),
            .in1(N__47342),
            .in2(_gnd_net_),
            .in3(N__72702),
            .lcout(REG_mem_4_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3719_3720_LC_9_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3719_3720_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3719_3720_LC_9_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3719_3720_LC_9_11_7  (
            .in0(N__47341),
            .in1(N__44451),
            .in2(_gnd_net_),
            .in3(N__59274),
            .lcout(REG_mem_38_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93276),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9832_3_lut_LC_9_12_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9832_3_lut_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9832_3_lut_LC_9_12_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9832_3_lut_LC_9_12_0  (
            .in0(N__42376),
            .in1(N__42220),
            .in2(_gnd_net_),
            .in3(N__44188),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11481_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.full_ext_r_117_LC_9_12_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.full_ext_r_117_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.full_ext_r_117_LC_9_12_1 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.full_ext_r_117_LC_9_12_1  (
            .in0(N__43673),
            .in1(N__42214),
            .in2(N__42223),
            .in3(N__49117),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.full_o ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93287),
            .ce(),
            .sr(N__73477));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9772_4_lut_LC_9_12_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9772_4_lut_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9772_4_lut_LC_9_12_2 .LUT_INIT=16'b1111100110011111;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9772_4_lut_LC_9_12_2  (
            .in0(N__43843),
            .in1(N__49028),
            .in2(N__50056),
            .in3(N__44052),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i11017_4_lut_LC_9_12_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i11017_4_lut_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i11017_4_lut_LC_9_12_3 .LUT_INIT=16'b0001001000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i11017_4_lut_LC_9_12_3  (
            .in0(N__44053),
            .in1(N__44233),
            .in2(N__49911),
            .in3(N__42205),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12527 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_6__I_0_2_lut_LC_9_12_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_6__I_0_2_lut_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_6__I_0_2_lut_LC_9_12_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_6__I_0_2_lut_LC_9_12_4  (
            .in0(N__49238),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52867),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.full_max_w_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5_4_lut_LC_9_12_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5_4_lut_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5_4_lut_LC_9_12_5 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5_4_lut_LC_9_12_5  (
            .in0(N__43729),
            .in1(N__48945),
            .in2(N__42208),
            .in3(N__43842),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6417_2_lut_LC_9_12_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6417_2_lut_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6417_2_lut_LC_9_12_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6417_2_lut_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__43672),
            .in2(_gnd_net_),
            .in3(N__43927),
            .lcout(n7596),
            .ltout(n7596_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i7_3_lut_LC_9_12_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i7_3_lut_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i7_3_lut_LC_9_12_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i7_3_lut_LC_9_12_7  (
            .in0(N__52435),
            .in1(_gnd_net_),
            .in2(N__42367),
            .in3(N__49239),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_w_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10182_3_lut_LC_9_13_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10182_3_lut_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10182_3_lut_LC_9_13_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10182_3_lut_LC_9_13_0  (
            .in0(N__43528),
            .in1(_gnd_net_),
            .in2(N__87354),
            .in3(N__45523),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11831 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2093_2094_LC_9_13_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2093_2094_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2093_2094_LC_9_13_1 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2093_2094_LC_9_13_1  (
            .in0(N__94328),
            .in1(N__47026),
            .in2(N__42345),
            .in3(N__76986),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93299),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3533_3534_LC_9_13_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3533_3534_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3533_3534_LC_9_13_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3533_3534_LC_9_13_2  (
            .in0(N__45975),
            .in1(_gnd_net_),
            .in2(N__47039),
            .in3(N__54093),
            .lcout(REG_mem_36_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93299),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i839_840_LC_9_13_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i839_840_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i839_840_LC_9_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i839_840_LC_9_13_3  (
            .in0(N__47458),
            .in1(N__42531),
            .in2(_gnd_net_),
            .in3(N__67326),
            .lcout(REG_mem_8_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93299),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4109_4110_LC_9_13_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4109_4110_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4109_4110_LC_9_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4109_4110_LC_9_13_4  (
            .in0(N__47030),
            .in1(N__42315),
            .in2(_gnd_net_),
            .in3(N__68000),
            .lcout(REG_mem_42_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93299),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3914_3915_LC_9_13_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3914_3915_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3914_3915_LC_9_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3914_3915_LC_9_13_5  (
            .in0(N__46349),
            .in1(N__42297),
            .in2(_gnd_net_),
            .in3(N__65892),
            .lcout(REG_mem_40_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93299),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1703_1704_LC_9_13_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1703_1704_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1703_1704_LC_9_13_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1703_1704_LC_9_13_6  (
            .in0(N__42276),
            .in1(N__47459),
            .in2(_gnd_net_),
            .in3(N__66586),
            .lcout(REG_mem_17_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93299),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4559_4560_LC_9_13_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4559_4560_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4559_4560_LC_9_13_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4559_4560_LC_9_13_7  (
            .in0(N__61291),
            .in1(N__42477),
            .in2(_gnd_net_),
            .in3(N__66251),
            .lcout(REG_mem_47_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93299),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1898_1899_LC_9_14_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1898_1899_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1898_1899_LC_9_14_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1898_1899_LC_9_14_0  (
            .in0(N__42465),
            .in1(N__46469),
            .in2(_gnd_net_),
            .in3(N__72075),
            .lcout(REG_mem_19_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4679_4680_LC_9_14_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4679_4680_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4679_4680_LC_9_14_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4679_4680_LC_9_14_1  (
            .in0(N__45840),
            .in1(_gnd_net_),
            .in2(N__47387),
            .in3(N__75568),
            .lcout(REG_mem_48_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4010_4011_LC_9_14_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4010_4011_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4010_4011_LC_9_14_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4010_4011_LC_9_14_2  (
            .in0(N__42438),
            .in1(N__46470),
            .in2(_gnd_net_),
            .in3(N__66017),
            .lcout(REG_mem_41_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1133_1134_LC_9_14_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1133_1134_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1133_1134_LC_9_14_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1133_1134_LC_9_14_3  (
            .in0(N__42420),
            .in1(_gnd_net_),
            .in2(N__47038),
            .in3(N__66812),
            .lcout(REG_mem_11_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i941_942_LC_9_14_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i941_942_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i941_942_LC_9_14_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i941_942_LC_9_14_4  (
            .in0(N__67196),
            .in1(N__42405),
            .in2(_gnd_net_),
            .in3(N__47020),
            .lcout(REG_mem_9_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4970_4971_LC_9_14_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4970_4971_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4970_4971_LC_9_14_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4970_4971_LC_9_14_5  (
            .in0(N__46468),
            .in1(N__42387),
            .in2(_gnd_net_),
            .in3(N__72247),
            .lcout(REG_mem_51_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9752_4_lut_4_lut_LC_9_14_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9752_4_lut_4_lut_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9752_4_lut_4_lut_LC_9_14_6 .LUT_INIT=16'b1111011010011111;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9752_4_lut_4_lut_LC_9_14_6  (
            .in0(N__44275),
            .in1(N__49782),
            .in2(N__49591),
            .in3(N__45946),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i935_936_LC_9_14_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i935_936_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i935_936_LC_9_14_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i935_936_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__42546),
            .in2(N__47388),
            .in3(N__67195),
            .lcout(REG_mem_9_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93313),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2279_2280_LC_9_15_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2279_2280_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2279_2280_LC_9_15_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2279_2280_LC_9_15_0  (
            .in0(N__42603),
            .in1(N__47437),
            .in2(_gnd_net_),
            .in3(N__75019),
            .lcout(REG_mem_23_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i1_LC_9_15_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i1_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i1_LC_9_15_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i1_LC_9_15_1  (
            .in0(N__73379),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42727),
            .lcout(rp_sync1_r_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i1_LC_9_15_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i1_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i1_LC_9_15_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i1_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__73381),
            .in2(_gnd_net_),
            .in3(N__42592),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i359_360_LC_9_15_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i359_360_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i359_360_LC_9_15_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i359_360_LC_9_15_3  (
            .in0(N__47436),
            .in1(N__94329),
            .in2(N__42582),
            .in3(N__83341),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_55_LC_9_15_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_55_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_55_LC_9_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_55_LC_9_15_4  (
            .in0(N__42558),
            .in1(N__42565),
            .in2(_gnd_net_),
            .in3(N__44044),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i0_LC_9_15_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i0_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i0_LC_9_15_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i0_LC_9_15_5  (
            .in0(N__73380),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42823),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93326),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_45_LC_9_15_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_45_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_45_LC_9_15_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_45_LC_9_15_6  (
            .in0(N__42559),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44045),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14402_bdd_4_lut_LC_9_15_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14402_bdd_4_lut_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14402_bdd_4_lut_LC_9_15_7 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14402_bdd_4_lut_LC_9_15_7  (
            .in0(N__42499),
            .in1(N__90705),
            .in2(N__42550),
            .in3(N__42535),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_LC_9_16_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_LC_9_16_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_LC_9_16_0  (
            .in0(N__91363),
            .in1(N__42490),
            .in2(N__42520),
            .in3(N__87063),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1031_1032_LC_9_16_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1031_1032_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1031_1032_LC_9_16_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1031_1032_LC_9_16_1  (
            .in0(N__42489),
            .in1(N__47416),
            .in2(_gnd_net_),
            .in3(N__66961),
            .lcout(REG_mem_10_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93339),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2189_2190_LC_9_16_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2189_2190_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2189_2190_LC_9_16_2 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2189_2190_LC_9_16_2  (
            .in0(N__47023),
            .in1(N__94766),
            .in2(N__42690),
            .in3(N__76332),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93339),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2855_2856_LC_9_16_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2855_2856_LC_9_16_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2855_2856_LC_9_16_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2855_2856_LC_9_16_3  (
            .in0(N__94763),
            .in1(N__47417),
            .in2(N__42637),
            .in3(N__70975),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93339),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14240_bdd_4_lut_LC_9_16_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14240_bdd_4_lut_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14240_bdd_4_lut_LC_9_16_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14240_bdd_4_lut_LC_9_16_4  (
            .in0(N__91362),
            .in1(N__44815),
            .in2(N__42775),
            .in3(N__42660),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12042 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i77_78_LC_9_16_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i77_78_LC_9_16_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i77_78_LC_9_16_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i77_78_LC_9_16_5  (
            .in0(N__94765),
            .in1(N__47025),
            .in2(N__42661),
            .in3(N__82927),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93339),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i365_366_LC_9_16_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i365_366_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i365_366_LC_9_16_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i365_366_LC_9_16_6  (
            .in0(N__47024),
            .in1(N__94767),
            .in2(N__42792),
            .in3(N__83339),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93339),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5927_5928_LC_9_16_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5927_5928_LC_9_16_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5927_5928_LC_9_16_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5927_5928_LC_9_16_7  (
            .in0(N__94764),
            .in1(N__47418),
            .in2(N__47589),
            .in3(N__70976),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93339),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3047_3048_LC_9_17_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3047_3048_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3047_3048_LC_9_17_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3047_3048_LC_9_17_0  (
            .in0(N__42648),
            .in1(N__47384),
            .in2(_gnd_net_),
            .in3(N__72550),
            .lcout(REG_mem_31_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93353),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12108_LC_9_17_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12108_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12108_LC_9_17_1 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12108_LC_9_17_1  (
            .in0(N__91353),
            .in1(N__86983),
            .in2(N__42754),
            .in3(N__42649),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13940_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13940_bdd_4_lut_LC_9_17_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13940_bdd_4_lut_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13940_bdd_4_lut_LC_9_17_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13940_bdd_4_lut_LC_9_17_2  (
            .in0(N__42765),
            .in1(N__91352),
            .in2(N__42640),
            .in3(N__42636),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13943 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12348_LC_9_17_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12348_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12348_LC_9_17_3 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12348_LC_9_17_3  (
            .in0(N__91354),
            .in1(N__44878),
            .in2(N__42793),
            .in3(N__86984),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2759_2760_LC_9_17_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2759_2760_LC_9_17_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2759_2760_LC_9_17_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2759_2760_LC_9_17_4  (
            .in0(N__95005),
            .in1(N__47385),
            .in2(N__42766),
            .in3(N__70631),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93353),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2951_2952_LC_9_17_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2951_2952_LC_9_17_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2951_2952_LC_9_17_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2951_2952_LC_9_17_5  (
            .in0(N__47383),
            .in1(N__95007),
            .in2(N__42753),
            .in3(N__77758),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93353),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5831_5832_LC_9_17_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5831_5832_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5831_5832_LC_9_17_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5831_5832_LC_9_17_6  (
            .in0(N__95006),
            .in1(N__47386),
            .in2(N__47616),
            .in3(N__70632),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93353),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i167_168_LC_9_17_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i167_168_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i167_168_LC_9_17_7 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i167_168_LC_9_17_7  (
            .in0(N__47382),
            .in1(N__42738),
            .in2(N__95299),
            .in3(N__80248),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93353),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i5_1_lut_LC_9_18_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i5_1_lut_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i5_1_lut_LC_9_18_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i5_1_lut_LC_9_18_0  (
            .in0(N__81191),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i1_LC_9_18_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i1_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i1_LC_9_18_1 .LUT_INIT=16'b0011011010011100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i1_LC_9_18_1  (
            .in0(N__52558),
            .in1(N__52644),
            .in2(N__84966),
            .in3(N__50750),
            .lcout(rd_grey_sync_r_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97352),
            .ce(),
            .sr(N__73457));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i2_LC_9_18_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i2_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i2_LC_9_18_2 .LUT_INIT=16'b0011100101101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i2_LC_9_18_2  (
            .in0(N__52562),
            .in1(N__42713),
            .in2(N__50755),
            .in3(N__84908),
            .lcout(rd_grey_sync_r_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97352),
            .ce(),
            .sr(N__73457));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i3_LC_9_18_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i3_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i3_LC_9_18_3 .LUT_INIT=16'b0001111010110100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i3_LC_9_18_3  (
            .in0(N__52559),
            .in1(N__81187),
            .in2(N__42718),
            .in3(N__50636),
            .lcout(rd_grey_sync_r_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97352),
            .ce(),
            .sr(N__73457));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i4_LC_9_18_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i4_LC_9_18_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i4_LC_9_18_4 .LUT_INIT=16'b0110011000111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i4_LC_9_18_4  (
            .in0(N__50637),
            .in1(N__42807),
            .in2(N__81233),
            .in3(N__52560),
            .lcout(rd_grey_sync_r_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97352),
            .ce(),
            .sr(N__73457));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i5_LC_9_18_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i5_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i5_LC_9_18_5 .LUT_INIT=16'b0010110101111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i5_LC_9_18_5  (
            .in0(N__52561),
            .in1(N__50791),
            .in2(N__42811),
            .in3(N__44386),
            .lcout(rd_grey_sync_r_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97352),
            .ce(),
            .sr(N__73457));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_i2_3_lut_LC_9_18_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_i2_3_lut_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_i2_3_lut_LC_9_18_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_6__I_0_i2_3_lut_LC_9_18_6  (
            .in0(N__50814),
            .in1(N__52556),
            .in2(_gnd_net_),
            .in3(N__91356),
            .lcout(rd_addr_nxt_c_6_N_465_1),
            .ltout(rd_addr_nxt_c_6_N_465_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i0_LC_9_18_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i0_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i0_LC_9_18_7 .LUT_INIT=16'b0001111010110100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_grey_sync_r__i0_LC_9_18_7  (
            .in0(N__52557),
            .in1(N__86866),
            .in2(N__42796),
            .in3(N__51129),
            .lcout(rd_grey_sync_r_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97352),
            .ce(),
            .sr(N__73457));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i0_LC_9_19_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i0_LC_9_19_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i0_LC_9_19_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i0_LC_9_19_0  (
            .in0(N__73459),
            .in1(N__86859),
            .in2(N__52578),
            .in3(N__51122),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i6_LC_9_19_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i6_LC_9_19_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i6_LC_9_19_1 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i6_LC_9_19_1  (
            .in0(N__50780),
            .in1(N__73462),
            .in2(N__44391),
            .in3(N__52572),
            .lcout(rd_addr_r_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i7_1_lut_LC_9_19_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i7_1_lut_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i7_1_lut_LC_9_19_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i7_1_lut_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__44385),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n2_adj_1149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i1_1_lut_LC_9_19_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i1_1_lut_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i1_1_lut_LC_9_19_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i1_1_lut_LC_9_19_3  (
            .in0(N__86860),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n8_adj_1152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i4_LC_9_19_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i4_LC_9_19_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i4_LC_9_19_4 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i4_LC_9_19_4  (
            .in0(N__73461),
            .in1(N__52573),
            .in2(N__81186),
            .in3(N__50624),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i2_LC_9_19_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i2_LC_9_19_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i2_LC_9_19_5 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i2_LC_9_19_5  (
            .in0(N__50741),
            .in1(N__73460),
            .in2(N__84965),
            .in3(N__52571),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12278_LC_9_19_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12278_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12278_LC_9_19_6 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12278_LC_9_19_6  (
            .in0(N__91502),
            .in1(N__86858),
            .in2(N__43774),
            .in3(N__42907),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i5_LC_9_19_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i5_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i5_LC_9_19_7 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i5_LC_9_19_7  (
            .in0(N__80866),
            .in1(N__73458),
            .in2(N__58354),
            .in3(N__65373),
            .lcout(fifo_data_out_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5735_5736_LC_9_20_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5735_5736_LC_9_20_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5735_5736_LC_9_20_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5735_5736_LC_9_20_0  (
            .in0(N__47340),
            .in1(N__95417),
            .in2(N__47721),
            .in3(N__79661),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93394),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12068_LC_9_20_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12068_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12068_LC_9_20_1 .LUT_INIT=16'b1010110011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12068_LC_9_20_1  (
            .in0(N__42843),
            .in1(N__44575),
            .in2(N__86982),
            .in3(N__91764),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13904_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13904_bdd_4_lut_LC_9_20_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13904_bdd_4_lut_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13904_bdd_4_lut_LC_9_20_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13904_bdd_4_lut_LC_9_20_2  (
            .in0(N__91763),
            .in1(N__42892),
            .in2(N__42871),
            .in3(N__42855),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12174 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3149_3150_LC_9_20_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3149_3150_LC_9_20_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3149_3150_LC_9_20_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3149_3150_LC_9_20_3  (
            .in0(N__95414),
            .in1(N__47009),
            .in2(N__42856),
            .in3(N__82949),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93394),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5159_5160_LC_9_20_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5159_5160_LC_9_20_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5159_5160_LC_9_20_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5159_5160_LC_9_20_4  (
            .in0(N__47339),
            .in1(N__95416),
            .in2(N__44832),
            .in3(N__77046),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93394),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3437_3438_LC_9_20_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3437_3438_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3437_3438_LC_9_20_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3437_3438_LC_9_20_5  (
            .in0(N__95415),
            .in1(N__47010),
            .in2(N__42844),
            .in3(N__83340),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93394),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i0_LC_9_20_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i0_LC_9_20_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i0_LC_9_20_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i0_LC_9_20_7  (
            .in0(N__42832),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73463),
            .lcout(rp_sync1_r_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93394),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i230_231_LC_10_1_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i230_231_LC_10_1_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i230_231_LC_10_1_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i230_231_LC_10_1_0  (
            .in0(N__71470),
            .in1(N__95553),
            .in2(N__43038),
            .in3(N__80527),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3347_3348_LC_10_1_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3347_3348_LC_10_1_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3347_3348_LC_10_1_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3347_3348_LC_10_1_1  (
            .in0(N__80526),
            .in1(N__42951),
            .in2(N__95706),
            .in3(N__62422),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3443_3444_LC_10_1_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3443_3444_LC_10_1_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3443_3444_LC_10_1_2 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3443_3444_LC_10_1_2  (
            .in0(N__62420),
            .in1(N__42960),
            .in2(N__83383),
            .in3(N__95555),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1871_1872_LC_10_1_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1871_1872_LC_10_1_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1871_1872_LC_10_1_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1871_1872_LC_10_1_3  (
            .in0(N__43011),
            .in1(N__61248),
            .in2(_gnd_net_),
            .in3(N__72109),
            .lcout(REG_mem_19_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i371_372_LC_10_1_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i371_372_LC_10_1_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i371_372_LC_10_1_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i371_372_LC_10_1_4  (
            .in0(N__62421),
            .in1(N__95554),
            .in2(N__44991),
            .in3(N__83357),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i257_258_LC_10_1_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i257_258_LC_10_1_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i257_258_LC_10_1_5 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i257_258_LC_10_1_5  (
            .in0(N__80525),
            .in1(N__42996),
            .in2(N__95705),
            .in3(N__56619),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93396),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10692_3_lut_LC_10_1_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10692_3_lut_LC_10_1_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10692_3_lut_LC_10_1_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10692_3_lut_LC_10_1_6  (
            .in0(N__88814),
            .in1(_gnd_net_),
            .in2(N__43000),
            .in3(N__42988),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10338_3_lut_LC_10_1_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10338_3_lut_LC_10_1_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10338_3_lut_LC_10_1_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10338_3_lut_LC_10_1_7  (
            .in0(N__42961),
            .in1(N__88813),
            .in2(_gnd_net_),
            .in3(N__42952),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11987 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11964_LC_10_2_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11964_LC_10_2_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11964_LC_10_2_0 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11964_LC_10_2_0  (
            .in0(N__85630),
            .in1(N__92583),
            .in2(N__42934),
            .in3(N__42919),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13682_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13682_bdd_4_lut_LC_10_2_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13682_bdd_4_lut_LC_10_2_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13682_bdd_4_lut_LC_10_2_1 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13682_bdd_4_lut_LC_10_2_1  (
            .in0(N__43117),
            .in1(N__85628),
            .in2(N__43108),
            .in3(N__43075),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13685 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1889_1890_LC_10_2_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1889_1890_LC_10_2_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1889_1890_LC_10_2_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1889_1890_LC_10_2_2  (
            .in0(N__43236),
            .in1(N__56408),
            .in2(_gnd_net_),
            .in3(N__72093),
            .lcout(REG_mem_19_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93382),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14132_bdd_4_lut_LC_10_2_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14132_bdd_4_lut_LC_10_2_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14132_bdd_4_lut_LC_10_2_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14132_bdd_4_lut_LC_10_2_3  (
            .in0(N__71080),
            .in1(N__85629),
            .in2(N__43105),
            .in3(N__43087),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12098 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4085_4086_LC_10_2_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4085_4086_LC_10_2_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4085_4086_LC_10_2_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4085_4086_LC_10_2_4  (
            .in0(N__44955),
            .in1(N__62612),
            .in2(_gnd_net_),
            .in3(N__68077),
            .lcout(REG_mem_42_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93382),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10323_3_lut_LC_10_2_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10323_3_lut_LC_10_2_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10323_3_lut_LC_10_2_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10323_3_lut_LC_10_2_5  (
            .in0(N__43069),
            .in1(N__88698),
            .in2(_gnd_net_),
            .in3(N__44935),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11972 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4934_4935_LC_10_2_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4934_4935_LC_10_2_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4934_4935_LC_10_2_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4934_4935_LC_10_2_7  (
            .in0(N__43068),
            .in1(N__71353),
            .in2(_gnd_net_),
            .in3(N__72228),
            .lcout(REG_mem_51_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93382),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10439_3_lut_LC_10_3_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10439_3_lut_LC_10_3_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10439_3_lut_LC_10_3_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10439_3_lut_LC_10_3_0  (
            .in0(N__43050),
            .in1(N__88670),
            .in2(_gnd_net_),
            .in3(N__43060),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12088 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3125_3126_LC_10_3_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3125_3126_LC_10_3_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3125_3126_LC_10_3_1 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3125_3126_LC_10_3_1  (
            .in0(N__43059),
            .in1(N__62810),
            .in2(N__95721),
            .in3(N__82919),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3221_3222_LC_10_3_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3221_3222_LC_10_3_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3221_3222_LC_10_3_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3221_3222_LC_10_3_2  (
            .in0(N__62809),
            .in1(N__95584),
            .in2(N__43051),
            .in3(N__80166),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i53_54_LC_10_3_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i53_54_LC_10_3_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i53_54_LC_10_3_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i53_54_LC_10_3_3  (
            .in0(N__48132),
            .in1(N__62811),
            .in2(N__95722),
            .in3(N__82920),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i149_150_LC_10_3_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i149_150_LC_10_3_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i149_150_LC_10_3_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i149_150_LC_10_3_4  (
            .in0(N__62808),
            .in1(N__95583),
            .in2(N__48156),
            .in3(N__80165),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i236_237_LC_10_3_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i236_237_LC_10_3_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i236_237_LC_10_3_5 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i236_237_LC_10_3_5  (
            .in0(N__80581),
            .in1(N__75975),
            .in2(N__47865),
            .in3(N__95594),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1862_1863_LC_10_3_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1862_1863_LC_10_3_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1862_1863_LC_10_3_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1862_1863_LC_10_3_6  (
            .in0(N__43185),
            .in1(N__71471),
            .in2(_gnd_net_),
            .in3(N__72092),
            .lcout(REG_mem_19_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3308_3309_LC_10_3_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3308_3309_LC_10_3_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3308_3309_LC_10_3_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3308_3309_LC_10_3_7  (
            .in0(N__80582),
            .in1(N__75976),
            .in2(N__95723),
            .in3(N__48234),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93369),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11515_LC_10_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11515_LC_10_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11515_LC_10_4_0 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11515_LC_10_4_0  (
            .in0(N__88447),
            .in1(N__92431),
            .in2(N__43129),
            .in3(N__43174),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13232 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i233_234_LC_10_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i233_234_LC_10_4_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i233_234_LC_10_4_1 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i233_234_LC_10_4_1  (
            .in0(N__96776),
            .in1(N__95294),
            .in2(N__51465),
            .in3(N__80471),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i806_807_LC_10_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i806_807_LC_10_4_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i806_807_LC_10_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i806_807_LC_10_4_2  (
            .in0(N__71399),
            .in1(N__51582),
            .in2(_gnd_net_),
            .in3(N__67312),
            .lcout(REG_mem_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1766_1767_LC_10_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1766_1767_LC_10_4_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1766_1767_LC_10_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1766_1767_LC_10_4_3  (
            .in0(N__43146),
            .in1(N__71400),
            .in2(_gnd_net_),
            .in3(N__67491),
            .lcout(REG_mem_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1025_1026_LC_10_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1025_1026_LC_10_4_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1025_1026_LC_10_4_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1025_1026_LC_10_4_4  (
            .in0(N__43125),
            .in1(N__56593),
            .in2(_gnd_net_),
            .in3(N__66984),
            .lcout(REG_mem_10_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11445_LC_10_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11445_LC_10_4_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11445_LC_10_4_5 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11445_LC_10_4_5  (
            .in0(N__92432),
            .in1(N__85504),
            .in2(N__48187),
            .in3(N__43342),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12908 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3014_3015_LC_10_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3014_3015_LC_10_4_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3014_3015_LC_10_4_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3014_3015_LC_10_4_6  (
            .in0(N__71398),
            .in1(_gnd_net_),
            .in2(N__43335),
            .in3(N__72539),
            .lcout(REG_mem_31_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1811_1812_LC_10_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1811_1812_LC_10_4_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1811_1812_LC_10_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1811_1812_LC_10_4_7  (
            .in0(N__43305),
            .in1(N__62412),
            .in2(_gnd_net_),
            .in3(N__67492),
            .lcout(REG_mem_18_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93355),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10712_3_lut_LC_10_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10712_3_lut_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10712_3_lut_LC_10_5_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10712_3_lut_LC_10_5_0  (
            .in0(N__43294),
            .in1(N__88444),
            .in2(_gnd_net_),
            .in3(N__43501),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2534_2535_LC_10_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2534_2535_LC_10_5_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2534_2535_LC_10_5_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2534_2535_LC_10_5_1  (
            .in0(N__70295),
            .in1(N__43269),
            .in2(_gnd_net_),
            .in3(N__71462),
            .lcout(REG_mem_26_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93340),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4769_4770_LC_10_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4769_4770_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4769_4770_LC_10_5_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4769_4770_LC_10_5_2  (
            .in0(N__43254),
            .in1(N__56594),
            .in2(_gnd_net_),
            .in3(N__62989),
            .lcout(REG_mem_49_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93340),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1190_1191_LC_10_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1190_1191_LC_10_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1190_1191_LC_10_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1190_1191_LC_10_5_3  (
            .in0(N__45060),
            .in1(N__71461),
            .in2(_gnd_net_),
            .in3(N__59653),
            .lcout(REG_mem_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93340),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10713_3_lut_LC_10_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10713_3_lut_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10713_3_lut_LC_10_5_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10713_3_lut_LC_10_5_4  (
            .in0(N__43243),
            .in1(N__88445),
            .in2(_gnd_net_),
            .in3(N__48436),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12362_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12908_bdd_4_lut_LC_10_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12908_bdd_4_lut_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12908_bdd_4_lut_LC_10_5_5 .LUT_INIT=16'b1010101011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12908_bdd_4_lut_LC_10_5_5  (
            .in0(N__43225),
            .in1(N__43219),
            .in2(N__43213),
            .in3(N__85431),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12911 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i929_930_LC_10_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i929_930_LC_10_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i929_930_LC_10_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i929_930_LC_10_5_6  (
            .in0(N__43476),
            .in1(N__56595),
            .in2(_gnd_net_),
            .in3(N__67155),
            .lcout(REG_mem_9_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93340),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3989_3990_LC_10_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3989_3990_LC_10_5_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3989_3990_LC_10_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3989_3990_LC_10_5_7  (
            .in0(N__47763),
            .in1(N__62817),
            .in2(_gnd_net_),
            .in3(N__66007),
            .lcout(REG_mem_41_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93340),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4193_4194_LC_10_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4193_4194_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4193_4194_LC_10_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4193_4194_LC_10_6_0  (
            .in0(N__43452),
            .in1(N__56592),
            .in2(_gnd_net_),
            .in3(N__68244),
            .lcout(REG_mem_43_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3539_3540_LC_10_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3539_3540_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3539_3540_LC_10_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3539_3540_LC_10_6_1  (
            .in0(N__43395),
            .in1(N__62378),
            .in2(_gnd_net_),
            .in3(N__54073),
            .lcout(REG_mem_36_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4979_4980_LC_10_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4979_4980_LC_10_6_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4979_4980_LC_10_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4979_4980_LC_10_6_2  (
            .in0(N__62376),
            .in1(N__43434),
            .in2(_gnd_net_),
            .in3(N__72203),
            .lcout(REG_mem_51_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i740_741_LC_10_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i740_741_LC_10_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i740_741_LC_10_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i740_741_LC_10_6_3  (
            .in0(N__43407),
            .in1(N__48768),
            .in2(_gnd_net_),
            .in3(N__89612),
            .lcout(REG_mem_7_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10346_3_lut_LC_10_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10346_3_lut_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10346_3_lut_LC_10_6_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10346_3_lut_LC_10_6_4  (
            .in0(N__88443),
            .in1(N__43396),
            .in2(_gnd_net_),
            .in3(N__45373),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11995 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i947_948_LC_10_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i947_948_LC_10_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i947_948_LC_10_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i947_948_LC_10_6_5  (
            .in0(N__43368),
            .in1(N__62379),
            .in2(_gnd_net_),
            .in3(N__67153),
            .lcout(REG_mem_9_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2459_2460_LC_10_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2459_2460_LC_10_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2459_2460_LC_10_6_6 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2459_2460_LC_10_6_6  (
            .in0(N__63338),
            .in1(N__43353),
            .in2(N__95617),
            .in3(N__96941),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1139_1140_LC_10_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1139_1140_LC_10_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1139_1140_LC_10_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1139_1140_LC_10_6_7  (
            .in0(N__43542),
            .in1(N__62377),
            .in2(_gnd_net_),
            .in3(N__66761),
            .lcout(REG_mem_11_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93327),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i83_2_lut_3_lut_LC_10_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i83_2_lut_3_lut_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i83_2_lut_3_lut_LC_10_7_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i83_2_lut_3_lut_LC_10_7_0  (
            .in0(N__94483),
            .in1(N__49592),
            .in2(_gnd_net_),
            .in3(N__43611),
            .lcout(n26),
            .ltout(n26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3791_3792_LC_10_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3791_3792_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3791_3792_LC_10_7_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3791_3792_LC_10_7_1  (
            .in0(_gnd_net_),
            .in1(N__43518),
            .in2(N__43531),
            .in3(N__61247),
            .lcout(REG_mem_39_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3803_3804_LC_10_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3803_3804_LC_10_7_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3803_3804_LC_10_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3803_3804_LC_10_7_2  (
            .in0(N__48255),
            .in1(N__63490),
            .in2(_gnd_net_),
            .in3(N__61828),
            .lcout(REG_mem_39_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i84_2_lut_3_lut_LC_10_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i84_2_lut_3_lut_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i84_2_lut_3_lut_LC_10_7_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i84_2_lut_3_lut_LC_10_7_3  (
            .in0(N__43612),
            .in1(N__94484),
            .in2(_gnd_net_),
            .in3(N__49593),
            .lcout(n58),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i905_906_LC_10_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i905_906_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i905_906_LC_10_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i905_906_LC_10_7_4  (
            .in0(N__51609),
            .in1(N__96817),
            .in2(_gnd_net_),
            .in3(N__67098),
            .lcout(REG_mem_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4748_4749_LC_10_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4748_4749_LC_10_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4748_4749_LC_10_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4748_4749_LC_10_7_5  (
            .in0(N__45120),
            .in1(N__75973),
            .in2(_gnd_net_),
            .in3(N__62962),
            .lcout(REG_mem_49_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1697_1698_LC_10_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1697_1698_LC_10_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1697_1698_LC_10_7_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1697_1698_LC_10_7_6  (
            .in0(N__43494),
            .in1(N__66490),
            .in2(_gnd_net_),
            .in3(N__56625),
            .lcout(REG_mem_17_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5804_5805_LC_10_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5804_5805_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5804_5805_LC_10_7_7 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5804_5805_LC_10_7_7  (
            .in0(N__56139),
            .in1(N__94485),
            .in2(N__70692),
            .in3(N__75974),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93314),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i16_2_lut_LC_10_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i16_2_lut_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i16_2_lut_LC_10_8_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i16_2_lut_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__50042),
            .in2(_gnd_net_),
            .in3(N__43713),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n16 ),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i104_2_lut_3_lut_4_lut_LC_10_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i104_2_lut_3_lut_4_lut_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i104_2_lut_3_lut_4_lut_LC_10_8_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i104_2_lut_3_lut_4_lut_LC_10_8_1  (
            .in0(N__94686),
            .in1(N__49527),
            .in2(N__43567),
            .in3(N__49815),
            .lcout(n48),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i87_2_lut_3_lut_4_lut_LC_10_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i87_2_lut_3_lut_4_lut_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i87_2_lut_3_lut_4_lut_LC_10_8_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i87_2_lut_3_lut_4_lut_LC_10_8_2  (
            .in0(N__43563),
            .in1(N__94681),
            .in2(N__49841),
            .in3(N__49570),
            .lcout(n24_adj_1185),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i88_2_lut_3_lut_4_lut_LC_10_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i88_2_lut_3_lut_4_lut_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i88_2_lut_3_lut_4_lut_LC_10_8_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i88_2_lut_3_lut_4_lut_LC_10_8_3  (
            .in0(N__49569),
            .in1(N__49811),
            .in2(N__95177),
            .in3(N__43564),
            .lcout(n56),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i107_2_lut_3_lut_4_lut_LC_10_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i107_2_lut_3_lut_4_lut_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i107_2_lut_3_lut_4_lut_LC_10_8_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i107_2_lut_3_lut_4_lut_LC_10_8_4  (
            .in0(N__49810),
            .in1(N__43627),
            .in2(N__49580),
            .in3(N__94685),
            .lcout(n14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i103_2_lut_3_lut_4_lut_LC_10_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i103_2_lut_3_lut_4_lut_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i103_2_lut_3_lut_4_lut_LC_10_8_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i103_2_lut_3_lut_4_lut_LC_10_8_5  (
            .in0(N__49568),
            .in1(N__49809),
            .in2(N__95176),
            .in3(N__43562),
            .lcout(n16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i47_2_lut_3_lut_4_lut_LC_10_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i47_2_lut_3_lut_4_lut_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i47_2_lut_3_lut_4_lut_LC_10_8_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i47_2_lut_3_lut_4_lut_LC_10_8_6  (
            .in0(N__49807),
            .in1(N__50043),
            .in2(N__49579),
            .in3(N__43714),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i55_2_lut_3_lut_4_lut_LC_10_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i55_2_lut_3_lut_4_lut_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i55_2_lut_3_lut_4_lut_LC_10_8_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i55_2_lut_3_lut_4_lut_LC_10_8_7  (
            .in0(N__43715),
            .in1(N__49523),
            .in2(N__50054),
            .in3(N__49808),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i108_2_lut_3_lut_4_lut_LC_10_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i108_2_lut_3_lut_4_lut_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i108_2_lut_3_lut_4_lut_LC_10_9_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i108_2_lut_3_lut_4_lut_LC_10_9_0  (
            .in0(N__49796),
            .in1(N__49553),
            .in2(N__95174),
            .in3(N__43625),
            .lcout(n46),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i20_2_lut_LC_10_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i20_2_lut_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i20_2_lut_LC_10_9_1 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i20_2_lut_LC_10_9_1  (
            .in0(N__50036),
            .in1(N__43586),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n20_adj_1160 ),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n20_adj_1160_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i91_2_lut_3_lut_4_lut_LC_10_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i91_2_lut_3_lut_4_lut_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i91_2_lut_3_lut_4_lut_LC_10_9_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i91_2_lut_3_lut_4_lut_LC_10_9_2  (
            .in0(N__94671),
            .in1(N__49816),
            .in2(N__43552),
            .in3(N__49554),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i12_2_lut_3_lut_4_lut_LC_10_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i12_2_lut_3_lut_4_lut_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i12_2_lut_3_lut_4_lut_LC_10_9_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i12_2_lut_3_lut_4_lut_LC_10_9_3  (
            .in0(N__50159),
            .in1(N__49020),
            .in2(N__43693),
            .in3(N__43941),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12_adj_1156 ),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12_adj_1156_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i15_2_lut_LC_10_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i15_2_lut_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i15_2_lut_LC_10_9_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i15_2_lut_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43630),
            .in3(N__50034),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i44_2_lut_3_lut_4_lut_LC_10_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i44_2_lut_3_lut_4_lut_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i44_2_lut_3_lut_4_lut_LC_10_9_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i44_2_lut_3_lut_4_lut_LC_10_9_5  (
            .in0(N__50037),
            .in1(N__43587),
            .in2(N__49589),
            .in3(N__49795),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i92_2_lut_3_lut_4_lut_LC_10_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i92_2_lut_3_lut_4_lut_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i92_2_lut_3_lut_4_lut_LC_10_9_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i92_2_lut_3_lut_4_lut_LC_10_9_6  (
            .in0(N__49797),
            .in1(N__49555),
            .in2(N__95175),
            .in3(N__43626),
            .lcout(n54),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i36_2_lut_3_lut_LC_10_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i36_2_lut_3_lut_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i36_2_lut_3_lut_LC_10_9_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i36_2_lut_3_lut_LC_10_9_7  (
            .in0(N__50035),
            .in1(N__43585),
            .in2(_gnd_net_),
            .in3(N__49794),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i11_2_lut_3_lut_4_lut_LC_10_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i11_2_lut_3_lut_4_lut_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i11_2_lut_3_lut_4_lut_LC_10_10_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i11_2_lut_3_lut_4_lut_LC_10_10_0  (
            .in0(N__43940),
            .in1(N__43685),
            .in2(N__49030),
            .in3(N__50158),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11 ),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i35_2_lut_3_lut_LC_10_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i35_2_lut_3_lut_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i35_2_lut_3_lut_LC_10_10_1 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i35_2_lut_3_lut_LC_10_10_1  (
            .in0(N__50039),
            .in1(N__49799),
            .in2(N__43570),
            .in3(_gnd_net_),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i17_2_lut_LC_10_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i17_2_lut_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i17_2_lut_LC_10_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i17_2_lut_LC_10_10_2  (
            .in0(N__43649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50038),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2270_2271_LC_10_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2270_2271_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2270_2271_LC_10_10_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2270_2271_LC_10_10_3  (
            .in0(N__72366),
            .in1(N__89519),
            .in2(_gnd_net_),
            .in3(N__74961),
            .lcout(REG_mem_23_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93269),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i40_2_lut_3_lut_4_lut_LC_10_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i40_2_lut_3_lut_4_lut_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i40_2_lut_3_lut_4_lut_LC_10_10_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i40_2_lut_3_lut_4_lut_LC_10_10_4  (
            .in0(N__50028),
            .in1(N__49519),
            .in2(N__49840),
            .in3(N__43716),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i9_2_lut_3_lut_4_lut_LC_10_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i9_2_lut_3_lut_4_lut_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i9_2_lut_3_lut_4_lut_LC_10_10_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i9_2_lut_3_lut_4_lut_LC_10_10_5  (
            .in0(N__50157),
            .in1(N__49016),
            .in2(N__43689),
            .in3(N__43939),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n9 ),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i25_2_lut_3_lut_LC_10_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i25_2_lut_3_lut_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i25_2_lut_3_lut_LC_10_10_6 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i25_2_lut_3_lut_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__49798),
            .in2(N__43657),
            .in3(N__50040),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i26_2_lut_3_lut_LC_10_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i26_2_lut_3_lut_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i26_2_lut_3_lut_LC_10_10_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i26_2_lut_3_lut_LC_10_10_7  (
            .in0(N__50041),
            .in1(N__49800),
            .in2(_gnd_net_),
            .in3(N__43648),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n26_adj_1146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.state_timeout_counter_i0_i2_LC_10_11_0 .C_ON=1'b0;
    defparam \usb3_if_inst.state_timeout_counter_i0_i2_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.state_timeout_counter_i0_i2_LC_10_11_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \usb3_if_inst.state_timeout_counter_i0_i2_LC_10_11_0  (
            .in0(N__64143),
            .in1(N__64313),
            .in2(N__57630),
            .in3(N__54541),
            .lcout(\usb3_if_inst.state_timeout_counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_timeout_counter_i0_i2C_net ),
            .ce(N__54493),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i7_4_lut_LC_10_11_1 .C_ON=1'b0;
    defparam \usb3_if_inst.i7_4_lut_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i7_4_lut_LC_10_11_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \usb3_if_inst.i7_4_lut_LC_10_11_1  (
            .in0(N__54577),
            .in1(N__54421),
            .in2(N__54448),
            .in3(N__54601),
            .lcout(\usb3_if_inst.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i106_2_lut_3_lut_LC_10_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i106_2_lut_3_lut_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i106_2_lut_3_lut_LC_10_11_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i106_2_lut_3_lut_LC_10_11_2  (
            .in0(N__45459),
            .in1(N__93968),
            .in2(_gnd_net_),
            .in3(N__49502),
            .lcout(n47),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i42_2_lut_LC_10_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i42_2_lut_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i42_2_lut_LC_10_11_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i42_2_lut_LC_10_11_3  (
            .in0(N__49501),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45458),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i121_2_lut_3_lut_LC_10_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i121_2_lut_3_lut_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i121_2_lut_3_lut_LC_10_11_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i121_2_lut_3_lut_LC_10_11_4  (
            .in0(N__93965),
            .in1(N__49509),
            .in2(_gnd_net_),
            .in3(N__43807),
            .lcout(n7_adj_1183),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i122_2_lut_3_lut_LC_10_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i122_2_lut_3_lut_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i122_2_lut_3_lut_LC_10_11_5 .LUT_INIT=16'b0010000000100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i122_2_lut_3_lut_LC_10_11_5  (
            .in0(N__43808),
            .in1(N__93966),
            .in2(N__49571),
            .in3(_gnd_net_),
            .lcout(n39),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i89_2_lut_3_lut_LC_10_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i89_2_lut_3_lut_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i89_2_lut_3_lut_LC_10_11_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i89_2_lut_3_lut_LC_10_11_6  (
            .in0(N__93964),
            .in1(N__49500),
            .in2(_gnd_net_),
            .in3(N__43809),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i90_2_lut_3_lut_LC_10_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i90_2_lut_3_lut_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i90_2_lut_3_lut_LC_10_11_7 .LUT_INIT=16'b0000001000000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i90_2_lut_3_lut_LC_10_11_7  (
            .in0(N__43810),
            .in1(N__93967),
            .in2(N__49572),
            .in3(_gnd_net_),
            .lcout(n55),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4571_4572_LC_10_12_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4571_4572_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4571_4572_LC_10_12_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4571_4572_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__63505),
            .in2(N__43791),
            .in3(N__66219),
            .lcout(REG_mem_47_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93300),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5351_5352_LC_10_12_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5351_5352_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5351_5352_LC_10_12_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5351_5352_LC_10_12_1  (
            .in0(N__47373),
            .in1(N__43764),
            .in2(_gnd_net_),
            .in3(N__77192),
            .lcout(REG_mem_55_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93300),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i749_750_LC_10_12_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i749_750_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i749_750_LC_10_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i749_750_LC_10_12_2  (
            .in0(N__44421),
            .in1(N__46929),
            .in2(_gnd_net_),
            .in3(N__89650),
            .lcout(REG_mem_7_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93300),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i1_LC_10_12_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i1_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i1_LC_10_12_3 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i1_LC_10_12_3  (
            .in0(N__50142),
            .in1(N__50084),
            .in2(N__73481),
            .in3(N__49118),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93300),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4562_4563_LC_10_12_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4562_4563_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4562_4563_LC_10_12_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4562_4563_LC_10_12_4  (
            .in0(N__57081),
            .in1(N__76751),
            .in2(_gnd_net_),
            .in3(N__66218),
            .lcout(REG_mem_47_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93300),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4577_4578_LC_10_12_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4577_4578_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4577_4578_LC_10_12_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4577_4578_LC_10_12_5  (
            .in0(N__66220),
            .in1(N__43740),
            .in2(_gnd_net_),
            .in3(N__56615),
            .lcout(REG_mem_47_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93300),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i6_LC_10_12_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i6_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i6_LC_10_12_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i6_LC_10_12_6  (
            .in0(N__49119),
            .in1(N__73456),
            .in2(N__52442),
            .in3(N__49240),
            .lcout(wr_grey_sync_r_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93300),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9799_4_lut_LC_10_12_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9799_4_lut_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9799_4_lut_LC_10_12_7 .LUT_INIT=16'b1110101111010111;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9799_4_lut_LC_10_12_7  (
            .in0(N__49296),
            .in1(N__44212),
            .in2(N__50090),
            .in3(N__45942),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.FT_RD_internal_75_LC_10_13_0 .C_ON=1'b0;
    defparam \usb3_if_inst.FT_RD_internal_75_LC_10_13_0 .SEQ_MODE=4'b1001;
    defparam \usb3_if_inst.FT_RD_internal_75_LC_10_13_0 .LUT_INIT=16'b1101110111010001;
    LogicCell40 \usb3_if_inst.FT_RD_internal_75_LC_10_13_0  (
            .in0(N__43869),
            .in1(N__64109),
            .in2(N__57599),
            .in3(N__64292),
            .lcout(DEBUG_3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.FT_RD_internal_75C_net ),
            .ce(),
            .sr(N__73709));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2_2_lut_LC_10_13_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2_2_lut_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2_2_lut_LC_10_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2_2_lut_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__44124),
            .in2(_gnd_net_),
            .in3(N__44112),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n6_adj_1172 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2_3_lut_LC_10_13_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2_3_lut_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2_3_lut_LC_10_13_2 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2_3_lut_LC_10_13_2  (
            .in0(N__44113),
            .in1(_gnd_net_),
            .in2(N__44128),
            .in3(N__43825),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10784_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9815_4_lut_LC_10_13_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9815_4_lut_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9815_4_lut_LC_10_13_3 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9815_4_lut_LC_10_13_3  (
            .in0(N__64293),
            .in1(N__44101),
            .in2(N__44020),
            .in3(N__44080),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11463 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i11082_3_lut_LC_10_13_4 .C_ON=1'b0;
    defparam \usb3_if_inst.i11082_3_lut_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i11082_3_lut_LC_10_13_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \usb3_if_inst.i11082_3_lut_LC_10_13_4  (
            .in0(N__57583),
            .in1(N__43881),
            .in2(_gnd_net_),
            .in3(N__43970),
            .lcout(afull_flag_impl_af_flag_p_w_N_603_3),
            .ltout(afull_flag_impl_af_flag_p_w_N_603_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_4_lut_adj_57_LC_10_13_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_4_lut_adj_57_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_4_lut_adj_57_LC_10_13_5 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_4_lut_adj_57_LC_10_13_5  (
            .in0(N__43824),
            .in1(N__44100),
            .in2(N__43906),
            .in3(N__43903),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n3_adj_1166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.FT_OE_internal_74_LC_10_13_6 .C_ON=1'b0;
    defparam \usb3_if_inst.FT_OE_internal_74_LC_10_13_6 .SEQ_MODE=4'b1001;
    defparam \usb3_if_inst.FT_OE_internal_74_LC_10_13_6 .LUT_INIT=16'b1100110100000001;
    LogicCell40 \usb3_if_inst.FT_OE_internal_74_LC_10_13_6  (
            .in0(N__43868),
            .in1(N__64108),
            .in2(N__57262),
            .in3(N__57517),
            .lcout(FT_OE_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.FT_RD_internal_75C_net ),
            .ce(),
            .sr(N__73709));
    defparam \usb3_if_inst.state_FSM_i6_LC_10_13_7 .C_ON=1'b0;
    defparam \usb3_if_inst.state_FSM_i6_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.state_FSM_i6_LC_10_13_7 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \usb3_if_inst.state_FSM_i6_LC_10_13_7  (
            .in0(N__64291),
            .in1(N__57584),
            .in2(N__64129),
            .in3(N__43870),
            .lcout(\usb3_if_inst.n550 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.FT_RD_internal_75C_net ),
            .ce(),
            .sr(N__73709));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_2_lut_LC_10_14_0 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_2_lut_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_2_lut_LC_10_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_2_lut_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__43836),
            .in2(N__49029),
            .in3(N__43813),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_sig_diff0_w_0 ),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10625 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_3_lut_LC_10_14_1 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_3_lut_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_3_lut_LC_10_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_3_lut_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__44204),
            .in2(N__50160),
            .in3(N__44116),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_sig_diff0_w_1 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10625 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10626 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_4_lut_LC_10_14_2 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_4_lut_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_4_lut_LC_10_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_4_lut_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__44046),
            .in2(N__50025),
            .in3(N__44104),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_sig_diff0_w_2 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10626 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10627 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_5_lut_LC_10_14_3 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_5_lut_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_5_lut_LC_10_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_5_lut_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(N__44026),
            .in2(N__49837),
            .in3(N__44092),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_sig_diff0_w_3 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10627 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10628 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_6_lut_LC_10_14_4 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_6_lut_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_6_lut_LC_10_14_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_6_lut_LC_10_14_4  (
            .in0(N__44089),
            .in1(N__45935),
            .in2(N__49590),
            .in3(N__44074),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11436 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10628 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10629 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_7_lut_LC_10_14_5 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_7_lut_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_7_lut_LC_10_14_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_add_2_7_lut_LC_10_14_5  (
            .in0(N__44071),
            .in1(N__94458),
            .in2(N__46105),
            .in3(N__44065),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11475 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10629 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10630 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.afull_flag_impl_af_flag_ext_r_121_LC_10_14_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.afull_flag_impl_af_flag_ext_r_121_LC_10_14_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.afull_flag_impl_af_flag_ext_r_121_LC_10_14_6 .LUT_INIT=16'b1110110111011110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.afull_flag_impl_af_flag_ext_r_121_LC_10_14_6  (
            .in0(N__52834),
            .in1(N__44062),
            .in2(N__52446),
            .in3(N__44056),
            .lcout(DEBUG_9_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93328),
            .ce(),
            .sr(N__73373));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_56_LC_10_15_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_56_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_56_LC_10_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_56_LC_10_15_0  (
            .in0(N__44273),
            .in1(N__44170),
            .in2(_gnd_net_),
            .in3(N__45933),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_LC_10_15_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_LC_10_15_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_LC_10_15_1  (
            .in0(N__45934),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44274),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_3 ),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9736_4_lut_LC_10_15_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9736_4_lut_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9736_4_lut_LC_10_15_2 .LUT_INIT=16'b1110101111010111;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9736_4_lut_LC_10_15_2  (
            .in0(N__49276),
            .in1(N__49631),
            .in2(N__44236),
            .in3(N__46091),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i746_747_LC_10_15_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i746_747_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i746_747_LC_10_15_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i746_747_LC_10_15_3  (
            .in0(N__46588),
            .in1(N__44304),
            .in2(_gnd_net_),
            .in3(N__89651),
            .lcout(REG_mem_7_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93341),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i2_LC_10_15_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i2_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i2_LC_10_15_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i2_LC_10_15_4  (
            .in0(N__44224),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73293),
            .lcout(rp_sync1_r_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93341),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9754_4_lut_LC_10_15_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9754_4_lut_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9754_4_lut_LC_10_15_5 .LUT_INIT=16'b1110110110110111;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9754_4_lut_LC_10_15_5  (
            .in0(N__94296),
            .in1(N__50155),
            .in2(N__46098),
            .in3(N__44208),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i2_LC_10_15_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i2_LC_10_15_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i2_LC_10_15_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i2_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__73295),
            .in2(_gnd_net_),
            .in3(N__44176),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93341),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i3_LC_10_15_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i3_LC_10_15_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i3_LC_10_15_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i3_LC_10_15_7  (
            .in0(N__73294),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44164),
            .lcout(rp_sync1_r_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93341),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i938_939_LC_10_16_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i938_939_LC_10_16_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i938_939_LC_10_16_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i938_939_LC_10_16_0  (
            .in0(N__44151),
            .in1(N__46584),
            .in2(_gnd_net_),
            .in3(N__67156),
            .lcout(REG_mem_9_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11675_LC_10_16_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11675_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11675_LC_10_16_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11675_LC_10_16_1  (
            .in0(N__90978),
            .in1(N__87466),
            .in2(N__44254),
            .in3(N__44335),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13430_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13430_bdd_4_lut_LC_10_16_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13430_bdd_4_lut_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13430_bdd_4_lut_LC_10_16_2 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13430_bdd_4_lut_LC_10_16_2  (
            .in0(N__44344),
            .in1(N__44152),
            .in2(N__44140),
            .in3(N__90977),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i842_843_LC_10_16_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i842_843_LC_10_16_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i842_843_LC_10_16_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i842_843_LC_10_16_3  (
            .in0(N__46582),
            .in1(N__44343),
            .in2(_gnd_net_),
            .in3(N__67344),
            .lcout(REG_mem_8_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1034_1035_LC_10_16_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1034_1035_LC_10_16_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1034_1035_LC_10_16_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1034_1035_LC_10_16_4  (
            .in0(N__44334),
            .in1(N__46583),
            .in2(_gnd_net_),
            .in3(N__66960),
            .lcout(REG_mem_10_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2567_2568_LC_10_16_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2567_2568_LC_10_16_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2567_2568_LC_10_16_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2567_2568_LC_10_16_5  (
            .in0(N__70294),
            .in1(N__44532),
            .in2(_gnd_net_),
            .in3(N__47431),
            .lcout(REG_mem_26_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4013_4014_LC_10_16_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4013_4014_LC_10_16_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4013_4014_LC_10_16_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4013_4014_LC_10_16_6  (
            .in0(N__44319),
            .in1(N__47012),
            .in2(_gnd_net_),
            .in3(N__66006),
            .lcout(REG_mem_41_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93356),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10650_3_lut_LC_10_16_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10650_3_lut_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10650_3_lut_LC_10_16_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10650_3_lut_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(N__87465),
            .in2(N__44308),
            .in3(N__46168),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3812_3813_LC_10_17_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3812_3813_LC_10_17_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3812_3813_LC_10_17_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3812_3813_LC_10_17_0  (
            .in0(N__50709),
            .in1(N__48895),
            .in2(_gnd_net_),
            .in3(N__61885),
            .lcout(REG_mem_39_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2663_2664_LC_10_17_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2663_2664_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2663_2664_LC_10_17_1 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2663_2664_LC_10_17_1  (
            .in0(N__47429),
            .in1(N__94771),
            .in2(N__44520),
            .in3(N__79795),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i3_LC_10_17_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i3_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i3_LC_10_17_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i3_LC_10_17_2  (
            .in0(N__73296),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44284),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1130_1131_LC_10_17_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1130_1131_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1130_1131_LC_10_17_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1130_1131_LC_10_17_3  (
            .in0(N__46581),
            .in1(N__44247),
            .in2(_gnd_net_),
            .in3(N__66827),
            .lcout(REG_mem_11_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1895_1896_LC_10_17_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1895_1896_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1895_1896_LC_10_17_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1895_1896_LC_10_17_4  (
            .in0(N__44496),
            .in1(N__47430),
            .in2(_gnd_net_),
            .in3(N__72105),
            .lcout(REG_mem_19_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4973_4974_LC_10_17_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4973_4974_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4973_4974_LC_10_17_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4973_4974_LC_10_17_5  (
            .in0(N__47004),
            .in1(N__44355),
            .in2(_gnd_net_),
            .in3(N__72262),
            .lcout(REG_mem_51_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i461_462_LC_10_17_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i461_462_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i461_462_LC_10_17_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i461_462_LC_10_17_6  (
            .in0(N__44484),
            .in1(N__47005),
            .in2(_gnd_net_),
            .in3(N__72730),
            .lcout(REG_mem_4_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93368),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14222_bdd_4_lut_LC_10_17_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14222_bdd_4_lut_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14222_bdd_4_lut_LC_10_17_7 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14222_bdd_4_lut_LC_10_17_7  (
            .in0(N__91347),
            .in1(N__44485),
            .in2(N__46156),
            .in3(N__44410),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12051 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11670_LC_10_18_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11670_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11670_LC_10_18_0 .LUT_INIT=16'b1100101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11670_LC_10_18_0  (
            .in0(N__44461),
            .in1(N__44404),
            .in2(N__87175),
            .in3(N__91349),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12343_LC_10_18_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12343_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12343_LC_10_18_1 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12343_LC_10_18_1  (
            .in0(N__91351),
            .in1(N__86989),
            .in2(N__46060),
            .in3(N__44425),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3815_3816_LC_10_18_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3815_3816_LC_10_18_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3815_3816_LC_10_18_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3815_3816_LC_10_18_2  (
            .in0(N__44403),
            .in1(N__47428),
            .in2(_gnd_net_),
            .in3(N__61893),
            .lcout(REG_mem_39_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93381),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i6_LC_10_18_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i6_LC_10_18_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i6_LC_10_18_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i6_LC_10_18_3  (
            .in0(N__44390),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73297),
            .lcout(rp_sync1_r_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93381),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4781_4782_LC_10_18_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4781_4782_LC_10_18_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4781_4782_LC_10_18_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4781_4782_LC_10_18_4  (
            .in0(N__44655),
            .in1(N__47016),
            .in2(_gnd_net_),
            .in3(N__63005),
            .lcout(REG_mem_49_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93381),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11809_LC_10_18_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11809_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11809_LC_10_18_5 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11809_LC_10_18_5  (
            .in0(N__91350),
            .in1(N__45826),
            .in2(N__44359),
            .in3(N__86988),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13592_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13592_bdd_4_lut_LC_10_18_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13592_bdd_4_lut_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13592_bdd_4_lut_LC_10_18_6 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13592_bdd_4_lut_LC_10_18_6  (
            .in0(N__44656),
            .in1(N__91348),
            .in2(N__44647),
            .in3(N__44644),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11565_LC_10_18_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11565_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11565_LC_10_18_7 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11565_LC_10_18_7  (
            .in0(N__89978),
            .in1(N__84934),
            .in2(N__44617),
            .in3(N__47497),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2087_2088_LC_10_19_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2087_2088_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2087_2088_LC_10_19_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2087_2088_LC_10_19_0  (
            .in0(N__77045),
            .in1(N__47453),
            .in2(N__44592),
            .in3(N__94770),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93395),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3341_3342_LC_10_19_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3341_3342_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3341_3342_LC_10_19_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3341_3342_LC_10_19_1  (
            .in0(N__94768),
            .in1(N__44574),
            .in2(N__47041),
            .in3(N__80512),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93395),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1802_1803_LC_10_19_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1802_1803_LC_10_19_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1802_1803_LC_10_19_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1802_1803_LC_10_19_2  (
            .in0(N__44553),
            .in1(N__46471),
            .in2(_gnd_net_),
            .in3(N__67460),
            .lcout(REG_mem_18_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93395),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12043_LC_10_19_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12043_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12043_LC_10_19_3 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12043_LC_10_19_3  (
            .in0(N__86862),
            .in1(N__91355),
            .in2(N__44542),
            .in3(N__44521),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13874 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2471_2472_LC_10_19_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2471_2472_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2471_2472_LC_10_19_4 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2471_2472_LC_10_19_4  (
            .in0(N__44763),
            .in1(N__47454),
            .in2(N__95298),
            .in3(N__96981),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93395),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5543_5544_LC_10_19_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5543_5544_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5543_5544_LC_10_19_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5543_5544_LC_10_19_5  (
            .in0(N__96980),
            .in1(N__47676),
            .in2(N__47461),
            .in3(N__94776),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93395),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i269_270_LC_10_19_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i269_270_LC_10_19_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i269_270_LC_10_19_6 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i269_270_LC_10_19_6  (
            .in0(N__47040),
            .in1(N__94769),
            .in2(N__80570),
            .in3(N__44874),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93395),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6023_6024_LC_10_19_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6023_6024_LC_10_19_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6023_6024_LC_10_19_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6023_6024_LC_10_19_7  (
            .in0(N__47452),
            .in1(N__94772),
            .in2(N__47637),
            .in3(N__77935),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93395),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14144_bdd_4_lut_LC_10_20_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14144_bdd_4_lut_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14144_bdd_4_lut_LC_10_20_0 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14144_bdd_4_lut_LC_10_20_0  (
            .in0(N__91236),
            .in1(N__44863),
            .in2(N__44857),
            .in3(N__44833),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i173_174_LC_10_20_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i173_174_LC_10_20_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i173_174_LC_10_20_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i173_174_LC_10_20_4  (
            .in0(N__47011),
            .in1(N__95418),
            .in2(N__44811),
            .in3(N__80299),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93407),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13874_bdd_4_lut_LC_10_20_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13874_bdd_4_lut_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13874_bdd_4_lut_LC_10_20_5 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13874_bdd_4_lut_LC_10_20_5  (
            .in0(N__44794),
            .in1(N__91235),
            .in2(N__44770),
            .in3(N__44752),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13877 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13040_bdd_4_lut_LC_11_1_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13040_bdd_4_lut_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13040_bdd_4_lut_LC_11_1_0 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13040_bdd_4_lut_LC_11_1_0  (
            .in0(N__92620),
            .in1(N__44737),
            .in2(N__44974),
            .in3(N__44716),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13043_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10409_3_lut_LC_11_1_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10409_3_lut_LC_11_1_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10409_3_lut_LC_11_1_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10409_3_lut_LC_11_1_1  (
            .in0(_gnd_net_),
            .in1(N__85631),
            .in2(N__44701),
            .in3(N__44662),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12058 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11256_LC_11_1_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11256_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11256_LC_11_1_2 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11256_LC_11_1_2  (
            .in0(N__92621),
            .in1(N__45334),
            .in2(N__88880),
            .in3(N__44944),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12926_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12926_bdd_4_lut_LC_11_1_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12926_bdd_4_lut_LC_11_1_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12926_bdd_4_lut_LC_11_1_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12926_bdd_4_lut_LC_11_1_3  (
            .in0(N__44965),
            .in1(N__92619),
            .in2(N__44680),
            .in3(N__44677),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12929 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11350_LC_11_1_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11350_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11350_LC_11_1_4 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11350_LC_11_1_4  (
            .in0(N__88818),
            .in1(N__92622),
            .in2(N__44995),
            .in3(N__53365),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13040 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i563_564_LC_11_1_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i563_564_LC_11_1_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i563_564_LC_11_1_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i563_564_LC_11_1_5  (
            .in0(N__44964),
            .in1(N__62423),
            .in2(_gnd_net_),
            .in3(N__67864),
            .lcout(REG_mem_5_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93408),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11934_LC_11_1_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11934_LC_11_1_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11934_LC_11_1_6 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11934_LC_11_1_6  (
            .in0(N__88819),
            .in1(N__92623),
            .in2(N__51772),
            .in3(N__44956),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13742 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i659_660_LC_11_1_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i659_660_LC_11_1_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i659_660_LC_11_1_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i659_660_LC_11_1_7  (
            .in0(N__44943),
            .in1(N__62424),
            .in2(_gnd_net_),
            .in3(N__66424),
            .lcout(REG_mem_6_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93408),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4361_4362_LC_11_2_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4361_4362_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4361_4362_LC_11_2_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4361_4362_LC_11_2_1  (
            .in0(N__47949),
            .in1(N__96709),
            .in2(_gnd_net_),
            .in3(N__71885),
            .lcout(REG_mem_45_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4838_4839_LC_11_2_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4838_4839_LC_11_2_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4838_4839_LC_11_2_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4838_4839_LC_11_2_2  (
            .in0(N__44934),
            .in1(N__71455),
            .in2(_gnd_net_),
            .in3(N__73046),
            .lcout(REG_mem_50_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.usb3_data_in_latched__i1_LC_11_2_3 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i1_LC_11_2_3 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i1_LC_11_2_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i1_LC_11_2_3  (
            .in0(_gnd_net_),
            .in1(N__73681),
            .in2(_gnd_net_),
            .in3(N__44920),
            .lcout(\usb3_if_inst.usb3_data_in_latched_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4553_4554_LC_11_2_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4553_4554_LC_11_2_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4553_4554_LC_11_2_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4553_4554_LC_11_2_4  (
            .in0(N__96710),
            .in1(N__47799),
            .in2(_gnd_net_),
            .in3(N__66268),
            .lcout(REG_mem_47_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4649_4650_LC_11_2_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4649_4650_LC_11_2_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4649_4650_LC_11_2_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4649_4650_LC_11_2_5  (
            .in0(N__47823),
            .in1(N__96711),
            .in2(_gnd_net_),
            .in3(N__75579),
            .lcout(REG_mem_48_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5531_5532_LC_11_2_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5531_5532_LC_11_2_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5531_5532_LC_11_2_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5531_5532_LC_11_2_6  (
            .in0(N__63163),
            .in1(N__95772),
            .in2(N__45081),
            .in3(N__96989),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4745_4746_LC_11_2_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4745_4746_LC_11_2_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4745_4746_LC_11_2_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4745_4746_LC_11_2_7  (
            .in0(N__47811),
            .in1(N__96712),
            .in2(_gnd_net_),
            .in3(N__62997),
            .lcout(REG_mem_49_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93397),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13832_bdd_4_lut_LC_11_3_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13832_bdd_4_lut_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13832_bdd_4_lut_LC_11_3_0 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13832_bdd_4_lut_LC_11_3_0  (
            .in0(N__45064),
            .in1(N__92617),
            .in2(N__45022),
            .in3(N__45013),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13835_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10389_3_lut_LC_11_3_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10389_3_lut_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10389_3_lut_LC_11_3_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10389_3_lut_LC_11_3_1  (
            .in0(N__85754),
            .in1(_gnd_net_),
            .in2(N__45049),
            .in3(N__51571),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12038 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4457_4458_LC_11_3_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4457_4458_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4457_4458_LC_11_3_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4457_4458_LC_11_3_2  (
            .in0(N__47788),
            .in1(N__96784),
            .in2(_gnd_net_),
            .in3(N__89122),
            .lcout(REG_mem_46_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93384),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10370_3_lut_LC_11_3_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10370_3_lut_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10370_3_lut_LC_11_3_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10370_3_lut_LC_11_3_3  (
            .in0(N__45271),
            .in1(N__88006),
            .in2(_gnd_net_),
            .in3(N__45256),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12019 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12008_LC_11_3_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12008_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12008_LC_11_3_4 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12008_LC_11_3_4  (
            .in0(N__88007),
            .in1(N__92618),
            .in2(N__45145),
            .in3(N__45004),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13832 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1286_1287_LC_11_3_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1286_1287_LC_11_3_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1286_1287_LC_11_3_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1286_1287_LC_11_3_5  (
            .in0(N__45012),
            .in1(N__71492),
            .in2(_gnd_net_),
            .in3(N__70113),
            .lcout(REG_mem_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93384),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2837_2838_LC_11_3_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2837_2838_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2837_2838_LC_11_3_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2837_2838_LC_11_3_6  (
            .in0(N__62796),
            .in1(N__95582),
            .in2(N__56187),
            .in3(N__70990),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93384),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1382_1383_LC_11_3_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1382_1383_LC_11_3_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1382_1383_LC_11_3_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1382_1383_LC_11_3_7  (
            .in0(N__45003),
            .in1(N__71493),
            .in2(_gnd_net_),
            .in3(N__74757),
            .lcout(REG_mem_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93384),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10365_3_lut_LC_11_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10365_3_lut_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10365_3_lut_LC_11_4_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10365_3_lut_LC_11_4_0  (
            .in0(N__88448),
            .in1(N__47938),
            .in2(_gnd_net_),
            .in3(N__45172),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12014 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4844_4845_LC_11_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4844_4845_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4844_4845_LC_11_4_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4844_4845_LC_11_4_1  (
            .in0(N__75955),
            .in1(N__45213),
            .in2(_gnd_net_),
            .in3(N__73025),
            .lcout(REG_mem_50_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93370),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4595_4596_LC_11_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4595_4596_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4595_4596_LC_11_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4595_4596_LC_11_4_2  (
            .in0(N__62374),
            .in1(N__45171),
            .in2(_gnd_net_),
            .in3(N__66259),
            .lcout(REG_mem_47_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93370),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4403_4404_LC_11_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4403_4404_LC_11_4_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4403_4404_LC_11_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4403_4404_LC_11_4_3  (
            .in0(N__45156),
            .in1(N__62375),
            .in2(_gnd_net_),
            .in3(N__71884),
            .lcout(REG_mem_45_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93370),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1685_1686_LC_11_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1685_1686_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1685_1686_LC_11_4_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1685_1686_LC_11_4_4  (
            .in0(N__55827),
            .in1(N__62801),
            .in2(_gnd_net_),
            .in3(N__66577),
            .lcout(REG_mem_17_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93370),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1478_1479_LC_11_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1478_1479_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1478_1479_LC_11_4_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1478_1479_LC_11_4_5  (
            .in0(N__45141),
            .in1(N__71494),
            .in2(_gnd_net_),
            .in3(N__64006),
            .lcout(REG_mem_15_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93370),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5324_5325_LC_11_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5324_5325_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5324_5325_LC_11_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5324_5325_LC_11_4_6  (
            .in0(N__75954),
            .in1(N__59097),
            .in2(_gnd_net_),
            .in3(N__77229),
            .lcout(REG_mem_55_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93370),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13976_bdd_4_lut_LC_11_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13976_bdd_4_lut_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13976_bdd_4_lut_LC_11_4_7 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13976_bdd_4_lut_LC_11_4_7  (
            .in0(N__90859),
            .in1(N__45196),
            .in2(N__45130),
            .in3(N__48058),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13979 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1043_1044_LC_11_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1043_1044_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1043_1044_LC_11_5_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1043_1044_LC_11_5_0  (
            .in0(N__66979),
            .in1(N__45102),
            .in2(_gnd_net_),
            .in3(N__62373),
            .lcout(REG_mem_10_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4787_4788_LC_11_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4787_4788_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4787_4788_LC_11_5_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4787_4788_LC_11_5_1  (
            .in0(N__62371),
            .in1(N__45267),
            .in2(_gnd_net_),
            .in3(N__62979),
            .lcout(REG_mem_49_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4691_4692_LC_11_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4691_4692_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4691_4692_LC_11_5_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4691_4692_LC_11_5_2  (
            .in0(N__45252),
            .in1(N__62372),
            .in2(_gnd_net_),
            .in3(N__75572),
            .lcout(REG_mem_48_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1493_1494_LC_11_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1493_1494_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1493_1494_LC_11_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1493_1494_LC_11_5_3  (
            .in0(N__58779),
            .in1(N__62813),
            .in2(_gnd_net_),
            .in3(N__63980),
            .lcout(REG_mem_15_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1589_1590_LC_11_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1589_1590_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1589_1590_LC_11_5_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1589_1590_LC_11_5_4  (
            .in0(N__65678),
            .in1(_gnd_net_),
            .in2(N__62854),
            .in3(N__55842),
            .lcout(REG_mem_16_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1001_1002_LC_11_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1001_1002_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1001_1002_LC_11_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1001_1002_LC_11_5_5  (
            .in0(N__48000),
            .in1(N__96773),
            .in2(_gnd_net_),
            .in3(N__66978),
            .lcout(REG_mem_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1781_1782_LC_11_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1781_1782_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1781_1782_LC_11_5_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1781_1782_LC_11_5_6  (
            .in0(N__62812),
            .in1(N__55980),
            .in2(_gnd_net_),
            .in3(N__67467),
            .lcout(REG_mem_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1577_1578_LC_11_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1577_1578_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1577_1578_LC_11_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1577_1578_LC_11_5_7  (
            .in0(N__55800),
            .in1(N__96774),
            .in2(_gnd_net_),
            .in3(N__65677),
            .lcout(REG_mem_16_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93357),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4391_4392_LC_11_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4391_4392_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4391_4392_LC_11_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4391_4392_LC_11_6_0  (
            .in0(N__45228),
            .in1(N__47180),
            .in2(_gnd_net_),
            .in3(N__71850),
            .lcout(REG_mem_45_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93342),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12128_LC_11_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12128_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12128_LC_11_6_1 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12128_LC_11_6_1  (
            .in0(N__92062),
            .in1(N__88446),
            .in2(N__45217),
            .in3(N__45319),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13976 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4757_4758_LC_11_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4757_4758_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4757_4758_LC_11_6_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4757_4758_LC_11_6_2  (
            .in0(N__62978),
            .in1(N__48345),
            .in2(_gnd_net_),
            .in3(N__62802),
            .lcout(REG_mem_49_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93342),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i755_756_LC_11_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i755_756_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i755_756_LC_11_6_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i755_756_LC_11_6_3  (
            .in0(N__89626),
            .in1(N__45330),
            .in2(_gnd_net_),
            .in3(N__62383),
            .lcout(REG_mem_7_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93342),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3785_3786_LC_11_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3785_3786_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3785_3786_LC_11_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3785_3786_LC_11_6_4  (
            .in0(N__53556),
            .in1(N__96775),
            .in2(_gnd_net_),
            .in3(N__61830),
            .lcout(REG_mem_39_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93342),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4940_4941_LC_11_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4940_4941_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4940_4941_LC_11_6_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4940_4941_LC_11_6_5  (
            .in0(N__75939),
            .in1(N__45318),
            .in2(_gnd_net_),
            .in3(N__72207),
            .lcout(REG_mem_51_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93342),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i716_717_LC_11_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i716_717_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i716_717_LC_11_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i716_717_LC_11_6_6  (
            .in0(N__47889),
            .in1(N__75940),
            .in2(_gnd_net_),
            .in3(N__89624),
            .lcout(REG_mem_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93342),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i725_726_LC_11_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i725_726_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i725_726_LC_11_6_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i725_726_LC_11_6_7  (
            .in0(N__89625),
            .in1(N__62803),
            .in2(_gnd_net_),
            .in3(N__51315),
            .lcout(REG_mem_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93342),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i722_723_LC_11_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i722_723_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i722_723_LC_11_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i722_723_LC_11_7_0  (
            .in0(N__62001),
            .in1(N__76744),
            .in2(_gnd_net_),
            .in3(N__89610),
            .lcout(REG_mem_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93329),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3782_3783_LC_11_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3782_3783_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3782_3783_LC_11_7_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3782_3783_LC_11_7_1  (
            .in0(N__53805),
            .in1(N__61827),
            .in2(_gnd_net_),
            .in3(N__71555),
            .lcout(REG_mem_39_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93329),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3713_3714_LC_11_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3713_3714_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3713_3714_LC_11_7_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3713_3714_LC_11_7_2  (
            .in0(N__56569),
            .in1(N__45300),
            .in2(_gnd_net_),
            .in3(N__59239),
            .lcout(REG_mem_38_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93329),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4001_4002_LC_11_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4001_4002_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4001_4002_LC_11_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4001_4002_LC_11_7_3  (
            .in0(N__66015),
            .in1(N__45282),
            .in2(_gnd_net_),
            .in3(N__56570),
            .lcout(REG_mem_41_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93329),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3635_3636_LC_11_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3635_3636_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3635_3636_LC_11_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3635_3636_LC_11_7_4  (
            .in0(N__45372),
            .in1(N__62414),
            .in2(_gnd_net_),
            .in3(N__63676),
            .lcout(REG_mem_37_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93329),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i731_732_LC_11_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i731_732_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i731_732_LC_11_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i731_732_LC_11_7_5  (
            .in0(N__89611),
            .in1(N__51975),
            .in2(_gnd_net_),
            .in3(N__63534),
            .lcout(REG_mem_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93329),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3998_3999_LC_11_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3998_3999_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3998_3999_LC_11_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3998_3999_LC_11_7_6  (
            .in0(N__85872),
            .in1(N__89527),
            .in2(_gnd_net_),
            .in3(N__66016),
            .lcout(REG_mem_41_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93329),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1094_1095_LC_11_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1094_1095_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1094_1095_LC_11_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1094_1095_LC_11_7_7  (
            .in0(N__51810),
            .in1(N__71554),
            .in2(_gnd_net_),
            .in3(N__66762),
            .lcout(REG_mem_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93329),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1598_1599_LC_11_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1598_1599_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1598_1599_LC_11_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1598_1599_LC_11_8_0  (
            .in0(N__89475),
            .in1(N__67524),
            .in2(_gnd_net_),
            .in3(N__65650),
            .lcout(REG_mem_16_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93316),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11485_LC_11_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11485_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11485_LC_11_8_1 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11485_LC_11_8_1  (
            .in0(N__91797),
            .in1(N__53842),
            .in2(N__48361),
            .in3(N__88148),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13202_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13202_bdd_4_lut_LC_11_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13202_bdd_4_lut_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13202_bdd_4_lut_LC_11_8_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13202_bdd_4_lut_LC_11_8_2  (
            .in0(N__48451),
            .in1(N__91796),
            .in2(N__45361),
            .in3(N__45343),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1217_1218_LC_11_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1217_1218_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1217_1218_LC_11_8_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1217_1218_LC_11_8_3  (
            .in0(N__45342),
            .in1(_gnd_net_),
            .in2(N__56606),
            .in3(N__59634),
            .lcout(REG_mem_12_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93316),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3902_3903_LC_11_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3902_3903_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3902_3903_LC_11_8_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3902_3903_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__85893),
            .in2(N__89518),
            .in3(N__65839),
            .lcout(REG_mem_40_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93316),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3608_3609_LC_11_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3608_3609_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3608_3609_LC_11_8_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3608_3609_LC_11_8_5  (
            .in0(N__53448),
            .in1(N__63636),
            .in2(_gnd_net_),
            .in3(N__96382),
            .lcout(REG_mem_37_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93316),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i545_546_LC_11_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i545_546_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i545_546_LC_11_8_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i545_546_LC_11_8_6  (
            .in0(N__45420),
            .in1(N__67799),
            .in2(_gnd_net_),
            .in3(N__56571),
            .lcout(REG_mem_5_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93316),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1691_1692_LC_11_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1691_1692_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1691_1692_LC_11_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1691_1692_LC_11_8_7  (
            .in0(N__52023),
            .in1(N__63544),
            .in2(_gnd_net_),
            .in3(N__66489),
            .lcout(REG_mem_17_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93316),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i79_2_lut_3_lut_4_lut_LC_11_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i79_2_lut_3_lut_4_lut_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i79_2_lut_3_lut_4_lut_LC_11_9_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i79_2_lut_3_lut_4_lut_LC_11_9_0  (
            .in0(N__45406),
            .in1(N__49581),
            .in2(N__94480),
            .in3(N__49783),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i80_2_lut_3_lut_4_lut_LC_11_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i80_2_lut_3_lut_4_lut_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i80_2_lut_3_lut_4_lut_LC_11_9_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i80_2_lut_3_lut_4_lut_LC_11_9_1  (
            .in0(N__49784),
            .in1(N__94048),
            .in2(N__49596),
            .in3(N__45407),
            .lcout(n60),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i95_2_lut_3_lut_4_lut_LC_11_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i95_2_lut_3_lut_4_lut_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i95_2_lut_3_lut_4_lut_LC_11_9_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i95_2_lut_3_lut_4_lut_LC_11_9_2  (
            .in0(N__45408),
            .in1(N__49582),
            .in2(N__94481),
            .in3(N__49792),
            .lcout(n20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i96_2_lut_3_lut_4_lut_LC_11_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i96_2_lut_3_lut_4_lut_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i96_2_lut_3_lut_4_lut_LC_11_9_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i96_2_lut_3_lut_4_lut_LC_11_9_3  (
            .in0(N__49785),
            .in1(N__94050),
            .in2(N__49597),
            .in3(N__45409),
            .lcout(n52),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i81_2_lut_3_lut_4_lut_LC_11_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i81_2_lut_3_lut_4_lut_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i81_2_lut_3_lut_4_lut_LC_11_9_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i81_2_lut_3_lut_4_lut_LC_11_9_4  (
            .in0(N__49448),
            .in1(N__49793),
            .in2(N__94482),
            .in3(N__45559),
            .lcout(n27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i82_2_lut_3_lut_4_lut_LC_11_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i82_2_lut_3_lut_4_lut_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i82_2_lut_3_lut_4_lut_LC_11_9_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i82_2_lut_3_lut_4_lut_LC_11_9_5  (
            .in0(N__45560),
            .in1(N__94049),
            .in2(N__49838),
            .in3(N__49446),
            .lcout(n59),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6116_6117_LC_11_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6116_6117_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6116_6117_LC_11_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6116_6117_LC_11_9_6  (
            .in0(N__48769),
            .in1(N__45384),
            .in2(_gnd_net_),
            .in3(N__67623),
            .lcout(REG_mem_63_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93301),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i98_2_lut_3_lut_4_lut_LC_11_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i98_2_lut_3_lut_4_lut_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i98_2_lut_3_lut_4_lut_LC_11_9_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i98_2_lut_3_lut_4_lut_LC_11_9_7  (
            .in0(N__45561),
            .in1(N__94051),
            .in2(N__49839),
            .in3(N__49447),
            .lcout(n51),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i100_2_lut_3_lut_LC_11_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i100_2_lut_3_lut_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i100_2_lut_3_lut_LC_11_10_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i100_2_lut_3_lut_LC_11_10_0  (
            .in0(N__49480),
            .in1(N__45472),
            .in2(_gnd_net_),
            .in3(N__93773),
            .lcout(n50),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i5_LC_11_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i5_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i5_LC_11_10_1 .LUT_INIT=16'b0001101111100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i5_LC_11_10_1  (
            .in0(N__49140),
            .in1(N__49275),
            .in2(N__94103),
            .in3(N__45490),
            .lcout(wr_grey_sync_r_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93279),
            .ce(),
            .sr(N__73464));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i5_3_lut_LC_11_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i5_3_lut_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i5_3_lut_LC_11_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_135_i5_3_lut_LC_11_10_2  (
            .in0(N__49481),
            .in1(N__49297),
            .in2(_gnd_net_),
            .in3(N__49138),
            .lcout(wr_addr_nxt_c_4),
            .ltout(wr_addr_nxt_c_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i4_LC_11_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i4_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i4_LC_11_10_3 .LUT_INIT=16'b0001111010110100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_grey_sync_r__i4_LC_11_10_3  (
            .in0(N__49139),
            .in1(N__49274),
            .in2(N__45478),
            .in3(N__93769),
            .lcout(wr_grey_sync_r_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93279),
            .ce(),
            .sr(N__73464));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i131_2_lut_3_lut_LC_11_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i131_2_lut_3_lut_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i131_2_lut_3_lut_LC_11_10_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i131_2_lut_3_lut_LC_11_10_4  (
            .in0(N__49477),
            .in1(N__45473),
            .in2(_gnd_net_),
            .in3(N__93771),
            .lcout(n2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i132_2_lut_3_lut_LC_11_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i132_2_lut_3_lut_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i132_2_lut_3_lut_LC_11_10_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i132_2_lut_3_lut_LC_11_10_5  (
            .in0(N__45474),
            .in1(N__93768),
            .in2(_gnd_net_),
            .in3(N__49476),
            .lcout(n34),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i99_2_lut_3_lut_LC_11_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i99_2_lut_3_lut_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i99_2_lut_3_lut_LC_11_10_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i99_2_lut_3_lut_LC_11_10_6  (
            .in0(N__49479),
            .in1(N__45475),
            .in2(_gnd_net_),
            .in3(N__93772),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i105_2_lut_3_lut_LC_11_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i105_2_lut_3_lut_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i105_2_lut_3_lut_LC_11_10_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i105_2_lut_3_lut_LC_11_10_7  (
            .in0(N__93770),
            .in1(N__49478),
            .in2(_gnd_net_),
            .in3(N__45460),
            .lcout(n15_adj_1184),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12433_LC_11_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12433_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12433_LC_11_11_0 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12433_LC_11_11_0  (
            .in0(N__49162),
            .in1(N__90858),
            .in2(N__45634),
            .in3(N__88070),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1391_1392_LC_11_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1391_1392_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1391_1392_LC_11_11_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1391_1392_LC_11_11_1  (
            .in0(N__45630),
            .in1(N__61307),
            .in2(_gnd_net_),
            .in3(N__74703),
            .lcout(REG_mem_14_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4871_4872_LC_11_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4871_4872_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4871_4872_LC_11_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4871_4872_LC_11_11_2  (
            .in0(N__47410),
            .in1(N__45864),
            .in2(_gnd_net_),
            .in3(N__72941),
            .lcout(REG_mem_50_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1295_1296_LC_11_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1295_1296_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1295_1296_LC_11_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1295_1296_LC_11_11_3  (
            .in0(N__45615),
            .in1(N__61306),
            .in2(_gnd_net_),
            .in3(N__70102),
            .lcout(REG_mem_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1517_1518_LC_11_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1517_1518_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1517_1518_LC_11_11_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1517_1518_LC_11_11_4  (
            .in0(N__45594),
            .in1(N__46901),
            .in2(_gnd_net_),
            .in3(N__63953),
            .lcout(REG_mem_15_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4205_4206_LC_11_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4205_4206_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4205_4206_LC_11_11_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4205_4206_LC_11_11_5  (
            .in0(N__46900),
            .in1(N__45573),
            .in2(_gnd_net_),
            .in3(N__68237),
            .lcout(REG_mem_43_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i97_2_lut_3_lut_4_lut_LC_11_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i97_2_lut_3_lut_4_lut_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i97_2_lut_3_lut_4_lut_LC_11_11_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.EnabledDecoder_2_i97_2_lut_3_lut_4_lut_LC_11_11_6  (
            .in0(N__49407),
            .in1(N__49701),
            .in2(N__94102),
            .in3(N__45562),
            .lcout(n19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4583_4584_LC_11_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4583_4584_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4583_4584_LC_11_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4583_4584_LC_11_11_7  (
            .in0(N__66183),
            .in1(N__45534),
            .in2(_gnd_net_),
            .in3(N__47411),
            .lcout(REG_mem_47_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93302),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3695_3696_LC_11_12_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3695_3696_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3695_3696_LC_11_12_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3695_3696_LC_11_12_0  (
            .in0(N__45513),
            .in1(N__61240),
            .in2(_gnd_net_),
            .in3(N__59243),
            .lcout(REG_mem_38_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93317),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11944_LC_11_12_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11944_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11944_LC_11_12_1 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11944_LC_11_12_1  (
            .in0(N__87527),
            .in1(N__90857),
            .in2(N__46033),
            .in3(N__45744),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13754 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1403_1404_LC_11_12_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1403_1404_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1403_1404_LC_11_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1403_1404_LC_11_12_2  (
            .in0(N__45777),
            .in1(N__63509),
            .in2(_gnd_net_),
            .in3(N__74704),
            .lcout(REG_mem_14_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93317),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4490_4491_LC_11_12_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4490_4491_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4490_4491_LC_11_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4490_4491_LC_11_12_3  (
            .in0(N__45759),
            .in1(N__46585),
            .in2(_gnd_net_),
            .in3(N__89011),
            .lcout(REG_mem_46_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93317),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3335_3336_LC_11_12_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3335_3336_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3335_3336_LC_11_12_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3335_3336_LC_11_12_4  (
            .in0(N__47412),
            .in1(N__93815),
            .in2(N__45745),
            .in3(N__80445),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93317),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5615_5616_LC_11_12_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5615_5616_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5615_5616_LC_11_12_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5615_5616_LC_11_12_5  (
            .in0(N__61239),
            .in1(N__45720),
            .in2(_gnd_net_),
            .in3(N__79911),
            .lcout(REG_mem_58_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93317),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3053_3054_LC_11_12_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3053_3054_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3053_3054_LC_11_12_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3053_3054_LC_11_12_6  (
            .in0(N__45699),
            .in1(N__46902),
            .in2(_gnd_net_),
            .in3(N__72491),
            .lcout(REG_mem_31_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93317),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4487_4488_LC_11_12_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4487_4488_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4487_4488_LC_11_12_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4487_4488_LC_11_12_7  (
            .in0(N__45681),
            .in1(_gnd_net_),
            .in2(N__47451),
            .in3(N__89010),
            .lcout(REG_mem_46_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93317),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1322_1323_LC_11_13_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1322_1323_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1322_1323_LC_11_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1322_1323_LC_11_13_0  (
            .in0(N__70100),
            .in1(N__45669),
            .in2(_gnd_net_),
            .in3(N__46568),
            .lcout(REG_mem_13_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11660_LC_11_13_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11660_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11660_LC_11_13_1 .LUT_INIT=16'b1011110010110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11660_LC_11_13_1  (
            .in0(N__45877),
            .in1(N__90856),
            .in2(N__87792),
            .in3(N__45886),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13412_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13412_bdd_4_lut_LC_11_13_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13412_bdd_4_lut_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13412_bdd_4_lut_LC_11_13_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13412_bdd_4_lut_LC_11_13_2  (
            .in0(N__90855),
            .in1(N__45670),
            .in2(N__45661),
            .in3(N__45643),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1226_1227_LC_11_13_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1226_1227_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1226_1227_LC_11_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1226_1227_LC_11_13_3  (
            .in0(N__45642),
            .in1(N__46565),
            .in2(_gnd_net_),
            .in3(N__59644),
            .lcout(REG_mem_12_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1418_1419_LC_11_13_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1418_1419_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1418_1419_LC_11_13_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1418_1419_LC_11_13_4  (
            .in0(N__45885),
            .in1(N__46567),
            .in2(_gnd_net_),
            .in3(N__74741),
            .lcout(REG_mem_14_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1514_1515_LC_11_13_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1514_1515_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1514_1515_LC_11_13_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1514_1515_LC_11_13_5  (
            .in0(N__45876),
            .in1(N__46566),
            .in2(_gnd_net_),
            .in3(N__63984),
            .lcout(REG_mem_15_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6119_6120_LC_11_13_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6119_6120_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6119_6120_LC_11_13_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6119_6120_LC_11_13_6  (
            .in0(N__47408),
            .in1(N__47655),
            .in2(_gnd_net_),
            .in3(N__67667),
            .lcout(REG_mem_63_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5639_5640_LC_11_13_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5639_5640_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5639_5640_LC_11_13_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5639_5640_LC_11_13_7  (
            .in0(N__79946),
            .in1(N__47736),
            .in2(_gnd_net_),
            .in3(N__47409),
            .lcout(REG_mem_58_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93330),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4775_4776_LC_11_14_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4775_4776_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4775_4776_LC_11_14_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4775_4776_LC_11_14_0  (
            .in0(N__45852),
            .in1(N__47435),
            .in2(_gnd_net_),
            .in3(N__62996),
            .lcout(REG_mem_49_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12318_LC_11_14_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12318_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12318_LC_11_14_1 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12318_LC_11_14_1  (
            .in0(N__90854),
            .in1(N__46042),
            .in2(N__87791),
            .in3(N__45868),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14204_bdd_4_lut_LC_11_14_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14204_bdd_4_lut_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14204_bdd_4_lut_LC_11_14_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14204_bdd_4_lut_LC_11_14_2  (
            .in0(N__45853),
            .in1(N__90853),
            .in2(N__45844),
            .in3(N__45841),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4877_4878_LC_11_14_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4877_4878_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4877_4878_LC_11_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4877_4878_LC_11_14_3  (
            .in0(N__47021),
            .in1(N__45819),
            .in2(_gnd_net_),
            .in3(N__72993),
            .lcout(REG_mem_50_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4589_4590_LC_11_14_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4589_4590_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4589_4590_LC_11_14_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4589_4590_LC_11_14_4  (
            .in0(N__45801),
            .in1(N__47022),
            .in2(_gnd_net_),
            .in3(N__66250),
            .lcout(REG_mem_47_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4967_4968_LC_11_14_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4967_4968_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4967_4968_LC_11_14_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4967_4968_LC_11_14_5  (
            .in0(N__47432),
            .in1(N__46041),
            .in2(_gnd_net_),
            .in3(N__72257),
            .lcout(REG_mem_51_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3431_3432_LC_11_14_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3431_3432_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3431_3432_LC_11_14_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3431_3432_LC_11_14_6  (
            .in0(N__94591),
            .in1(N__47434),
            .in2(N__46026),
            .in3(N__83328),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i551_552_LC_11_14_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i551_552_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i551_552_LC_11_14_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i551_552_LC_11_14_7  (
            .in0(N__47433),
            .in1(N__46002),
            .in2(_gnd_net_),
            .in3(N__67846),
            .lcout(REG_mem_5_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93343),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3629_3630_LC_11_15_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3629_3630_LC_11_15_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3629_3630_LC_11_15_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3629_3630_LC_11_15_0  (
            .in0(N__46995),
            .in1(N__45990),
            .in2(_gnd_net_),
            .in3(N__63677),
            .lcout(REG_mem_37_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93358),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12018_LC_11_15_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12018_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12018_LC_11_15_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12018_LC_11_15_1  (
            .in0(N__45910),
            .in1(N__90635),
            .in2(N__45901),
            .in3(N__87334),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13838_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13838_bdd_4_lut_LC_11_15_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13838_bdd_4_lut_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13838_bdd_4_lut_LC_11_15_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13838_bdd_4_lut_LC_11_15_2  (
            .in0(N__90634),
            .in1(N__45991),
            .in2(N__45982),
            .in3(N__45979),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12189 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2_3_lut_adj_46_LC_11_15_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2_3_lut_adj_46_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2_3_lut_adj_46_LC_11_15_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2_3_lut_adj_46_LC_11_15_3  (
            .in0(N__52852),
            .in1(N__46123),
            .in2(_gnd_net_),
            .in3(N__46116),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3725_3726_LC_11_15_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3725_3726_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3725_3726_LC_11_15_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3725_3726_LC_11_15_4  (
            .in0(N__46996),
            .in1(N__45909),
            .in2(_gnd_net_),
            .in3(N__59273),
            .lcout(REG_mem_38_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93358),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3821_3822_LC_11_15_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3821_3822_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3821_3822_LC_11_15_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3821_3822_LC_11_15_5  (
            .in0(N__45897),
            .in1(N__46997),
            .in2(_gnd_net_),
            .in3(N__61894),
            .lcout(REG_mem_39_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93358),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4874_4875_LC_11_15_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4874_4875_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4874_4875_LC_11_15_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4874_4875_LC_11_15_6  (
            .in0(N__46599),
            .in1(_gnd_net_),
            .in2(N__46586),
            .in3(N__72994),
            .lcout(REG_mem_50_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93358),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i650_651_LC_11_15_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i650_651_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i650_651_LC_11_15_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i650_651_LC_11_15_7  (
            .in0(N__66412),
            .in1(N__46167),
            .in2(_gnd_net_),
            .in3(N__46569),
            .lcout(REG_mem_6_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93358),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i557_558_LC_11_16_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i557_558_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i557_558_LC_11_16_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i557_558_LC_11_16_0  (
            .in0(N__46152),
            .in1(N__46998),
            .in2(_gnd_net_),
            .in3(N__67847),
            .lcout(REG_mem_5_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i4_LC_11_16_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i4_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i4_LC_11_16_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i4_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__73465),
            .in2(_gnd_net_),
            .in3(N__46141),
            .lcout(rp_sync1_r_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i4_LC_11_16_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i4_LC_11_16_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i4_LC_11_16_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i4_LC_11_16_2  (
            .in0(N__73467),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46129),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i5_LC_11_16_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i5_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i5_LC_11_16_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i5_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__73468),
            .in2(_gnd_net_),
            .in3(N__46066),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_6__I_0_136_i1_2_lut_LC_11_16_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_6__I_0_136_i1_2_lut_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_6__I_0_136_i1_2_lut_LC_11_16_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_6__I_0_136_i1_2_lut_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__52853),
            .in2(_gnd_net_),
            .in3(N__46117),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync_w_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i5_LC_11_16_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i5_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i5_LC_11_16_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync1_r__i5_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__73466),
            .in2(_gnd_net_),
            .in3(N__46078),
            .lcout(rp_sync1_r_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i653_654_LC_11_16_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i653_654_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i653_654_LC_11_16_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i653_654_LC_11_16_6  (
            .in0(N__66402),
            .in1(N__46053),
            .in2(_gnd_net_),
            .in3(N__46999),
            .lcout(REG_mem_6_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i6_LC_11_16_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i6_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i6_LC_11_16_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r__i6_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__73469),
            .in2(_gnd_net_),
            .in3(N__47518),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rp_sync2_r_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93371),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1319_1320_LC_11_17_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1319_1320_LC_11_17_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1319_1320_LC_11_17_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1319_1320_LC_11_17_0  (
            .in0(N__70101),
            .in1(_gnd_net_),
            .in2(N__47460),
            .in3(N__47508),
            .lcout(REG_mem_13_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93383),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12478_LC_11_17_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12478_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12478_LC_11_17_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12478_LC_11_17_1  (
            .in0(N__47482),
            .in1(N__91111),
            .in2(N__47473),
            .in3(N__87259),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14396_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14396_bdd_4_lut_LC_11_17_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14396_bdd_4_lut_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14396_bdd_4_lut_LC_11_17_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14396_bdd_4_lut_LC_11_17_2  (
            .in0(N__91110),
            .in1(N__47509),
            .in2(N__47500),
            .in3(N__47491),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1223_1224_LC_11_17_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1223_1224_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1223_1224_LC_11_17_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1223_1224_LC_11_17_3  (
            .in0(N__47490),
            .in1(N__47446),
            .in2(_gnd_net_),
            .in3(N__59657),
            .lcout(REG_mem_12_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93383),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1415_1416_LC_11_17_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1415_1416_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1415_1416_LC_11_17_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1415_1416_LC_11_17_4  (
            .in0(N__47444),
            .in1(N__47481),
            .in2(_gnd_net_),
            .in3(N__74763),
            .lcout(REG_mem_14_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93383),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1511_1512_LC_11_17_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1511_1512_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1511_1512_LC_11_17_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1511_1512_LC_11_17_5  (
            .in0(N__47469),
            .in1(N__47447),
            .in2(_gnd_net_),
            .in3(N__63985),
            .lcout(REG_mem_15_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93383),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i647_648_LC_11_17_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i647_648_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i647_648_LC_11_17_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i647_648_LC_11_17_6  (
            .in0(N__47445),
            .in1(N__47052),
            .in2(_gnd_net_),
            .in3(N__66423),
            .lcout(REG_mem_6_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93383),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4397_4398_LC_11_17_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4397_4398_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4397_4398_LC_11_17_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4397_4398_LC_11_17_7  (
            .in0(N__46620),
            .in1(N__47000),
            .in2(_gnd_net_),
            .in3(N__71878),
            .lcout(REG_mem_45_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93383),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.counter_1109__i0_LC_11_18_0 .C_ON=1'b1;
    defparam \spi0.counter_1109__i0_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \spi0.counter_1109__i0_LC_11_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.counter_1109__i0_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__50935),
            .in2(_gnd_net_),
            .in3(N__47545),
            .lcout(\spi0.counter_0 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\spi0.n10694 ),
            .clk(N__97363),
            .ce(N__52945),
            .sr(N__53032));
    defparam \spi0.counter_1109__i1_LC_11_18_1 .C_ON=1'b1;
    defparam \spi0.counter_1109__i1_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \spi0.counter_1109__i1_LC_11_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.counter_1109__i1_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__50980),
            .in2(N__86655),
            .in3(N__47542),
            .lcout(\spi0.counter_1 ),
            .ltout(),
            .carryin(\spi0.n10694 ),
            .carryout(\spi0.n10695 ),
            .clk(N__97363),
            .ce(N__52945),
            .sr(N__53032));
    defparam \spi0.counter_1109__i2_LC_11_18_2 .C_ON=1'b1;
    defparam \spi0.counter_1109__i2_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \spi0.counter_1109__i2_LC_11_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.counter_1109__i2_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__50959),
            .in2(N__86659),
            .in3(N__47539),
            .lcout(\spi0.counter_2 ),
            .ltout(),
            .carryin(\spi0.n10695 ),
            .carryout(\spi0.n10696 ),
            .clk(N__97363),
            .ce(N__52945),
            .sr(N__53032));
    defparam \spi0.counter_1109__i3_LC_11_18_3 .C_ON=1'b1;
    defparam \spi0.counter_1109__i3_LC_11_18_3 .SEQ_MODE=4'b1000;
    defparam \spi0.counter_1109__i3_LC_11_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.counter_1109__i3_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__50998),
            .in2(N__86656),
            .in3(N__47536),
            .lcout(\spi0.counter_3 ),
            .ltout(),
            .carryin(\spi0.n10696 ),
            .carryout(\spi0.n10697 ),
            .clk(N__97363),
            .ce(N__52945),
            .sr(N__53032));
    defparam \spi0.counter_1109__i4_LC_11_18_4 .C_ON=1'b1;
    defparam \spi0.counter_1109__i4_LC_11_18_4 .SEQ_MODE=4'b1000;
    defparam \spi0.counter_1109__i4_LC_11_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.counter_1109__i4_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__52793),
            .in2(N__86660),
            .in3(N__47533),
            .lcout(\spi0.counter_4 ),
            .ltout(),
            .carryin(\spi0.n10697 ),
            .carryout(\spi0.n10698 ),
            .clk(N__97363),
            .ce(N__52945),
            .sr(N__53032));
    defparam \spi0.counter_1109__i5_LC_11_18_5 .C_ON=1'b1;
    defparam \spi0.counter_1109__i5_LC_11_18_5 .SEQ_MODE=4'b1000;
    defparam \spi0.counter_1109__i5_LC_11_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.counter_1109__i5_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__51063),
            .in2(N__86657),
            .in3(N__47530),
            .lcout(\spi0.counter_5 ),
            .ltout(),
            .carryin(\spi0.n10698 ),
            .carryout(\spi0.n10699 ),
            .clk(N__97363),
            .ce(N__52945),
            .sr(N__53032));
    defparam \spi0.counter_1109__i6_LC_11_18_6 .C_ON=1'b1;
    defparam \spi0.counter_1109__i6_LC_11_18_6 .SEQ_MODE=4'b1000;
    defparam \spi0.counter_1109__i6_LC_11_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.counter_1109__i6_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__51024),
            .in2(N__86661),
            .in3(N__47527),
            .lcout(\spi0.counter_6 ),
            .ltout(),
            .carryin(\spi0.n10699 ),
            .carryout(\spi0.n10700 ),
            .clk(N__97363),
            .ce(N__52945),
            .sr(N__53032));
    defparam \spi0.counter_1109__i7_LC_11_18_7 .C_ON=1'b1;
    defparam \spi0.counter_1109__i7_LC_11_18_7 .SEQ_MODE=4'b1000;
    defparam \spi0.counter_1109__i7_LC_11_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.counter_1109__i7_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__51012),
            .in2(N__86658),
            .in3(N__47524),
            .lcout(\spi0.counter_7 ),
            .ltout(),
            .carryin(\spi0.n10700 ),
            .carryout(\spi0.n10701 ),
            .clk(N__97363),
            .ce(N__52945),
            .sr(N__53032));
    defparam \spi0.counter_1109__i8_LC_11_19_0 .C_ON=1'b1;
    defparam \spi0.counter_1109__i8_LC_11_19_0 .SEQ_MODE=4'b1001;
    defparam \spi0.counter_1109__i8_LC_11_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.counter_1109__i8_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__51036),
            .in2(N__86662),
            .in3(N__47521),
            .lcout(\spi0.counter_8 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\spi0.n10702 ),
            .clk(N__97371),
            .ce(N__52938),
            .sr(N__53031));
    defparam \spi0.counter_1109__i9_LC_11_19_1 .C_ON=1'b0;
    defparam \spi0.counter_1109__i9_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \spi0.counter_1109__i9_LC_11_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi0.counter_1109__i9_LC_11_19_1  (
            .in0(N__51051),
            .in1(N__86645),
            .in2(_gnd_net_),
            .in3(N__47746),
            .lcout(\spi0.counter_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97371),
            .ce(N__52938),
            .sr(N__53031));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11939_LC_11_20_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11939_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11939_LC_11_20_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11939_LC_11_20_0  (
            .in0(N__90872),
            .in1(N__47743),
            .in2(N__47725),
            .in3(N__87217),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13748_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13748_bdd_4_lut_LC_11_20_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13748_bdd_4_lut_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13748_bdd_4_lut_LC_11_20_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13748_bdd_4_lut_LC_11_20_1  (
            .in0(N__90870),
            .in1(N__47704),
            .in2(N__47680),
            .in3(N__47677),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13751 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11839_LC_11_20_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11839_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11839_LC_11_20_2 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11839_LC_11_20_2  (
            .in0(N__90871),
            .in1(N__87216),
            .in2(N__47665),
            .in3(N__47638),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13616_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13616_bdd_4_lut_LC_11_20_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13616_bdd_4_lut_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13616_bdd_4_lut_LC_11_20_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13616_bdd_4_lut_LC_11_20_3  (
            .in0(N__90869),
            .in1(N__47620),
            .in2(N__47599),
            .in3(N__47596),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13619_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12423_LC_11_20_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12423_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12423_LC_11_20_4 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12423_LC_11_20_4  (
            .in0(N__85075),
            .in1(N__89906),
            .in2(N__47572),
            .in3(N__47569),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14324_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14324_bdd_4_lut_LC_11_20_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14324_bdd_4_lut_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14324_bdd_4_lut_LC_11_20_5 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14324_bdd_4_lut_LC_11_20_5  (
            .in0(N__47563),
            .in1(N__89905),
            .in2(N__47557),
            .in3(N__47554),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14120_bdd_4_lut_LC_12_1_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14120_bdd_4_lut_LC_12_1_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14120_bdd_4_lut_LC_12_1_0 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14120_bdd_4_lut_LC_12_1_0  (
            .in0(N__51730),
            .in1(N__92625),
            .in2(N__51925),
            .in3(N__47848),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14123_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10697_3_lut_LC_12_1_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10697_3_lut_LC_12_1_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10697_3_lut_LC_12_1_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10697_3_lut_LC_12_1_1  (
            .in0(N__47875),
            .in1(_gnd_net_),
            .in2(N__47899),
            .in3(N__85846),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12058_LC_12_1_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12058_LC_12_1_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12058_LC_12_1_2 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12058_LC_12_1_2  (
            .in0(N__47989),
            .in1(N__92626),
            .in2(N__88588),
            .in3(N__47896),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13886_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13886_bdd_4_lut_LC_12_1_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13886_bdd_4_lut_LC_12_1_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13886_bdd_4_lut_LC_12_1_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13886_bdd_4_lut_LC_12_1_3  (
            .in0(N__92624),
            .in1(N__47833),
            .in2(N__47878),
            .in3(N__47842),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13889 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12248_LC_12_1_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12248_LC_12_1_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12248_LC_12_1_4 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12248_LC_12_1_4  (
            .in0(N__88330),
            .in1(N__47869),
            .in2(N__53161),
            .in3(N__92627),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i524_525_LC_12_1_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i524_525_LC_12_1_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i524_525_LC_12_1_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i524_525_LC_12_1_5  (
            .in0(N__75956),
            .in1(N__47841),
            .in2(_gnd_net_),
            .in3(N__67883),
            .lcout(REG_mem_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93416),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i428_429_LC_12_1_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i428_429_LC_12_1_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i428_429_LC_12_1_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i428_429_LC_12_1_6  (
            .in0(N__47832),
            .in1(N__75957),
            .in2(_gnd_net_),
            .in3(N__72724),
            .lcout(REG_mem_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93416),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10070_3_lut_LC_12_2_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10070_3_lut_LC_12_2_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10070_3_lut_LC_12_2_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10070_3_lut_LC_12_2_0  (
            .in0(N__47824),
            .in1(N__87998),
            .in2(_gnd_net_),
            .in3(N__47812),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11719 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10065_3_lut_LC_12_2_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10065_3_lut_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10065_3_lut_LC_12_2_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10065_3_lut_LC_12_2_1  (
            .in0(N__87997),
            .in1(N__47800),
            .in2(_gnd_net_),
            .in3(N__47787),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13742_bdd_4_lut_LC_12_2_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13742_bdd_4_lut_LC_12_2_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13742_bdd_4_lut_LC_12_2_2 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13742_bdd_4_lut_LC_12_2_2  (
            .in0(N__92616),
            .in1(N__47923),
            .in2(N__47773),
            .in3(N__47752),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i620_621_LC_12_2_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i620_621_LC_12_2_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i620_621_LC_12_2_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i620_621_LC_12_2_3  (
            .in0(N__47988),
            .in1(N__75864),
            .in2(_gnd_net_),
            .in3(N__66415),
            .lcout(REG_mem_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93409),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10656_3_lut_LC_12_2_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10656_3_lut_LC_12_2_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10656_3_lut_LC_12_2_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10656_3_lut_LC_12_2_5  (
            .in0(N__87999),
            .in1(N__47977),
            .in2(_gnd_net_),
            .in3(N__47911),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10064_3_lut_LC_12_2_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10064_3_lut_LC_12_2_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10064_3_lut_LC_12_2_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10064_3_lut_LC_12_2_6  (
            .in0(N__47950),
            .in1(N__87996),
            .in2(_gnd_net_),
            .in3(N__51496),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11713 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2729_2730_LC_12_2_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2729_2730_LC_12_2_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2729_2730_LC_12_2_7 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2729_2730_LC_12_2_7  (
            .in0(N__96664),
            .in1(N__94139),
            .in2(N__58635),
            .in3(N__70719),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93409),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3701_3702_LC_12_3_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3701_3702_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3701_3702_LC_12_3_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3701_3702_LC_12_3_1  (
            .in0(N__51369),
            .in1(N__62780),
            .in2(_gnd_net_),
            .in3(N__59283),
            .lcout(REG_mem_38_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93398),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4499_4500_LC_12_3_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4499_4500_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4499_4500_LC_12_3_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4499_4500_LC_12_3_2  (
            .in0(N__62367),
            .in1(N__47934),
            .in2(_gnd_net_),
            .in3(N__89123),
            .lcout(REG_mem_46_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93398),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2261_2262_LC_12_3_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2261_2262_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2261_2262_LC_12_3_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2261_2262_LC_12_3_3  (
            .in0(N__55962),
            .in1(N__62779),
            .in2(_gnd_net_),
            .in3(N__75064),
            .lcout(REG_mem_23_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93398),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3893_3894_LC_12_3_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3893_3894_LC_12_3_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3893_3894_LC_12_3_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3893_3894_LC_12_3_4  (
            .in0(N__62777),
            .in1(N__47922),
            .in2(_gnd_net_),
            .in3(N__65901),
            .lcout(REG_mem_40_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93398),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4169_4170_LC_12_3_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4169_4170_LC_12_3_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4169_4170_LC_12_3_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4169_4170_LC_12_3_5  (
            .in0(N__51213),
            .in1(N__96783),
            .in2(_gnd_net_),
            .in3(N__68295),
            .lcout(REG_mem_43_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93398),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5333_5334_LC_12_3_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5333_5334_LC_12_3_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5333_5334_LC_12_3_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5333_5334_LC_12_3_6  (
            .in0(N__62778),
            .in1(N__47910),
            .in2(_gnd_net_),
            .in3(N__77232),
            .lcout(REG_mem_55_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93398),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10859_3_lut_LC_12_3_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10859_3_lut_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10859_3_lut_LC_12_3_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10859_3_lut_LC_12_3_7  (
            .in0(N__48160),
            .in1(N__48139),
            .in2(_gnd_net_),
            .in3(N__88008),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10007_3_lut_LC_12_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10007_3_lut_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10007_3_lut_LC_12_4_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10007_3_lut_LC_12_4_0  (
            .in0(N__48106),
            .in1(N__88581),
            .in2(_gnd_net_),
            .in3(N__48121),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i812_813_LC_12_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i812_813_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i812_813_LC_12_4_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i812_813_LC_12_4_1  (
            .in0(N__66648),
            .in1(N__75942),
            .in2(_gnd_net_),
            .in3(N__67336),
            .lcout(REG_mem_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93385),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i521_522_LC_12_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i521_522_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i521_522_LC_12_4_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i521_522_LC_12_4_2  (
            .in0(N__48105),
            .in1(N__96730),
            .in2(_gnd_net_),
            .in3(N__67869),
            .lcout(REG_mem_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93385),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10481_3_lut_LC_12_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10481_3_lut_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10481_3_lut_LC_12_4_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10481_3_lut_LC_12_4_3  (
            .in0(N__88583),
            .in1(N__53647),
            .in2(_gnd_net_),
            .in3(N__48097),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5126_5127_LC_12_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5126_5127_LC_12_4_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5126_5127_LC_12_4_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5126_5127_LC_12_4_4  (
            .in0(N__71457),
            .in1(N__95773),
            .in2(N__48075),
            .in3(N__77003),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93385),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4652_4653_LC_12_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4652_4653_LC_12_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4652_4653_LC_12_4_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4652_4653_LC_12_4_5  (
            .in0(N__48057),
            .in1(N__75941),
            .in2(_gnd_net_),
            .in3(N__75577),
            .lcout(REG_mem_48_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93385),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12238_LC_12_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12238_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12238_LC_12_4_6 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12238_LC_12_4_6  (
            .in0(N__48046),
            .in1(N__90232),
            .in2(N__48031),
            .in3(N__81510),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14078 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10011_3_lut_LC_12_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10011_3_lut_LC_12_4_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10011_3_lut_LC_12_4_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10011_3_lut_LC_12_4_7  (
            .in0(N__88582),
            .in1(N__52012),
            .in2(_gnd_net_),
            .in3(N__48001),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11660 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4853_4854_LC_12_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4853_4854_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4853_4854_LC_12_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4853_4854_LC_12_5_0  (
            .in0(N__48300),
            .in1(N__62799),
            .in2(_gnd_net_),
            .in3(N__73032),
            .lcout(REG_mem_50_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12388_LC_12_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12388_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12388_LC_12_5_1 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12388_LC_12_5_1  (
            .in0(N__92449),
            .in1(N__51744),
            .in2(N__48244),
            .in3(N__87666),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2165_2166_LC_12_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2165_2166_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2165_2166_LC_12_5_2 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2165_2166_LC_12_5_2  (
            .in0(N__62797),
            .in1(N__95685),
            .in2(N__55947),
            .in3(N__76345),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2069_2070_LC_12_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2069_2070_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2069_2070_LC_12_5_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2069_2070_LC_12_5_3  (
            .in0(N__95683),
            .in1(N__62798),
            .in2(N__55926),
            .in3(N__76943),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5141_5142_LC_12_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5141_5142_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5141_5142_LC_12_5_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5141_5142_LC_12_5_4  (
            .in0(N__76945),
            .in1(N__62800),
            .in2(N__48216),
            .in3(N__95686),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2081_2082_LC_12_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2081_2082_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2081_2082_LC_12_5_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2081_2082_LC_12_5_5  (
            .in0(N__95684),
            .in1(N__56511),
            .in2(N__48199),
            .in3(N__76944),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10733_3_lut_LC_12_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10733_3_lut_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10733_3_lut_LC_12_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10733_3_lut_LC_12_5_6  (
            .in0(N__87665),
            .in1(N__48198),
            .in2(_gnd_net_),
            .in3(N__48171),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1985_1986_LC_12_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1985_1986_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1985_1986_LC_12_5_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1985_1986_LC_12_5_7  (
            .in0(N__95682),
            .in1(N__56510),
            .in2(N__48172),
            .in3(N__77464),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93372),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i824_825_LC_12_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i824_825_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i824_825_LC_12_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i824_825_LC_12_6_0  (
            .in0(N__70164),
            .in1(N__96315),
            .in2(_gnd_net_),
            .in3(N__67340),
            .lcout(REG_mem_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93359),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10646_3_lut_LC_12_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10646_3_lut_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10646_3_lut_LC_12_6_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10646_3_lut_LC_12_6_1  (
            .in0(N__48271),
            .in1(N__88301),
            .in2(_gnd_net_),
            .in3(N__48346),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11495_LC_12_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11495_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11495_LC_12_6_2 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11495_LC_12_6_2  (
            .in0(N__85823),
            .in1(N__92448),
            .in2(N__48334),
            .in3(N__48322),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13214_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13214_bdd_4_lut_LC_12_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13214_bdd_4_lut_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13214_bdd_4_lut_LC_12_6_3 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13214_bdd_4_lut_LC_12_6_3  (
            .in0(N__48313),
            .in1(N__85822),
            .in2(N__48307),
            .in3(N__48277),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4949_4950_LC_12_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4949_4950_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4949_4950_LC_12_6_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4949_4950_LC_12_6_4  (
            .in0(N__62823),
            .in1(N__48288),
            .in2(_gnd_net_),
            .in3(N__72243),
            .lcout(REG_mem_51_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93359),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10647_3_lut_LC_12_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10647_3_lut_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10647_3_lut_LC_12_6_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10647_3_lut_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__88302),
            .in2(N__48304),
            .in3(N__48289),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4661_4662_LC_12_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4661_4662_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4661_4662_LC_12_6_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4661_4662_LC_12_6_6  (
            .in0(N__62822),
            .in1(N__48270),
            .in2(_gnd_net_),
            .in3(N__75567),
            .lcout(REG_mem_48_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93359),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10113_3_lut_LC_12_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10113_3_lut_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10113_3_lut_LC_12_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10113_3_lut_LC_12_6_7  (
            .in0(N__48373),
            .in1(N__51685),
            .in2(_gnd_net_),
            .in3(N__88300),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11762 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3611_3612_LC_12_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3611_3612_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3611_3612_LC_12_7_0 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3611_3612_LC_12_7_0  (
            .in0(N__63685),
            .in1(_gnd_net_),
            .in2(N__48418),
            .in3(N__63526),
            .lcout(REG_mem_37_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12033_LC_12_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12033_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12033_LC_12_7_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12033_LC_12_7_1  (
            .in0(N__92040),
            .in1(N__88619),
            .in2(N__48262),
            .in3(N__51646),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13862_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13862_bdd_4_lut_LC_12_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13862_bdd_4_lut_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13862_bdd_4_lut_LC_12_7_2 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13862_bdd_4_lut_LC_12_7_2  (
            .in0(N__48417),
            .in1(N__48403),
            .in2(N__48406),
            .in3(N__92039),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3515_3516_LC_12_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3515_3516_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3515_3516_LC_12_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3515_3516_LC_12_7_3  (
            .in0(N__63525),
            .in1(N__48402),
            .in2(_gnd_net_),
            .in3(N__54082),
            .lcout(REG_mem_36_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11869_LC_12_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11869_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11869_LC_12_7_4 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11869_LC_12_7_4  (
            .in0(N__85721),
            .in1(N__48391),
            .in2(N__51874),
            .in3(N__92041),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i710_711_LC_12_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i710_711_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i710_711_LC_12_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i710_711_LC_12_7_5  (
            .in0(N__48372),
            .in1(N__71600),
            .in2(_gnd_net_),
            .in3(N__89642),
            .lcout(REG_mem_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4274_4275_LC_12_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4274_4275_LC_12_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4274_4275_LC_12_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4274_4275_LC_12_7_6  (
            .in0(N__57024),
            .in1(N__76703),
            .in2(_gnd_net_),
            .in3(N__71739),
            .lcout(REG_mem_44_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3593_3594_LC_12_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3593_3594_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3593_3594_LC_12_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3593_3594_LC_12_7_7  (
            .in0(N__96731),
            .in1(N__53208),
            .in2(_gnd_net_),
            .in3(N__63684),
            .lcout(REG_mem_37_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93344),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1397_1398_LC_12_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1397_1398_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1397_1398_LC_12_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1397_1398_LC_12_8_0  (
            .in0(N__62821),
            .in1(N__58752),
            .in2(_gnd_net_),
            .in3(N__74679),
            .lcout(REG_mem_14_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i518_519_LC_12_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i518_519_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i518_519_LC_12_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i518_519_LC_12_8_1  (
            .in0(N__51885),
            .in1(N__71545),
            .in2(_gnd_net_),
            .in3(N__67800),
            .lcout(REG_mem_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3881_3882_LC_12_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3881_3882_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3881_3882_LC_12_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3881_3882_LC_12_8_2  (
            .in0(N__51414),
            .in1(N__96733),
            .in2(_gnd_net_),
            .in3(N__65876),
            .lcout(REG_mem_40_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1409_1410_LC_12_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1409_1410_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1409_1410_LC_12_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1409_1410_LC_12_8_3  (
            .in0(N__74680),
            .in1(N__48357),
            .in2(_gnd_net_),
            .in3(N__56508),
            .lcout(REG_mem_14_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3689_3690_LC_12_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3689_3690_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3689_3690_LC_12_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3689_3690_LC_12_8_4  (
            .in0(N__53571),
            .in1(N__96732),
            .in2(_gnd_net_),
            .in3(N__59206),
            .lcout(REG_mem_38_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3590_3591_LC_12_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3590_3591_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3590_3591_LC_12_8_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3590_3591_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(N__71544),
            .in2(N__53790),
            .in3(N__63648),
            .lcout(REG_mem_37_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i923_924_LC_12_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i923_924_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i923_924_LC_12_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i923_924_LC_12_8_6  (
            .in0(N__63527),
            .in1(N__48462),
            .in2(_gnd_net_),
            .in3(N__67133),
            .lcout(REG_mem_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1313_1314_LC_12_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1313_1314_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1313_1314_LC_12_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1313_1314_LC_12_8_7  (
            .in0(N__48447),
            .in1(N__56507),
            .in2(_gnd_net_),
            .in3(N__70079),
            .lcout(REG_mem_13_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93331),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i59_60_LC_12_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i59_60_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i59_60_LC_12_9_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i59_60_LC_12_9_0  (
            .in0(N__63540),
            .in1(N__94101),
            .in2(N__54252),
            .in3(N__82817),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1793_1794_LC_12_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1793_1794_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1793_1794_LC_12_9_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1793_1794_LC_12_9_1  (
            .in0(N__48429),
            .in1(N__56509),
            .in2(_gnd_net_),
            .in3(N__67490),
            .lcout(REG_mem_18_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3692_3693_LC_12_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3692_3693_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3692_3693_LC_12_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3692_3693_LC_12_9_2  (
            .in0(N__61935),
            .in1(N__75987),
            .in2(_gnd_net_),
            .in3(N__59199),
            .lcout(REG_mem_38_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i443_444_LC_12_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i443_444_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i443_444_LC_12_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i443_444_LC_12_9_3  (
            .in0(N__51951),
            .in1(N__63541),
            .in2(_gnd_net_),
            .in3(N__72720),
            .lcout(REG_mem_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5810_5811_LC_12_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5810_5811_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5810_5811_LC_12_9_4 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5810_5811_LC_12_9_4  (
            .in0(N__59907),
            .in1(N__94100),
            .in2(N__70714),
            .in3(N__76761),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i539_540_LC_12_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i539_540_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i539_540_LC_12_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i539_540_LC_12_9_5  (
            .in0(N__51936),
            .in1(N__63542),
            .in2(_gnd_net_),
            .in3(N__67798),
            .lcout(REG_mem_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4370_4371_LC_12_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4370_4371_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4370_4371_LC_12_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4370_4371_LC_12_9_6  (
            .in0(N__57042),
            .in1(N__76760),
            .in2(_gnd_net_),
            .in3(N__71809),
            .lcout(REG_mem_45_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i635_636_LC_12_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i635_636_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i635_636_LC_12_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i635_636_LC_12_9_7  (
            .in0(N__51963),
            .in1(N__63543),
            .in2(_gnd_net_),
            .in3(N__66348),
            .lcout(REG_mem_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93318),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5429_5430_LC_12_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5429_5430_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5429_5430_LC_12_10_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5429_5430_LC_12_10_0  (
            .in0(N__62855),
            .in1(N__93811),
            .in2(N__53415),
            .in3(N__95997),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93291),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1523_1524_LC_12_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1523_1524_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1523_1524_LC_12_10_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1523_1524_LC_12_10_1  (
            .in0(N__48909),
            .in1(N__63952),
            .in2(_gnd_net_),
            .in3(N__62413),
            .lcout(REG_mem_15_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93291),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3602_3603_LC_12_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3602_3603_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3602_3603_LC_12_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3602_3603_LC_12_10_2  (
            .in0(N__56940),
            .in1(N__76753),
            .in2(_gnd_net_),
            .in3(N__63649),
            .lcout(REG_mem_37_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93291),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4556_4557_LC_12_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4556_4557_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4556_4557_LC_12_10_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4556_4557_LC_12_10_3  (
            .in0(N__75986),
            .in1(N__56679),
            .in2(_gnd_net_),
            .in3(N__66181),
            .lcout(REG_mem_47_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93291),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4082_4083_LC_12_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4082_4083_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4082_4083_LC_12_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4082_4083_LC_12_10_4  (
            .in0(N__57003),
            .in1(N__76754),
            .in2(_gnd_net_),
            .in3(N__68034),
            .lcout(REG_mem_42_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93291),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5822_5823_LC_12_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5822_5823_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5822_5823_LC_12_10_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5822_5823_LC_12_10_5  (
            .in0(N__70662),
            .in1(N__67557),
            .in2(N__94140),
            .in3(N__89515),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93291),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4580_4581_LC_12_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4580_4581_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4580_4581_LC_12_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4580_4581_LC_12_10_6  (
            .in0(N__66182),
            .in1(N__48489),
            .in2(_gnd_net_),
            .in3(N__48891),
            .lcout(REG_mem_47_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93291),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5906_5907_LC_12_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5906_5907_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5906_5907_LC_12_10_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5906_5907_LC_12_10_7  (
            .in0(N__93810),
            .in1(N__59925),
            .in2(N__76762),
            .in3(N__70915),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93291),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i5_LC_12_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i5_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i5_LC_12_11_0 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i5_LC_12_11_0  (
            .in0(N__49270),
            .in1(N__93805),
            .in2(N__73475),
            .in3(N__49149),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93319),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1490_1491_LC_12_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1490_1491_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1490_1491_LC_12_11_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1490_1491_LC_12_11_1  (
            .in0(N__76745),
            .in1(N__52287),
            .in2(_gnd_net_),
            .in3(N__63955),
            .lcout(REG_mem_15_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93319),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i0_LC_12_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i0_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i0_LC_12_11_2 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i0_LC_12_11_2  (
            .in0(N__48938),
            .in1(N__49006),
            .in2(N__73473),
            .in3(N__49150),
            .lcout(wr_addr_r_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93319),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1487_1488_LC_12_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1487_1488_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1487_1488_LC_12_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1487_1488_LC_12_11_3  (
            .in0(N__49161),
            .in1(N__61221),
            .in2(_gnd_net_),
            .in3(N__63954),
            .lcout(REG_mem_15_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93319),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i3_LC_12_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i3_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i3_LC_12_11_4 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i3_LC_12_11_4  (
            .in0(N__49702),
            .in1(N__49619),
            .in2(N__73474),
            .in3(N__49148),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93319),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i2_LC_12_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i2_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i2_LC_12_11_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i2_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__73436),
            .in2(_gnd_net_),
            .in3(N__49072),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93319),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i4_LC_12_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i4_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i4_LC_12_11_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r__i4_LC_12_11_6  (
            .in0(N__73440),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49047),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93319),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i251_252_LC_12_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i251_252_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i251_252_LC_12_11_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i251_252_LC_12_11_7  (
            .in0(N__93804),
            .in1(N__63539),
            .in2(N__54291),
            .in3(N__80508),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93319),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_2_lut_LC_12_12_0 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_2_lut_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_2_lut_LC_12_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_2_lut_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__48982),
            .in2(_gnd_net_),
            .in3(N__50167),
            .lcout(wr_addr_p1_w_0),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10631 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_3_lut_LC_12_12_1 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_3_lut_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_3_lut_LC_12_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_3_lut_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__50156),
            .in2(_gnd_net_),
            .in3(N__50059),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_1 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10631 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10632 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_4_lut_LC_12_12_2 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_4_lut_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_4_lut_LC_12_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_4_lut_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__49941),
            .in2(_gnd_net_),
            .in3(N__49888),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_2 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10632 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10633 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_5_lut_LC_12_12_3 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_5_lut_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_5_lut_LC_12_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_5_lut_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__49679),
            .in2(_gnd_net_),
            .in3(N__49600),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_3 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10633 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10634 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_6_lut_LC_12_12_4 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_6_lut_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_6_lut_LC_12_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_6_lut_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__49341),
            .in2(_gnd_net_),
            .in3(N__49279),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_4 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10634 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10635 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_7_lut_LC_12_12_5 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_7_lut_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_7_lut_LC_12_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_7_lut_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__93618),
            .in2(_gnd_net_),
            .in3(N__49246),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_p1_w_5 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10635 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10636 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_8_lut_LC_12_12_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_8_lut_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_8_lut_LC_12_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_141_8_lut_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__52434),
            .in2(_gnd_net_),
            .in3(N__49243),
            .lcout(wr_addr_p1_w_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i11_LC_12_13_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i11_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i11_LC_12_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i11_LC_12_13_0  (
            .in0(N__81050),
            .in1(N__49222),
            .in2(_gnd_net_),
            .in3(N__49207),
            .lcout(REG_out_raw_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97346),
            .ce(N__80816),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12428_LC_12_13_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12428_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12428_LC_12_13_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12428_LC_12_13_1  (
            .in0(N__49189),
            .in1(N__81056),
            .in2(N__49180),
            .in3(N__81305),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14318_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i12_LC_12_13_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i12_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i12_LC_12_13_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i12_LC_12_13_2  (
            .in0(N__81051),
            .in1(N__50344),
            .in2(N__50326),
            .in3(N__50323),
            .lcout(REG_out_raw_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97346),
            .ce(N__80816),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i2_LC_12_13_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i2_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i2_LC_12_13_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i2_LC_12_13_3  (
            .in0(N__53503),
            .in1(N__81055),
            .in2(_gnd_net_),
            .in3(N__51280),
            .lcout(REG_out_raw_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97346),
            .ce(N__80816),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i16_LC_12_13_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i16_LC_12_13_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i16_LC_12_13_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i16_LC_12_13_4  (
            .in0(N__81053),
            .in1(_gnd_net_),
            .in2(N__50308),
            .in3(N__50287),
            .lcout(REG_out_raw_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97346),
            .ce(N__80816),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i1_LC_12_13_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i1_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i1_LC_12_13_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i1_LC_12_13_5  (
            .in0(N__50275),
            .in1(N__50263),
            .in2(_gnd_net_),
            .in3(N__81054),
            .lcout(REG_out_raw_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97346),
            .ce(N__80816),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i10_LC_12_13_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i10_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i10_LC_12_13_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i10_LC_12_13_6  (
            .in0(N__81049),
            .in1(N__50248),
            .in2(_gnd_net_),
            .in3(N__50230),
            .lcout(REG_out_raw_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97346),
            .ce(N__80816),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i15_LC_12_13_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i15_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i15_LC_12_13_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i15_LC_12_13_7  (
            .in0(N__50218),
            .in1(N__50200),
            .in2(_gnd_net_),
            .in3(N__81052),
            .lcout(REG_out_raw_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97346),
            .ce(N__80816),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i1_LC_12_14_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i1_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i1_LC_12_14_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i1_LC_12_14_0  (
            .in0(N__73419),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50188),
            .lcout(wp_sync1_r_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97348),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i10_LC_12_14_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i10_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i10_LC_12_14_1 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i10_LC_12_14_1  (
            .in0(N__50173),
            .in1(N__80729),
            .in2(N__58101),
            .in3(N__73418),
            .lcout(fifo_data_out_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97348),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i4_LC_12_14_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i4_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i4_LC_12_14_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i4_LC_12_14_2  (
            .in0(N__73424),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50392),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97348),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i4_LC_12_14_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i4_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i4_LC_12_14_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i4_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__50404),
            .in2(_gnd_net_),
            .in3(N__73421),
            .lcout(wp_sync1_r_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97348),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i3_LC_12_14_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i3_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i3_LC_12_14_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i3_LC_12_14_4  (
            .in0(N__73423),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50371),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97348),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i5_LC_12_14_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i5_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i5_LC_12_14_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i5_LC_12_14_5  (
            .in0(N__50353),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73425),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97348),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i3_LC_12_14_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i3_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i3_LC_12_14_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i3_LC_12_14_6  (
            .in0(N__73420),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50386),
            .lcout(wp_sync1_r_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97348),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i5_LC_12_14_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i5_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i5_LC_12_14_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i5_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__50365),
            .in2(_gnd_net_),
            .in3(N__73422),
            .lcout(wp_sync1_r_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97348),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_LC_12_15_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_LC_12_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_LC_12_15_0  (
            .in0(N__52386),
            .in1(N__50532),
            .in2(_gnd_net_),
            .in3(N__50546),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_4 ),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_53_LC_12_15_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_53_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_53_LC_12_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_53_LC_12_15_1  (
            .in0(N__50518),
            .in1(_gnd_net_),
            .in2(N__50347),
            .in3(N__50508),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_143_i1_2_lut_LC_12_15_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_143_i1_2_lut_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_143_i1_2_lut_LC_12_15_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_143_i1_2_lut_LC_12_15_2  (
            .in0(N__52388),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50548),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i2_LC_12_15_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i2_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i2_LC_12_15_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i2_LC_12_15_3  (
            .in0(N__73427),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52342),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97353),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i1_LC_12_15_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i1_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i1_LC_12_15_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i1_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__50587),
            .in2(_gnd_net_),
            .in3(N__73426),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97353),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_47_LC_12_15_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_47_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_47_LC_12_15_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_47_LC_12_15_5  (
            .in0(N__50547),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52387),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n4027 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_4_lut_LC_12_15_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_4_lut_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_4_lut_LC_12_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_4_lut_LC_12_15_6  (
            .in0(N__52385),
            .in1(N__50545),
            .in2(N__50533),
            .in3(N__50517),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_3 ),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_54_LC_12_15_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_54_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_54_LC_12_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_3_lut_adj_54_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__50509),
            .in2(N__50500),
            .in3(N__50497),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_2_lut_LC_12_16_0 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_2_lut_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_2_lut_LC_12_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_2_lut_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__52662),
            .in2(N__50491),
            .in3(N__50476),
            .lcout(rd_sig_diff0_w_0),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10619 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_3_lut_LC_12_16_1 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_3_lut_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_3_lut_LC_12_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_3_lut_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__52633),
            .in2(N__52704),
            .in3(N__50473),
            .lcout(rd_sig_diff0_w_1),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10619 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10620 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_4_lut_LC_12_16_2 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_4_lut_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_4_lut_LC_12_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_4_lut_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__52743),
            .in2(N__50470),
            .in3(N__50452),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_sig_diff0_w_2 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10620 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10621 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_5_lut_LC_12_16_3 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_5_lut_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_5_lut_LC_12_16_3 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_5_lut_LC_12_16_3  (
            .in0(N__50827),
            .in1(N__50436),
            .in2(N__50425),
            .in3(N__50407),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n8 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10621 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10622 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_6_lut_LC_12_16_4 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_6_lut_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_6_lut_LC_12_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_6_lut_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__50649),
            .in2(N__50905),
            .in3(N__50890),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_sig_diff0_w_4 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10622 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10623 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_7_lut_LC_12_16_5 .C_ON=1'b1;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_7_lut_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_7_lut_LC_12_16_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_7_lut_LC_12_16_5  (
            .in0(N__50887),
            .in1(N__50878),
            .in2(N__50863),
            .in3(N__50854),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7 ),
            .ltout(),
            .carryin(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10623 ),
            .carryout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10624 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_8_lut_LC_12_16_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_8_lut_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_8_lut_LC_12_16_6 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_add_2_8_lut_LC_12_16_6  (
            .in0(N__52389),
            .in1(N__50851),
            .in2(N__50839),
            .in3(N__50830),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_4_lut_LC_12_17_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_4_lut_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_4_lut_LC_12_17_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_4_lut_LC_12_17_0  (
            .in0(N__52705),
            .in1(N__52393),
            .in2(N__50821),
            .in3(N__50790),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n8_adj_1157_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6_4_lut_LC_12_17_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6_4_lut_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6_4_lut_LC_12_17_1 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6_4_lut_LC_12_17_1  (
            .in0(N__50754),
            .in1(N__52747),
            .in2(N__50719),
            .in3(N__51094),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n10760 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9797_4_lut_LC_12_17_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9797_4_lut_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9797_4_lut_LC_12_17_2 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9797_4_lut_LC_12_17_2  (
            .in0(N__50656),
            .in1(N__87335),
            .in2(N__81293),
            .in3(N__52669),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9936_3_lut_LC_12_17_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9936_3_lut_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9936_3_lut_LC_12_17_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9936_3_lut_LC_12_17_3  (
            .in0(N__87336),
            .in1(_gnd_net_),
            .in2(N__50716),
            .in3(N__50698),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11585 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_49_LC_12_17_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_49_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_49_LC_12_17_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_49_LC_12_17_4  (
            .in0(N__50655),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50638),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n4025_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5_4_lut_adj_50_LC_12_17_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5_4_lut_adj_50_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5_4_lut_adj_50_LC_12_17_5 .LUT_INIT=16'b1111110111111110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5_4_lut_adj_50_LC_12_17_5  (
            .in0(N__52668),
            .in1(N__50602),
            .in2(N__51133),
            .in3(N__51130),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12_adj_1158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i0_LC_12_17_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i0_LC_12_17_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i0_LC_12_17_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i0_LC_12_17_6  (
            .in0(N__73429),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51070),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97364),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i0_LC_12_17_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i0_LC_12_17_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i0_LC_12_17_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i0_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__51088),
            .in2(_gnd_net_),
            .in3(N__73428),
            .lcout(wp_sync1_r_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97364),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_2_lut_4_lut_adj_37_LC_12_18_0 .C_ON=1'b0;
    defparam \spi0.i1_2_lut_4_lut_adj_37_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_2_lut_4_lut_adj_37_LC_12_18_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \spi0.i1_2_lut_4_lut_adj_37_LC_12_18_0  (
            .in0(N__50999),
            .in1(N__50981),
            .in2(N__50965),
            .in3(N__50936),
            .lcout(\spi0.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i3_4_lut_adj_27_LC_12_18_1 .C_ON=1'b0;
    defparam \spi0.i3_4_lut_adj_27_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \spi0.i3_4_lut_adj_27_LC_12_18_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \spi0.i3_4_lut_adj_27_LC_12_18_1  (
            .in0(N__50983),
            .in1(N__51001),
            .in2(N__50941),
            .in3(N__50963),
            .lcout(\spi0.n11317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i6_4_lut_LC_12_18_2 .C_ON=1'b0;
    defparam \spi0.i6_4_lut_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \spi0.i6_4_lut_LC_12_18_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \spi0.i6_4_lut_LC_12_18_2  (
            .in0(N__51064),
            .in1(N__51052),
            .in2(N__51040),
            .in3(N__51025),
            .lcout(\spi0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_2_lut_adj_29_LC_12_18_3 .C_ON=1'b0;
    defparam \spi0.i1_2_lut_adj_29_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_2_lut_adj_29_LC_12_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \spi0.i1_2_lut_adj_29_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__51013),
            .in2(_gnd_net_),
            .in3(N__52794),
            .lcout(\spi0.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i2_3_lut_adj_28_LC_12_18_4 .C_ON=1'b0;
    defparam \spi0.i2_3_lut_adj_28_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \spi0.i2_3_lut_adj_28_LC_12_18_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \spi0.i2_3_lut_adj_28_LC_12_18_4  (
            .in0(N__51000),
            .in1(N__50982),
            .in2(_gnd_net_),
            .in3(N__50964),
            .lcout(),
            .ltout(\spi0.n3909_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i7_4_lut_LC_12_18_5 .C_ON=1'b0;
    defparam \spi0.i7_4_lut_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \spi0.i7_4_lut_LC_12_18_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \spi0.i7_4_lut_LC_12_18_5  (
            .in0(N__50940),
            .in1(N__50920),
            .in2(N__50914),
            .in3(N__50911),
            .lcout(\spi0.n19 ),
            .ltout(\spi0.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i106_2_lut_LC_12_18_6 .C_ON=1'b0;
    defparam \spi0.i106_2_lut_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \spi0.i106_2_lut_LC_12_18_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \spi0.i106_2_lut_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51190),
            .in3(N__55047),
            .lcout(\spi0.n88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i2318_4_lut_4_lut_LC_12_18_7 .C_ON=1'b0;
    defparam \spi0.i2318_4_lut_4_lut_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \spi0.i2318_4_lut_4_lut_LC_12_18_7 .LUT_INIT=16'b1111001011101111;
    LogicCell40 \spi0.i2318_4_lut_4_lut_LC_12_18_7  (
            .in0(N__55048),
            .in1(N__55251),
            .in2(N__55498),
            .in3(N__55588),
            .lcout(\spi0.n4409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i11041_4_lut_LC_12_19_0 .C_ON=1'b0;
    defparam \spi0.i11041_4_lut_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \spi0.i11041_4_lut_LC_12_19_0 .LUT_INIT=16'b1100000010001100;
    LogicCell40 \spi0.i11041_4_lut_LC_12_19_0  (
            .in0(N__51178),
            .in1(N__55599),
            .in2(N__55252),
            .in3(N__55070),
            .lcout(\spi0.n12566 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i8592_4_lut_LC_12_19_1 .C_ON=1'b0;
    defparam \spi0.i8592_4_lut_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \spi0.i8592_4_lut_LC_12_19_1 .LUT_INIT=16'b1000101011001110;
    LogicCell40 \spi0.i8592_4_lut_LC_12_19_1  (
            .in0(N__55218),
            .in1(N__55483),
            .in2(N__51187),
            .in3(N__55767),
            .lcout(\spi0.n10106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i2_3_lut_4_lut_adj_35_LC_12_19_2 .C_ON=1'b0;
    defparam \spi0.i2_3_lut_4_lut_adj_35_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \spi0.i2_3_lut_4_lut_adj_35_LC_12_19_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \spi0.i2_3_lut_4_lut_adj_35_LC_12_19_2  (
            .in0(N__55482),
            .in1(N__55603),
            .in2(N__55253),
            .in3(N__55072),
            .lcout(\spi0.n11351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i11020_2_lut_4_lut_LC_12_19_3 .C_ON=1'b0;
    defparam \spi0.i11020_2_lut_4_lut_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \spi0.i11020_2_lut_4_lut_LC_12_19_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \spi0.i11020_2_lut_4_lut_LC_12_19_3  (
            .in0(N__55069),
            .in1(N__51177),
            .in2(N__55612),
            .in3(N__55210),
            .lcout(),
            .ltout(\spi0.n12567_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_4_lut_LC_12_19_4 .C_ON=1'b0;
    defparam \spi0.i1_4_lut_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_4_lut_LC_12_19_4 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \spi0.i1_4_lut_LC_12_19_4  (
            .in0(N__55480),
            .in1(N__51169),
            .in2(N__51163),
            .in3(N__52796),
            .lcout(\spi0.SCLK_N_977 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i2_3_lut_4_lut_LC_12_19_5 .C_ON=1'b0;
    defparam \spi0.i2_3_lut_4_lut_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \spi0.i2_3_lut_4_lut_LC_12_19_5 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \spi0.i2_3_lut_4_lut_LC_12_19_5  (
            .in0(N__55071),
            .in1(N__55481),
            .in2(N__55613),
            .in3(N__55214),
            .lcout(),
            .ltout(\spi0.n2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_4_lut_adj_23_LC_12_19_6 .C_ON=1'b0;
    defparam \spi0.i1_4_lut_adj_23_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_4_lut_adj_23_LC_12_19_6 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \spi0.i1_4_lut_adj_23_LC_12_19_6  (
            .in0(N__52818),
            .in1(N__51142),
            .in2(N__51136),
            .in3(N__52797),
            .lcout(n1928),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i11112_3_lut_LC_12_19_7 .C_ON=1'b0;
    defparam \spi0.i11112_3_lut_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \spi0.i11112_3_lut_LC_12_19_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi0.i11112_3_lut_LC_12_19_7  (
            .in0(N__52795),
            .in1(N__51295),
            .in2(_gnd_net_),
            .in3(N__52817),
            .lcout(n4093),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13970_bdd_4_lut_LC_13_1_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13970_bdd_4_lut_LC_13_1_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13970_bdd_4_lut_LC_13_1_0 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13970_bdd_4_lut_LC_13_1_0  (
            .in0(N__51202),
            .in1(N__85848),
            .in2(N__51244),
            .in3(N__51403),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11750 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12208_LC_13_1_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12208_LC_13_1_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12208_LC_13_1_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12208_LC_13_1_1  (
            .in0(N__81289),
            .in1(N__90388),
            .in2(N__58822),
            .in3(N__55654),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13844_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13844_bdd_4_lut_LC_13_1_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13844_bdd_4_lut_LC_13_1_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13844_bdd_4_lut_LC_13_1_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13844_bdd_4_lut_LC_13_1_2  (
            .in0(N__51223),
            .in1(N__81288),
            .in2(N__51289),
            .in3(N__51286),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13847 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12133_LC_13_1_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12133_LC_13_1_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12133_LC_13_1_3 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12133_LC_13_1_3  (
            .in0(N__85850),
            .in1(N__92580),
            .in2(N__51265),
            .in3(N__51250),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13970 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11615_LC_13_1_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11615_LC_13_1_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11615_LC_13_1_4 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11615_LC_13_1_4  (
            .in0(N__53197),
            .in1(N__85849),
            .in2(N__92664),
            .in3(N__53545),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13358_bdd_4_lut_LC_13_1_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13358_bdd_4_lut_LC_13_1_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13358_bdd_4_lut_LC_13_1_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13358_bdd_4_lut_LC_13_1_5  (
            .in0(N__85847),
            .in1(N__51235),
            .in2(N__51226),
            .in3(N__53179),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10056_3_lut_LC_13_1_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10056_3_lut_LC_13_1_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10056_3_lut_LC_13_1_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10056_3_lut_LC_13_1_6  (
            .in0(N__51217),
            .in1(N__53596),
            .in2(_gnd_net_),
            .in3(N__88587),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9840_3_lut_LC_13_2_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9840_3_lut_LC_13_2_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9840_3_lut_LC_13_2_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9840_3_lut_LC_13_2_1  (
            .in0(N__85851),
            .in1(N__51196),
            .in2(_gnd_net_),
            .in3(N__51535),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11489_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14258_bdd_4_lut_LC_13_2_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14258_bdd_4_lut_LC_13_2_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14258_bdd_4_lut_LC_13_2_2 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14258_bdd_4_lut_LC_13_2_2  (
            .in0(N__51331),
            .in1(N__81511),
            .in2(N__51394),
            .in3(N__51376),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12393_LC_13_2_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12393_LC_13_2_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12393_LC_13_2_3 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_12393_LC_13_2_3  (
            .in0(N__81512),
            .in1(N__90387),
            .in2(N__51391),
            .in3(N__53239),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1385_1386_LC_13_2_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1385_1386_LC_13_2_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1385_1386_LC_13_2_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1385_1386_LC_13_2_4  (
            .in0(N__53271),
            .in1(N__96639),
            .in2(_gnd_net_),
            .in3(N__74769),
            .lcout(REG_mem_14_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93417),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10482_3_lut_LC_13_2_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10482_3_lut_LC_13_2_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10482_3_lut_LC_13_2_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10482_3_lut_LC_13_2_5  (
            .in0(N__51370),
            .in1(N__88318),
            .in2(_gnd_net_),
            .in3(N__59131),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12131_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11196_LC_13_2_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11196_LC_13_2_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11196_LC_13_2_6 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11196_LC_13_2_6  (
            .in0(N__91221),
            .in1(N__85853),
            .in2(N__51358),
            .in3(N__51355),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12818_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12818_bdd_4_lut_LC_13_2_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12818_bdd_4_lut_LC_13_2_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12818_bdd_4_lut_LC_13_2_7 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12818_bdd_4_lut_LC_13_2_7  (
            .in0(N__85852),
            .in1(N__51346),
            .in2(N__51334),
            .in3(N__53107),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12821 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9858_3_lut_LC_13_3_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9858_3_lut_LC_13_3_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9858_3_lut_LC_13_3_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9858_3_lut_LC_13_3_0  (
            .in0(N__88321),
            .in1(_gnd_net_),
            .in2(N__51325),
            .in3(N__51673),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11507_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12378_LC_13_3_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12378_LC_13_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12378_LC_13_3_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12378_LC_13_3_1  (
            .in0(N__85827),
            .in1(N__92027),
            .in2(N__51304),
            .in3(N__51301),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9857_3_lut_LC_13_3_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9857_3_lut_LC_13_3_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9857_3_lut_LC_13_3_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9857_3_lut_LC_13_3_2  (
            .in0(N__88320),
            .in1(_gnd_net_),
            .in2(N__53932),
            .in3(N__51901),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10860_3_lut_LC_13_3_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10860_3_lut_LC_13_3_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10860_3_lut_LC_13_3_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10860_3_lut_LC_13_3_3  (
            .in0(N__51477),
            .in1(N__88319),
            .in2(_gnd_net_),
            .in3(N__53137),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12509_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14276_bdd_4_lut_LC_13_3_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14276_bdd_4_lut_LC_13_3_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14276_bdd_4_lut_LC_13_3_4 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14276_bdd_4_lut_LC_13_3_4  (
            .in0(N__51514),
            .in1(N__85826),
            .in2(N__51508),
            .in3(N__51505),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4265_4266_LC_13_3_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4265_4266_LC_13_3_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4265_4266_LC_13_3_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4265_4266_LC_13_3_5  (
            .in0(N__51489),
            .in1(N__96750),
            .in2(_gnd_net_),
            .in3(N__71762),
            .lcout(REG_mem_44_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93410),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2357_2358_LC_13_3_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2357_2358_LC_13_3_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2357_2358_LC_13_3_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2357_2358_LC_13_3_6  (
            .in0(N__62781),
            .in1(N__95762),
            .in2(N__53332),
            .in3(N__96011),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93410),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i245_246_LC_13_3_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i245_246_LC_13_3_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i245_246_LC_13_3_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i245_246_LC_13_3_7  (
            .in0(N__95761),
            .in1(N__62782),
            .in2(N__51478),
            .in3(N__80577),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93410),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2924_2925_LC_13_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2924_2925_LC_13_4_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2924_2925_LC_13_4_0 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2924_2925_LC_13_4_0  (
            .in0(N__95774),
            .in1(N__75919),
            .in2(N__61647),
            .in3(N__77964),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10005_3_lut_LC_13_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10005_3_lut_LC_13_4_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10005_3_lut_LC_13_4_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10005_3_lut_LC_13_4_1  (
            .in0(N__51466),
            .in1(N__88584),
            .in2(_gnd_net_),
            .in3(N__51448),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11654 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10055_3_lut_LC_13_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10055_3_lut_LC_13_4_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10055_3_lut_LC_13_4_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10055_3_lut_LC_13_4_2  (
            .in0(N__88586),
            .in1(_gnd_net_),
            .in2(N__51424),
            .in3(N__53872),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2453_2454_LC_13_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2453_2454_LC_13_4_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2453_2454_LC_13_4_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2453_2454_LC_13_4_3  (
            .in0(N__62790),
            .in1(N__95775),
            .in2(N__53347),
            .in3(N__97049),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2456_2457_LC_13_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2456_2457_LC_13_4_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2456_2457_LC_13_4_4 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2456_2457_LC_13_4_4  (
            .in0(N__97048),
            .in1(N__96157),
            .in2(N__95779),
            .in3(N__69807),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i809_810_LC_13_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i809_810_LC_13_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i809_810_LC_13_4_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i809_810_LC_13_4_5  (
            .in0(N__51633),
            .in1(N__96740),
            .in2(_gnd_net_),
            .in3(N__67337),
            .lcout(REG_mem_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3497_3498_LC_13_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3497_3498_LC_13_4_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3497_3498_LC_13_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3497_3498_LC_13_4_6  (
            .in0(N__96739),
            .in1(N__53229),
            .in2(_gnd_net_),
            .in3(N__54108),
            .lcout(REG_mem_36_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93399),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10010_3_lut_LC_13_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10010_3_lut_LC_13_4_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10010_3_lut_LC_13_4_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10010_3_lut_LC_13_4_7  (
            .in0(N__51634),
            .in1(N__88585),
            .in2(_gnd_net_),
            .in3(N__51622),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14288_bdd_4_lut_LC_13_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14288_bdd_4_lut_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14288_bdd_4_lut_LC_13_5_0 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14288_bdd_4_lut_LC_13_5_0  (
            .in0(N__92352),
            .in1(N__51705),
            .in2(N__51598),
            .in3(N__51525),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12030 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13856_bdd_4_lut_LC_13_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13856_bdd_4_lut_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13856_bdd_4_lut_LC_13_5_1 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13856_bdd_4_lut_LC_13_5_1  (
            .in0(N__51589),
            .in1(N__92351),
            .in2(N__51865),
            .in3(N__51781),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13859 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13574_bdd_4_lut_LC_13_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13574_bdd_4_lut_LC_13_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13574_bdd_4_lut_LC_13_5_2 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13574_bdd_4_lut_LC_13_5_2  (
            .in0(N__92350),
            .in1(N__51691),
            .in2(N__51559),
            .in3(N__53467),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3116_3117_LC_13_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3116_3117_LC_13_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3116_3117_LC_13_5_3 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3116_3117_LC_13_5_3  (
            .in0(N__75928),
            .in1(N__94582),
            .in2(N__51526),
            .in3(N__82921),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93386),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2156_2157_LC_13_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2156_2157_LC_13_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2156_2157_LC_13_5_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2156_2157_LC_13_5_4  (
            .in0(N__94581),
            .in1(N__75931),
            .in2(N__58992),
            .in3(N__76346),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93386),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3404_3405_LC_13_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3404_3405_LC_13_5_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3404_3405_LC_13_5_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3404_3405_LC_13_5_5  (
            .in0(N__75929),
            .in1(N__94583),
            .in2(N__51748),
            .in3(N__83361),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93386),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i140_141_LC_13_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i140_141_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i140_141_LC_13_5_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i140_141_LC_13_5_6  (
            .in0(N__94580),
            .in1(N__75930),
            .in2(N__51729),
            .in3(N__80283),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93386),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5528_5529_LC_13_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5528_5529_LC_13_5_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5528_5529_LC_13_5_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5528_5529_LC_13_5_7  (
            .in0(N__96229),
            .in1(N__94584),
            .in2(N__76056),
            .in3(N__96990),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93386),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3212_3213_LC_13_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3212_3213_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3212_3213_LC_13_6_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3212_3213_LC_13_6_0  (
            .in0(N__75971),
            .in1(N__94579),
            .in2(N__51706),
            .in3(N__80232),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93373),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11799_LC_13_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11799_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11799_LC_13_6_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11799_LC_13_6_1  (
            .in0(N__91662),
            .in1(N__88303),
            .in2(N__51658),
            .in3(N__51826),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13574 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i614_615_LC_13_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i614_615_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i614_615_LC_13_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i614_615_LC_13_6_2  (
            .in0(N__71596),
            .in1(N__51684),
            .in2(_gnd_net_),
            .in3(N__66413),
            .lcout(REG_mem_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93373),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1109_1110_LC_13_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1109_1110_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1109_1110_LC_13_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1109_1110_LC_13_6_3  (
            .in0(N__56109),
            .in1(N__62843),
            .in2(_gnd_net_),
            .in3(N__66804),
            .lcout(REG_mem_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93373),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i629_630_LC_13_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i629_630_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i629_630_LC_13_6_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i629_630_LC_13_6_4  (
            .in0(N__62842),
            .in1(N__51669),
            .in2(_gnd_net_),
            .in3(N__66414),
            .lcout(REG_mem_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93373),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4565_4566_LC_13_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4565_4566_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4565_4566_LC_13_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4565_4566_LC_13_6_5  (
            .in0(N__51654),
            .in1(N__62844),
            .in2(_gnd_net_),
            .in3(N__66270),
            .lcout(REG_mem_47_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93373),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3707_3708_LC_13_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3707_3708_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3707_3708_LC_13_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3707_3708_LC_13_6_6  (
            .in0(N__51645),
            .in1(N__63258),
            .in2(_gnd_net_),
            .in3(N__59280),
            .lcout(REG_mem_38_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93373),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i44_45_LC_13_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i44_45_LC_13_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i44_45_LC_13_6_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i44_45_LC_13_6_7  (
            .in0(N__94578),
            .in1(N__75972),
            .in2(N__51918),
            .in3(N__82898),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93373),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i998_999_LC_13_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i998_999_LC_13_7_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i998_999_LC_13_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i998_999_LC_13_7_0  (
            .in0(N__71602),
            .in1(N__51792),
            .in2(_gnd_net_),
            .in3(N__66985),
            .lcout(REG_mem_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i533_534_LC_13_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i533_534_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i533_534_LC_13_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i533_534_LC_13_7_1  (
            .in0(N__51897),
            .in1(N__62835),
            .in2(_gnd_net_),
            .in3(N__67868),
            .lcout(REG_mem_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10112_3_lut_LC_13_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10112_3_lut_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10112_3_lut_LC_13_7_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10112_3_lut_LC_13_7_2  (
            .in0(N__53701),
            .in1(N__88473),
            .in2(_gnd_net_),
            .in3(N__51886),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i902_903_LC_13_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i902_903_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i902_903_LC_13_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i902_903_LC_13_7_3  (
            .in0(N__51858),
            .in1(N__71601),
            .in2(_gnd_net_),
            .in3(N__67163),
            .lcout(REG_mem_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1907_1908_LC_13_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1907_1908_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1907_1908_LC_13_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1907_1908_LC_13_7_4  (
            .in0(N__62444),
            .in1(N__51837),
            .in2(_gnd_net_),
            .in3(N__72065),
            .lcout(REG_mem_19_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4469_4470_LC_13_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4469_4470_LC_13_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4469_4470_LC_13_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4469_4470_LC_13_7_5  (
            .in0(N__51825),
            .in1(N__62834),
            .in2(_gnd_net_),
            .in3(N__89102),
            .lcout(REG_mem_46_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12028_LC_13_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12028_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12028_LC_13_7_6 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12028_LC_13_7_6  (
            .in0(N__51814),
            .in1(N__91242),
            .in2(N__51796),
            .in3(N__88474),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13856 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4181_4182_LC_13_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4181_4182_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4181_4182_LC_13_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4181_4182_LC_13_7_7  (
            .in0(N__51759),
            .in1(N__62833),
            .in2(_gnd_net_),
            .in3(N__68274),
            .lcout(REG_mem_43_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93360),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13982_bdd_4_lut_LC_13_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13982_bdd_4_lut_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13982_bdd_4_lut_LC_13_8_0 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13982_bdd_4_lut_LC_13_8_0  (
            .in0(N__56782),
            .in1(N__91239),
            .in2(N__52033),
            .in3(N__51994),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1097_1098_LC_13_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1097_1098_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1097_1098_LC_13_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1097_1098_LC_13_8_1  (
            .in0(N__52005),
            .in1(N__96778),
            .in2(_gnd_net_),
            .in3(N__66803),
            .lcout(REG_mem_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93345),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3890_3891_LC_13_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3890_3891_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3890_3891_LC_13_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3890_3891_LC_13_8_2  (
            .in0(N__56982),
            .in1(N__76707),
            .in2(_gnd_net_),
            .in3(N__65877),
            .lcout(REG_mem_40_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93345),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1595_1596_LC_13_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1595_1596_LC_13_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1595_1596_LC_13_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1595_1596_LC_13_8_3  (
            .in0(N__51993),
            .in1(N__63528),
            .in2(_gnd_net_),
            .in3(N__65676),
            .lcout(REG_mem_16_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93345),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4658_4659_LC_13_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4658_4659_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4658_4659_LC_13_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4658_4659_LC_13_8_4  (
            .in0(N__63018),
            .in1(N__76708),
            .in2(_gnd_net_),
            .in3(N__75559),
            .lcout(REG_mem_48_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93345),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12213_LC_13_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12213_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12213_LC_13_8_5 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12213_LC_13_8_5  (
            .in0(N__91241),
            .in1(N__87977),
            .in2(N__51985),
            .in3(N__51964),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14072_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14072_bdd_4_lut_LC_13_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14072_bdd_4_lut_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14072_bdd_4_lut_LC_13_8_6 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14072_bdd_4_lut_LC_13_8_6  (
            .in0(N__51952),
            .in1(N__91240),
            .in2(N__51940),
            .in3(N__51937),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1883_1884_LC_13_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1883_1884_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1883_1884_LC_13_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1883_1884_LC_13_8_7  (
            .in0(N__56793),
            .in1(N__63529),
            .in2(_gnd_net_),
            .in3(N__72085),
            .lcout(REG_mem_19_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93345),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13718_bdd_4_lut_LC_13_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13718_bdd_4_lut_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13718_bdd_4_lut_LC_13_9_0 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13718_bdd_4_lut_LC_13_9_0  (
            .in0(N__52105),
            .in1(N__91238),
            .in2(N__52096),
            .in3(N__59824),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5033_5034_LC_13_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5033_5034_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5033_5034_LC_13_9_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5033_5034_LC_13_9_1  (
            .in0(N__94121),
            .in1(N__96806),
            .in2(N__52122),
            .in3(N__77418),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5339_5340_LC_13_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5339_5340_LC_13_9_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5339_5340_LC_13_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5339_5340_LC_13_9_2  (
            .in0(N__59835),
            .in1(N__63341),
            .in2(_gnd_net_),
            .in3(N__77210),
            .lcout(REG_mem_55_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5147_5148_LC_13_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5147_5148_LC_13_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5147_5148_LC_13_9_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5147_5148_LC_13_9_3  (
            .in0(N__94122),
            .in1(N__52104),
            .in2(N__63441),
            .in3(N__76927),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5051_5052_LC_13_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5051_5052_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5051_5052_LC_13_9_4 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5051_5052_LC_13_9_4  (
            .in0(N__52092),
            .in1(N__63343),
            .in2(N__95009),
            .in3(N__77417),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3518_3519_LC_13_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3518_3519_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3518_3519_LC_13_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3518_3519_LC_13_9_5  (
            .in0(N__67032),
            .in1(N__89526),
            .in2(_gnd_net_),
            .in3(N__54080),
            .lcout(REG_mem_36_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1979_1980_LC_13_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1979_1980_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1979_1980_LC_13_9_6 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1979_1980_LC_13_9_6  (
            .in0(N__54186),
            .in1(N__63342),
            .in2(N__95008),
            .in3(N__77416),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i347_348_LC_13_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i347_348_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i347_348_LC_13_9_7 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i347_348_LC_13_9_7  (
            .in0(N__94120),
            .in1(N__54270),
            .in2(N__63440),
            .in3(N__83291),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93332),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13478_bdd_4_lut_LC_13_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13478_bdd_4_lut_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13478_bdd_4_lut_LC_13_10_0 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13478_bdd_4_lut_LC_13_10_0  (
            .in0(N__90252),
            .in1(N__52084),
            .in2(N__54175),
            .in3(N__52069),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12282 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13316_bdd_4_lut_LC_13_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13316_bdd_4_lut_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13316_bdd_4_lut_LC_13_10_1 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13316_bdd_4_lut_LC_13_10_1  (
            .in0(N__52060),
            .in1(N__90250),
            .in2(N__52045),
            .in3(N__59437),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12330_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_11680_LC_13_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_11680_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_11680_LC_13_10_2 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_11680_LC_13_10_2  (
            .in0(N__81063),
            .in1(N__81239),
            .in2(N__52258),
            .in3(N__52228),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13466_bdd_4_lut_LC_13_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13466_bdd_4_lut_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13466_bdd_4_lut_LC_13_10_3 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13466_bdd_4_lut_LC_13_10_3  (
            .in0(N__52165),
            .in1(N__90251),
            .in2(N__52255),
            .in3(N__52240),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13580_bdd_4_lut_LC_13_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13580_bdd_4_lut_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13580_bdd_4_lut_LC_13_10_4 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13580_bdd_4_lut_LC_13_10_4  (
            .in0(N__90253),
            .in1(N__52222),
            .in2(N__52207),
            .in3(N__54235),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12258_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i8_LC_13_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i8_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i8_LC_13_10_5 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i8_LC_13_10_5  (
            .in0(N__52195),
            .in1(N__81062),
            .in2(N__52189),
            .in3(N__52186),
            .lcout(REG_out_raw_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97347),
            .ce(N__80854),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3227_3228_LC_13_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3227_3228_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3227_3228_LC_13_11_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3227_3228_LC_13_11_0  (
            .in0(N__80201),
            .in1(N__63449),
            .in2(N__52180),
            .in3(N__93809),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12048_LC_13_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12048_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12048_LC_13_11_1 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12048_LC_13_11_1  (
            .in0(N__52299),
            .in1(N__52147),
            .in2(N__91237),
            .in3(N__88243),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13880_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13880_bdd_4_lut_LC_13_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13880_bdd_4_lut_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13880_bdd_4_lut_LC_13_11_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13880_bdd_4_lut_LC_13_11_2  (
            .in0(N__52179),
            .in1(N__90878),
            .in2(N__52168),
            .in3(N__52158),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3131_3132_LC_13_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3131_3132_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3131_3132_LC_13_11_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3131_3132_LC_13_11_3  (
            .in0(N__93806),
            .in1(N__63447),
            .in2(N__52159),
            .in3(N__82897),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3323_3324_LC_13_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3323_3324_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3323_3324_LC_13_11_4 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3323_3324_LC_13_11_4  (
            .in0(N__63446),
            .in1(N__52143),
            .in2(N__94590),
            .in3(N__80507),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3419_3420_LC_13_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3419_3420_LC_13_11_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3419_3420_LC_13_11_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3419_3420_LC_13_11_5  (
            .in0(N__93807),
            .in1(N__63448),
            .in2(N__52300),
            .in3(N__83343),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2075_2076_LC_13_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2075_2076_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2075_2076_LC_13_11_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2075_2076_LC_13_11_6  (
            .in0(N__63445),
            .in1(N__93808),
            .in2(N__54205),
            .in3(N__76985),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93333),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9990_3_lut_LC_13_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9990_3_lut_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9990_3_lut_LC_13_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9990_3_lut_LC_13_11_7  (
            .in0(N__52288),
            .in1(N__53722),
            .in2(_gnd_net_),
            .in3(N__88242),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11639 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i1726_4_lut_LC_13_12_0 .C_ON=1'b0;
    defparam \usb3_if_inst.i1726_4_lut_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i1726_4_lut_LC_13_12_0 .LUT_INIT=16'b1100010111000000;
    LogicCell40 \usb3_if_inst.i1726_4_lut_LC_13_12_0  (
            .in0(N__52264),
            .in1(N__52270),
            .in2(N__64080),
            .in3(N__57205),
            .lcout(),
            .ltout(\usb3_if_inst.n2912_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.state_timeout_counter_i0_i1_LC_13_12_1 .C_ON=1'b0;
    defparam \usb3_if_inst.state_timeout_counter_i0_i1_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.state_timeout_counter_i0_i1_LC_13_12_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \usb3_if_inst.state_timeout_counter_i0_i1_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__64142),
            .in2(N__52276),
            .in3(N__64345),
            .lcout(\usb3_if_inst.state_timeout_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_timeout_counter_i0_i1C_net ),
            .ce(N__54482),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i3_4_lut_LC_13_12_2 .C_ON=1'b0;
    defparam \usb3_if_inst.i3_4_lut_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i3_4_lut_LC_13_12_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \usb3_if_inst.i3_4_lut_LC_13_12_2  (
            .in0(N__57491),
            .in1(N__54348),
            .in2(N__54513),
            .in3(N__54322),
            .lcout(\usb3_if_inst.n7 ),
            .ltout(\usb3_if_inst.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.mux_40_i2_3_lut_4_lut_LC_13_12_3 .C_ON=1'b0;
    defparam \usb3_if_inst.mux_40_i2_3_lut_4_lut_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.mux_40_i2_3_lut_4_lut_LC_13_12_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \usb3_if_inst.mux_40_i2_3_lut_4_lut_LC_13_12_3  (
            .in0(N__57731),
            .in1(N__54328),
            .in2(N__52273),
            .in3(N__54352),
            .lcout(\usb3_if_inst.n137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i1_2_lut_LC_13_12_4 .C_ON=1'b0;
    defparam \usb3_if_inst.i1_2_lut_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i1_2_lut_LC_13_12_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \usb3_if_inst.i1_2_lut_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__54349),
            .in2(_gnd_net_),
            .in3(N__54323),
            .lcout(\usb3_if_inst.n3684 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.mux_40_i1_4_lut_LC_13_12_5 .C_ON=1'b0;
    defparam \usb3_if_inst.mux_40_i1_4_lut_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.mux_40_i1_4_lut_LC_13_12_5 .LUT_INIT=16'b0100010001110100;
    LogicCell40 \usb3_if_inst.mux_40_i1_4_lut_LC_13_12_5  (
            .in0(N__54324),
            .in1(N__57397),
            .in2(N__57748),
            .in3(N__64516),
            .lcout(),
            .ltout(\usb3_if_inst.n138_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i1555_4_lut_LC_13_12_6 .C_ON=1'b0;
    defparam \usb3_if_inst.i1555_4_lut_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i1555_4_lut_LC_13_12_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \usb3_if_inst.i1555_4_lut_LC_13_12_6  (
            .in0(N__64072),
            .in1(N__54325),
            .in2(N__52453),
            .in3(N__57204),
            .lcout(),
            .ltout(\usb3_if_inst.n2739_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.state_timeout_counter_i0_i0_LC_13_12_7 .C_ON=1'b0;
    defparam \usb3_if_inst.state_timeout_counter_i0_i0_LC_13_12_7 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.state_timeout_counter_i0_i0_LC_13_12_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \usb3_if_inst.state_timeout_counter_i0_i0_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__64141),
            .in2(N__52450),
            .in3(N__64344),
            .lcout(\usb3_if_inst.state_timeout_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_timeout_counter_i0_i1C_net ),
            .ce(N__54482),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.genblk16_rd_prev_r_132_LC_13_13_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.genblk16_rd_prev_r_132_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.genblk16_rd_prev_r_132_LC_13_13_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.genblk16_rd_prev_r_132_LC_13_13_0  (
            .in0(N__57711),
            .in1(N__73200),
            .in2(_gnd_net_),
            .in3(N__69046),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.genblk16_rd_prev_r ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97349),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i6_LC_13_13_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i6_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i6_LC_13_13_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i6_LC_13_13_1  (
            .in0(N__73202),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52447),
            .lcout(wp_sync1_r_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97349),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i6_LC_13_13_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i6_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i6_LC_13_13_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r__i6_LC_13_13_2  (
            .in0(N__52399),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73203),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97349),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i2_LC_13_13_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i2_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i2_LC_13_13_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync1_r__i2_LC_13_13_3  (
            .in0(N__73201),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52360),
            .lcout(wp_sync1_r_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97349),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i7_LC_13_13_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i7_LC_13_13_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i7_LC_13_13_4 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i7_LC_13_13_4  (
            .in0(N__80735),
            .in1(N__73199),
            .in2(N__65043),
            .in3(N__52333),
            .lcout(fifo_data_out_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97349),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i14_LC_13_13_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i14_LC_13_13_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i14_LC_13_13_5 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i14_LC_13_13_5  (
            .in0(N__73197),
            .in1(N__80733),
            .in2(N__68931),
            .in3(N__52324),
            .lcout(fifo_data_out_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97349),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i13_LC_13_13_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i13_LC_13_13_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i13_LC_13_13_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i13_LC_13_13_6  (
            .in0(N__80732),
            .in1(N__73196),
            .in2(N__52318),
            .in3(N__68496),
            .lcout(fifo_data_out_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97349),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i4_LC_13_13_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i4_LC_13_13_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i4_LC_13_13_7 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i4_LC_13_13_7  (
            .in0(N__73198),
            .in1(N__80734),
            .in2(N__64989),
            .in3(N__73108),
            .lcout(fifo_data_out_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97349),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.empty_o_I_0_1_lut_LC_13_14_0 .C_ON=1'b0;
    defparam \usb3_if_inst.empty_o_I_0_1_lut_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.empty_o_I_0_1_lut_LC_13_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \usb3_if_inst.empty_o_I_0_1_lut_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57709),
            .lcout(\usb3_if_inst.empty_o_N_599 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9834_3_lut_LC_13_14_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9834_3_lut_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9834_3_lut_LC_13_14_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9834_3_lut_LC_13_14_1  (
            .in0(N__52615),
            .in1(N__52606),
            .in2(_gnd_net_),
            .in3(N__52726),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11483_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.empty_ext_r_124_LC_13_14_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.empty_ext_r_124_LC_13_14_2 .SEQ_MODE=4'b1001;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.empty_ext_r_124_LC_13_14_2 .LUT_INIT=16'b0000110000101110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.empty_ext_r_124_LC_13_14_2  (
            .in0(N__69037),
            .in1(N__57706),
            .in2(N__52591),
            .in3(N__52588),
            .lcout(DEBUG_5_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97354),
            .ce(),
            .sr(N__73413));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_52_LC_13_14_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_52_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_52_LC_13_14_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_52_LC_13_14_3  (
            .in0(N__57707),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69038),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_fifo_en_w ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4_2_lut_LC_13_14_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4_2_lut_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4_2_lut_LC_13_14_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4_2_lut_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(N__52498),
            .in2(_gnd_net_),
            .in3(N__52489),
            .lcout(),
            .ltout(n5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.aempty_flag_impl_ae_flag_ext_r_130_LC_13_14_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.aempty_flag_impl_ae_flag_ext_r_130_LC_13_14_5 .SEQ_MODE=4'b1011;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.aempty_flag_impl_ae_flag_ext_r_130_LC_13_14_5 .LUT_INIT=16'b0000011100000011;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.aempty_flag_impl_ae_flag_ext_r_130_LC_13_14_5  (
            .in0(N__52480),
            .in1(N__52471),
            .in2(N__52462),
            .in3(N__69036),
            .lcout(dc32_fifo_almost_empty),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97354),
            .ce(),
            .sr(N__73413));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_fifo_en_w_I_0_158_2_lut_3_lut_LC_13_14_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_fifo_en_w_I_0_158_2_lut_3_lut_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_fifo_en_w_I_0_158_2_lut_3_lut_LC_13_14_6 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_fifo_en_w_I_0_158_2_lut_3_lut_LC_13_14_6  (
            .in0(N__69039),
            .in1(N__57708),
            .in2(_gnd_net_),
            .in3(N__52459),
            .lcout(t_rd_fifo_en_w),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i163_2_lut_2_lut_LC_13_14_7 .C_ON=1'b0;
    defparam \usb3_if_inst.i163_2_lut_2_lut_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i163_2_lut_2_lut_LC_13_14_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \usb3_if_inst.i163_2_lut_2_lut_LC_13_14_7  (
            .in0(N__57710),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57385),
            .lcout(\usb3_if_inst.n534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i11_LC_13_15_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i11_LC_13_15_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i11_LC_13_15_0 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i11_LC_13_15_0  (
            .in0(N__73415),
            .in1(N__80730),
            .in2(N__52759),
            .in3(N__58146),
            .lcout(fifo_data_out_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97358),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9782_4_lut_LC_13_15_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9782_4_lut_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9782_4_lut_LC_13_15_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9782_4_lut_LC_13_15_1  (
            .in0(N__52697),
            .in1(N__52742),
            .in2(N__85302),
            .in3(N__90527),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i2_LC_13_15_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i2_LC_13_15_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i2_LC_13_15_2 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i2_LC_13_15_2  (
            .in0(N__73416),
            .in1(N__80731),
            .in2(N__61549),
            .in3(N__65475),
            .lcout(fifo_data_out_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97358),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i0_LC_13_15_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i0_LC_13_15_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i0_LC_13_15_3 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i0_LC_13_15_3  (
            .in0(N__57315),
            .in1(N__80728),
            .in2(N__52720),
            .in3(N__73414),
            .lcout(fifo_data_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97358),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_48_LC_13_15_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_48_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_48_LC_13_15_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1_2_lut_adj_48_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__52696),
            .in2(_gnd_net_),
            .in3(N__52678),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync_w_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i1_LC_13_15_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i1_LC_13_15_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i1_LC_13_15_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r__i1_LC_13_15_6  (
            .in0(N__73417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52651),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97358),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i2_1_lut_LC_13_15_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i2_1_lut_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i2_1_lut_LC_13_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wp_sync2_r_6__I_0_149_inv_0_i2_1_lut_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90528),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n7_adj_1151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i1_LC_13_16_0 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i1_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i1_LC_13_16_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \spi0.tx_shift_reg_i0_i1_LC_13_16_0  (
            .in0(N__57891),
            .in1(N__57949),
            .in2(_gnd_net_),
            .in3(N__54793),
            .lcout(\spi0.tx_shift_reg_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97365),
            .ce(N__57962),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i2_LC_13_16_1 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i2_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i2_LC_13_16_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.tx_shift_reg_i0_i2_LC_13_16_1  (
            .in0(N__52627),
            .in1(N__58228),
            .in2(_gnd_net_),
            .in3(N__57892),
            .lcout(\spi0.tx_shift_reg_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97365),
            .ce(N__57962),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i3_LC_13_16_2 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i3_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i3_LC_13_16_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \spi0.tx_shift_reg_i0_i3_LC_13_16_2  (
            .in0(N__57893),
            .in1(N__52621),
            .in2(_gnd_net_),
            .in3(N__54845),
            .lcout(\spi0.tx_shift_reg_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97365),
            .ce(N__57962),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i4_LC_13_16_3 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i4_LC_13_16_3 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i4_LC_13_16_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.tx_shift_reg_i0_i4_LC_13_16_3  (
            .in0(N__52885),
            .in1(N__69443),
            .in2(_gnd_net_),
            .in3(N__57894),
            .lcout(\spi0.tx_shift_reg_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97365),
            .ce(N__57962),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i5_LC_13_16_4 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i5_LC_13_16_4 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i5_LC_13_16_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi0.tx_shift_reg_i0_i5_LC_13_16_4  (
            .in0(N__57895),
            .in1(N__54870),
            .in2(_gnd_net_),
            .in3(N__52879),
            .lcout(\spi0.tx_shift_reg_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97365),
            .ce(N__57962),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i6_LC_13_16_5 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i6_LC_13_16_5 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i6_LC_13_16_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.tx_shift_reg_i0_i6_LC_13_16_5  (
            .in0(N__52873),
            .in1(N__54816),
            .in2(_gnd_net_),
            .in3(N__57896),
            .lcout(\spi0.tx_shift_reg_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97365),
            .ce(N__57962),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_inv_0_i7_1_lut_LC_13_16_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_inv_0_i7_1_lut_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_inv_0_i7_1_lut_LC_13_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.wr_addr_r_6__I_0_inv_0_i7_1_lut_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52863),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6205_1_lut_LC_13_16_7.C_ON=1'b0;
    defparam i6205_1_lut_LC_13_16_7.SEQ_MODE=4'b0000;
    defparam i6205_1_lut_LC_13_16_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 i6205_1_lut_LC_13_16_7 (
            .in0(N__84712),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n7383),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_4_lut_adj_24_LC_13_17_0 .C_ON=1'b0;
    defparam \spi0.i1_4_lut_adj_24_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_4_lut_adj_24_LC_13_17_0 .LUT_INIT=16'b1110111000001110;
    LogicCell40 \spi0.i1_4_lut_adj_24_LC_13_17_0  (
            .in0(N__55487),
            .in1(N__55585),
            .in2(N__52822),
            .in3(N__52804),
            .lcout(\spi0.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i30_4_lut_LC_13_17_1 .C_ON=1'b0;
    defparam \spi0.i30_4_lut_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \spi0.i30_4_lut_LC_13_17_1 .LUT_INIT=16'b1111101001010001;
    LogicCell40 \spi0.i30_4_lut_LC_13_17_1  (
            .in0(N__55586),
            .in1(N__58479),
            .in2(N__55269),
            .in3(N__55489),
            .lcout(),
            .ltout(\spi0.n24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i11115_3_lut_4_lut_LC_13_17_2 .C_ON=1'b0;
    defparam \spi0.i11115_3_lut_4_lut_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \spi0.i11115_3_lut_4_lut_LC_13_17_2 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \spi0.i11115_3_lut_4_lut_LC_13_17_2  (
            .in0(N__55260),
            .in1(N__55008),
            .in2(N__52768),
            .in3(N__52765),
            .lcout(n4070),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i8605_3_lut_3_lut_LC_13_17_3 .C_ON=1'b0;
    defparam \spi0.i8605_3_lut_3_lut_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \spi0.i8605_3_lut_3_lut_LC_13_17_3 .LUT_INIT=16'b0000101001011010;
    LogicCell40 \spi0.i8605_3_lut_3_lut_LC_13_17_3  (
            .in0(N__55011),
            .in1(_gnd_net_),
            .in2(N__55270),
            .in3(N__55493),
            .lcout(\spi0.n10119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i4_4_lut_LC_13_17_4 .C_ON=1'b0;
    defparam \spi0.i4_4_lut_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \spi0.i4_4_lut_LC_13_17_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \spi0.i4_4_lut_LC_13_17_4  (
            .in0(N__58480),
            .in1(N__55265),
            .in2(N__55497),
            .in3(N__55105),
            .lcout(\spi0.n4105 ),
            .ltout(\spi0.n4105_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_2_lut_4_lut_LC_13_17_5 .C_ON=1'b0;
    defparam \spi0.i1_2_lut_4_lut_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_2_lut_4_lut_LC_13_17_5 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \spi0.i1_2_lut_4_lut_LC_13_17_5  (
            .in0(N__55009),
            .in1(N__55261),
            .in2(N__52918),
            .in3(N__52978),
            .lcout(\spi0.n11345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_rep_17_2_lut_LC_13_17_6 .C_ON=1'b0;
    defparam \spi0.i1_rep_17_2_lut_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_rep_17_2_lut_LC_13_17_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \spi0.i1_rep_17_2_lut_LC_13_17_6  (
            .in0(N__55488),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55010),
            .lcout(\spi0.n14442 ),
            .ltout(\spi0.n14442_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.state_i2_LC_13_17_7 .C_ON=1'b0;
    defparam \spi0.state_i2_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \spi0.state_i2_LC_13_17_7 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \spi0.state_i2_LC_13_17_7  (
            .in0(N__55587),
            .in1(N__54769),
            .in2(N__52915),
            .in3(N__52912),
            .lcout(\spi0.state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97372),
            .ce(N__52906),
            .sr(_gnd_net_));
    defparam \spi0.i11033_3_lut_LC_13_18_0 .C_ON=1'b0;
    defparam \spi0.i11033_3_lut_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \spi0.i11033_3_lut_LC_13_18_0 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \spi0.i11033_3_lut_LC_13_18_0  (
            .in0(N__55012),
            .in1(N__55233),
            .in2(_gnd_net_),
            .in3(N__54926),
            .lcout(),
            .ltout(\spi0.n12594_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.state_i1_LC_13_18_1 .C_ON=1'b0;
    defparam \spi0.state_i1_LC_13_18_1 .SEQ_MODE=4'b1000;
    defparam \spi0.state_i1_LC_13_18_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \spi0.state_i1_LC_13_18_1  (
            .in0(N__54763),
            .in1(N__55466),
            .in2(N__52897),
            .in3(N__55579),
            .lcout(\spi0.state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97379),
            .ce(N__52891),
            .sr(_gnd_net_));
    defparam \spi0.i2103_2_lut_LC_13_18_2 .C_ON=1'b0;
    defparam \spi0.i2103_2_lut_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \spi0.i2103_2_lut_LC_13_18_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \spi0.i2103_2_lut_LC_13_18_2  (
            .in0(N__55577),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55234),
            .lcout(),
            .ltout(\spi0.n3295_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_4_lut_adj_34_LC_13_18_3 .C_ON=1'b0;
    defparam \spi0.i1_4_lut_adj_34_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_4_lut_adj_34_LC_13_18_3 .LUT_INIT=16'b0101011100000000;
    LogicCell40 \spi0.i1_4_lut_adj_34_LC_13_18_3  (
            .in0(N__55463),
            .in1(N__55014),
            .in2(N__52894),
            .in3(N__52963),
            .lcout(\spi0.n11346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i2_3_lut_adj_26_LC_13_18_4 .C_ON=1'b0;
    defparam \spi0.i2_3_lut_adj_26_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \spi0.i2_3_lut_adj_26_LC_13_18_4 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \spi0.i2_3_lut_adj_26_LC_13_18_4  (
            .in0(N__55015),
            .in1(N__52977),
            .in2(_gnd_net_),
            .in3(N__55235),
            .lcout(\spi0.n4260 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i2_3_lut_LC_13_18_5 .C_ON=1'b0;
    defparam \spi0.i2_3_lut_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \spi0.i2_3_lut_LC_13_18_5 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \spi0.i2_3_lut_LC_13_18_5  (
            .in0(N__54927),
            .in1(N__55464),
            .in2(_gnd_net_),
            .in3(N__55578),
            .lcout(\spi0.n11311 ),
            .ltout(\spi0.n11311_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_3_lut_LC_13_18_6 .C_ON=1'b0;
    defparam \spi0.i1_3_lut_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_3_lut_LC_13_18_6 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \spi0.i1_3_lut_LC_13_18_6  (
            .in0(N__55013),
            .in1(_gnd_net_),
            .in2(N__52966),
            .in3(N__52956),
            .lcout(\spi0.n11344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i2_4_lut_LC_13_18_7 .C_ON=1'b0;
    defparam \spi0.i2_4_lut_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \spi0.i2_4_lut_LC_13_18_7 .LUT_INIT=16'b1010001010101010;
    LogicCell40 \spi0.i2_4_lut_LC_13_18_7  (
            .in0(N__52957),
            .in1(N__54928),
            .in2(N__55259),
            .in3(N__55465),
            .lcout(\spi0.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i11024_3_lut_4_lut_LC_13_19_0 .C_ON=1'b0;
    defparam \spi0.i11024_3_lut_4_lut_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \spi0.i11024_3_lut_4_lut_LC_13_19_0 .LUT_INIT=16'b0101011101010101;
    LogicCell40 \spi0.i11024_3_lut_4_lut_LC_13_19_0  (
            .in0(N__55436),
            .in1(N__55061),
            .in2(N__55231),
            .in3(N__55740),
            .lcout(),
            .ltout(\spi0.n12607_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i8614_4_lut_LC_13_19_1 .C_ON=1'b0;
    defparam \spi0.i8614_4_lut_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \spi0.i8614_4_lut_LC_13_19_1 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \spi0.i8614_4_lut_LC_13_19_1  (
            .in0(N__55064),
            .in1(N__55584),
            .in2(N__52948),
            .in3(N__52924),
            .lcout(\spi0.n4120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i11053_2_lut_LC_13_19_2 .C_ON=1'b0;
    defparam \spi0.i11053_2_lut_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \spi0.i11053_2_lut_LC_13_19_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \spi0.i11053_2_lut_LC_13_19_2  (
            .in0(N__55438),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55184),
            .lcout(\spi0.n12702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.byte_recv_92_i3_LC_13_19_3 .C_ON=1'b0;
    defparam \spi0.byte_recv_92_i3_LC_13_19_3 .SEQ_MODE=4'b1000;
    defparam \spi0.byte_recv_92_i3_LC_13_19_3 .LUT_INIT=16'b0000010000100000;
    LogicCell40 \spi0.byte_recv_92_i3_LC_13_19_3  (
            .in0(N__55059),
            .in1(N__55435),
            .in2(N__55230),
            .in3(N__55580),
            .lcout(spi_rx_byte_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97386),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i2026_4_lut_4_lut_LC_13_19_4 .C_ON=1'b0;
    defparam \spi0.i2026_4_lut_4_lut_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \spi0.i2026_4_lut_4_lut_LC_13_19_4 .LUT_INIT=16'b1111111010111111;
    LogicCell40 \spi0.i2026_4_lut_4_lut_LC_13_19_4  (
            .in0(N__55583),
            .in1(N__55446),
            .in2(N__55232),
            .in3(N__55063),
            .lcout(n3204),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i10998_2_lut_3_lut_LC_13_19_5 .C_ON=1'b0;
    defparam \spi0.i10998_2_lut_3_lut_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \spi0.i10998_2_lut_3_lut_LC_13_19_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \spi0.i10998_2_lut_3_lut_LC_13_19_5  (
            .in0(N__55060),
            .in1(N__55581),
            .in2(_gnd_net_),
            .in3(N__55185),
            .lcout(\spi0.n12586 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i11039_3_lut_LC_13_19_6 .C_ON=1'b0;
    defparam \spi0.i11039_3_lut_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \spi0.i11039_3_lut_LC_13_19_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \spi0.i11039_3_lut_LC_13_19_6  (
            .in0(N__55437),
            .in1(N__55183),
            .in2(_gnd_net_),
            .in3(N__55062),
            .lcout(),
            .ltout(\spi0.n12598_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_4_lut_adj_32_LC_13_19_7 .C_ON=1'b0;
    defparam \spi0.i1_4_lut_adj_32_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_4_lut_adj_32_LC_13_19_7 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \spi0.i1_4_lut_adj_32_LC_13_19_7  (
            .in0(N__53065),
            .in1(N__55582),
            .in2(N__53059),
            .in3(N__53056),
            .lcout(\spi0.CS_N_974 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i8568_4_lut_LC_13_20_0 .C_ON=1'b0;
    defparam \spi0.i8568_4_lut_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \spi0.i8568_4_lut_LC_13_20_0 .LUT_INIT=16'b1100000011001010;
    LogicCell40 \spi0.i8568_4_lut_LC_13_20_0  (
            .in0(N__55178),
            .in1(N__53005),
            .in2(N__55615),
            .in3(N__52984),
            .lcout(\spi0.n10082 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_2_lut_LC_13_20_1 .C_ON=1'b0;
    defparam \spi0.i1_2_lut_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_2_lut_LC_13_20_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \spi0.i1_2_lut_LC_13_20_1  (
            .in0(N__55459),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55065),
            .lcout(\spi0.n11350 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i8562_4_lut_4_lut_LC_13_20_2 .C_ON=1'b0;
    defparam \spi0.i8562_4_lut_4_lut_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \spi0.i8562_4_lut_4_lut_LC_13_20_2 .LUT_INIT=16'b0110001001110011;
    LogicCell40 \spi0.i8562_4_lut_4_lut_LC_13_20_2  (
            .in0(N__55067),
            .in1(N__55461),
            .in2(N__55768),
            .in3(N__54949),
            .lcout(),
            .ltout(\spi0.n10076_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i8567_3_lut_LC_13_20_3 .C_ON=1'b0;
    defparam \spi0.i8567_3_lut_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \spi0.i8567_3_lut_LC_13_20_3 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \spi0.i8567_3_lut_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(N__55177),
            .in2(N__53008),
            .in3(N__52999),
            .lcout(\spi0.n10081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i9750_3_lut_LC_13_20_4 .C_ON=1'b0;
    defparam \spi0.i9750_3_lut_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \spi0.i9750_3_lut_LC_13_20_4 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \spi0.i9750_3_lut_LC_13_20_4  (
            .in0(N__55068),
            .in1(N__55462),
            .in2(_gnd_net_),
            .in3(N__54950),
            .lcout(\spi0.n11398 ),
            .ltout(\spi0.n11398_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_4_lut_adj_36_LC_13_20_5 .C_ON=1'b0;
    defparam \spi0.i1_4_lut_adj_36_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_4_lut_adj_36_LC_13_20_5 .LUT_INIT=16'b0000110010001000;
    LogicCell40 \spi0.i1_4_lut_adj_36_LC_13_20_5  (
            .in0(N__52993),
            .in1(N__55608),
            .in2(N__52987),
            .in3(N__55176),
            .lcout(\spi0.n4281 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1_2_lut_adj_25_LC_13_20_6 .C_ON=1'b0;
    defparam \spi0.i1_2_lut_adj_25_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \spi0.i1_2_lut_adj_25_LC_13_20_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \spi0.i1_2_lut_adj_25_LC_13_20_6  (
            .in0(N__55066),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55460),
            .lcout(\spi0.n81 ),
            .ltout(\spi0.n81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.state_i0_LC_13_20_7 .C_ON=1'b0;
    defparam \spi0.state_i0_LC_13_20_7 .SEQ_MODE=4'b1000;
    defparam \spi0.state_i0_LC_13_20_7 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \spi0.state_i0_LC_13_20_7  (
            .in0(N__54739),
            .in1(_gnd_net_),
            .in2(N__53182),
            .in3(N__55179),
            .lcout(\spi0.state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97395),
            .ce(N__55081),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10050_3_lut_LC_14_1_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10050_3_lut_LC_14_1_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10050_3_lut_LC_14_1_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10050_3_lut_LC_14_1_0  (
            .in0(N__53896),
            .in1(N__53172),
            .in2(_gnd_net_),
            .in3(N__88845),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11699 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3401_3402_LC_14_1_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3401_3402_LC_14_1_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3401_3402_LC_14_1_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3401_3402_LC_14_1_1  (
            .in0(N__83379),
            .in1(N__96729),
            .in2(N__53173),
            .in3(N__95728),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93430),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i332_333_LC_14_1_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i332_333_LC_14_1_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i332_333_LC_14_1_2 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i332_333_LC_14_1_2  (
            .in0(N__95725),
            .in1(N__75932),
            .in2(N__53154),
            .in3(N__83381),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93430),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i341_342_LC_14_1_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i341_342_LC_14_1_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i341_342_LC_14_1_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i341_342_LC_14_1_3  (
            .in0(N__83380),
            .in1(N__62845),
            .in2(N__53133),
            .in3(N__95729),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93430),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3413_3414_LC_14_1_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3413_3414_LC_14_1_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3413_3414_LC_14_1_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3413_3414_LC_14_1_4  (
            .in0(N__95726),
            .in1(N__53115),
            .in2(N__62863),
            .in3(N__83382),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93430),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10440_3_lut_LC_14_1_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10440_3_lut_LC_14_1_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10440_3_lut_LC_14_1_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10440_3_lut_LC_14_1_5  (
            .in0(N__53116),
            .in1(_gnd_net_),
            .in2(N__88887),
            .in3(N__53101),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12089 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3317_3318_LC_14_1_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3317_3318_LC_14_1_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3317_3318_LC_14_1_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3317_3318_LC_14_1_6  (
            .in0(N__95724),
            .in1(N__53100),
            .in2(N__62862),
            .in3(N__80571),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93430),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i134_135_LC_14_1_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i134_135_LC_14_1_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i134_135_LC_14_1_7 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i134_135_LC_14_1_7  (
            .in0(N__71540),
            .in1(N__95727),
            .in2(N__53082),
            .in3(N__80317),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93430),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4937_4938_LC_14_2_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4937_4938_LC_14_2_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4937_4938_LC_14_2_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4937_4938_LC_14_2_0  (
            .in0(N__55632),
            .in1(N__96638),
            .in2(_gnd_net_),
            .in3(N__72261),
            .lcout(REG_mem_51_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93424),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10023_3_lut_LC_14_2_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10023_3_lut_LC_14_2_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10023_3_lut_LC_14_2_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10023_3_lut_LC_14_2_1  (
            .in0(N__53827),
            .in1(N__88881),
            .in2(_gnd_net_),
            .in3(N__53272),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11672 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1769_1770_LC_14_2_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1769_1770_LC_14_2_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1769_1770_LC_14_2_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1769_1770_LC_14_2_2  (
            .in0(N__53259),
            .in1(N__96635),
            .in2(_gnd_net_),
            .in3(N__67510),
            .lcout(REG_mem_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93424),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10029_3_lut_LC_14_2_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10029_3_lut_LC_14_2_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10029_3_lut_LC_14_2_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10029_3_lut_LC_14_2_3  (
            .in0(N__53260),
            .in1(N__53248),
            .in2(_gnd_net_),
            .in3(N__88882),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11678 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1865_1866_LC_14_2_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1865_1866_LC_14_2_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1865_1866_LC_14_2_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1865_1866_LC_14_2_4  (
            .in0(N__53247),
            .in1(N__96636),
            .in2(_gnd_net_),
            .in3(N__72112),
            .lcout(REG_mem_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93424),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2537_2538_LC_14_2_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2537_2538_LC_14_2_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2537_2538_LC_14_2_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2537_2538_LC_14_2_5  (
            .in0(N__96637),
            .in1(N__58914),
            .in2(_gnd_net_),
            .in3(N__70391),
            .lcout(REG_mem_26_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93424),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9906_3_lut_LC_14_2_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9906_3_lut_LC_14_2_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9906_3_lut_LC_14_2_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9906_3_lut_LC_14_2_6  (
            .in0(N__56884),
            .in1(N__85626),
            .in2(_gnd_net_),
            .in3(N__53398),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11555 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10052_3_lut_LC_14_2_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10052_3_lut_LC_14_2_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10052_3_lut_LC_14_2_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10052_3_lut_LC_14_2_7  (
            .in0(N__53233),
            .in1(N__88883),
            .in2(_gnd_net_),
            .in3(N__53218),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5621_5622_LC_14_3_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5621_5622_LC_14_3_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5621_5622_LC_14_3_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5621_5622_LC_14_3_0  (
            .in0(N__53190),
            .in1(_gnd_net_),
            .in2(N__62807),
            .in3(N__79967),
            .lcout(REG_mem_58_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11630_LC_14_3_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11630_LC_14_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11630_LC_14_3_1 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11630_LC_14_3_1  (
            .in0(N__92031),
            .in1(N__53191),
            .in2(N__53380),
            .in3(N__88821),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13340_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13340_bdd_4_lut_LC_14_3_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13340_bdd_4_lut_LC_14_3_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13340_bdd_4_lut_LC_14_3_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13340_bdd_4_lut_LC_14_3_2  (
            .in0(N__92028),
            .in1(N__53391),
            .in2(N__53425),
            .in3(N__53422),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5525_5526_LC_14_3_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5525_5526_LC_14_3_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5525_5526_LC_14_3_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5525_5526_LC_14_3_3  (
            .in0(N__95730),
            .in1(N__62718),
            .in2(N__53392),
            .in3(N__97035),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4190_4191_LC_14_3_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4190_4191_LC_14_3_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4190_4191_LC_14_3_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4190_4191_LC_14_3_4  (
            .in0(N__89439),
            .in1(N__85935),
            .in2(_gnd_net_),
            .in3(N__68297),
            .lcout(REG_mem_43_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5717_5718_LC_14_3_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5717_5718_LC_14_3_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5717_5718_LC_14_3_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5717_5718_LC_14_3_5  (
            .in0(N__95731),
            .in1(N__62719),
            .in2(N__53379),
            .in3(N__79658),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i275_276_LC_14_3_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i275_276_LC_14_3_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i275_276_LC_14_3_6 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i275_276_LC_14_3_6  (
            .in0(N__62353),
            .in1(N__53358),
            .in2(N__95770),
            .in3(N__80602),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93418),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10331_3_lut_LC_14_3_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10331_3_lut_LC_14_3_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10331_3_lut_LC_14_3_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10331_3_lut_LC_14_3_7  (
            .in0(N__53346),
            .in1(N__88820),
            .in2(_gnd_net_),
            .in3(N__53331),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11980 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11605_LC_14_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11605_LC_14_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11605_LC_14_4_0 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11605_LC_14_4_0  (
            .in0(N__85655),
            .in1(N__92029),
            .in2(N__53317),
            .in3(N__59005),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13346_bdd_4_lut_LC_14_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13346_bdd_4_lut_LC_14_4_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13346_bdd_4_lut_LC_14_4_1 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13346_bdd_4_lut_LC_14_4_1  (
            .in0(N__53305),
            .in1(N__53299),
            .in2(N__53284),
            .in3(N__85652),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12253_LC_14_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12253_LC_14_4_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12253_LC_14_4_2 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12253_LC_14_4_2  (
            .in0(N__85656),
            .in1(N__53281),
            .in2(N__53629),
            .in3(N__92030),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13994_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13994_bdd_4_lut_LC_14_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13994_bdd_4_lut_LC_14_4_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13994_bdd_4_lut_LC_14_4_3 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13994_bdd_4_lut_LC_14_4_3  (
            .in0(N__53533),
            .in1(N__53521),
            .in2(N__53515),
            .in3(N__85654),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11744_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13376_bdd_4_lut_LC_14_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13376_bdd_4_lut_LC_14_4_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13376_bdd_4_lut_LC_14_4_4 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13376_bdd_4_lut_LC_14_4_4  (
            .in0(N__53473),
            .in1(N__81448),
            .in2(N__53512),
            .in3(N__53509),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13352_bdd_4_lut_LC_14_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13352_bdd_4_lut_LC_14_4_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13352_bdd_4_lut_LC_14_4_5 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13352_bdd_4_lut_LC_14_4_5  (
            .in0(N__53485),
            .in1(N__85653),
            .in2(N__66106),
            .in3(N__55774),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11834_LC_14_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11834_LC_14_4_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11834_LC_14_4_6 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11834_LC_14_4_6  (
            .in0(N__90362),
            .in1(N__81449),
            .in2(N__53476),
            .in3(N__58726),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4373_4374_LC_14_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4373_4374_LC_14_5_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4373_4374_LC_14_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4373_4374_LC_14_5_0  (
            .in0(N__53466),
            .in1(N__62724),
            .in2(_gnd_net_),
            .in3(N__71887),
            .lcout(REG_mem_45_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11784_LC_14_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11784_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11784_LC_14_5_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11784_LC_14_5_1  (
            .in0(N__53668),
            .in1(N__91812),
            .in2(N__53659),
            .in3(N__88598),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13550_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13550_bdd_4_lut_LC_14_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13550_bdd_4_lut_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13550_bdd_4_lut_LC_14_5_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13550_bdd_4_lut_LC_14_5_2  (
            .in0(N__91811),
            .in1(N__53455),
            .in2(N__53437),
            .in3(N__53434),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11838 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3512_3513_LC_14_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3512_3513_LC_14_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3512_3513_LC_14_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3512_3513_LC_14_5_3  (
            .in0(N__53433),
            .in1(N__96368),
            .in2(_gnd_net_),
            .in3(N__54086),
            .lcout(REG_mem_36_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3704_3705_LC_14_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3704_3705_LC_14_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3704_3705_LC_14_5_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3704_3705_LC_14_5_4  (
            .in0(N__96366),
            .in1(N__53667),
            .in2(_gnd_net_),
            .in3(N__59272),
            .lcout(REG_mem_38_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3800_3801_LC_14_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3800_3801_LC_14_5_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3800_3801_LC_14_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3800_3801_LC_14_5_5  (
            .in0(N__53655),
            .in1(N__96369),
            .in2(_gnd_net_),
            .in3(N__61878),
            .lcout(REG_mem_39_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3605_3606_LC_14_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3605_3606_LC_14_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3605_3606_LC_14_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3605_3606_LC_14_5_6  (
            .in0(N__53640),
            .in1(N__62723),
            .in2(_gnd_net_),
            .in3(N__63717),
            .lcout(REG_mem_37_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1112_1113_LC_14_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1112_1113_LC_14_5_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1112_1113_LC_14_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1112_1113_LC_14_5_7  (
            .in0(N__66057),
            .in1(N__96367),
            .in2(_gnd_net_),
            .in3(N__66828),
            .lcout(REG_mem_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93400),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10022_3_lut_LC_14_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10022_3_lut_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10022_3_lut_LC_14_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10022_3_lut_LC_14_6_0  (
            .in0(N__53617),
            .in1(N__53608),
            .in2(_gnd_net_),
            .in3(N__88596),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1193_1194_LC_14_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1193_1194_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1193_1194_LC_14_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1193_1194_LC_14_6_1  (
            .in0(N__96695),
            .in1(N__53616),
            .in2(_gnd_net_),
            .in3(N__59658),
            .lcout(REG_mem_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1289_1290_LC_14_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1289_1290_LC_14_6_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1289_1290_LC_14_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1289_1290_LC_14_6_2  (
            .in0(N__53607),
            .in1(N__96696),
            .in2(_gnd_net_),
            .in3(N__70132),
            .lcout(REG_mem_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4073_4074_LC_14_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4073_4074_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4073_4074_LC_14_6_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4073_4074_LC_14_6_3  (
            .in0(N__96699),
            .in1(N__53589),
            .in2(_gnd_net_),
            .in3(N__68078),
            .lcout(REG_mem_42_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1673_1674_LC_14_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1673_1674_LC_14_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1673_1674_LC_14_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1673_1674_LC_14_6_4  (
            .in0(N__55785),
            .in1(N__96698),
            .in2(_gnd_net_),
            .in3(N__66580),
            .lcout(REG_mem_17_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10053_3_lut_LC_14_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10053_3_lut_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10053_3_lut_LC_14_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10053_3_lut_LC_14_6_5  (
            .in0(N__88597),
            .in1(N__53578),
            .in2(_gnd_net_),
            .in3(N__53560),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1481_1482_LC_14_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1481_1482_LC_14_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1481_1482_LC_14_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1481_1482_LC_14_6_6  (
            .in0(N__53820),
            .in1(N__96697),
            .in2(_gnd_net_),
            .in3(N__64005),
            .lcout(REG_mem_15_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3596_3597_LC_14_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3596_3597_LC_14_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3596_3597_LC_14_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3596_3597_LC_14_6_7  (
            .in0(N__61494),
            .in1(N__75988),
            .in2(_gnd_net_),
            .in3(N__63711),
            .lcout(REG_mem_37_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93387),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3794_3795_LC_14_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3794_3795_LC_14_7_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3794_3795_LC_14_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3794_3795_LC_14_7_0  (
            .in0(N__76691),
            .in1(N__59307),
            .in2(_gnd_net_),
            .in3(N__61891),
            .lcout(REG_mem_39_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11330_LC_14_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11330_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11330_LC_14_7_1 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11330_LC_14_7_1  (
            .in0(N__91643),
            .in1(N__88475),
            .in2(N__53734),
            .in3(N__53809),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13016_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13016_bdd_4_lut_LC_14_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13016_bdd_4_lut_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13016_bdd_4_lut_LC_14_7_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13016_bdd_4_lut_LC_14_7_2  (
            .in0(N__53794),
            .in1(N__91642),
            .in2(N__53773),
            .in3(N__53770),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13019 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3686_3687_LC_14_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3686_3687_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3686_3687_LC_14_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3686_3687_LC_14_7_3  (
            .in0(N__53730),
            .in1(N__71552),
            .in2(_gnd_net_),
            .in3(N__59275),
            .lcout(REG_mem_38_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1394_1395_LC_14_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1394_1395_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1394_1395_LC_14_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1394_1395_LC_14_7_4  (
            .in0(N__76690),
            .in1(N__53712),
            .in2(_gnd_net_),
            .in3(N__74753),
            .lcout(REG_mem_14_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i422_423_LC_14_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i422_423_LC_14_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i422_423_LC_14_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i422_423_LC_14_7_5  (
            .in0(N__53700),
            .in1(N__71553),
            .in2(_gnd_net_),
            .in3(N__72728),
            .lcout(REG_mem_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4454_4455_LC_14_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4454_4455_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4454_4455_LC_14_7_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4454_4455_LC_14_7_6  (
            .in0(N__71551),
            .in1(N__53679),
            .in2(_gnd_net_),
            .in3(N__89103),
            .lcout(REG_mem_46_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3305_3306_LC_14_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3305_3306_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3305_3306_LC_14_7_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3305_3306_LC_14_7_7  (
            .in0(N__96771),
            .in1(N__94577),
            .in2(N__53889),
            .in3(N__80547),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93374),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3977_3978_LC_14_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3977_3978_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3977_3978_LC_14_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3977_3978_LC_14_8_0  (
            .in0(N__53865),
            .in1(N__96770),
            .in2(_gnd_net_),
            .in3(N__66004),
            .lcout(REG_mem_41_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93361),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12308_LC_14_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12308_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12308_LC_14_8_1 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12308_LC_14_8_1  (
            .in0(N__91405),
            .in1(N__59737),
            .in2(N__88737),
            .in3(N__53851),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14192_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14192_bdd_4_lut_LC_14_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14192_bdd_4_lut_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14192_bdd_4_lut_LC_14_8_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14192_bdd_4_lut_LC_14_8_2  (
            .in0(N__53944),
            .in1(N__91404),
            .in2(N__53854),
            .in3(N__53911),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4766_4767_LC_14_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4766_4767_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4766_4767_LC_14_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4766_4767_LC_14_8_3  (
            .in0(N__89398),
            .in1(N__59694),
            .in2(_gnd_net_),
            .in3(N__62986),
            .lcout(REG_mem_49_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93361),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1406_1407_LC_14_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1406_1407_LC_14_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1406_1407_LC_14_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1406_1407_LC_14_8_4  (
            .in0(N__53850),
            .in1(N__89400),
            .in2(_gnd_net_),
            .in3(N__74745),
            .lcout(REG_mem_14_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93361),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1505_1506_LC_14_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1505_1506_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1505_1506_LC_14_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1505_1506_LC_14_8_5  (
            .in0(N__53838),
            .in1(N__56613),
            .in2(_gnd_net_),
            .in3(N__64010),
            .lcout(REG_mem_15_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93361),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1022_1023_LC_14_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1022_1023_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1022_1023_LC_14_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1022_1023_LC_14_8_6  (
            .in0(N__59385),
            .in1(N__89399),
            .in2(_gnd_net_),
            .in3(N__66980),
            .lcout(REG_mem_10_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93361),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1676_1677_LC_14_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1676_1677_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1676_1677_LC_14_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1676_1677_LC_14_8_7  (
            .in0(N__66529),
            .in1(N__56085),
            .in2(_gnd_net_),
            .in3(N__75998),
            .lcout(REG_mem_17_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93361),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10347_3_lut_LC_14_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10347_3_lut_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10347_3_lut_LC_14_9_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10347_3_lut_LC_14_9_0  (
            .in0(N__54127),
            .in1(N__88511),
            .in2(_gnd_net_),
            .in3(N__54118),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11996 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3731_3732_LC_14_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3731_3732_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3731_3732_LC_14_9_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3731_3732_LC_14_9_1  (
            .in0(N__59247),
            .in1(N__54126),
            .in2(_gnd_net_),
            .in3(N__62446),
            .lcout(REG_mem_38_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3827_3828_LC_14_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3827_3828_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3827_3828_LC_14_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3827_3828_LC_14_9_2  (
            .in0(N__62445),
            .in1(N__54117),
            .in2(_gnd_net_),
            .in3(N__61879),
            .lcout(REG_mem_39_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3506_3507_LC_14_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3506_3507_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3506_3507_LC_14_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3506_3507_LC_14_9_3  (
            .in0(N__56955),
            .in1(N__76702),
            .in2(_gnd_net_),
            .in3(N__54081),
            .lcout(REG_mem_36_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1310_1311_LC_14_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1310_1311_LC_14_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1310_1311_LC_14_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1310_1311_LC_14_9_4  (
            .in0(N__53943),
            .in1(N__89522),
            .in2(_gnd_net_),
            .in3(N__70109),
            .lcout(REG_mem_13_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2750_2751_LC_14_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2750_2751_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2750_2751_LC_14_9_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2750_2751_LC_14_9_5  (
            .in0(N__89521),
            .in1(N__94473),
            .in2(N__92694),
            .in3(N__70680),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i437_438_LC_14_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i437_438_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i437_438_LC_14_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i437_438_LC_14_9_6  (
            .in0(N__53922),
            .in1(N__62860),
            .in2(_gnd_net_),
            .in3(N__72687),
            .lcout(REG_mem_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1214_1215_LC_14_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1214_1215_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1214_1215_LC_14_9_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1214_1215_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(N__59611),
            .in2(N__89530),
            .in3(N__53907),
            .lcout(REG_mem_12_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93347),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2171_2172_LC_14_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2171_2172_LC_14_10_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2171_2172_LC_14_10_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2171_2172_LC_14_10_0  (
            .in0(N__63339),
            .in1(N__94471),
            .in2(N__54229),
            .in3(N__76235),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93321),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2267_2268_LC_14_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2267_2268_LC_14_10_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2267_2268_LC_14_10_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2267_2268_LC_14_10_1  (
            .in0(N__54213),
            .in1(N__63340),
            .in2(_gnd_net_),
            .in3(N__75002),
            .lcout(REG_mem_23_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93321),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2840_2841_LC_14_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2840_2841_LC_14_10_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2840_2841_LC_14_10_2 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2840_2841_LC_14_10_2  (
            .in0(N__96365),
            .in1(N__94472),
            .in2(N__69846),
            .in3(N__70964),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93321),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12223_LC_14_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12223_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12223_LC_14_10_3 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12223_LC_14_10_3  (
            .in0(N__54295),
            .in1(N__54274),
            .in2(N__91730),
            .in3(N__88510),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14090_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14090_bdd_4_lut_LC_14_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14090_bdd_4_lut_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14090_bdd_4_lut_LC_14_10_4 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14090_bdd_4_lut_LC_14_10_4  (
            .in0(N__63568),
            .in1(N__91283),
            .in2(N__54259),
            .in3(N__54256),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12123_LC_14_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12123_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12123_LC_14_10_5 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12123_LC_14_10_5  (
            .in0(N__91284),
            .in1(N__54228),
            .in2(N__54217),
            .in3(N__88509),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13964_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13964_bdd_4_lut_LC_14_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13964_bdd_4_lut_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13964_bdd_4_lut_LC_14_10_6 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13964_bdd_4_lut_LC_14_10_6  (
            .in0(N__54204),
            .in1(N__91282),
            .in2(N__54190),
            .in3(N__54187),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3059_3060_LC_14_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3059_3060_LC_14_10_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3059_3060_LC_14_10_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3059_3060_LC_14_10_7  (
            .in0(N__54156),
            .in1(N__62354),
            .in2(_gnd_net_),
            .in3(N__72501),
            .lcout(REG_mem_31_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93321),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1106_1107_LC_14_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1106_1107_LC_14_11_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1106_1107_LC_14_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1106_1107_LC_14_11_0  (
            .in0(N__76712),
            .in1(N__56922),
            .in2(_gnd_net_),
            .in3(N__66808),
            .lcout(REG_mem_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93348),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12053_LC_14_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12053_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12053_LC_14_11_1 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12053_LC_14_11_1  (
            .in0(N__85406),
            .in1(N__63829),
            .in2(N__91403),
            .in3(N__64027),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13796 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10014_3_lut_LC_14_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10014_3_lut_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10014_3_lut_LC_14_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10014_3_lut_LC_14_11_2  (
            .in0(N__88245),
            .in1(N__54385),
            .in2(_gnd_net_),
            .in3(N__54394),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11663 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1778_1779_LC_14_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1778_1779_LC_14_11_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1778_1779_LC_14_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1778_1779_LC_14_11_3  (
            .in0(N__54393),
            .in1(N__76716),
            .in2(_gnd_net_),
            .in3(N__67486),
            .lcout(REG_mem_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93348),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1874_1875_LC_14_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1874_1875_LC_14_11_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1874_1875_LC_14_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1874_1875_LC_14_11_4  (
            .in0(N__76714),
            .in1(N__54384),
            .in2(_gnd_net_),
            .in3(N__72100),
            .lcout(REG_mem_19_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93348),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10013_3_lut_LC_14_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10013_3_lut_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10013_3_lut_LC_14_11_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10013_3_lut_LC_14_11_5  (
            .in0(N__54364),
            .in1(N__88244),
            .in2(_gnd_net_),
            .in3(N__54375),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1586_1587_LC_14_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1586_1587_LC_14_11_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1586_1587_LC_14_11_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1586_1587_LC_14_11_6  (
            .in0(N__76713),
            .in1(_gnd_net_),
            .in2(N__54376),
            .in3(N__65687),
            .lcout(REG_mem_16_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93348),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1682_1683_LC_14_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1682_1683_LC_14_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1682_1683_LC_14_11_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1682_1683_LC_14_11_7  (
            .in0(N__54363),
            .in1(N__76715),
            .in2(_gnd_net_),
            .in3(N__66581),
            .lcout(REG_mem_17_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93348),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i1_3_lut_4_lut_adj_21_LC_14_12_0 .C_ON=1'b0;
    defparam \usb3_if_inst.i1_3_lut_4_lut_adj_21_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i1_3_lut_4_lut_adj_21_LC_14_12_0 .LUT_INIT=16'b0000111100011110;
    LogicCell40 \usb3_if_inst.i1_3_lut_4_lut_adj_21_LC_14_12_0  (
            .in0(N__57501),
            .in1(N__54351),
            .in2(N__54514),
            .in3(N__54327),
            .lcout(\usb3_if_inst.n3686 ),
            .ltout(\usb3_if_inst.n3686_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.mux_40_i4_4_lut_LC_14_12_1 .C_ON=1'b0;
    defparam \usb3_if_inst.mux_40_i4_4_lut_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.mux_40_i4_4_lut_LC_14_12_1 .LUT_INIT=16'b0100111000001010;
    LogicCell40 \usb3_if_inst.mux_40_i4_4_lut_LC_14_12_1  (
            .in0(N__57393),
            .in1(N__64517),
            .in2(N__54355),
            .in3(N__57753),
            .lcout(\usb3_if_inst.n135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i1277_2_lut_LC_14_12_2 .C_ON=1'b0;
    defparam \usb3_if_inst.i1277_2_lut_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i1277_2_lut_LC_14_12_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \usb3_if_inst.i1277_2_lut_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__54350),
            .in2(_gnd_net_),
            .in3(N__54326),
            .lcout(\usb3_if_inst.n4 ),
            .ltout(\usb3_if_inst.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.mux_40_i3_3_lut_4_lut_LC_14_12_3 .C_ON=1'b0;
    defparam \usb3_if_inst.mux_40_i3_3_lut_4_lut_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.mux_40_i3_3_lut_4_lut_LC_14_12_3 .LUT_INIT=16'b0100111011100100;
    LogicCell40 \usb3_if_inst.mux_40_i3_3_lut_4_lut_LC_14_12_3  (
            .in0(N__57392),
            .in1(N__57752),
            .in2(N__54298),
            .in3(N__57500),
            .lcout(),
            .ltout(\usb3_if_inst.n4403_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i5710_4_lut_LC_14_12_4 .C_ON=1'b0;
    defparam \usb3_if_inst.i5710_4_lut_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i5710_4_lut_LC_14_12_4 .LUT_INIT=16'b0000101001001110;
    LogicCell40 \usb3_if_inst.i5710_4_lut_LC_14_12_4  (
            .in0(N__64071),
            .in1(N__57223),
            .in2(N__54544),
            .in3(N__57454),
            .lcout(\usb3_if_inst.n6904 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.state_timeout_counter_i0_i3_LC_14_12_5 .C_ON=1'b0;
    defparam \usb3_if_inst.state_timeout_counter_i0_i3_LC_14_12_5 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.state_timeout_counter_i0_i3_LC_14_12_5 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \usb3_if_inst.state_timeout_counter_i0_i3_LC_14_12_5  (
            .in0(N__64070),
            .in1(N__54529),
            .in2(N__54523),
            .in3(N__57203),
            .lcout(\usb3_if_inst.state_timeout_counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_timeout_counter_i0_i3C_net ),
            .ce(N__54492),
            .sr(N__57178));
    defparam \usb3_if_inst.i10966_2_lut_LC_14_12_6 .C_ON=1'b0;
    defparam \usb3_if_inst.i10966_2_lut_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i10966_2_lut_LC_14_12_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \usb3_if_inst.i10966_2_lut_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(N__64069),
            .in2(_gnd_net_),
            .in3(N__57222),
            .lcout(),
            .ltout(\usb3_if_inst.n12582_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i1_4_lut_LC_14_12_7 .C_ON=1'b0;
    defparam \usb3_if_inst.i1_4_lut_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i1_4_lut_LC_14_12_7 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \usb3_if_inst.i1_4_lut_LC_14_12_7  (
            .in0(N__64149),
            .in1(N__73718),
            .in2(N__54496),
            .in3(N__57513),
            .lcout(\usb3_if_inst.n4061 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.num_lines_clocked_out_i0_LC_14_13_0 .C_ON=1'b1;
    defparam \usb3_if_inst.num_lines_clocked_out_i0_LC_14_13_0 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.num_lines_clocked_out_i0_LC_14_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \usb3_if_inst.num_lines_clocked_out_i0_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__54441),
            .in2(N__54457),
            .in3(N__54427),
            .lcout(\usb3_if_inst.num_lines_clocked_out_0 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\usb3_if_inst.n10660 ),
            .clk(\INVusb3_if_inst.num_lines_clocked_out_i0C_net ),
            .ce(N__57334),
            .sr(N__73656));
    defparam \usb3_if_inst.num_lines_clocked_out_i1_LC_14_13_1 .C_ON=1'b1;
    defparam \usb3_if_inst.num_lines_clocked_out_i1_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.num_lines_clocked_out_i1_LC_14_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \usb3_if_inst.num_lines_clocked_out_i1_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__64821),
            .in2(N__86571),
            .in3(N__54424),
            .lcout(\usb3_if_inst.num_lines_clocked_out_1 ),
            .ltout(),
            .carryin(\usb3_if_inst.n10660 ),
            .carryout(\usb3_if_inst.n10661 ),
            .clk(\INVusb3_if_inst.num_lines_clocked_out_i0C_net ),
            .ce(N__57334),
            .sr(N__73656));
    defparam \usb3_if_inst.num_lines_clocked_out_i2_LC_14_13_2 .C_ON=1'b1;
    defparam \usb3_if_inst.num_lines_clocked_out_i2_LC_14_13_2 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.num_lines_clocked_out_i2_LC_14_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \usb3_if_inst.num_lines_clocked_out_i2_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__86484),
            .in2(N__54420),
            .in3(N__54400),
            .lcout(\usb3_if_inst.num_lines_clocked_out_2 ),
            .ltout(),
            .carryin(\usb3_if_inst.n10661 ),
            .carryout(\usb3_if_inst.n10662 ),
            .clk(\INVusb3_if_inst.num_lines_clocked_out_i0C_net ),
            .ce(N__57334),
            .sr(N__73656));
    defparam \usb3_if_inst.num_lines_clocked_out_i3_LC_14_13_3 .C_ON=1'b1;
    defparam \usb3_if_inst.num_lines_clocked_out_i3_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.num_lines_clocked_out_i3_LC_14_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \usb3_if_inst.num_lines_clocked_out_i3_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__64629),
            .in2(N__86572),
            .in3(N__54397),
            .lcout(\usb3_if_inst.num_lines_clocked_out_3 ),
            .ltout(),
            .carryin(\usb3_if_inst.n10662 ),
            .carryout(\usb3_if_inst.n10663 ),
            .clk(\INVusb3_if_inst.num_lines_clocked_out_i0C_net ),
            .ce(N__57334),
            .sr(N__73656));
    defparam \usb3_if_inst.num_lines_clocked_out_i4_LC_14_13_4 .C_ON=1'b1;
    defparam \usb3_if_inst.num_lines_clocked_out_i4_LC_14_13_4 .SEQ_MODE=4'b1001;
    defparam \usb3_if_inst.num_lines_clocked_out_i4_LC_14_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \usb3_if_inst.num_lines_clocked_out_i4_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__86488),
            .in2(N__64542),
            .in3(N__54610),
            .lcout(\usb3_if_inst.num_lines_clocked_out_4 ),
            .ltout(),
            .carryin(\usb3_if_inst.n10663 ),
            .carryout(\usb3_if_inst.n10664 ),
            .clk(\INVusb3_if_inst.num_lines_clocked_out_i0C_net ),
            .ce(N__57334),
            .sr(N__73656));
    defparam \usb3_if_inst.num_lines_clocked_out_i5_LC_14_13_5 .C_ON=1'b1;
    defparam \usb3_if_inst.num_lines_clocked_out_i5_LC_14_13_5 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.num_lines_clocked_out_i5_LC_14_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \usb3_if_inst.num_lines_clocked_out_i5_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__64839),
            .in2(N__86573),
            .in3(N__54607),
            .lcout(\usb3_if_inst.num_lines_clocked_out_5 ),
            .ltout(),
            .carryin(\usb3_if_inst.n10664 ),
            .carryout(\usb3_if_inst.n10665 ),
            .clk(\INVusb3_if_inst.num_lines_clocked_out_i0C_net ),
            .ce(N__57334),
            .sr(N__73656));
    defparam \usb3_if_inst.num_lines_clocked_out_i6_LC_14_13_6 .C_ON=1'b1;
    defparam \usb3_if_inst.num_lines_clocked_out_i6_LC_14_13_6 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.num_lines_clocked_out_i6_LC_14_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \usb3_if_inst.num_lines_clocked_out_i6_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__86492),
            .in2(N__64614),
            .in3(N__54604),
            .lcout(\usb3_if_inst.num_lines_clocked_out_6 ),
            .ltout(),
            .carryin(\usb3_if_inst.n10665 ),
            .carryout(\usb3_if_inst.n10666 ),
            .clk(\INVusb3_if_inst.num_lines_clocked_out_i0C_net ),
            .ce(N__57334),
            .sr(N__73656));
    defparam \usb3_if_inst.num_lines_clocked_out_i7_LC_14_13_7 .C_ON=1'b1;
    defparam \usb3_if_inst.num_lines_clocked_out_i7_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.num_lines_clocked_out_i7_LC_14_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \usb3_if_inst.num_lines_clocked_out_i7_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(N__54597),
            .in2(N__86574),
            .in3(N__54583),
            .lcout(\usb3_if_inst.num_lines_clocked_out_7 ),
            .ltout(),
            .carryin(\usb3_if_inst.n10666 ),
            .carryout(\usb3_if_inst.n10667 ),
            .clk(\INVusb3_if_inst.num_lines_clocked_out_i0C_net ),
            .ce(N__57334),
            .sr(N__73656));
    defparam \usb3_if_inst.num_lines_clocked_out_i8_LC_14_14_0 .C_ON=1'b1;
    defparam \usb3_if_inst.num_lines_clocked_out_i8_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.num_lines_clocked_out_i8_LC_14_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \usb3_if_inst.num_lines_clocked_out_i8_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__64557),
            .in2(N__86575),
            .in3(N__54580),
            .lcout(\usb3_if_inst.num_lines_clocked_out_8 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\usb3_if_inst.n10668 ),
            .clk(\INVusb3_if_inst.num_lines_clocked_out_i8C_net ),
            .ce(N__57333),
            .sr(N__73704));
    defparam \usb3_if_inst.num_lines_clocked_out_i9_LC_14_14_1 .C_ON=1'b1;
    defparam \usb3_if_inst.num_lines_clocked_out_i9_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.num_lines_clocked_out_i9_LC_14_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \usb3_if_inst.num_lines_clocked_out_i9_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__86500),
            .in2(N__54576),
            .in3(N__54556),
            .lcout(\usb3_if_inst.num_lines_clocked_out_9 ),
            .ltout(),
            .carryin(\usb3_if_inst.n10668 ),
            .carryout(\usb3_if_inst.n10669 ),
            .clk(\INVusb3_if_inst.num_lines_clocked_out_i8C_net ),
            .ce(N__57333),
            .sr(N__73704));
    defparam \usb3_if_inst.num_lines_clocked_out_i10_LC_14_14_2 .C_ON=1'b0;
    defparam \usb3_if_inst.num_lines_clocked_out_i10_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.num_lines_clocked_out_i10_LC_14_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \usb3_if_inst.num_lines_clocked_out_i10_LC_14_14_2  (
            .in0(N__86496),
            .in1(N__64587),
            .in2(_gnd_net_),
            .in3(N__54553),
            .lcout(\usb3_if_inst.num_lines_clocked_out_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.num_lines_clocked_out_i8C_net ),
            .ce(N__57333),
            .sr(N__73704));
    defparam \spi0.tx_shift_reg_i0_i9_LC_14_15_0 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i9_LC_14_15_0 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i9_LC_14_15_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi0.tx_shift_reg_i0_i9_LC_14_15_0  (
            .in0(N__57924),
            .in1(N__54730),
            .in2(_gnd_net_),
            .in3(N__54640),
            .lcout(\spi0.tx_shift_reg_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97366),
            .ce(N__57980),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i10_LC_14_15_1 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i10_LC_14_15_1 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i10_LC_14_15_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.tx_shift_reg_i0_i10_LC_14_15_1  (
            .in0(N__54550),
            .in1(N__58198),
            .in2(_gnd_net_),
            .in3(N__57917),
            .lcout(\spi0.tx_shift_reg_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97366),
            .ce(N__57980),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i11_LC_14_15_2 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i11_LC_14_15_2 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i11_LC_14_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \spi0.tx_shift_reg_i0_i11_LC_14_15_2  (
            .in0(N__57918),
            .in1(N__54667),
            .in2(_gnd_net_),
            .in3(N__54889),
            .lcout(\spi0.tx_shift_reg_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97366),
            .ce(N__57980),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i12_LC_14_15_3 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i12_LC_14_15_3 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i12_LC_14_15_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.tx_shift_reg_i0_i12_LC_14_15_3  (
            .in0(N__54661),
            .in1(N__69319),
            .in2(_gnd_net_),
            .in3(N__57919),
            .lcout(\spi0.tx_shift_reg_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97366),
            .ce(N__57980),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i13_LC_14_15_4 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i13_LC_14_15_4 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i13_LC_14_15_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi0.tx_shift_reg_i0_i13_LC_14_15_4  (
            .in0(N__57920),
            .in1(N__54622),
            .in2(_gnd_net_),
            .in3(N__54655),
            .lcout(\spi0.tx_shift_reg_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97366),
            .ce(N__57980),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i14_LC_14_15_5 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i14_LC_14_15_5 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i14_LC_14_15_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.tx_shift_reg_i0_i14_LC_14_15_5  (
            .in0(N__54646),
            .in1(N__54706),
            .in2(_gnd_net_),
            .in3(N__57921),
            .lcout(\spi0.tx_shift_reg_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97366),
            .ce(N__57980),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i8_LC_14_15_6 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i8_LC_14_15_6 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i8_LC_14_15_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi0.tx_shift_reg_i0_i8_LC_14_15_6  (
            .in0(N__57923),
            .in1(N__54682),
            .in2(_gnd_net_),
            .in3(N__54628),
            .lcout(\spi0.tx_shift_reg_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97366),
            .ce(N__57980),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i7_LC_14_15_7 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i7_LC_14_15_7 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i7_LC_14_15_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.tx_shift_reg_i0_i7_LC_14_15_7  (
            .in0(N__54634),
            .in1(N__58451),
            .in2(_gnd_net_),
            .in3(N__57922),
            .lcout(\spi0.tx_shift_reg_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97366),
            .ce(N__57980),
            .sr(_gnd_net_));
    defparam tx_data_byte_r_i0_i5_LC_14_16_0.C_ON=1'b0;
    defparam tx_data_byte_r_i0_i5_LC_14_16_0.SEQ_MODE=4'b1000;
    defparam tx_data_byte_r_i0_i5_LC_14_16_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 tx_data_byte_r_i0_i5_LC_14_16_0 (
            .in0(N__54869),
            .in1(N__54717),
            .in2(_gnd_net_),
            .in3(N__69407),
            .lcout(tx_data_byte_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97373),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_Rx_Byte_i7_LC_14_16_1 .C_ON=1'b0;
    defparam \pc_rx.r_Rx_Byte_i7_LC_14_16_1 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Rx_Byte_i7_LC_14_16_1 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \pc_rx.r_Rx_Byte_i7_LC_14_16_1  (
            .in0(N__60726),
            .in1(N__60175),
            .in2(N__57820),
            .in3(N__58305),
            .lcout(pc_data_rx_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97373),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_addr_byte_r_i0_i5_LC_14_16_2.C_ON=1'b0;
    defparam tx_addr_byte_r_i0_i5_LC_14_16_2.SEQ_MODE=4'b1000;
    defparam tx_addr_byte_r_i0_i5_LC_14_16_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 tx_addr_byte_r_i0_i5_LC_14_16_2 (
            .in0(N__54868),
            .in1(N__69404),
            .in2(_gnd_net_),
            .in3(N__54621),
            .lcout(tx_addr_byte_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97373),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_addr_byte_r_i0_i1_LC_14_16_3.C_ON=1'b0;
    defparam tx_addr_byte_r_i0_i1_LC_14_16_3.SEQ_MODE=4'b1000;
    defparam tx_addr_byte_r_i0_i1_LC_14_16_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 tx_addr_byte_r_i0_i1_LC_14_16_3 (
            .in0(N__54792),
            .in1(N__69403),
            .in2(_gnd_net_),
            .in3(N__54729),
            .lcout(tx_addr_byte_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97373),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_data_byte_r_i0_i3_LC_14_16_4.C_ON=1'b0;
    defparam tx_data_byte_r_i0_i3_LC_14_16_4.SEQ_MODE=4'b1000;
    defparam tx_data_byte_r_i0_i3_LC_14_16_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 tx_data_byte_r_i0_i3_LC_14_16_4 (
            .in0(N__60136),
            .in1(N__69406),
            .in2(_gnd_net_),
            .in3(N__54844),
            .lcout(tx_data_byte_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97373),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_Rx_Byte_i5_LC_14_16_5 .C_ON=1'b0;
    defparam \pc_rx.r_Rx_Byte_i5_LC_14_16_5 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Rx_Byte_i5_LC_14_16_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \pc_rx.r_Rx_Byte_i5_LC_14_16_5  (
            .in0(N__60725),
            .in1(N__60174),
            .in2(N__54718),
            .in3(N__58336),
            .lcout(pc_data_rx_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97373),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_data_byte_r_i0_i6_LC_14_16_6.C_ON=1'b0;
    defparam tx_data_byte_r_i0_i6_LC_14_16_6.SEQ_MODE=4'b1000;
    defparam tx_data_byte_r_i0_i6_LC_14_16_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 tx_data_byte_r_i0_i6_LC_14_16_6 (
            .in0(N__54815),
            .in1(N__69408),
            .in2(_gnd_net_),
            .in3(N__58240),
            .lcout(tx_data_byte_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97373),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_addr_byte_r_i0_i6_LC_14_16_7.C_ON=1'b0;
    defparam tx_addr_byte_r_i0_i6_LC_14_16_7.SEQ_MODE=4'b1000;
    defparam tx_addr_byte_r_i0_i6_LC_14_16_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 tx_addr_byte_r_i0_i6_LC_14_16_7 (
            .in0(N__69405),
            .in1(N__54814),
            .in2(_gnd_net_),
            .in3(N__54705),
            .lcout(tx_addr_byte_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97373),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i3_4_lut_LC_14_17_0 .C_ON=1'b0;
    defparam \pc_rx.i3_4_lut_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i3_4_lut_LC_14_17_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \pc_rx.i3_4_lut_LC_14_17_0  (
            .in0(N__60385),
            .in1(N__60796),
            .in2(N__58324),
            .in3(N__60082),
            .lcout(),
            .ltout(n10847_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_Rx_Byte_i0_LC_14_17_1 .C_ON=1'b0;
    defparam \pc_rx.r_Rx_Byte_i0_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Rx_Byte_i0_LC_14_17_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \pc_rx.r_Rx_Byte_i0_LC_14_17_1  (
            .in0(N__54690),
            .in1(_gnd_net_),
            .in2(N__54694),
            .in3(N__60733),
            .lcout(pc_data_rx_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97380),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_data_byte_r_i0_i0_LC_14_17_2.C_ON=1'b0;
    defparam tx_data_byte_r_i0_i0_LC_14_17_2.SEQ_MODE=4'b1000;
    defparam tx_data_byte_r_i0_i0_LC_14_17_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 tx_data_byte_r_i0_i0_LC_14_17_2 (
            .in0(N__58019),
            .in1(N__69377),
            .in2(_gnd_net_),
            .in3(N__54691),
            .lcout(tx_data_byte_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97380),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_addr_byte_r_i0_i0_LC_14_17_3.C_ON=1'b0;
    defparam tx_addr_byte_r_i0_i0_LC_14_17_3.SEQ_MODE=4'b1000;
    defparam tx_addr_byte_r_i0_i0_LC_14_17_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 tx_addr_byte_r_i0_i0_LC_14_17_3 (
            .in0(N__69375),
            .in1(N__58018),
            .in2(_gnd_net_),
            .in3(N__54678),
            .lcout(tx_addr_byte_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97380),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i1_2_lut_3_lut_LC_14_17_4 .C_ON=1'b0;
    defparam \pc_rx.i1_2_lut_3_lut_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i1_2_lut_3_lut_LC_14_17_4 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \pc_rx.i1_2_lut_3_lut_LC_14_17_4  (
            .in0(N__60384),
            .in1(N__60795),
            .in2(_gnd_net_),
            .in3(N__60081),
            .lcout(n3997),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_addr_byte_r_i0_i3_LC_14_17_5.C_ON=1'b0;
    defparam tx_addr_byte_r_i0_i3_LC_14_17_5.SEQ_MODE=4'b1000;
    defparam tx_addr_byte_r_i0_i3_LC_14_17_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 tx_addr_byte_r_i0_i3_LC_14_17_5 (
            .in0(N__69376),
            .in1(N__54846),
            .in2(_gnd_net_),
            .in3(N__54885),
            .lcout(tx_addr_byte_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97380),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_data_byte_r_i0_i2_LC_14_17_6.C_ON=1'b0;
    defparam tx_data_byte_r_i0_i2_LC_14_17_6.SEQ_MODE=4'b1000;
    defparam tx_data_byte_r_i0_i2_LC_14_17_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 tx_data_byte_r_i0_i2_LC_14_17_6 (
            .in0(N__58219),
            .in1(N__69378),
            .in2(_gnd_net_),
            .in3(N__58173),
            .lcout(tx_data_byte_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97380),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_data_byte_r_i0_i1_LC_14_17_7.C_ON=1'b0;
    defparam tx_data_byte_r_i0_i1_LC_14_17_7.SEQ_MODE=4'b1000;
    defparam tx_data_byte_r_i0_i1_LC_14_17_7.LUT_INIT=16'b1110111000100010;
    LogicCell40 tx_data_byte_r_i0_i1_LC_14_17_7 (
            .in0(N__54790),
            .in1(N__69379),
            .in2(_gnd_net_),
            .in3(N__58414),
            .lcout(tx_data_byte_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97380),
            .ce(),
            .sr(_gnd_net_));
    defparam i9764_2_lut_LC_14_18_0.C_ON=1'b0;
    defparam i9764_2_lut_LC_14_18_0.SEQ_MODE=4'b0000;
    defparam i9764_2_lut_LC_14_18_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 i9764_2_lut_LC_14_18_0 (
            .in0(N__58459),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54874),
            .lcout(),
            .ltout(n11412_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9823_4_lut_LC_14_18_1.C_ON=1'b0;
    defparam i9823_4_lut_LC_14_18_1.SEQ_MODE=4'b0000;
    defparam i9823_4_lut_LC_14_18_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 i9823_4_lut_LC_14_18_1 (
            .in0(N__69444),
            .in1(N__54850),
            .in2(N__54823),
            .in3(N__58227),
            .lcout(),
            .ltout(n11471_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam multi_byte_spi_trans_flag_r_86_LC_14_18_2.C_ON=1'b0;
    defparam multi_byte_spi_trans_flag_r_86_LC_14_18_2.SEQ_MODE=4'b1000;
    defparam multi_byte_spi_trans_flag_r_86_LC_14_18_2.LUT_INIT=16'b0000000000010000;
    LogicCell40 multi_byte_spi_trans_flag_r_86_LC_14_18_2 (
            .in0(N__58020),
            .in1(N__54820),
            .in2(N__54796),
            .in3(N__54791),
            .lcout(multi_byte_spi_trans_flag_r),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97387),
            .ce(),
            .sr(N__58501));
    defparam \spi0.i10988_3_lut_4_lut_LC_14_18_3 .C_ON=1'b0;
    defparam \spi0.i10988_3_lut_4_lut_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \spi0.i10988_3_lut_4_lut_LC_14_18_3 .LUT_INIT=16'b0101010100010000;
    LogicCell40 \spi0.i10988_3_lut_4_lut_LC_14_18_3  (
            .in0(N__55254),
            .in1(N__55439),
            .in2(N__54756),
            .in3(N__55049),
            .lcout(\spi0.n12605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i8576_4_lut_4_lut_LC_14_18_4 .C_ON=1'b0;
    defparam \spi0.i8576_4_lut_4_lut_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \spi0.i8576_4_lut_4_lut_LC_14_18_4 .LUT_INIT=16'b1111010100000100;
    LogicCell40 \spi0.i8576_4_lut_4_lut_LC_14_18_4  (
            .in0(N__55051),
            .in1(N__54752),
            .in2(N__55478),
            .in3(N__55257),
            .lcout(\spi0.n10090 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i8618_4_lut_LC_14_18_5 .C_ON=1'b0;
    defparam \spi0.i8618_4_lut_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \spi0.i8618_4_lut_LC_14_18_5 .LUT_INIT=16'b1000100101000101;
    LogicCell40 \spi0.i8618_4_lut_LC_14_18_5  (
            .in0(N__55258),
            .in1(N__55590),
            .in2(N__54757),
            .in3(N__54945),
            .lcout(\spi0.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i11009_4_lut_LC_14_18_6 .C_ON=1'b0;
    defparam \spi0.i11009_4_lut_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \spi0.i11009_4_lut_LC_14_18_6 .LUT_INIT=16'b1111110000010000;
    LogicCell40 \spi0.i11009_4_lut_LC_14_18_6  (
            .in0(N__55050),
            .in1(N__55479),
            .in2(N__54951),
            .in3(N__55255),
            .lcout(),
            .ltout(\spi0.n12576_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i42_4_lut_LC_14_18_7 .C_ON=1'b0;
    defparam \spi0.i42_4_lut_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \spi0.i42_4_lut_LC_14_18_7 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \spi0.i42_4_lut_LC_14_18_7  (
            .in0(N__55256),
            .in1(N__55589),
            .in2(N__55114),
            .in3(N__54898),
            .lcout(\spi0.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i11110_3_lut_LC_14_19_0 .C_ON=1'b0;
    defparam \spi0.i11110_3_lut_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \spi0.i11110_3_lut_LC_14_19_0 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \spi0.i11110_3_lut_LC_14_19_0  (
            .in0(N__55111),
            .in1(N__55430),
            .in2(_gnd_net_),
            .in3(N__55073),
            .lcout(\spi0.n19_adj_1139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i1584_2_lut_LC_14_19_1 .C_ON=1'b0;
    defparam \spi0.i1584_2_lut_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \spi0.i1584_2_lut_LC_14_19_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \spi0.i1584_2_lut_LC_14_19_1  (
            .in0(N__55074),
            .in1(_gnd_net_),
            .in2(N__55614),
            .in3(_gnd_net_),
            .lcout(\spi0.n2768 ),
            .ltout(\spi0.n2768_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i3_4_lut_LC_14_19_2 .C_ON=1'b0;
    defparam \spi0.i3_4_lut_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \spi0.i3_4_lut_LC_14_19_2 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \spi0.i3_4_lut_LC_14_19_2  (
            .in0(N__55096),
            .in1(N__55432),
            .in2(N__55090),
            .in3(N__55087),
            .lcout(\spi0.n14414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i3253_2_lut_LC_14_19_3 .C_ON=1'b0;
    defparam \spi0.i3253_2_lut_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \spi0.i3253_2_lut_LC_14_19_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \spi0.i3253_2_lut_LC_14_19_3  (
            .in0(N__55431),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55701),
            .lcout(\spi0.n4455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i44_4_lut_LC_14_19_4 .C_ON=1'b0;
    defparam \spi0.i44_4_lut_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \spi0.i44_4_lut_LC_14_19_4 .LUT_INIT=16'b1111000000010001;
    LogicCell40 \spi0.i44_4_lut_LC_14_19_4  (
            .in0(N__58470),
            .in1(N__55075),
            .in2(N__54955),
            .in3(N__55433),
            .lcout(\spi0.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i2_2_lut_LC_14_19_5 .C_ON=1'b0;
    defparam \spi0.i2_2_lut_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \spi0.i2_2_lut_LC_14_19_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \spi0.i2_2_lut_LC_14_19_5  (
            .in0(N__55306),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55327),
            .lcout(),
            .ltout(\spi0.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i7_4_lut_adj_31_LC_14_19_6 .C_ON=1'b0;
    defparam \spi0.i7_4_lut_adj_31_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \spi0.i7_4_lut_adj_31_LC_14_19_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \spi0.i7_4_lut_adj_31_LC_14_19_6  (
            .in0(N__55288),
            .in1(N__74068),
            .in2(N__54892),
            .in3(N__55342),
            .lcout(\spi0.n1979 ),
            .ltout(\spi0.n1979_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.state_i3_LC_14_19_7 .C_ON=1'b0;
    defparam \spi0.state_i3_LC_14_19_7 .SEQ_MODE=4'b1000;
    defparam \spi0.state_i3_LC_14_19_7 .LUT_INIT=16'b1111011110100010;
    LogicCell40 \spi0.state_i3_LC_14_19_7  (
            .in0(N__55434),
            .in1(N__55607),
            .in2(N__55507),
            .in3(N__55504),
            .lcout(\spi0.state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97396),
            .ce(N__55351),
            .sr(_gnd_net_));
    defparam \spi0.multi_byte_counter_i0_LC_14_20_0 .C_ON=1'b1;
    defparam \spi0.multi_byte_counter_i0_LC_14_20_0 .SEQ_MODE=4'b1000;
    defparam \spi0.multi_byte_counter_i0_LC_14_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.multi_byte_counter_i0_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__55341),
            .in2(N__55763),
            .in3(_gnd_net_),
            .lcout(\spi0.multi_byte_counter_0 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\spi0.n10653 ),
            .clk(N__97404),
            .ce(N__55702),
            .sr(N__55687));
    defparam \spi0.multi_byte_counter_i1_LC_14_20_1 .C_ON=1'b1;
    defparam \spi0.multi_byte_counter_i1_LC_14_20_1 .SEQ_MODE=4'b1000;
    defparam \spi0.multi_byte_counter_i1_LC_14_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.multi_byte_counter_i1_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__55744),
            .in2(N__74085),
            .in3(N__55330),
            .lcout(\spi0.multi_byte_counter_1 ),
            .ltout(),
            .carryin(\spi0.n10653 ),
            .carryout(\spi0.n10654 ),
            .clk(N__97404),
            .ce(N__55702),
            .sr(N__55687));
    defparam \spi0.multi_byte_counter_i2_LC_14_20_2 .C_ON=1'b1;
    defparam \spi0.multi_byte_counter_i2_LC_14_20_2 .SEQ_MODE=4'b1000;
    defparam \spi0.multi_byte_counter_i2_LC_14_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.multi_byte_counter_i2_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__55323),
            .in2(N__55764),
            .in3(N__55312),
            .lcout(\spi0.multi_byte_counter_2 ),
            .ltout(),
            .carryin(\spi0.n10654 ),
            .carryout(\spi0.n10655 ),
            .clk(N__97404),
            .ce(N__55702),
            .sr(N__55687));
    defparam \spi0.multi_byte_counter_i3_LC_14_20_3 .C_ON=1'b1;
    defparam \spi0.multi_byte_counter_i3_LC_14_20_3 .SEQ_MODE=4'b1000;
    defparam \spi0.multi_byte_counter_i3_LC_14_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.multi_byte_counter_i3_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__55748),
            .in2(N__74109),
            .in3(N__55309),
            .lcout(\spi0.multi_byte_counter_3 ),
            .ltout(),
            .carryin(\spi0.n10655 ),
            .carryout(\spi0.n10656 ),
            .clk(N__97404),
            .ce(N__55702),
            .sr(N__55687));
    defparam \spi0.multi_byte_counter_i4_LC_14_20_4 .C_ON=1'b1;
    defparam \spi0.multi_byte_counter_i4_LC_14_20_4 .SEQ_MODE=4'b1000;
    defparam \spi0.multi_byte_counter_i4_LC_14_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.multi_byte_counter_i4_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__55305),
            .in2(N__55765),
            .in3(N__55294),
            .lcout(\spi0.multi_byte_counter_4 ),
            .ltout(),
            .carryin(\spi0.n10656 ),
            .carryout(\spi0.n10657 ),
            .clk(N__97404),
            .ce(N__55702),
            .sr(N__55687));
    defparam \spi0.multi_byte_counter_i5_LC_14_20_5 .C_ON=1'b1;
    defparam \spi0.multi_byte_counter_i5_LC_14_20_5 .SEQ_MODE=4'b1001;
    defparam \spi0.multi_byte_counter_i5_LC_14_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.multi_byte_counter_i5_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__55752),
            .in2(N__74133),
            .in3(N__55291),
            .lcout(\spi0.multi_byte_counter_5 ),
            .ltout(),
            .carryin(\spi0.n10657 ),
            .carryout(\spi0.n10658 ),
            .clk(N__97404),
            .ce(N__55702),
            .sr(N__55687));
    defparam \spi0.multi_byte_counter_i6_LC_14_20_6 .C_ON=1'b1;
    defparam \spi0.multi_byte_counter_i6_LC_14_20_6 .SEQ_MODE=4'b1000;
    defparam \spi0.multi_byte_counter_i6_LC_14_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \spi0.multi_byte_counter_i6_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(N__55284),
            .in2(N__55766),
            .in3(N__55273),
            .lcout(\spi0.multi_byte_counter_6 ),
            .ltout(),
            .carryin(\spi0.n10658 ),
            .carryout(\spi0.n10659 ),
            .clk(N__97404),
            .ce(N__55702),
            .sr(N__55687));
    defparam \spi0.multi_byte_counter_i7_LC_14_20_7 .C_ON=1'b0;
    defparam \spi0.multi_byte_counter_i7_LC_14_20_7 .SEQ_MODE=4'b1001;
    defparam \spi0.multi_byte_counter_i7_LC_14_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi0.multi_byte_counter_i7_LC_14_20_7  (
            .in0(N__74151),
            .in1(N__55756),
            .in2(_gnd_net_),
            .in3(N__55705),
            .lcout(\spi0.multi_byte_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97404),
            .ce(N__55702),
            .sr(N__55687));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13364_bdd_4_lut_LC_15_1_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13364_bdd_4_lut_LC_15_1_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13364_bdd_4_lut_LC_15_1_3 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13364_bdd_4_lut_LC_15_1_3  (
            .in0(N__85660),
            .in1(N__55678),
            .in2(N__55669),
            .in3(N__55621),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2825_2826_LC_15_2_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2825_2826_LC_15_2_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2825_2826_LC_15_2_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2825_2826_LC_15_2_0  (
            .in0(N__96582),
            .in1(N__95743),
            .in2(N__58654),
            .in3(N__71007),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93431),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4841_4842_LC_15_2_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4841_4842_LC_15_2_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4841_4842_LC_15_2_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4841_4842_LC_15_2_1  (
            .in0(N__55644),
            .in1(N__96580),
            .in2(_gnd_net_),
            .in3(N__73053),
            .lcout(REG_mem_50_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93431),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10851_3_lut_LC_15_2_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10851_3_lut_LC_15_2_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10851_3_lut_LC_15_2_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10851_3_lut_LC_15_2_2  (
            .in0(N__85659),
            .in1(N__58660),
            .in2(_gnd_net_),
            .in3(N__56002),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6089_6090_LC_15_2_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6089_6090_LC_15_2_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6089_6090_LC_15_2_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6089_6090_LC_15_2_3  (
            .in0(N__58593),
            .in1(N__96581),
            .in2(_gnd_net_),
            .in3(N__67715),
            .lcout(REG_mem_63_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93431),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10071_3_lut_LC_15_2_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10071_3_lut_LC_15_2_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10071_3_lut_LC_15_2_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10071_3_lut_LC_15_2_4  (
            .in0(N__88849),
            .in1(N__55645),
            .in2(_gnd_net_),
            .in3(N__55636),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11720 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5993_5994_LC_15_2_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5993_5994_LC_15_2_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5993_5994_LC_15_2_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5993_5994_LC_15_2_5  (
            .in0(N__95742),
            .in1(N__96584),
            .in2(N__58582),
            .in3(N__77897),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93431),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5897_5898_LC_15_2_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5897_5898_LC_15_2_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5897_5898_LC_15_2_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5897_5898_LC_15_2_6  (
            .in0(N__96583),
            .in1(N__95744),
            .in2(N__58609),
            .in3(N__71008),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93431),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13850_bdd_4_lut_LC_15_3_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13850_bdd_4_lut_LC_15_3_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13850_bdd_4_lut_LC_15_3_0 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13850_bdd_4_lut_LC_15_3_0  (
            .in0(N__92610),
            .in1(N__56098),
            .in2(N__56050),
            .in3(N__56065),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13853 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11744_LC_15_3_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11744_LC_15_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11744_LC_15_3_1 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11744_LC_15_3_1  (
            .in0(N__88885),
            .in1(N__92612),
            .in2(N__55996),
            .in3(N__58879),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11211_LC_15_3_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11211_LC_15_3_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11211_LC_15_3_2 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11211_LC_15_3_2  (
            .in0(N__92611),
            .in1(N__88884),
            .in2(N__55969),
            .in3(N__55951),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12872_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12872_bdd_4_lut_LC_15_3_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12872_bdd_4_lut_LC_15_3_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12872_bdd_4_lut_LC_15_3_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12872_bdd_4_lut_LC_15_3_3  (
            .in0(N__55930),
            .in1(N__92609),
            .in2(N__55909),
            .in3(N__55906),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12875_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10862_3_lut_LC_15_3_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10862_3_lut_LC_15_3_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10862_3_lut_LC_15_3_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10862_3_lut_LC_15_3_4  (
            .in0(N__85842),
            .in1(_gnd_net_),
            .in2(N__55882),
            .in3(N__55816),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12511_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11560_LC_15_3_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11560_LC_15_3_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11560_LC_15_3_5 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11560_LC_15_3_5  (
            .in0(N__56011),
            .in1(N__81514),
            .in2(N__55879),
            .in3(N__90301),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13250_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13250_bdd_4_lut_LC_15_3_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13250_bdd_4_lut_LC_15_3_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13250_bdd_4_lut_LC_15_3_6 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13250_bdd_4_lut_LC_15_3_6  (
            .in0(N__55876),
            .in1(N__81513),
            .in2(N__55870),
            .in3(N__55867),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13253 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13514_bdd_4_lut_LC_15_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13514_bdd_4_lut_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13514_bdd_4_lut_LC_15_4_0 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13514_bdd_4_lut_LC_15_4_0  (
            .in0(N__92176),
            .in1(N__55858),
            .in2(N__55852),
            .in3(N__55831),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10028_3_lut_LC_15_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10028_3_lut_LC_15_4_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10028_3_lut_LC_15_4_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10028_3_lut_LC_15_4_1  (
            .in0(N__55810),
            .in1(N__55789),
            .in2(_gnd_net_),
            .in3(N__88602),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12023_LC_15_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12023_LC_15_4_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12023_LC_15_4_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12023_LC_15_4_2  (
            .in0(N__88603),
            .in1(N__56116),
            .in2(N__92430),
            .in3(N__56035),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13850 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13280_bdd_4_lut_LC_15_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13280_bdd_4_lut_LC_15_4_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13280_bdd_4_lut_LC_15_4_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13280_bdd_4_lut_LC_15_4_3  (
            .in0(N__56092),
            .in1(N__92175),
            .in2(N__58957),
            .in3(N__56074),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1580_1581_LC_15_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1580_1581_LC_15_4_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1580_1581_LC_15_4_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1580_1581_LC_15_4_4  (
            .in0(N__56073),
            .in1(N__75896),
            .in2(_gnd_net_),
            .in3(N__65688),
            .lcout(REG_mem_16_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93419),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i917_918_LC_15_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i917_918_LC_15_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i917_918_LC_15_4_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i917_918_LC_15_4_5  (
            .in0(N__56061),
            .in1(N__62635),
            .in2(_gnd_net_),
            .in3(N__67188),
            .lcout(REG_mem_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93419),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i821_822_LC_15_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i821_822_LC_15_4_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i821_822_LC_15_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i821_822_LC_15_4_6  (
            .in0(N__62633),
            .in1(N__56046),
            .in2(_gnd_net_),
            .in3(N__67338),
            .lcout(REG_mem_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93419),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1013_1014_LC_15_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1013_1014_LC_15_4_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1013_1014_LC_15_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1013_1014_LC_15_4_7  (
            .in0(N__56034),
            .in1(N__62634),
            .in2(_gnd_net_),
            .in3(N__66996),
            .lcout(REG_mem_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93419),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10377_3_lut_LC_15_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10377_3_lut_LC_15_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10377_3_lut_LC_15_5_0 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10377_3_lut_LC_15_5_0  (
            .in0(N__88728),
            .in1(_gnd_net_),
            .in2(N__62470),
            .in3(N__56701),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12026_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12418_LC_15_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12418_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12418_LC_15_5_1 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12418_LC_15_5_1  (
            .in0(N__85658),
            .in1(N__56170),
            .in2(N__56026),
            .in3(N__92492),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14282_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14282_bdd_4_lut_LC_15_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14282_bdd_4_lut_LC_15_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14282_bdd_4_lut_LC_15_5_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14282_bdd_4_lut_LC_15_5_2  (
            .in0(N__56023),
            .in1(N__85657),
            .in2(N__56014),
            .in3(N__56632),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12512 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2549_2550_LC_15_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2549_2550_LC_15_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2549_2550_LC_15_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2549_2550_LC_15_5_3  (
            .in0(N__56643),
            .in1(N__62677),
            .in2(_gnd_net_),
            .in3(N__70387),
            .lcout(REG_mem_26_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93411),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i617_618_LC_15_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i617_618_LC_15_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i617_618_LC_15_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i617_618_LC_15_5_4  (
            .in0(N__59016),
            .in1(N__96694),
            .in2(_gnd_net_),
            .in3(N__66420),
            .lcout(REG_mem_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93411),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10332_3_lut_LC_15_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10332_3_lut_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10332_3_lut_LC_15_5_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10332_3_lut_LC_15_5_5  (
            .in0(N__56724),
            .in1(N__56644),
            .in2(_gnd_net_),
            .in3(N__88726),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11981 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i641_642_LC_15_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i641_642_LC_15_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i641_642_LC_15_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i641_642_LC_15_5_6  (
            .in0(N__56202),
            .in1(N__56614),
            .in2(_gnd_net_),
            .in3(N__66421),
            .lcout(REG_mem_6_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93411),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10376_3_lut_LC_15_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10376_3_lut_LC_15_5_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10376_3_lut_LC_15_5_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10376_3_lut_LC_15_5_7  (
            .in0(N__56836),
            .in1(N__88727),
            .in2(_gnd_net_),
            .in3(N__56191),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12025 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6092_6093_LC_15_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6092_6093_LC_15_6_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6092_6093_LC_15_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6092_6093_LC_15_6_0  (
            .in0(N__56160),
            .in1(N__75865),
            .in2(_gnd_net_),
            .in3(N__67700),
            .lcout(REG_mem_63_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93401),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11824_LC_15_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11824_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11824_LC_15_6_1 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11824_LC_15_6_1  (
            .in0(N__91680),
            .in1(N__56161),
            .in2(N__88773),
            .in3(N__56710),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13604_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13604_bdd_4_lut_LC_15_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13604_bdd_4_lut_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13604_bdd_4_lut_LC_15_6_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13604_bdd_4_lut_LC_15_6_2  (
            .in0(N__56128),
            .in1(N__91679),
            .in2(N__56152),
            .in3(N__56149),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5900_5901_LC_15_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5900_5901_LC_15_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5900_5901_LC_15_6_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5900_5901_LC_15_6_3  (
            .in0(N__95746),
            .in1(N__56127),
            .in2(N__75959),
            .in3(N__70999),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93401),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2645_2646_LC_15_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2645_2646_LC_15_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2645_2646_LC_15_6_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2645_2646_LC_15_6_4  (
            .in0(N__62853),
            .in1(N__95748),
            .in2(N__56725),
            .in3(N__79785),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93401),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5996_5997_LC_15_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5996_5997_LC_15_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5996_5997_LC_15_6_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5996_5997_LC_15_6_5  (
            .in0(N__95747),
            .in1(N__56709),
            .in2(N__75960),
            .in3(N__77973),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93401),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2732_2733_LC_15_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2732_2733_LC_15_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2732_2733_LC_15_6_6 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2732_2733_LC_15_6_6  (
            .in0(N__61665),
            .in1(N__95749),
            .in2(N__70720),
            .in3(N__75875),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93401),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2828_2829_LC_15_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2828_2829_LC_15_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2828_2829_LC_15_6_7 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2828_2829_LC_15_6_7  (
            .in0(N__95745),
            .in1(N__61680),
            .in2(N__75958),
            .in3(N__70998),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93401),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4268_4269_LC_15_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4268_4269_LC_15_7_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4268_4269_LC_15_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4268_4269_LC_15_7_0  (
            .in0(N__56667),
            .in1(N__75966),
            .in2(_gnd_net_),
            .in3(N__71740),
            .lcout(REG_mem_44_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93389),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3029_3030_LC_15_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3029_3030_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3029_3030_LC_15_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3029_3030_LC_15_7_1  (
            .in0(N__56697),
            .in1(N__62717),
            .in2(_gnd_net_),
            .in3(N__72535),
            .lcout(REG_mem_31_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93389),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12218_LC_15_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12218_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12218_LC_15_7_2 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12218_LC_15_7_2  (
            .in0(N__92216),
            .in1(N__88776),
            .in2(N__56656),
            .in3(N__56686),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14084_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14084_bdd_4_lut_LC_15_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14084_bdd_4_lut_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14084_bdd_4_lut_LC_15_7_3 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14084_bdd_4_lut_LC_15_7_3  (
            .in0(N__56815),
            .in1(N__56668),
            .in2(N__56659),
            .in3(N__92213),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4460_4461_LC_15_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4460_4461_LC_15_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4460_4461_LC_15_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4460_4461_LC_15_7_4  (
            .in0(N__56652),
            .in1(N__75967),
            .in2(_gnd_net_),
            .in3(N__89104),
            .lcout(REG_mem_46_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93389),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14168_bdd_4_lut_LC_15_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14168_bdd_4_lut_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14168_bdd_4_lut_LC_15_7_5 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14168_bdd_4_lut_LC_15_7_5  (
            .in0(N__56764),
            .in1(N__92214),
            .in2(N__56752),
            .in3(N__56770),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12078 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6101_6102_LC_15_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6101_6102_LC_15_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6101_6102_LC_15_7_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6101_6102_LC_15_7_6  (
            .in0(N__62716),
            .in1(N__56898),
            .in2(_gnd_net_),
            .in3(N__67696),
            .lcout(REG_mem_63_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93389),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12143_LC_15_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12143_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12143_LC_15_7_7 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12143_LC_15_7_7  (
            .in0(N__88775),
            .in1(N__92215),
            .in2(N__63085),
            .in3(N__56800),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13982 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4859_4860_LC_15_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4859_4860_LC_15_8_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4859_4860_LC_15_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4859_4860_LC_15_8_0  (
            .in0(N__59460),
            .in1(N__63377),
            .in2(_gnd_net_),
            .in3(N__73033),
            .lcout(REG_mem_50_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12288_LC_15_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12288_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12288_LC_15_8_1 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12288_LC_15_8_1  (
            .in0(N__56736),
            .in1(N__91886),
            .in2(N__61705),
            .in3(N__88354),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3980_3981_LC_15_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3980_3981_LC_15_8_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3980_3981_LC_15_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3980_3981_LC_15_8_2  (
            .in0(N__56763),
            .in1(N__75964),
            .in2(_gnd_net_),
            .in3(N__66005),
            .lcout(REG_mem_41_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3884_3885_LC_15_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3884_3885_LC_15_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3884_3885_LC_15_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3884_3885_LC_15_8_3  (
            .in0(N__75961),
            .in1(N__56748),
            .in2(_gnd_net_),
            .in3(N__65878),
            .lcout(REG_mem_40_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4574_4575_LC_15_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4574_4575_LC_15_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4574_4575_LC_15_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4574_4575_LC_15_8_4  (
            .in0(N__84837),
            .in1(N__89458),
            .in2(_gnd_net_),
            .in3(N__66266),
            .lcout(REG_mem_47_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4172_4173_LC_15_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4172_4173_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4172_4173_LC_15_8_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4172_4173_LC_15_8_5  (
            .in0(N__75962),
            .in1(_gnd_net_),
            .in2(N__56737),
            .in3(N__68278),
            .lcout(REG_mem_43_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1388_1389_LC_15_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1388_1389_LC_15_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1388_1389_LC_15_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1388_1389_LC_15_8_6  (
            .in0(N__72285),
            .in1(N__75963),
            .in2(_gnd_net_),
            .in3(N__74764),
            .lcout(REG_mem_14_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4760_4761_LC_15_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4760_4761_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4760_4761_LC_15_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4760_4761_LC_15_8_7  (
            .in0(N__75168),
            .in1(N__96370),
            .in2(_gnd_net_),
            .in3(N__62987),
            .lcout(REG_mem_49_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93376),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3710_3711_LC_15_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3710_3711_LC_15_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3710_3711_LC_15_9_0 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3710_3711_LC_15_9_0  (
            .in0(N__89454),
            .in1(_gnd_net_),
            .in2(N__63750),
            .in3(N__59248),
            .lcout(REG_mem_38_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93363),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11306_LC_15_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11306_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11306_LC_15_9_1 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11306_LC_15_9_1  (
            .in0(N__56847),
            .in1(N__56902),
            .in2(N__92212),
            .in3(N__88514),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12986_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12986_bdd_4_lut_LC_15_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12986_bdd_4_lut_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12986_bdd_4_lut_LC_15_9_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12986_bdd_4_lut_LC_15_9_2  (
            .in0(N__56859),
            .in1(N__91879),
            .in2(N__56887),
            .in3(N__56871),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12989 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5909_5910_LC_15_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5909_5910_LC_15_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5909_5910_LC_15_9_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5909_5910_LC_15_9_3  (
            .in0(N__62856),
            .in1(N__95095),
            .in2(N__56872),
            .in3(N__70977),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93363),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5813_5814_LC_15_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5813_5814_LC_15_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5813_5814_LC_15_9_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5813_5814_LC_15_9_4  (
            .in0(N__95094),
            .in1(N__62859),
            .in2(N__56860),
            .in3(N__70572),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93363),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6005_6006_LC_15_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6005_6006_LC_15_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6005_6006_LC_15_9_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6005_6006_LC_15_9_5  (
            .in0(N__62857),
            .in1(N__95096),
            .in2(N__56848),
            .in3(N__77934),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93363),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2741_2742_LC_15_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2741_2742_LC_15_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2741_2742_LC_15_9_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2741_2742_LC_15_9_6  (
            .in0(N__95093),
            .in1(N__62858),
            .in2(N__56832),
            .in3(N__70571),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93363),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4364_4365_LC_15_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4364_4365_LC_15_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4364_4365_LC_15_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4364_4365_LC_15_9_7  (
            .in0(N__75965),
            .in1(N__56811),
            .in2(_gnd_net_),
            .in3(N__71863),
            .lcout(REG_mem_45_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93363),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11311_LC_15_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11311_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11311_LC_15_10_0 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11311_LC_15_10_0  (
            .in0(N__91291),
            .in1(N__88512),
            .in2(N__57094),
            .in3(N__57070),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12992_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12992_bdd_4_lut_LC_15_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12992_bdd_4_lut_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12992_bdd_4_lut_LC_15_10_1 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12992_bdd_4_lut_LC_15_10_1  (
            .in0(N__57049),
            .in1(N__91288),
            .in2(N__57031),
            .in3(N__57028),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12995 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11415_LC_15_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11415_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11415_LC_15_10_2 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11415_LC_15_10_2  (
            .in0(N__91292),
            .in1(N__88513),
            .in2(N__57010),
            .in3(N__68149),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13118_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13118_bdd_4_lut_LC_15_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13118_bdd_4_lut_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13118_bdd_4_lut_LC_15_10_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13118_bdd_4_lut_LC_15_10_3  (
            .in0(N__61912),
            .in1(N__91289),
            .in2(N__56992),
            .in3(N__56989),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13121_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12098_LC_15_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12098_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12098_LC_15_10_4 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12098_LC_15_10_4  (
            .in0(N__56971),
            .in1(N__90343),
            .in2(N__56965),
            .in3(N__85540),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13622_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13622_bdd_4_lut_LC_15_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13622_bdd_4_lut_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13622_bdd_4_lut_LC_15_10_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13622_bdd_4_lut_LC_15_10_5  (
            .in0(N__90342),
            .in1(N__64228),
            .in2(N__56962),
            .in3(N__56929),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13178_bdd_4_lut_LC_15_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13178_bdd_4_lut_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13178_bdd_4_lut_LC_15_10_6 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13178_bdd_4_lut_LC_15_10_6  (
            .in0(N__91290),
            .in1(N__59296),
            .in2(N__56959),
            .in3(N__56944),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9903_3_lut_LC_15_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9903_3_lut_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9903_3_lut_LC_15_11_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9903_3_lut_LC_15_11_0  (
            .in0(N__88247),
            .in1(N__56923),
            .in2(_gnd_net_),
            .in3(N__57157),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11552 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12118_LC_15_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12118_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12118_LC_15_11_1 .LUT_INIT=16'b1011110010110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12118_LC_15_11_1  (
            .in0(N__56911),
            .in1(N__85523),
            .in2(N__91878),
            .in3(N__59503),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13934_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13934_bdd_4_lut_LC_15_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13934_bdd_4_lut_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13934_bdd_4_lut_LC_15_11_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13934_bdd_4_lut_LC_15_11_2  (
            .in0(N__85522),
            .in1(N__57127),
            .in2(N__57166),
            .in3(N__57163),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13937 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1010_1011_LC_15_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1010_1011_LC_15_11_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1010_1011_LC_15_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1010_1011_LC_15_11_3  (
            .in0(N__57156),
            .in1(N__76710),
            .in2(_gnd_net_),
            .in3(N__66915),
            .lcout(REG_mem_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93364),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13796_bdd_4_lut_LC_15_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13796_bdd_4_lut_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13796_bdd_4_lut_LC_15_11_4 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13796_bdd_4_lut_LC_15_11_4  (
            .in0(N__85521),
            .in1(N__57148),
            .in2(N__57142),
            .in3(N__57133),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13799 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9902_3_lut_LC_15_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9902_3_lut_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9902_3_lut_LC_15_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9902_3_lut_LC_15_11_5  (
            .in0(N__57121),
            .in1(N__57112),
            .in2(_gnd_net_),
            .in3(N__88246),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i818_819_LC_15_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i818_819_LC_15_11_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i818_819_LC_15_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i818_819_LC_15_11_6  (
            .in0(N__76709),
            .in1(N__57120),
            .in2(_gnd_net_),
            .in3(N__67339),
            .lcout(REG_mem_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93364),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i914_915_LC_15_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i914_915_LC_15_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i914_915_LC_15_11_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i914_915_LC_15_11_7  (
            .in0(N__57111),
            .in1(N__76711),
            .in2(_gnd_net_),
            .in3(N__67187),
            .lcout(REG_mem_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93364),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i1571_3_lut_4_lut_LC_15_12_0 .C_ON=1'b0;
    defparam \usb3_if_inst.i1571_3_lut_4_lut_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i1571_3_lut_4_lut_LC_15_12_0 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \usb3_if_inst.i1571_3_lut_4_lut_LC_15_12_0  (
            .in0(N__57225),
            .in1(N__57388),
            .in2(N__57646),
            .in3(N__64360),
            .lcout(),
            .ltout(\usb3_if_inst.n2755_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i1_4_lut_adj_17_LC_15_12_1 .C_ON=1'b0;
    defparam \usb3_if_inst.i1_4_lut_adj_17_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i1_4_lut_adj_17_LC_15_12_1 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \usb3_if_inst.i1_4_lut_adj_17_LC_15_12_1  (
            .in0(N__64361),
            .in1(N__57637),
            .in2(N__57100),
            .in3(N__64144),
            .lcout(),
            .ltout(\usb3_if_inst.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.state_FSM_i2_LC_15_12_2 .C_ON=1'b0;
    defparam \usb3_if_inst.state_FSM_i2_LC_15_12_2 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.state_FSM_i2_LC_15_12_2 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \usb3_if_inst.state_FSM_i2_LC_15_12_2  (
            .in0(N__57655),
            .in1(N__57187),
            .in2(N__57097),
            .in3(N__64519),
            .lcout(\usb3_if_inst.n554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_FSM_i2C_net ),
            .ce(),
            .sr(N__73689));
    defparam \usb3_if_inst.state_FSM_i4_LC_15_12_3 .C_ON=1'b0;
    defparam \usb3_if_inst.state_FSM_i4_LC_15_12_3 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.state_FSM_i4_LC_15_12_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \usb3_if_inst.state_FSM_i4_LC_15_12_3  (
            .in0(N__64362),
            .in1(N__57638),
            .in2(N__57399),
            .in3(N__57226),
            .lcout(\usb3_if_inst.n552 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_FSM_i2C_net ),
            .ce(),
            .sr(N__73689));
    defparam \usb3_if_inst.i1612_2_lut_3_lut_4_lut_LC_15_12_4 .C_ON=1'b0;
    defparam \usb3_if_inst.i1612_2_lut_3_lut_4_lut_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i1612_2_lut_3_lut_4_lut_LC_15_12_4 .LUT_INIT=16'b1000100010001010;
    LogicCell40 \usb3_if_inst.i1612_2_lut_3_lut_4_lut_LC_15_12_4  (
            .in0(N__57224),
            .in1(N__57386),
            .in2(N__57647),
            .in3(N__64359),
            .lcout(\usb3_if_inst.n2798 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i2_3_lut_LC_15_12_5 .C_ON=1'b0;
    defparam \usb3_if_inst.i2_3_lut_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i2_3_lut_LC_15_12_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \usb3_if_inst.i2_3_lut_LC_15_12_5  (
            .in0(N__57387),
            .in1(N__57751),
            .in2(_gnd_net_),
            .in3(N__64076),
            .lcout(\usb3_if_inst.n3973 ),
            .ltout(\usb3_if_inst.n3973_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.state_FSM_i1_LC_15_12_6 .C_ON=1'b0;
    defparam \usb3_if_inst.state_FSM_i1_LC_15_12_6 .SEQ_MODE=4'b1001;
    defparam \usb3_if_inst.state_FSM_i1_LC_15_12_6 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \usb3_if_inst.state_FSM_i1_LC_15_12_6  (
            .in0(N__57775),
            .in1(N__57667),
            .in2(N__57181),
            .in3(N__64518),
            .lcout(\usb3_if_inst.n555 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_FSM_i2C_net ),
            .ce(),
            .sr(N__73689));
    defparam \usb3_if_inst.i2_3_lut_4_lut_adj_20_LC_15_12_7 .C_ON=1'b0;
    defparam \usb3_if_inst.i2_3_lut_4_lut_adj_20_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i2_3_lut_4_lut_adj_20_LC_15_12_7 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \usb3_if_inst.i2_3_lut_4_lut_adj_20_LC_15_12_7  (
            .in0(N__64358),
            .in1(N__73690),
            .in2(N__57648),
            .in3(N__64145),
            .lcout(\usb3_if_inst.n10751 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.state_timeout_counter_i0_i2_LC_15_13_0 .C_ON=1'b0;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i2_LC_15_13_0 .SEQ_MODE=4'b1001;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i2_LC_15_13_0 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \bluejay_data_inst.state_timeout_counter_i0_i2_LC_15_13_0  (
            .in0(N__59857),
            .in1(_gnd_net_),
            .in2(N__68598),
            .in3(N__64681),
            .lcout(\bluejay_data_inst.state_timeout_counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97359),
            .ce(N__69170),
            .sr(N__58159));
    defparam \bluejay_data_inst.i1_2_lut_adj_66_LC_15_13_1 .C_ON=1'b0;
    defparam \bluejay_data_inst.i1_2_lut_adj_66_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i1_2_lut_adj_66_LC_15_13_1 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \bluejay_data_inst.i1_2_lut_adj_66_LC_15_13_1  (
            .in0(N__59953),
            .in1(N__60001),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\bluejay_data_inst.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i4_4_lut_LC_15_13_2 .C_ON=1'b0;
    defparam \bluejay_data_inst.i4_4_lut_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i4_4_lut_LC_15_13_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \bluejay_data_inst.i4_4_lut_LC_15_13_2  (
            .in0(N__59868),
            .in1(N__59980),
            .in2(N__57169),
            .in3(N__59893),
            .lcout(\bluejay_data_inst.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i1_2_lut_LC_15_13_3 .C_ON=1'b0;
    defparam \bluejay_data_inst.i1_2_lut_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i1_2_lut_LC_15_13_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \bluejay_data_inst.i1_2_lut_LC_15_13_3  (
            .in0(N__73538),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68575),
            .lcout(\bluejay_data_inst.n11177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i2_3_lut_adj_14_LC_15_13_4 .C_ON=1'b0;
    defparam \usb3_if_inst.i2_3_lut_adj_14_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i2_3_lut_adj_14_LC_15_13_4 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \usb3_if_inst.i2_3_lut_adj_14_LC_15_13_4  (
            .in0(N__68579),
            .in1(N__57749),
            .in2(_gnd_net_),
            .in3(N__57625),
            .lcout(\usb3_if_inst.n10869 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i3_4_lut_adj_18_LC_15_13_5 .C_ON=1'b0;
    defparam \usb3_if_inst.i3_4_lut_adj_18_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i3_4_lut_adj_18_LC_15_13_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \usb3_if_inst.i3_4_lut_adj_18_LC_15_13_5  (
            .in0(N__57750),
            .in1(N__68580),
            .in2(N__57645),
            .in3(N__57666),
            .lcout(\usb3_if_inst.n10746 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i6182_2_lut_LC_15_13_6 .C_ON=1'b0;
    defparam \usb3_if_inst.i6182_2_lut_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i6182_2_lut_LC_15_13_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \usb3_if_inst.i6182_2_lut_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__57629),
            .in2(_gnd_net_),
            .in3(N__64353),
            .lcout(\usb3_if_inst.n7360 ),
            .ltout(\usb3_if_inst.n7360_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i6327_2_lut_3_lut_4_lut_LC_15_13_7 .C_ON=1'b0;
    defparam \usb3_if_inst.i6327_2_lut_3_lut_4_lut_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i6327_2_lut_3_lut_4_lut_LC_15_13_7 .LUT_INIT=16'b0110011000000110;
    LogicCell40 \usb3_if_inst.i6327_2_lut_3_lut_4_lut_LC_15_13_7  (
            .in0(N__57502),
            .in1(N__57463),
            .in2(N__57457),
            .in3(N__57398),
            .lcout(\usb3_if_inst.n7505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i16_LC_15_14_0 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i16_LC_15_14_0 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i16_LC_15_14_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i16_LC_15_14_0  (
            .in0(N__68988),
            .in1(N__68906),
            .in2(_gnd_net_),
            .in3(N__58252),
            .lcout(DATA15_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i16C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i1_2_lut_adj_67_LC_15_14_1 .C_ON=1'b0;
    defparam \bluejay_data_inst.i1_2_lut_adj_67_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i1_2_lut_adj_67_LC_15_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \bluejay_data_inst.i1_2_lut_adj_67_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__68991),
            .in2(_gnd_net_),
            .in3(N__68904),
            .lcout(\bluejay_data_inst.valid_N_707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i1_3_lut_LC_15_14_2 .C_ON=1'b0;
    defparam \usb3_if_inst.i1_3_lut_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i1_3_lut_LC_15_14_2 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \usb3_if_inst.i1_3_lut_LC_15_14_2  (
            .in0(N__73691),
            .in1(N__64081),
            .in2(_gnd_net_),
            .in3(N__57400),
            .lcout(\usb3_if_inst.n4178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i1_LC_15_14_3 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i1_LC_15_14_3 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i1_LC_15_14_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i1_LC_15_14_3  (
            .in0(N__57322),
            .in1(N__68989),
            .in2(_gnd_net_),
            .in3(N__68903),
            .lcout(DATA16_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i16C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i1_2_lut_adj_58_LC_15_14_4 .C_ON=1'b0;
    defparam \bluejay_data_inst.i1_2_lut_adj_58_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i1_2_lut_adj_58_LC_15_14_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \bluejay_data_inst.i1_2_lut_adj_58_LC_15_14_4  (
            .in0(N__68990),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69155),
            .lcout(\bluejay_data_inst.n4522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i12_LC_15_14_5 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i12_LC_15_14_5 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i12_LC_15_14_5 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i12_LC_15_14_5  (
            .in0(N__58153),
            .in1(N__68987),
            .in2(_gnd_net_),
            .in3(N__68902),
            .lcout(DATA11_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i16C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i11_LC_15_14_6 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i11_LC_15_14_6 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i11_LC_15_14_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i11_LC_15_14_6  (
            .in0(N__68986),
            .in1(N__68905),
            .in2(_gnd_net_),
            .in3(N__58102),
            .lcout(DATA10_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i16C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i10_LC_15_14_7 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i10_LC_15_14_7 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i10_LC_15_14_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i10_LC_15_14_7  (
            .in0(N__57789),
            .in1(N__68985),
            .in2(_gnd_net_),
            .in3(N__68901),
            .lcout(DATA9_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i16C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.tx_shift_reg_i0_i0_LC_15_15_0 .C_ON=1'b0;
    defparam \spi0.tx_shift_reg_i0_i0_LC_15_15_0 .SEQ_MODE=4'b1000;
    defparam \spi0.tx_shift_reg_i0_i0_LC_15_15_0 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \spi0.tx_shift_reg_i0_i0_LC_15_15_0  (
            .in0(N__58024),
            .in1(N__57942),
            .in2(N__57987),
            .in3(N__57931),
            .lcout(tx_shift_reg_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97374),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.mux_946_i16_3_lut_LC_15_15_1 .C_ON=1'b0;
    defparam \spi0.mux_946_i16_3_lut_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \spi0.mux_946_i16_3_lut_LC_15_15_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi0.mux_946_i16_3_lut_LC_15_15_1  (
            .in0(N__57930),
            .in1(N__58432),
            .in2(_gnd_net_),
            .in3(N__57862),
            .lcout(\spi0.n1930 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i12_LC_15_15_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i12_LC_15_15_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i12_LC_15_15_2 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i12_LC_15_15_2  (
            .in0(N__80826),
            .in1(N__73298),
            .in2(N__57835),
            .in3(N__68433),
            .lcout(fifo_data_out_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97374),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_data_byte_r_i0_i7_LC_15_15_3.C_ON=1'b0;
    defparam tx_data_byte_r_i0_i7_LC_15_15_3.SEQ_MODE=4'b1000;
    defparam tx_data_byte_r_i0_i7_LC_15_15_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 tx_data_byte_r_i0_i7_LC_15_15_3 (
            .in0(N__69402),
            .in1(N__58450),
            .in2(_gnd_net_),
            .in3(N__57819),
            .lcout(tx_data_byte_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97374),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i9_LC_15_15_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i9_LC_15_15_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i9_LC_15_15_4 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i9_LC_15_15_4  (
            .in0(N__80830),
            .in1(N__73302),
            .in2(N__57793),
            .in3(N__57805),
            .lcout(fifo_data_out_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97374),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i3_LC_15_15_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i3_LC_15_15_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i3_LC_15_15_5 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i3_LC_15_15_5  (
            .in0(N__73300),
            .in1(N__80828),
            .in2(N__58285),
            .in3(N__65532),
            .lcout(fifo_data_out_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97374),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i8_LC_15_15_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i8_LC_15_15_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i8_LC_15_15_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i8_LC_15_15_6  (
            .in0(N__80829),
            .in1(N__73301),
            .in2(N__80902),
            .in3(N__65088),
            .lcout(fifo_data_out_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97374),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i15_LC_15_15_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i15_LC_15_15_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i15_LC_15_15_7 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i15_LC_15_15_7  (
            .in0(N__73299),
            .in1(N__80827),
            .in2(N__58267),
            .in3(N__58251),
            .lcout(fifo_data_out_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97374),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_Rx_Byte_i6_LC_15_16_0 .C_ON=1'b0;
    defparam \pc_rx.r_Rx_Byte_i6_LC_15_16_0 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Rx_Byte_i6_LC_15_16_0 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \pc_rx.r_Rx_Byte_i6_LC_15_16_0  (
            .in0(N__60701),
            .in1(N__58239),
            .in2(N__58306),
            .in3(N__58186),
            .lcout(pc_data_rx_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97381),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_Rx_Byte_i4_LC_15_16_1 .C_ON=1'b0;
    defparam \pc_rx.r_Rx_Byte_i4_LC_15_16_1 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Rx_Byte_i4_LC_15_16_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \pc_rx.r_Rx_Byte_i4_LC_15_16_1  (
            .in0(N__58185),
            .in1(N__60700),
            .in2(N__58401),
            .in3(N__58335),
            .lcout(pc_data_rx_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97381),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_addr_byte_r_i0_i2_LC_15_16_2.C_ON=1'b0;
    defparam tx_addr_byte_r_i0_i2_LC_15_16_2.SEQ_MODE=4'b1000;
    defparam tx_addr_byte_r_i0_i2_LC_15_16_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 tx_addr_byte_r_i0_i2_LC_15_16_2 (
            .in0(N__58226),
            .in1(N__69400),
            .in2(_gnd_net_),
            .in3(N__58197),
            .lcout(tx_addr_byte_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97381),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.Rx_Recv_Byte_i4_LC_15_16_3 .C_ON=1'b0;
    defparam \spi0.Rx_Recv_Byte_i4_LC_15_16_3 .SEQ_MODE=4'b1000;
    defparam \spi0.Rx_Recv_Byte_i4_LC_15_16_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.Rx_Recv_Byte_i4_LC_15_16_3  (
            .in0(N__69749),
            .in1(N__64945),
            .in2(_gnd_net_),
            .in3(N__65161),
            .lcout(rx_buf_byte_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97381),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_Rx_Byte_i2_LC_15_16_4 .C_ON=1'b0;
    defparam \pc_rx.r_Rx_Byte_i2_LC_15_16_4 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Rx_Byte_i2_LC_15_16_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \pc_rx.r_Rx_Byte_i2_LC_15_16_4  (
            .in0(N__60699),
            .in1(N__60147),
            .in2(N__58174),
            .in3(N__58184),
            .lcout(pc_data_rx_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97381),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.buffer_switch_done_latched_81_LC_15_16_5 .C_ON=1'b0;
    defparam \usb3_if_inst.buffer_switch_done_latched_81_LC_15_16_5 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.buffer_switch_done_latched_81_LC_15_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.buffer_switch_done_latched_81_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73558),
            .lcout(buffer_switch_done_latched),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97381),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_Rx_Byte_i1_LC_15_16_6 .C_ON=1'b0;
    defparam \pc_rx.r_Rx_Byte_i1_LC_15_16_6 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Rx_Byte_i1_LC_15_16_6 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \pc_rx.r_Rx_Byte_i1_LC_15_16_6  (
            .in0(N__60698),
            .in1(N__58413),
            .in2(N__60168),
            .in3(N__58320),
            .lcout(pc_data_rx_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97381),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_data_byte_r_i0_i4_LC_15_16_7.C_ON=1'b0;
    defparam tx_data_byte_r_i0_i4_LC_15_16_7.SEQ_MODE=4'b1000;
    defparam tx_data_byte_r_i0_i4_LC_15_16_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 tx_data_byte_r_i0_i4_LC_15_16_7 (
            .in0(N__69401),
            .in1(_gnd_net_),
            .in2(N__58402),
            .in3(N__69433),
            .lcout(tx_data_byte_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97381),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i6_LC_15_17_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i6_LC_15_17_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i6_LC_15_17_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i6_LC_15_17_0  (
            .in0(N__58387),
            .in1(N__81037),
            .in2(_gnd_net_),
            .in3(N__58366),
            .lcout(REG_out_raw_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97388),
            .ce(N__80835),
            .sr(_gnd_net_));
    defparam \pc_rx.i5315_3_lut_LC_15_17_1 .C_ON=1'b0;
    defparam \pc_rx.i5315_3_lut_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i5315_3_lut_LC_15_17_1 .LUT_INIT=16'b0110011000100010;
    LogicCell40 \pc_rx.i5315_3_lut_LC_15_17_1  (
            .in0(N__60780),
            .in1(N__60229),
            .in2(_gnd_net_),
            .in3(N__58291),
            .lcout(\pc_rx.n6515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.equal_137_i4_2_lut_LC_15_17_2 .C_ON=1'b0;
    defparam \pc_rx.equal_137_i4_2_lut_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \pc_rx.equal_137_i4_2_lut_LC_15_17_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \pc_rx.equal_137_i4_2_lut_LC_15_17_2  (
            .in0(N__60102),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60039),
            .lcout(n4_adj_1205),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.equal_140_i4_2_lut_LC_15_17_3 .C_ON=1'b0;
    defparam \pc_rx.equal_140_i4_2_lut_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \pc_rx.equal_140_i4_2_lut_LC_15_17_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \pc_rx.equal_140_i4_2_lut_LC_15_17_3  (
            .in0(N__60040),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60103),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.equal_142_i4_2_lut_LC_15_17_4 .C_ON=1'b0;
    defparam \pc_rx.equal_142_i4_2_lut_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \pc_rx.equal_142_i4_2_lut_LC_15_17_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \pc_rx.equal_142_i4_2_lut_LC_15_17_4  (
            .in0(N__60104),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60041),
            .lcout(n4_adj_1206),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i6277_2_lut_LC_15_17_5 .C_ON=1'b0;
    defparam \pc_rx.i6277_2_lut_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i6277_2_lut_LC_15_17_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pc_rx.i6277_2_lut_LC_15_17_5  (
            .in0(N__60043),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60106),
            .lcout(n7455),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i2_2_lut_3_lut_LC_15_17_6 .C_ON=1'b0;
    defparam \pc_rx.i2_2_lut_3_lut_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i2_2_lut_3_lut_LC_15_17_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pc_rx.i2_2_lut_3_lut_LC_15_17_6  (
            .in0(N__60105),
            .in1(N__60072),
            .in2(_gnd_net_),
            .in3(N__60042),
            .lcout(\pc_rx.n149 ),
            .ltout(\pc_rx.n149_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i3268_3_lut_LC_15_17_7 .C_ON=1'b0;
    defparam \pc_rx.i3268_3_lut_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i3268_3_lut_LC_15_17_7 .LUT_INIT=16'b1111001100000000;
    LogicCell40 \pc_rx.i3268_3_lut_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__60356),
            .in2(N__58522),
            .in3(N__60407),
            .lcout(\pc_rx.n4470 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i5281_4_lut_4_lut_LC_15_18_0 .C_ON=1'b0;
    defparam \pc_rx.i5281_4_lut_4_lut_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i5281_4_lut_4_lut_LC_15_18_0 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \pc_rx.i5281_4_lut_4_lut_LC_15_18_0  (
            .in0(N__60300),
            .in1(N__60225),
            .in2(N__60649),
            .in3(N__60351),
            .lcout(\pc_rx.n6481 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_Rx_DV_52_LC_15_18_1 .C_ON=1'b0;
    defparam \pc_rx.r_Rx_DV_52_LC_15_18_1 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Rx_DV_52_LC_15_18_1 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \pc_rx.r_Rx_DV_52_LC_15_18_1  (
            .in0(N__58517),
            .in1(N__60301),
            .in2(N__60424),
            .in3(N__60352),
            .lcout(debug_led3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97397),
            .ce(),
            .sr(_gnd_net_));
    defparam uart_rx_complete_prev_83_LC_15_18_2.C_ON=1'b0;
    defparam uart_rx_complete_prev_83_LC_15_18_2.SEQ_MODE=4'b1000;
    defparam uart_rx_complete_prev_83_LC_15_18_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 uart_rx_complete_prev_83_LC_15_18_2 (
            .in0(_gnd_net_),
            .in1(N__58518),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uart_rx_complete_prev),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97397),
            .ce(),
            .sr(_gnd_net_));
    defparam uart_rx_complete_rising_edge_82_LC_15_18_3.C_ON=1'b0;
    defparam uart_rx_complete_rising_edge_82_LC_15_18_3.SEQ_MODE=4'b1000;
    defparam uart_rx_complete_rising_edge_82_LC_15_18_3.LUT_INIT=16'b0000000010101010;
    LogicCell40 uart_rx_complete_rising_edge_82_LC_15_18_3 (
            .in0(N__58519),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58507),
            .lcout(uart_rx_complete_rising_edge),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97397),
            .ce(),
            .sr(_gnd_net_));
    defparam even_byte_flag_89_LC_15_18_4.C_ON=1'b0;
    defparam even_byte_flag_89_LC_15_18_4.SEQ_MODE=4'b1000;
    defparam even_byte_flag_89_LC_15_18_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 even_byte_flag_89_LC_15_18_4 (
            .in0(_gnd_net_),
            .in1(N__69366),
            .in2(_gnd_net_),
            .in3(N__58490),
            .lcout(even_byte_flag),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97397),
            .ce(),
            .sr(_gnd_net_));
    defparam i3241_1_lut_2_lut_LC_15_18_5.C_ON=1'b0;
    defparam i3241_1_lut_2_lut_LC_15_18_5.SEQ_MODE=4'b0000;
    defparam i3241_1_lut_2_lut_LC_15_18_5.LUT_INIT=16'b0101111101011111;
    LogicCell40 i3241_1_lut_2_lut_LC_15_18_5 (
            .in0(N__69367),
            .in1(_gnd_net_),
            .in2(N__58495),
            .in3(_gnd_net_),
            .lcout(n4443),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam spi_start_transfer_r_84_LC_15_18_6.C_ON=1'b0;
    defparam spi_start_transfer_r_84_LC_15_18_6.SEQ_MODE=4'b1000;
    defparam spi_start_transfer_r_84_LC_15_18_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 spi_start_transfer_r_84_LC_15_18_6 (
            .in0(_gnd_net_),
            .in1(N__69368),
            .in2(_gnd_net_),
            .in3(N__58494),
            .lcout(spi_start_transfer_r),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97397),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_addr_byte_r_i0_i7_LC_15_18_7.C_ON=1'b0;
    defparam tx_addr_byte_r_i0_i7_LC_15_18_7.SEQ_MODE=4'b1000;
    defparam tx_addr_byte_r_i0_i7_LC_15_18_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 tx_addr_byte_r_i0_i7_LC_15_18_7 (
            .in0(N__69369),
            .in1(N__58458),
            .in2(_gnd_net_),
            .in3(N__58425),
            .lcout(tx_addr_byte_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97397),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_Clock_Count_1111__i0_LC_15_19_0 .C_ON=1'b1;
    defparam \pc_rx.r_Clock_Count_1111__i0_LC_15_19_0 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Clock_Count_1111__i0_LC_15_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_rx.r_Clock_Count_1111__i0_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__60515),
            .in2(_gnd_net_),
            .in3(N__58552),
            .lcout(\pc_rx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\pc_rx.n10703 ),
            .clk(N__97405),
            .ce(N__60435),
            .sr(N__58713));
    defparam \pc_rx.r_Clock_Count_1111__i1_LC_15_19_1 .C_ON=1'b1;
    defparam \pc_rx.r_Clock_Count_1111__i1_LC_15_19_1 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Clock_Count_1111__i1_LC_15_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_rx.r_Clock_Count_1111__i1_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__60533),
            .in2(_gnd_net_),
            .in3(N__58549),
            .lcout(\pc_rx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\pc_rx.n10703 ),
            .carryout(\pc_rx.n10704 ),
            .clk(N__97405),
            .ce(N__60435),
            .sr(N__58713));
    defparam \pc_rx.r_Clock_Count_1111__i2_LC_15_19_2 .C_ON=1'b1;
    defparam \pc_rx.r_Clock_Count_1111__i2_LC_15_19_2 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Clock_Count_1111__i2_LC_15_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_rx.r_Clock_Count_1111__i2_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__60473),
            .in2(_gnd_net_),
            .in3(N__58546),
            .lcout(\pc_rx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\pc_rx.n10704 ),
            .carryout(\pc_rx.n10705 ),
            .clk(N__97405),
            .ce(N__60435),
            .sr(N__58713));
    defparam \pc_rx.r_Clock_Count_1111__i3_LC_15_19_3 .C_ON=1'b1;
    defparam \pc_rx.r_Clock_Count_1111__i3_LC_15_19_3 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Clock_Count_1111__i3_LC_15_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_rx.r_Clock_Count_1111__i3_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(N__60500),
            .in2(_gnd_net_),
            .in3(N__58543),
            .lcout(\pc_rx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\pc_rx.n10705 ),
            .carryout(\pc_rx.n10706 ),
            .clk(N__97405),
            .ce(N__60435),
            .sr(N__58713));
    defparam \pc_rx.r_Clock_Count_1111__i4_LC_15_19_4 .C_ON=1'b1;
    defparam \pc_rx.r_Clock_Count_1111__i4_LC_15_19_4 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Clock_Count_1111__i4_LC_15_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_rx.r_Clock_Count_1111__i4_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__60548),
            .in2(_gnd_net_),
            .in3(N__58540),
            .lcout(\pc_rx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\pc_rx.n10706 ),
            .carryout(\pc_rx.n10707 ),
            .clk(N__97405),
            .ce(N__60435),
            .sr(N__58713));
    defparam \pc_rx.r_Clock_Count_1111__i5_LC_15_19_5 .C_ON=1'b1;
    defparam \pc_rx.r_Clock_Count_1111__i5_LC_15_19_5 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Clock_Count_1111__i5_LC_15_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_rx.r_Clock_Count_1111__i5_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__60243),
            .in2(_gnd_net_),
            .in3(N__58537),
            .lcout(\pc_rx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\pc_rx.n10707 ),
            .carryout(\pc_rx.n10708 ),
            .clk(N__97405),
            .ce(N__60435),
            .sr(N__58713));
    defparam \pc_rx.r_Clock_Count_1111__i6_LC_15_19_6 .C_ON=1'b1;
    defparam \pc_rx.r_Clock_Count_1111__i6_LC_15_19_6 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Clock_Count_1111__i6_LC_15_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_rx.r_Clock_Count_1111__i6_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(N__60255),
            .in2(_gnd_net_),
            .in3(N__58534),
            .lcout(\pc_rx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\pc_rx.n10708 ),
            .carryout(\pc_rx.n10709 ),
            .clk(N__97405),
            .ce(N__60435),
            .sr(N__58713));
    defparam \pc_rx.r_Clock_Count_1111__i7_LC_15_19_7 .C_ON=1'b1;
    defparam \pc_rx.r_Clock_Count_1111__i7_LC_15_19_7 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Clock_Count_1111__i7_LC_15_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_rx.r_Clock_Count_1111__i7_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__60567),
            .in2(_gnd_net_),
            .in3(N__58531),
            .lcout(\pc_rx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(\pc_rx.n10709 ),
            .carryout(\pc_rx.n10710 ),
            .clk(N__97405),
            .ce(N__60435),
            .sr(N__58713));
    defparam \pc_rx.r_Clock_Count_1111__i8_LC_15_20_0 .C_ON=1'b1;
    defparam \pc_rx.r_Clock_Count_1111__i8_LC_15_20_0 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Clock_Count_1111__i8_LC_15_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_rx.r_Clock_Count_1111__i8_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(N__60579),
            .in2(_gnd_net_),
            .in3(N__58528),
            .lcout(\pc_rx.r_Clock_Count_8 ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\pc_rx.n10711 ),
            .clk(N__97417),
            .ce(N__60442),
            .sr(N__58714));
    defparam \pc_rx.r_Clock_Count_1111__i9_LC_15_20_1 .C_ON=1'b0;
    defparam \pc_rx.r_Clock_Count_1111__i9_LC_15_20_1 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Clock_Count_1111__i9_LC_15_20_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pc_rx.r_Clock_Count_1111__i9_LC_15_20_1  (
            .in0(N__60270),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58525),
            .lcout(\pc_rx.r_Clock_Count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97417),
            .ce(N__60442),
            .sr(N__58714));
    defparam \usb3_if_inst.usb3_data_in_latched__i8_LC_16_1_2 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i8_LC_16_1_2 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i8_LC_16_1_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i8_LC_16_1_2  (
            .in0(N__58696),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\usb3_if_inst.usb3_data_in_latched_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93446),
            .ce(),
            .sr(N__73711));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14018_bdd_4_lut_LC_16_2_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14018_bdd_4_lut_LC_16_2_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14018_bdd_4_lut_LC_16_2_0 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14018_bdd_4_lut_LC_16_2_0  (
            .in0(N__58684),
            .in1(N__92581),
            .in2(N__58741),
            .in3(N__59716),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14021 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10046_3_lut_LC_16_2_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10046_3_lut_LC_16_2_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10046_3_lut_LC_16_2_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10046_3_lut_LC_16_2_1  (
            .in0(N__58653),
            .in1(N__88853),
            .in2(_gnd_net_),
            .in3(N__58639),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11695 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10047_3_lut_LC_16_2_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10047_3_lut_LC_16_2_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10047_3_lut_LC_16_2_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10047_3_lut_LC_16_2_2  (
            .in0(N__88854),
            .in1(_gnd_net_),
            .in2(N__58567),
            .in3(N__58936),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11696_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12138_LC_16_2_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12138_LC_16_2_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12138_LC_16_2_3 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12138_LC_16_2_3  (
            .in0(N__85861),
            .in1(N__58618),
            .in2(N__58612),
            .in3(N__92582),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13988 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10091_3_lut_LC_16_2_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10091_3_lut_LC_16_2_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10091_3_lut_LC_16_2_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10091_3_lut_LC_16_2_4  (
            .in0(N__88855),
            .in1(N__58608),
            .in2(_gnd_net_),
            .in3(N__58860),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11740 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10092_3_lut_LC_16_2_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10092_3_lut_LC_16_2_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10092_3_lut_LC_16_2_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10092_3_lut_LC_16_2_5  (
            .in0(N__58594),
            .in1(N__58581),
            .in2(_gnd_net_),
            .in3(N__88856),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2921_2922_LC_16_2_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2921_2922_LC_16_2_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2921_2922_LC_16_2_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2921_2922_LC_16_2_6  (
            .in0(N__96573),
            .in1(N__95752),
            .in2(N__58566),
            .in3(N__77937),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93437),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5801_5802_LC_16_2_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5801_5802_LC_16_2_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5801_5802_LC_16_2_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5801_5802_LC_16_2_7  (
            .in0(N__95751),
            .in1(N__96574),
            .in2(N__58861),
            .in3(N__70718),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93437),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10077_3_lut_LC_16_3_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10077_3_lut_LC_16_3_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10077_3_lut_LC_16_3_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10077_3_lut_LC_16_3_0  (
            .in0(N__58797),
            .in1(N__88325),
            .in2(_gnd_net_),
            .in3(N__58807),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11726 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12088_LC_16_3_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12088_LC_16_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12088_LC_16_3_1 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_12088_LC_16_3_1  (
            .in0(N__92107),
            .in1(N__85845),
            .in2(N__58849),
            .in3(N__58840),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13892_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13892_bdd_4_lut_LC_16_3_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13892_bdd_4_lut_LC_16_3_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13892_bdd_4_lut_LC_16_3_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13892_bdd_4_lut_LC_16_3_2  (
            .in0(N__85843),
            .in1(N__58831),
            .in2(N__58825),
            .in3(N__86758),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5609_5610_LC_16_3_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5609_5610_LC_16_3_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5609_5610_LC_16_3_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5609_5610_LC_16_3_3  (
            .in0(N__58806),
            .in1(N__96528),
            .in2(_gnd_net_),
            .in3(N__79996),
            .lcout(REG_mem_58_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93432),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5705_5706_LC_16_3_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5705_5706_LC_16_3_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5705_5706_LC_16_3_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5705_5706_LC_16_3_4  (
            .in0(N__95707),
            .in1(N__96576),
            .in2(N__58798),
            .in3(N__79660),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93432),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2633_2634_LC_16_3_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2633_2634_LC_16_3_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2633_2634_LC_16_3_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2633_2634_LC_16_3_5  (
            .in0(N__96575),
            .in1(N__95708),
            .in2(N__58903),
            .in3(N__79659),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93432),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12163_LC_16_3_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12163_LC_16_3_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12163_LC_16_3_6 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12163_LC_16_3_6  (
            .in0(N__58786),
            .in1(N__92106),
            .in2(N__58768),
            .in3(N__88326),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14018 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13988_bdd_4_lut_LC_16_3_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13988_bdd_4_lut_LC_16_3_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13988_bdd_4_lut_LC_16_3_7 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13988_bdd_4_lut_LC_16_3_7  (
            .in0(N__58888),
            .in1(N__85844),
            .in2(N__88969),
            .in3(N__58732),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10008_3_lut_LC_16_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10008_3_lut_LC_16_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10008_3_lut_LC_16_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10008_3_lut_LC_16_4_0  (
            .in0(N__88756),
            .in1(N__89551),
            .in2(_gnd_net_),
            .in3(N__59017),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11657 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2060_2061_LC_16_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2060_2061_LC_16_4_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2060_2061_LC_16_4_1 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2060_2061_LC_16_4_1  (
            .in0(N__75897),
            .in1(N__95092),
            .in2(N__58975),
            .in3(N__77039),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93425),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11370_LC_16_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11370_LC_16_4_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11370_LC_16_4_2 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11370_LC_16_4_2  (
            .in0(N__88758),
            .in1(N__58996),
            .in2(N__92398),
            .in3(N__58945),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13064_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13064_bdd_4_lut_LC_16_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13064_bdd_4_lut_LC_16_4_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13064_bdd_4_lut_LC_16_4_3 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13064_bdd_4_lut_LC_16_4_3  (
            .in0(N__59058),
            .in1(N__58974),
            .in2(N__58960),
            .in3(N__92097),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13067 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11580_LC_16_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11580_LC_16_4_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11580_LC_16_4_4 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11580_LC_16_4_4  (
            .in0(N__88759),
            .in1(N__61756),
            .in2(N__92399),
            .in3(N__61735),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2252_2253_LC_16_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2252_2253_LC_16_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2252_2253_LC_16_4_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2252_2253_LC_16_4_5  (
            .in0(N__58944),
            .in1(N__75819),
            .in2(_gnd_net_),
            .in3(N__75048),
            .lcout(REG_mem_23_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93425),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3017_3018_LC_16_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3017_3018_LC_16_4_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3017_3018_LC_16_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3017_3018_LC_16_4_6  (
            .in0(N__96665),
            .in1(N__58932),
            .in2(_gnd_net_),
            .in3(N__72568),
            .lcout(REG_mem_31_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93425),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10035_3_lut_LC_16_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10035_3_lut_LC_16_4_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10035_3_lut_LC_16_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10035_3_lut_LC_16_4_7  (
            .in0(N__58921),
            .in1(N__58902),
            .in2(_gnd_net_),
            .in3(N__88757),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11684 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1877_1878_LC_16_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1877_1878_LC_16_5_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1877_1878_LC_16_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1877_1878_LC_16_5_0  (
            .in0(N__58872),
            .in1(N__62676),
            .in2(_gnd_net_),
            .in3(N__72110),
            .lcout(REG_mem_19_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12073_LC_16_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12073_LC_16_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12073_LC_16_5_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12073_LC_16_5_1  (
            .in0(N__59070),
            .in1(N__92494),
            .in2(N__59110),
            .in3(N__88545),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13910_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13910_bdd_4_lut_LC_16_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13910_bdd_4_lut_LC_16_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13910_bdd_4_lut_LC_16_5_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13910_bdd_4_lut_LC_16_5_2  (
            .in0(N__59082),
            .in1(N__92493),
            .in2(N__59086),
            .in3(N__66046),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13913 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1208_1209_LC_16_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1208_1209_LC_16_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1208_1209_LC_16_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1208_1209_LC_16_5_3  (
            .in0(N__74841),
            .in1(N__96189),
            .in2(_gnd_net_),
            .in3(N__59662),
            .lcout(REG_mem_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5036_5037_LC_16_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5036_5037_LC_16_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5036_5037_LC_16_5_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5036_5037_LC_16_5_4  (
            .in0(N__75904),
            .in1(N__95494),
            .in2(N__59083),
            .in3(N__77475),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5228_5229_LC_16_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5228_5229_LC_16_5_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5228_5229_LC_16_5_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5228_5229_LC_16_5_5  (
            .in0(N__95492),
            .in1(N__75905),
            .in2(N__59071),
            .in3(N__76354),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1964_1965_LC_16_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1964_1965_LC_16_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1964_1965_LC_16_5_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1964_1965_LC_16_5_6  (
            .in0(N__75903),
            .in1(N__95493),
            .in2(N__59059),
            .in3(N__77474),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93420),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10727_3_lut_LC_16_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10727_3_lut_LC_16_5_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10727_3_lut_LC_16_5_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10727_3_lut_LC_16_5_7  (
            .in0(N__85854),
            .in1(N__59044),
            .in2(_gnd_net_),
            .in3(N__59038),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2546_2547_LC_16_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2546_2547_LC_16_6_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2546_2547_LC_16_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2546_2547_LC_16_6_0  (
            .in0(N__76600),
            .in1(N__59025),
            .in2(_gnd_net_),
            .in3(N__70392),
            .lcout(REG_mem_26_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12038_LC_16_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12038_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12038_LC_16_6_1 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12038_LC_16_6_1  (
            .in0(N__59346),
            .in1(N__91699),
            .in2(N__59029),
            .in3(N__88540),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13868_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13868_bdd_4_lut_LC_16_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13868_bdd_4_lut_LC_16_6_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13868_bdd_4_lut_LC_16_6_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13868_bdd_4_lut_LC_16_6_2  (
            .in0(N__59358),
            .in1(N__92491),
            .in2(N__59374),
            .in3(N__59370),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13871 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2450_2451_LC_16_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2450_2451_LC_16_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2450_2451_LC_16_6_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2450_2451_LC_16_6_3  (
            .in0(N__95087),
            .in1(N__76602),
            .in2(N__59371),
            .in3(N__97021),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2354_2355_LC_16_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2354_2355_LC_16_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2354_2355_LC_16_6_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2354_2355_LC_16_6_4  (
            .in0(N__76601),
            .in1(N__95090),
            .in2(N__59359),
            .in3(N__96012),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2642_2643_LC_16_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2642_2643_LC_16_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2642_2643_LC_16_6_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2642_2643_LC_16_6_5  (
            .in0(N__95088),
            .in1(N__76603),
            .in2(N__59347),
            .in3(N__79759),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3206_3207_LC_16_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3206_3207_LC_16_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3206_3207_LC_16_6_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3206_3207_LC_16_6_6  (
            .in0(N__71569),
            .in1(N__95091),
            .in2(N__59328),
            .in3(N__80289),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5522_5523_LC_16_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5522_5523_LC_16_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5522_5523_LC_16_6_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5522_5523_LC_16_6_7  (
            .in0(N__95089),
            .in1(N__76604),
            .in2(N__61428),
            .in3(N__97022),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93412),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11465_LC_16_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11465_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11465_LC_16_7_0 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11465_LC_16_7_0  (
            .in0(N__88701),
            .in1(N__59146),
            .in2(N__92113),
            .in3(N__59311),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3698_3699_LC_16_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3698_3699_LC_16_7_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3698_3699_LC_16_7_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3698_3699_LC_16_7_1  (
            .in0(N__76605),
            .in1(N__59142),
            .in2(_gnd_net_),
            .in3(N__59284),
            .lcout(REG_mem_38_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93402),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3806_3807_LC_16_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3806_3807_LC_16_7_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3806_3807_LC_16_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3806_3807_LC_16_7_2  (
            .in0(N__61889),
            .in1(N__63765),
            .in2(_gnd_net_),
            .in3(N__89456),
            .lcout(REG_mem_39_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93402),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3797_3798_LC_16_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3797_3798_LC_16_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3797_3798_LC_16_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3797_3798_LC_16_7_3  (
            .in0(N__59121),
            .in1(N__62678),
            .in2(_gnd_net_),
            .in3(N__61890),
            .lcout(REG_mem_39_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93402),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1202_1203_LC_16_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1202_1203_LC_16_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1202_1203_LC_16_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1202_1203_LC_16_7_4  (
            .in0(N__59514),
            .in1(N__76606),
            .in2(_gnd_net_),
            .in3(N__59652),
            .lcout(REG_mem_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93402),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9989_3_lut_LC_16_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9989_3_lut_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9989_3_lut_LC_16_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9989_3_lut_LC_16_7_5  (
            .in0(N__63583),
            .in1(N__59515),
            .in2(_gnd_net_),
            .in3(N__88700),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1118_1119_LC_16_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1118_1119_LC_16_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1118_1119_LC_16_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1118_1119_LC_16_7_6  (
            .in0(N__59406),
            .in1(N__89455),
            .in2(_gnd_net_),
            .in3(N__66825),
            .lcout(REG_mem_11_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93402),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10208_3_lut_LC_16_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10208_3_lut_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10208_3_lut_LC_16_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10208_3_lut_LC_16_7_7  (
            .in0(N__59491),
            .in1(N__88699),
            .in2(_gnd_net_),
            .in3(N__63793),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11857 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4763_4764_LC_16_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4763_4764_LC_16_8_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4763_4764_LC_16_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4763_4764_LC_16_8_0  (
            .in0(N__62988),
            .in1(N__59448),
            .in2(_gnd_net_),
            .in3(N__63276),
            .lcout(REG_mem_49_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93390),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11954_LC_16_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11954_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11954_LC_16_8_1 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11954_LC_16_8_1  (
            .in0(N__59746),
            .in1(N__91417),
            .in2(N__59467),
            .in3(N__88254),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13760_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13760_bdd_4_lut_LC_16_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13760_bdd_4_lut_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13760_bdd_4_lut_LC_16_8_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13760_bdd_4_lut_LC_16_8_2  (
            .in0(N__91416),
            .in1(N__59449),
            .in2(N__59440),
            .in3(N__59419),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4667_4668_LC_16_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4667_4668_LC_16_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4667_4668_LC_16_8_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4667_4668_LC_16_8_3  (
            .in0(N__59418),
            .in1(_gnd_net_),
            .in2(N__63378),
            .in3(N__75580),
            .lcout(REG_mem_48_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93390),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12363_LC_16_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12363_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12363_LC_16_8_4 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12363_LC_16_8_4  (
            .in0(N__91418),
            .in1(N__59410),
            .in2(N__88538),
            .in3(N__59395),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4955_4956_LC_16_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4955_4956_LC_16_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4955_4956_LC_16_8_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4955_4956_LC_16_8_5  (
            .in0(N__59745),
            .in1(_gnd_net_),
            .in2(N__63379),
            .in3(N__72229),
            .lcout(REG_mem_51_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93390),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5426_5427_LC_16_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5426_5427_LC_16_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5426_5427_LC_16_8_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5426_5427_LC_16_8_6  (
            .in0(N__76610),
            .in1(N__95750),
            .in2(N__61449),
            .in3(N__95930),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93390),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1502_1503_LC_16_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1502_1503_LC_16_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1502_1503_LC_16_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1502_1503_LC_16_8_7  (
            .in0(N__59727),
            .in1(N__89457),
            .in2(_gnd_net_),
            .in3(N__64012),
            .lcout(REG_mem_15_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93390),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1301_1302_LC_16_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1301_1302_LC_16_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1301_1302_LC_16_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1301_1302_LC_16_9_0  (
            .in0(N__62861),
            .in1(N__59712),
            .in2(_gnd_net_),
            .in3(N__70122),
            .lcout(REG_mem_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11769_LC_16_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11769_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11769_LC_16_9_1 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11769_LC_16_9_1  (
            .in0(N__59671),
            .in1(N__91884),
            .in2(N__72898),
            .in3(N__88536),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13532_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13532_bdd_4_lut_LC_16_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13532_bdd_4_lut_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13532_bdd_4_lut_LC_16_9_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13532_bdd_4_lut_LC_16_9_2  (
            .in0(N__91883),
            .in1(N__59701),
            .in2(N__59683),
            .in3(N__59680),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11841 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4670_4671_LC_16_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4670_4671_LC_16_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4670_4671_LC_16_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4670_4671_LC_16_9_3  (
            .in0(N__59679),
            .in1(N__89452),
            .in2(_gnd_net_),
            .in3(N__75589),
            .lcout(REG_mem_48_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4382_4383_LC_16_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4382_4383_LC_16_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4382_4383_LC_16_9_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4382_4383_LC_16_9_4  (
            .in0(N__89451),
            .in1(_gnd_net_),
            .in2(N__89694),
            .in3(N__71864),
            .lcout(REG_mem_45_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4958_4959_LC_16_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4958_4959_LC_16_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4958_4959_LC_16_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4958_4959_LC_16_9_5  (
            .in0(N__59670),
            .in1(N__89453),
            .in2(_gnd_net_),
            .in3(N__72264),
            .lcout(REG_mem_51_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2153_2154_LC_16_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2153_2154_LC_16_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2153_2154_LC_16_9_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2153_2154_LC_16_9_6  (
            .in0(N__96769),
            .in1(N__95101),
            .in2(N__66126),
            .in3(N__76337),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93378),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11914_LC_16_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11914_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11914_LC_16_9_7 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11914_LC_16_9_7  (
            .in0(N__59845),
            .in1(N__91885),
            .in2(N__59809),
            .in3(N__88537),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5243_5244_LC_16_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5243_5244_LC_16_10_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5243_5244_LC_16_10_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5243_5244_LC_16_10_0  (
            .in0(N__63353),
            .in1(N__95100),
            .in2(N__59805),
            .in3(N__76236),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93349),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11929_LC_16_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11929_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11929_LC_16_10_1 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11929_LC_16_10_1  (
            .in0(N__91295),
            .in1(N__88253),
            .in2(N__59761),
            .in3(N__70414),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13736_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13736_bdd_4_lut_LC_16_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13736_bdd_4_lut_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13736_bdd_4_lut_LC_16_10_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13736_bdd_4_lut_LC_16_10_2  (
            .in0(N__59772),
            .in1(N__91293),
            .in2(N__59788),
            .in3(N__59784),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13739 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2834_2835_LC_16_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2834_2835_LC_16_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2834_2835_LC_16_10_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2834_2835_LC_16_10_3  (
            .in0(N__95097),
            .in1(N__76721),
            .in2(N__59785),
            .in3(N__70965),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93349),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2738_2739_LC_16_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2738_2739_LC_16_10_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2738_2739_LC_16_10_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2738_2739_LC_16_10_4  (
            .in0(N__76720),
            .in1(N__95099),
            .in2(N__59773),
            .in3(N__70721),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93349),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2930_2931_LC_16_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2930_2931_LC_16_10_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2930_2931_LC_16_10_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2930_2931_LC_16_10_5  (
            .in0(N__95098),
            .in1(N__76722),
            .in2(N__59760),
            .in3(N__77930),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93349),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6098_6099_LC_16_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6098_6099_LC_16_10_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6098_6099_LC_16_10_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6098_6099_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__63060),
            .in2(N__76752),
            .in3(N__67673),
            .lcout(REG_mem_63_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93349),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14138_bdd_4_lut_LC_16_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14138_bdd_4_lut_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14138_bdd_4_lut_LC_16_10_7 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14138_bdd_4_lut_LC_16_10_7  (
            .in0(N__91294),
            .in1(N__63049),
            .in2(N__59932),
            .in3(N__59914),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12093 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.state_timeout_counter_i0_i0_LC_16_11_0 .C_ON=1'b1;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i0_LC_16_11_0 .SEQ_MODE=4'b1001;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i0_LC_16_11_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \bluejay_data_inst.state_timeout_counter_i0_i0_LC_16_11_0  (
            .in0(N__78032),
            .in1(N__64473),
            .in2(_gnd_net_),
            .in3(N__59896),
            .lcout(\bluejay_data_inst.state_timeout_counter_0 ),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\bluejay_data_inst.n10581 ),
            .clk(N__97351),
            .ce(N__69171),
            .sr(N__69073));
    defparam \bluejay_data_inst.state_timeout_counter_i0_i1_LC_16_11_1 .C_ON=1'b1;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i1_LC_16_11_1 .SEQ_MODE=4'b1001;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i1_LC_16_11_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \bluejay_data_inst.state_timeout_counter_i0_i1_LC_16_11_1  (
            .in0(N__78034),
            .in1(N__59886),
            .in2(N__86586),
            .in3(N__59875),
            .lcout(\bluejay_data_inst.state_timeout_counter_1 ),
            .ltout(),
            .carryin(\bluejay_data_inst.n10581 ),
            .carryout(\bluejay_data_inst.n10582 ),
            .clk(N__97351),
            .ce(N__69171),
            .sr(N__69073));
    defparam \bluejay_data_inst.sub_116_add_2_4_lut_LC_16_11_2 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_4_lut_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_4_lut_LC_16_11_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_4_lut_LC_16_11_2  (
            .in0(N__78033),
            .in1(N__59872),
            .in2(N__86587),
            .in3(N__59848),
            .lcout(\bluejay_data_inst.n86 ),
            .ltout(),
            .carryin(\bluejay_data_inst.n10582 ),
            .carryout(\bluejay_data_inst.n10583 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_0_LC_16_11_3 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_0_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_0_LC_16_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_0_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__86530),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10583 ),
            .carryout(\bluejay_data_inst.n10583_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_1_LC_16_11_4 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_1_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_1_LC_16_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_1_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__86528),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10583_THRU_CRY_0_THRU_CO ),
            .carryout(\bluejay_data_inst.n10583_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_2_LC_16_11_5 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_2_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_2_LC_16_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_2_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(N__86531),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10583_THRU_CRY_1_THRU_CO ),
            .carryout(\bluejay_data_inst.n10583_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_3_LC_16_11_6 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_3_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_3_LC_16_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_3_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__86529),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10583_THRU_CRY_2_THRU_CO ),
            .carryout(\bluejay_data_inst.n10583_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_4_LC_16_11_7 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_4_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_4_LC_16_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_4_THRU_CRY_4_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__86532),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10583_THRU_CRY_3_THRU_CO ),
            .carryout(\bluejay_data_inst.n10583_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.state_timeout_counter_i0_i3_LC_16_12_0 .C_ON=1'b1;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i3_LC_16_12_0 .SEQ_MODE=4'b1001;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i3_LC_16_12_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \bluejay_data_inst.state_timeout_counter_i0_i3_LC_16_12_0  (
            .in0(N__78047),
            .in1(N__64415),
            .in2(N__86427),
            .in3(N__59938),
            .lcout(state_timeout_counter_3),
            .ltout(),
            .carryin(bfn_16_12_0_),
            .carryout(\bluejay_data_inst.n10584 ),
            .clk(N__97360),
            .ce(N__69175),
            .sr(N__64663));
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_0_LC_16_12_1 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_0_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_0_LC_16_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_0_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__86305),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10584 ),
            .carryout(\bluejay_data_inst.n10584_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_1_LC_16_12_2 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_1_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_1_LC_16_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_1_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__86428),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10584_THRU_CRY_0_THRU_CO ),
            .carryout(\bluejay_data_inst.n10584_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_2_LC_16_12_3 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_2_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_2_LC_16_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_2_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(N__86309),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10584_THRU_CRY_1_THRU_CO ),
            .carryout(\bluejay_data_inst.n10584_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_3_LC_16_12_4 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_3_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_3_LC_16_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_3_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__86429),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10584_THRU_CRY_2_THRU_CO ),
            .carryout(\bluejay_data_inst.n10584_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_4_LC_16_12_5 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_4_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_4_LC_16_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_4_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__86313),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10584_THRU_CRY_3_THRU_CO ),
            .carryout(\bluejay_data_inst.n10584_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_5_LC_16_12_6 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_5_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_5_LC_16_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_5_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__86430),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10584_THRU_CRY_4_THRU_CO ),
            .carryout(\bluejay_data_inst.n10584_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_6_LC_16_12_7 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_6_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_6_LC_16_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_5_THRU_CRY_6_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(N__86317),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10584_THRU_CRY_5_THRU_CO ),
            .carryout(\bluejay_data_inst.n10584_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.state_timeout_counter_i0_i4_LC_16_13_0 .C_ON=1'b1;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i4_LC_16_13_0 .SEQ_MODE=4'b1001;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i4_LC_16_13_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \bluejay_data_inst.state_timeout_counter_i0_i4_LC_16_13_0  (
            .in0(N__78054),
            .in1(N__64456),
            .in2(N__86588),
            .in3(N__59935),
            .lcout(\bluejay_data_inst.state_timeout_counter_4 ),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(\bluejay_data_inst.n10585 ),
            .clk(N__97368),
            .ce(N__69169),
            .sr(N__59965));
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_0_LC_16_13_1 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_0_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_0_LC_16_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_0_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__86539),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10585 ),
            .carryout(\bluejay_data_inst.n10585_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_1_LC_16_13_2 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_1_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_1_LC_16_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_1_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__86543),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10585_THRU_CRY_0_THRU_CO ),
            .carryout(\bluejay_data_inst.n10585_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_2_LC_16_13_3 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_2_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_2_LC_16_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_2_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(N__86540),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10585_THRU_CRY_1_THRU_CO ),
            .carryout(\bluejay_data_inst.n10585_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_3_LC_16_13_4 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_3_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_3_LC_16_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_3_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(N__86544),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10585_THRU_CRY_2_THRU_CO ),
            .carryout(\bluejay_data_inst.n10585_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_4_LC_16_13_5 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_4_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_4_LC_16_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_4_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(N__86541),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10585_THRU_CRY_3_THRU_CO ),
            .carryout(\bluejay_data_inst.n10585_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_5_LC_16_13_6 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_5_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_5_LC_16_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_5_LC_16_13_6  (
            .in0(_gnd_net_),
            .in1(N__86545),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10585_THRU_CRY_4_THRU_CO ),
            .carryout(\bluejay_data_inst.n10585_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_6_LC_16_13_7 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_6_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_6_LC_16_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_6_THRU_CRY_6_LC_16_13_7  (
            .in0(_gnd_net_),
            .in1(N__86542),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10585_THRU_CRY_5_THRU_CO ),
            .carryout(\bluejay_data_inst.n10585_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.state_timeout_counter_i0_i5_LC_16_14_0 .C_ON=1'b1;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i5_LC_16_14_0 .SEQ_MODE=4'b1001;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i5_LC_16_14_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \bluejay_data_inst.state_timeout_counter_i0_i5_LC_16_14_0  (
            .in0(N__78055),
            .in1(N__59952),
            .in2(N__86589),
            .in3(N__59941),
            .lcout(\bluejay_data_inst.state_timeout_counter_5 ),
            .ltout(),
            .carryin(bfn_16_14_0_),
            .carryout(\bluejay_data_inst.n10586 ),
            .clk(N__97375),
            .ce(N__69152),
            .sr(N__64656));
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_0_LC_16_14_1 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_0_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_0_LC_16_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_0_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__86549),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10586 ),
            .carryout(\bluejay_data_inst.n10586_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_1_LC_16_14_2 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_1_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_1_LC_16_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_1_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(N__86553),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10586_THRU_CRY_0_THRU_CO ),
            .carryout(\bluejay_data_inst.n10586_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_2_LC_16_14_3 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_2_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_2_LC_16_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_2_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(N__86550),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10586_THRU_CRY_1_THRU_CO ),
            .carryout(\bluejay_data_inst.n10586_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_3_LC_16_14_4 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_3_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_3_LC_16_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_3_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(N__86554),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10586_THRU_CRY_2_THRU_CO ),
            .carryout(\bluejay_data_inst.n10586_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_4_LC_16_14_5 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_4_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_4_LC_16_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_4_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(N__86551),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10586_THRU_CRY_3_THRU_CO ),
            .carryout(\bluejay_data_inst.n10586_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_5_LC_16_14_6 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_5_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_5_LC_16_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_5_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__86555),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10586_THRU_CRY_4_THRU_CO ),
            .carryout(\bluejay_data_inst.n10586_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_6_LC_16_14_7 .C_ON=1'b1;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_6_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_6_LC_16_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \bluejay_data_inst.sub_116_add_2_7_THRU_CRY_6_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(N__86552),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\bluejay_data_inst.n10586_THRU_CRY_5_THRU_CO ),
            .carryout(\bluejay_data_inst.n10586_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.state_timeout_counter_i0_i6_LC_16_15_0 .C_ON=1'b1;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i6_LC_16_15_0 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i6_LC_16_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \bluejay_data_inst.state_timeout_counter_i0_i6_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__59997),
            .in2(N__86590),
            .in3(N__59986),
            .lcout(\bluejay_data_inst.state_timeout_counter_6 ),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\bluejay_data_inst.n10587 ),
            .clk(N__97382),
            .ce(N__69168),
            .sr(N__69187));
    defparam \bluejay_data_inst.state_timeout_counter_i0_i7_LC_16_15_1 .C_ON=1'b0;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i7_LC_16_15_1 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.state_timeout_counter_i0_i7_LC_16_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \bluejay_data_inst.state_timeout_counter_i0_i7_LC_16_15_1  (
            .in0(N__86559),
            .in1(N__59976),
            .in2(_gnd_net_),
            .in3(N__59983),
            .lcout(\bluejay_data_inst.state_timeout_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97382),
            .ce(N__69168),
            .sr(N__69187));
    defparam \pc_rx.r_Bit_Index_i0_LC_16_16_1 .C_ON=1'b0;
    defparam \pc_rx.r_Bit_Index_i0_LC_16_16_1 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Bit_Index_i0_LC_16_16_1 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \pc_rx.r_Bit_Index_i0_LC_16_16_1  (
            .in0(N__60069),
            .in1(N__60358),
            .in2(_gnd_net_),
            .in3(N__60415),
            .lcout(\pc_rx.r_Bit_Index_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97389),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_SM_Main_i2_LC_16_16_2 .C_ON=1'b0;
    defparam \pc_rx.r_SM_Main_i2_LC_16_16_2 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_SM_Main_i2_LC_16_16_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pc_rx.r_SM_Main_i2_LC_16_16_2  (
            .in0(N__60794),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60378),
            .lcout(\pc_rx.r_SM_Main_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97389),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_Rx_Data_50_LC_16_16_3 .C_ON=1'b0;
    defparam \pc_rx.r_Rx_Data_50_LC_16_16_3 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Rx_Data_50_LC_16_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pc_rx.r_Rx_Data_50_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60199),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97389),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i1_2_lut_3_lut_adj_38_LC_16_16_4 .C_ON=1'b0;
    defparam \pc_rx.i1_2_lut_3_lut_adj_38_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i1_2_lut_3_lut_adj_38_LC_16_16_4 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \pc_rx.i1_2_lut_3_lut_adj_38_LC_16_16_4  (
            .in0(N__60793),
            .in1(N__60068),
            .in2(_gnd_net_),
            .in3(N__60377),
            .lcout(n4002),
            .ltout(n4002_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_Rx_Byte_i3_LC_16_16_5 .C_ON=1'b0;
    defparam \pc_rx.r_Rx_Byte_i3_LC_16_16_5 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Rx_Byte_i3_LC_16_16_5 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \pc_rx.r_Rx_Byte_i3_LC_16_16_5  (
            .in0(N__60132),
            .in1(N__60697),
            .in2(N__60151),
            .in3(N__60148),
            .lcout(pc_data_rx_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97389),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i1_LC_16_16_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i1_LC_16_16_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i1_LC_16_16_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i1_LC_16_16_6  (
            .in0(N__80831),
            .in1(N__73303),
            .in2(N__60121),
            .in3(N__65424),
            .lcout(fifo_data_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97389),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_Bit_Index_i2_LC_16_17_0 .C_ON=1'b0;
    defparam \pc_rx.r_Bit_Index_i2_LC_16_17_0 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Bit_Index_i2_LC_16_17_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \pc_rx.r_Bit_Index_i2_LC_16_17_0  (
            .in0(N__60038),
            .in1(N__60071),
            .in2(_gnd_net_),
            .in3(N__60101),
            .lcout(\pc_rx.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97398),
            .ce(N__60414),
            .sr(N__60016));
    defparam \pc_rx.r_Bit_Index_i1_LC_16_17_1 .C_ON=1'b0;
    defparam \pc_rx.r_Bit_Index_i1_LC_16_17_1 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_Bit_Index_i1_LC_16_17_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pc_rx.r_Bit_Index_i1_LC_16_17_1  (
            .in0(N__60070),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60037),
            .lcout(\pc_rx.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97398),
            .ce(N__60414),
            .sr(N__60016));
    defparam \pc_rx.i1_2_lut_adj_39_LC_16_18_0 .C_ON=1'b0;
    defparam \pc_rx.i1_2_lut_adj_39_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i1_2_lut_adj_39_LC_16_18_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pc_rx.i1_2_lut_adj_39_LC_16_18_0  (
            .in0(N__60767),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60223),
            .lcout(),
            .ltout(\pc_rx.n55_adj_1144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_SM_Main_i1_LC_16_18_1 .C_ON=1'b0;
    defparam \pc_rx.r_SM_Main_i1_LC_16_18_1 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_SM_Main_i1_LC_16_18_1 .LUT_INIT=16'b0001101100001010;
    LogicCell40 \pc_rx.r_SM_Main_i1_LC_16_18_1  (
            .in0(N__60350),
            .in1(N__60722),
            .in2(N__60004),
            .in3(N__60451),
            .lcout(\pc_rx.r_SM_Main_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97406),
            .ce(),
            .sr(N__60295));
    defparam \pc_rx.i1_2_lut_adj_42_LC_16_18_2 .C_ON=1'b0;
    defparam \pc_rx.i1_2_lut_adj_42_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i1_2_lut_adj_42_LC_16_18_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \pc_rx.i1_2_lut_adj_42_LC_16_18_2  (
            .in0(N__60768),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60660),
            .lcout(\pc_rx.n145 ),
            .ltout(\pc_rx.n145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i11078_4_lut_LC_16_18_3 .C_ON=1'b0;
    defparam \pc_rx.i11078_4_lut_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i11078_4_lut_LC_16_18_3 .LUT_INIT=16'b0000000010111111;
    LogicCell40 \pc_rx.i11078_4_lut_LC_16_18_3  (
            .in0(N__60343),
            .in1(N__60721),
            .in2(N__60445),
            .in3(N__60296),
            .lcout(\pc_rx.n6490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i13_4_lut_4_lut_LC_16_18_4 .C_ON=1'b0;
    defparam \pc_rx.i13_4_lut_4_lut_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i13_4_lut_4_lut_LC_16_18_4 .LUT_INIT=16'b0100001100000011;
    LogicCell40 \pc_rx.i13_4_lut_4_lut_LC_16_18_4  (
            .in0(N__60297),
            .in1(N__60344),
            .in2(N__60781),
            .in3(N__60221),
            .lcout(\pc_rx.n4081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i2_4_lut_LC_16_18_5 .C_ON=1'b0;
    defparam \pc_rx.i2_4_lut_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i2_4_lut_LC_16_18_5 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \pc_rx.i2_4_lut_LC_16_18_5  (
            .in0(N__60224),
            .in1(N__60299),
            .in2(N__60357),
            .in3(N__60769),
            .lcout(\pc_rx.n4140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i1_2_lut_3_lut_adj_40_LC_16_18_6 .C_ON=1'b0;
    defparam \pc_rx.i1_2_lut_3_lut_adj_40_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i1_2_lut_3_lut_adj_40_LC_16_18_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \pc_rx.i1_2_lut_3_lut_adj_40_LC_16_18_6  (
            .in0(N__60298),
            .in1(N__60345),
            .in2(_gnd_net_),
            .in3(N__60222),
            .lcout(\pc_rx.n151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.r_SM_Main_i0_LC_16_18_7 .C_ON=1'b0;
    defparam \pc_rx.r_SM_Main_i0_LC_16_18_7 .SEQ_MODE=4'b1000;
    defparam \pc_rx.r_SM_Main_i0_LC_16_18_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pc_rx.r_SM_Main_i0_LC_16_18_7  (
            .in0(N__60349),
            .in1(N__60307),
            .in2(_gnd_net_),
            .in3(N__60457),
            .lcout(\pc_rx.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97406),
            .ce(),
            .sr(N__60295));
    defparam \pc_rx.i4_4_lut_LC_16_19_0 .C_ON=1'b0;
    defparam \pc_rx.i4_4_lut_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i4_4_lut_LC_16_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pc_rx.i4_4_lut_LC_16_19_0  (
            .in0(N__60556),
            .in1(N__60271),
            .in2(N__60259),
            .in3(N__60244),
            .lcout(\pc_rx.n140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i1_3_lut_adj_44_LC_16_19_1 .C_ON=1'b0;
    defparam \pc_rx.i1_3_lut_adj_44_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i1_3_lut_adj_44_LC_16_19_1 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \pc_rx.i1_3_lut_adj_44_LC_16_19_1  (
            .in0(N__60534),
            .in1(N__60516),
            .in2(_gnd_net_),
            .in3(N__60474),
            .lcout(),
            .ltout(\pc_rx.n4_adj_1145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i1_4_lut_LC_16_19_2 .C_ON=1'b0;
    defparam \pc_rx.i1_4_lut_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i1_4_lut_LC_16_19_2 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \pc_rx.i1_4_lut_LC_16_19_2  (
            .in0(N__60549),
            .in1(N__60501),
            .in2(N__60232),
            .in3(N__60486),
            .lcout(\pc_rx.r_SM_Main_2_N_732_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i1_2_lut_adj_43_LC_16_19_3 .C_ON=1'b0;
    defparam \pc_rx.i1_2_lut_adj_43_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i1_2_lut_adj_43_LC_16_19_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \pc_rx.i1_2_lut_adj_43_LC_16_19_3  (
            .in0(N__60580),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60568),
            .lcout(\pc_rx.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i3_4_lut_adj_41_LC_16_19_4 .C_ON=1'b0;
    defparam \pc_rx.i3_4_lut_adj_41_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i3_4_lut_adj_41_LC_16_19_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \pc_rx.i3_4_lut_adj_41_LC_16_19_4  (
            .in0(N__60550),
            .in1(N__60535),
            .in2(N__60520),
            .in3(N__60502),
            .lcout(),
            .ltout(\pc_rx.n8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i4_3_lut_LC_16_19_5 .C_ON=1'b0;
    defparam \pc_rx.i4_3_lut_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i4_3_lut_LC_16_19_5 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \pc_rx.i4_3_lut_LC_16_19_5  (
            .in0(N__60487),
            .in1(_gnd_net_),
            .in2(N__60478),
            .in3(N__60475),
            .lcout(\pc_rx.n13 ),
            .ltout(\pc_rx.n13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i5300_4_lut_3_lut_LC_16_19_6 .C_ON=1'b0;
    defparam \pc_rx.i5300_4_lut_3_lut_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i5300_4_lut_3_lut_LC_16_19_6 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \pc_rx.i5300_4_lut_3_lut_LC_16_19_6  (
            .in0(N__60723),
            .in1(_gnd_net_),
            .in2(N__60460),
            .in3(N__60770),
            .lcout(\pc_rx.n6500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_all_w_I_0_1_lut_LC_16_19_7.C_ON=1'b0;
    defparam reset_all_w_I_0_1_lut_LC_16_19_7.SEQ_MODE=4'b0000;
    defparam reset_all_w_I_0_1_lut_LC_16_19_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 reset_all_w_I_0_1_lut_LC_16_19_7 (
            .in0(N__78365),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESET_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_clk_counter_i3_1107__i1_LC_16_20_0.C_ON=1'b0;
    defparam reset_clk_counter_i3_1107__i1_LC_16_20_0.SEQ_MODE=4'b1000;
    defparam reset_clk_counter_i3_1107__i1_LC_16_20_0.LUT_INIT=16'b1001100111001100;
    LogicCell40 reset_clk_counter_i3_1107__i1_LC_16_20_0 (
            .in0(N__60818),
            .in1(N__60888),
            .in2(_gnd_net_),
            .in3(N__60834),
            .lcout(reset_clk_counter_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97426),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_clk_counter_i3_1107__i2_LC_16_20_1.C_ON=1'b0;
    defparam reset_clk_counter_i3_1107__i2_LC_16_20_1.SEQ_MODE=4'b1000;
    defparam reset_clk_counter_i3_1107__i2_LC_16_20_1.LUT_INIT=16'b1100110010011100;
    LogicCell40 reset_clk_counter_i3_1107__i2_LC_16_20_1 (
            .in0(N__60889),
            .in1(N__60857),
            .in2(N__60838),
            .in3(N__60819),
            .lcout(reset_clk_counter_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97426),
            .ce(),
            .sr(_gnd_net_));
    defparam i9054_2_lut_3_lut_LC_16_20_2.C_ON=1'b0;
    defparam i9054_2_lut_3_lut_LC_16_20_2.SEQ_MODE=4'b0000;
    defparam i9054_2_lut_3_lut_LC_16_20_2.LUT_INIT=16'b1110111011111111;
    LogicCell40 i9054_2_lut_3_lut_LC_16_20_2 (
            .in0(N__60813),
            .in1(N__60886),
            .in2(_gnd_net_),
            .in3(N__60833),
            .lcout(),
            .ltout(n10562_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_clk_counter_i3_1107__i3_LC_16_20_3.C_ON=1'b0;
    defparam reset_clk_counter_i3_1107__i3_LC_16_20_3.SEQ_MODE=4'b1000;
    defparam reset_clk_counter_i3_1107__i3_LC_16_20_3.LUT_INIT=16'b1100110011000011;
    LogicCell40 reset_clk_counter_i3_1107__i3_LC_16_20_3 (
            .in0(_gnd_net_),
            .in1(N__60871),
            .in2(N__60892),
            .in3(N__60858),
            .lcout(reset_clk_counter_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97426),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_all_r_77_LC_16_20_4.C_ON=1'b0;
    defparam reset_all_r_77_LC_16_20_4.SEQ_MODE=4'b1000;
    defparam reset_all_r_77_LC_16_20_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 reset_all_r_77_LC_16_20_4 (
            .in0(N__60870),
            .in1(N__60856),
            .in2(N__60820),
            .in3(N__60887),
            .lcout(reset_all_w),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97426),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_16_20_5.C_ON=1'b0;
    defparam i3_4_lut_LC_16_20_5.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_16_20_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i3_4_lut_LC_16_20_5 (
            .in0(N__60885),
            .in1(N__60869),
            .in2(N__60859),
            .in3(N__60812),
            .lcout(reset_all_w_N_61),
            .ltout(reset_all_w_N_61_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_clk_counter_i3_1107__i0_LC_16_20_6.C_ON=1'b0;
    defparam reset_clk_counter_i3_1107__i0_LC_16_20_6.SEQ_MODE=4'b1000;
    defparam reset_clk_counter_i3_1107__i0_LC_16_20_6.LUT_INIT=16'b0101101001011010;
    LogicCell40 reset_clk_counter_i3_1107__i0_LC_16_20_6 (
            .in0(N__60817),
            .in1(_gnd_net_),
            .in2(N__60823),
            .in3(_gnd_net_),
            .lcout(reset_clk_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97426),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_rx.i1_3_lut_LC_16_20_7 .C_ON=1'b0;
    defparam \pc_rx.i1_3_lut_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \pc_rx.i1_3_lut_LC_16_20_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \pc_rx.i1_3_lut_LC_16_20_7  (
            .in0(N__60787),
            .in1(N__60724),
            .in2(_gnd_net_),
            .in3(N__60661),
            .lcout(\pc_rx.n125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.usb3_data_in_latched__i5_LC_17_1_2 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i5_LC_17_1_2 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i5_LC_17_1_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i5_LC_17_1_2  (
            .in0(N__60637),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\usb3_if_inst.usb3_data_in_latched_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93451),
            .ce(),
            .sr(N__73712));
    defparam \usb3_if_inst.usb3_data_in_latched__i6_LC_17_1_3 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i6_LC_17_1_3 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i6_LC_17_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i6_LC_17_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60625),
            .lcout(\usb3_if_inst.usb3_data_in_latched_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93451),
            .ce(),
            .sr(N__73712));
    defparam \usb3_if_inst.usb3_data_in_latched__i7_LC_17_1_5 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i7_LC_17_1_5 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i7_LC_17_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i7_LC_17_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60613),
            .lcout(\usb3_if_inst.usb3_data_in_latched_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93451),
            .ce(),
            .sr(N__73712));
    defparam \usb3_if_inst.usb3_data_in_latched__i4_LC_17_1_6 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i4_LC_17_1_6 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i4_LC_17_1_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i4_LC_17_1_6  (
            .in0(N__60595),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\usb3_if_inst.usb3_data_in_latched_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93451),
            .ce(),
            .sr(N__73712));
    defparam \usb3_if_inst.dc32_fifo_data_in_i2_LC_17_2_1 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i2_LC_17_2_1 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i2_LC_17_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i2_LC_17_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65716),
            .lcout(dc32_fifo_data_in_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.dc32_fifo_data_in_i2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.dc32_fifo_data_in_i3_LC_17_2_2 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i3_LC_17_2_2 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i3_LC_17_2_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i3_LC_17_2_2  (
            .in0(N__65737),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(dc32_fifo_data_in_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.dc32_fifo_data_in_i2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.dc32_fifo_data_in_i4_LC_17_2_3 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i4_LC_17_2_3 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i4_LC_17_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i4_LC_17_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61411),
            .lcout(dc32_fifo_data_in_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.dc32_fifo_data_in_i2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.dc32_fifo_data_in_i5_LC_17_2_4 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i5_LC_17_2_4 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i5_LC_17_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i5_LC_17_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60967),
            .lcout(dc32_fifo_data_in_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.dc32_fifo_data_in_i2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.dc32_fifo_data_in_i6_LC_17_2_5 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i6_LC_17_2_5 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i6_LC_17_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i6_LC_17_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60961),
            .lcout(dc32_fifo_data_in_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.dc32_fifo_data_in_i2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.dc32_fifo_data_in_i7_LC_17_2_6 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i7_LC_17_2_6 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i7_LC_17_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i7_LC_17_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60955),
            .lcout(dc32_fifo_data_in_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.dc32_fifo_data_in_i2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.dc32_fifo_data_in_i8_LC_17_2_7 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i8_LC_17_2_7 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i8_LC_17_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i8_LC_17_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60949),
            .lcout(dc32_fifo_data_in_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.dc32_fifo_data_in_i2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12944_bdd_4_lut_LC_17_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12944_bdd_4_lut_LC_17_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12944_bdd_4_lut_LC_17_4_0 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12944_bdd_4_lut_LC_17_4_0  (
            .in0(N__90389),
            .in1(N__60898),
            .in2(N__60943),
            .in3(N__61483),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12947 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11286_LC_17_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11286_LC_17_4_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11286_LC_17_4_1 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11286_LC_17_4_1  (
            .in0(N__60925),
            .in1(N__90391),
            .in2(N__60913),
            .in3(N__85856),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12944 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_LC_17_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_LC_17_4_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_LC_17_4_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_LC_17_4_2  (
            .in0(N__85857),
            .in1(N__61594),
            .in2(N__90399),
            .in3(N__75235),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14408_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14408_bdd_4_lut_LC_17_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14408_bdd_4_lut_LC_17_4_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14408_bdd_4_lut_LC_17_4_3 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14408_bdd_4_lut_LC_17_4_3  (
            .in0(N__61579),
            .in1(N__90390),
            .in2(N__61570),
            .in3(N__61567),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9849_3_lut_LC_17_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9849_3_lut_LC_17_4_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9849_3_lut_LC_17_4_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i9849_3_lut_LC_17_4_4  (
            .in0(_gnd_net_),
            .in1(N__81495),
            .in2(N__61561),
            .in3(N__61558),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11498_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i3_LC_17_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i3_LC_17_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i3_LC_17_4_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i3_LC_17_4_5  (
            .in0(N__61951),
            .in1(_gnd_net_),
            .in2(N__61552),
            .in3(N__81093),
            .lcout(REG_out_raw_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97418),
            .ce(N__80881),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14210_bdd_4_lut_LC_17_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14210_bdd_4_lut_LC_17_4_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14210_bdd_4_lut_LC_17_4_6 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14210_bdd_4_lut_LC_17_4_6  (
            .in0(N__61525),
            .in1(N__92191),
            .in2(N__61924),
            .in3(N__61501),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12057 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5714_5715_LC_17_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5714_5715_LC_17_5_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5714_5715_LC_17_5_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5714_5715_LC_17_5_0  (
            .in0(N__79771),
            .in1(N__61461),
            .in2(N__95625),
            .in3(N__76621),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93426),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5618_5619_LC_17_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5618_5619_LC_17_5_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5618_5619_LC_17_5_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5618_5619_LC_17_5_1  (
            .in0(N__61473),
            .in1(N__76513),
            .in2(_gnd_net_),
            .in3(N__79995),
            .lcout(REG_mem_58_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93426),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12313_LC_17_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12313_LC_17_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12313_LC_17_5_2 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12313_LC_17_5_2  (
            .in0(N__88760),
            .in1(N__92105),
            .in2(N__61477),
            .in3(N__61462),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14198_bdd_4_lut_LC_17_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14198_bdd_4_lut_LC_17_5_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14198_bdd_4_lut_LC_17_5_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14198_bdd_4_lut_LC_17_5_3  (
            .in0(N__92104),
            .in1(N__61453),
            .in2(N__61432),
            .in3(N__61429),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12066 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4076_4077_LC_17_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4076_4077_LC_17_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4076_4077_LC_17_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4076_4077_LC_17_5_4  (
            .in0(N__61695),
            .in1(N__75805),
            .in2(_gnd_net_),
            .in3(N__68088),
            .lcout(REG_mem_42_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93426),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2636_2637_LC_17_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2636_2637_LC_17_5_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2636_2637_LC_17_5_5 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2636_2637_LC_17_5_5  (
            .in0(N__75804),
            .in1(N__61617),
            .in2(N__79798),
            .in3(N__95326),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93426),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2648_2649_LC_17_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2648_2649_LC_17_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2648_2649_LC_17_5_6 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2648_2649_LC_17_5_6  (
            .in0(N__79770),
            .in1(N__69822),
            .in2(N__95624),
            .in3(N__96231),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93426),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5720_5721_LC_17_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5720_5721_LC_17_5_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5720_5721_LC_17_5_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5720_5721_LC_17_5_7  (
            .in0(N__96230),
            .in1(N__95325),
            .in2(N__71142),
            .in3(N__79792),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93426),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14360_bdd_4_lut_LC_17_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14360_bdd_4_lut_LC_17_6_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14360_bdd_4_lut_LC_17_6_0 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14360_bdd_4_lut_LC_17_6_0  (
            .in0(N__61684),
            .in1(N__91834),
            .in2(N__61630),
            .in3(N__61669),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12453_LC_17_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12453_LC_17_6_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12453_LC_17_6_1 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12453_LC_17_6_1  (
            .in0(N__91836),
            .in1(N__61654),
            .in2(N__88748),
            .in3(N__63042),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11191_LC_17_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11191_LC_17_6_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11191_LC_17_6_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11191_LC_17_6_2  (
            .in0(N__61717),
            .in1(N__91835),
            .in2(N__61621),
            .in3(N__88541),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12848_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12848_bdd_4_lut_LC_17_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12848_bdd_4_lut_LC_17_6_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12848_bdd_4_lut_LC_17_6_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12848_bdd_4_lut_LC_17_6_3  (
            .in0(N__91833),
            .in1(N__71113),
            .in2(N__61606),
            .in3(N__75610),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12851_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10728_3_lut_LC_17_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10728_3_lut_LC_17_6_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10728_3_lut_LC_17_6_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10728_3_lut_LC_17_6_4  (
            .in0(N__85855),
            .in1(_gnd_net_),
            .in2(N__61603),
            .in3(N__61600),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12377_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11455_LC_17_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11455_LC_17_6_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11455_LC_17_6_5 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_3__bdd_4_lut_11455_LC_17_6_5  (
            .in0(N__81474),
            .in1(N__90369),
            .in2(N__61978),
            .in3(N__61975),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13010_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13010_bdd_4_lut_LC_17_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13010_bdd_4_lut_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13010_bdd_4_lut_LC_17_6_6 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13010_bdd_4_lut_LC_17_6_6  (
            .in0(N__61969),
            .in1(N__81473),
            .in2(N__61954),
            .in3(N__67003),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13013 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12323_LC_17_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12323_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12323_LC_17_7_0 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12323_LC_17_7_0  (
            .in0(N__61942),
            .in1(N__91743),
            .in2(N__88834),
            .in3(N__61765),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3986_3987_LC_17_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3986_3987_LC_17_7_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3986_3987_LC_17_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3986_3987_LC_17_7_1  (
            .in0(N__61905),
            .in1(N__76611),
            .in2(_gnd_net_),
            .in3(N__66026),
            .lcout(REG_mem_41_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93413),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3788_3789_LC_17_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3788_3789_LC_17_7_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3788_3789_LC_17_7_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3788_3789_LC_17_7_2  (
            .in0(N__75924),
            .in1(N__61764),
            .in2(_gnd_net_),
            .in3(N__61892),
            .lcout(REG_mem_39_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93413),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1484_1485_LC_17_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1484_1485_LC_17_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1484_1485_LC_17_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1484_1485_LC_17_7_3  (
            .in0(N__72300),
            .in1(N__75925),
            .in2(_gnd_net_),
            .in3(N__64009),
            .lcout(REG_mem_15_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93413),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1772_1773_LC_17_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1772_1773_LC_17_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1772_1773_LC_17_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1772_1773_LC_17_7_4  (
            .in0(N__75922),
            .in1(N__61746),
            .in2(_gnd_net_),
            .in3(N__67513),
            .lcout(REG_mem_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93413),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1868_1869_LC_17_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1868_1869_LC_17_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1868_1869_LC_17_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1868_1869_LC_17_7_5  (
            .in0(N__61728),
            .in1(N__75926),
            .in2(_gnd_net_),
            .in3(N__72101),
            .lcout(REG_mem_19_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93413),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2540_2541_LC_17_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2540_2541_LC_17_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2540_2541_LC_17_7_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2540_2541_LC_17_7_6  (
            .in0(N__75923),
            .in1(N__61716),
            .in2(_gnd_net_),
            .in3(N__70386),
            .lcout(REG_mem_26_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93413),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3020_3021_LC_17_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3020_3021_LC_17_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3020_3021_LC_17_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3020_3021_LC_17_7_7  (
            .in0(N__63043),
            .in1(N__75927),
            .in2(_gnd_net_),
            .in3(N__72560),
            .lcout(REG_mem_31_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93413),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14348_bdd_4_lut_LC_17_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14348_bdd_4_lut_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14348_bdd_4_lut_LC_17_8_0 .LUT_INIT=16'b1111101000001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14348_bdd_4_lut_LC_17_8_0  (
            .in0(N__62872),
            .in1(N__63028),
            .in2(N__91813),
            .in3(N__66595),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12006 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i908_909_LC_17_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i908_909_LC_17_8_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i908_909_LC_17_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i908_909_LC_17_8_1  (
            .in0(N__66636),
            .in1(N__75820),
            .in2(_gnd_net_),
            .in3(N__67192),
            .lcout(REG_mem_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4754_4755_LC_17_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4754_4755_LC_17_8_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4754_4755_LC_17_8_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4754_4755_LC_17_8_2  (
            .in0(N__62871),
            .in1(N__62985),
            .in2(_gnd_net_),
            .in3(N__76619),
            .lcout(REG_mem_49_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2933_2934_LC_17_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2933_2934_LC_17_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2933_2934_LC_17_8_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2933_2934_LC_17_8_3  (
            .in0(N__94825),
            .in1(N__62679),
            .in2(N__62463),
            .in3(N__77957),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4850_4851_LC_17_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4850_4851_LC_17_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4850_4851_LC_17_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4850_4851_LC_17_8_4  (
            .in0(N__66615),
            .in1(N__76617),
            .in2(_gnd_net_),
            .in3(N__73050),
            .lcout(REG_mem_50_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2579_2580_LC_17_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2579_2580_LC_17_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2579_2580_LC_17_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2579_2580_LC_17_8_5  (
            .in0(N__62019),
            .in1(N__62419),
            .in2(_gnd_net_),
            .in3(N__70385),
            .lcout(REG_mem_26_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i626_627_LC_17_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i626_627_LC_17_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i626_627_LC_17_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i626_627_LC_17_8_6  (
            .in0(N__61986),
            .in1(N__76618),
            .in2(_gnd_net_),
            .in3(N__66422),
            .lcout(REG_mem_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93403),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10872_3_lut_LC_17_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10872_3_lut_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10872_3_lut_LC_17_8_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10872_3_lut_LC_17_8_7  (
            .in0(N__88264),
            .in1(N__62008),
            .in2(_gnd_net_),
            .in3(N__61987),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12521 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1292_1293_LC_17_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1292_1293_LC_17_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1292_1293_LC_17_9_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1292_1293_LC_17_9_0  (
            .in0(N__63786),
            .in1(N__75821),
            .in2(_gnd_net_),
            .in3(N__70121),
            .lcout(REG_mem_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11988_LC_17_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11988_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11988_LC_17_9_1 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11988_LC_17_9_1  (
            .in0(N__91739),
            .in1(N__63775),
            .in2(N__88539),
            .in3(N__63754),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3614_3615_LC_17_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3614_3615_LC_17_9_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3614_3615_LC_17_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3614_3615_LC_17_9_2  (
            .in0(N__67056),
            .in1(N__89435),
            .in2(_gnd_net_),
            .in3(N__63689),
            .lcout(REG_mem_37_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1298_1299_LC_17_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1298_1299_LC_17_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1298_1299_LC_17_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1298_1299_LC_17_9_3  (
            .in0(N__70120),
            .in1(N__76620),
            .in2(_gnd_net_),
            .in3(N__63579),
            .lcout(REG_mem_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i155_156_LC_17_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i155_156_LC_17_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i155_156_LC_17_9_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i155_156_LC_17_9_4  (
            .in0(N__63380),
            .in1(N__95173),
            .in2(N__63561),
            .in3(N__80268),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1787_1788_LC_17_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1787_1788_LC_17_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1787_1788_LC_17_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1787_1788_LC_17_9_5  (
            .in0(N__63075),
            .in1(N__63381),
            .in2(_gnd_net_),
            .in3(N__67505),
            .lcout(REG_mem_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i638_639_LC_17_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i638_639_LC_17_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i638_639_LC_17_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i638_639_LC_17_9_6  (
            .in0(N__83076),
            .in1(N__89436),
            .in2(_gnd_net_),
            .in3(N__66387),
            .lcout(REG_mem_6_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i734_735_LC_17_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i734_735_LC_17_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i734_735_LC_17_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i734_735_LC_17_9_7  (
            .in0(N__89434),
            .in1(N__83061),
            .in2(_gnd_net_),
            .in3(N__89670),
            .lcout(REG_mem_7_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93391),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12263_LC_17_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12263_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12263_LC_17_10_0 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12263_LC_17_10_0  (
            .in0(N__88263),
            .in1(N__75145),
            .in2(N__63064),
            .in3(N__91731),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10106_3_lut_LC_17_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10106_3_lut_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10106_3_lut_LC_17_10_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10106_3_lut_LC_17_10_1  (
            .in0(N__63855),
            .in1(N__88261),
            .in2(_gnd_net_),
            .in3(N__77269),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1496_1497_LC_17_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1496_1497_LC_17_10_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1496_1497_LC_17_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1496_1497_LC_17_10_2  (
            .in0(N__74802),
            .in1(N__96260),
            .in2(_gnd_net_),
            .in3(N__63998),
            .lcout(REG_mem_15_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93365),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3410_3411_LC_17_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3410_3411_LC_17_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3410_3411_LC_17_10_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3410_3411_LC_17_10_3  (
            .in0(N__94823),
            .in1(N__76736),
            .in2(N__63808),
            .in3(N__83378),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93365),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2066_2067_LC_17_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2066_2067_LC_17_10_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2066_2067_LC_17_10_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2066_2067_LC_17_10_4  (
            .in0(N__76733),
            .in1(N__94824),
            .in2(N__63859),
            .in3(N__77019),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93365),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2162_2163_LC_17_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2162_2163_LC_17_10_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2162_2163_LC_17_10_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2162_2163_LC_17_10_5  (
            .in0(N__94822),
            .in1(N__76735),
            .in2(N__63841),
            .in3(N__76237),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93365),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10107_3_lut_LC_17_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10107_3_lut_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10107_3_lut_LC_17_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10107_3_lut_LC_17_10_6  (
            .in0(N__88262),
            .in1(N__63840),
            .in2(_gnd_net_),
            .in3(N__63817),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11756 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2258_2259_LC_17_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2258_2259_LC_17_10_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2258_2259_LC_17_10_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2258_2259_LC_17_10_7  (
            .in0(N__63816),
            .in1(N__76734),
            .in2(_gnd_net_),
            .in3(N__75012),
            .lcout(REG_mem_23_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93365),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3218_3219_LC_17_11_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3218_3219_LC_17_11_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3218_3219_LC_17_11_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3218_3219_LC_17_11_0  (
            .in0(N__76613),
            .in1(N__93926),
            .in2(N__64243),
            .in3(N__80267),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93392),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11665_LC_17_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11665_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11665_LC_17_11_1 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11665_LC_17_11_1  (
            .in0(N__91927),
            .in1(N__63807),
            .in2(N__64204),
            .in3(N__88342),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13418_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13418_bdd_4_lut_LC_17_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13418_bdd_4_lut_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13418_bdd_4_lut_LC_17_11_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13418_bdd_4_lut_LC_17_11_2  (
            .in0(N__64242),
            .in1(N__91926),
            .in2(N__64231),
            .in3(N__64215),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13421 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3122_3123_LC_17_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3122_3123_LC_17_11_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3122_3123_LC_17_11_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3122_3123_LC_17_11_3  (
            .in0(N__93923),
            .in1(N__76615),
            .in2(N__64216),
            .in3(N__82934),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93392),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3314_3315_LC_17_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3314_3315_LC_17_11_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3314_3315_LC_17_11_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3314_3315_LC_17_11_4  (
            .in0(N__76614),
            .in1(N__93927),
            .in2(N__64203),
            .in3(N__80569),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93392),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i50_51_LC_17_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i50_51_LC_17_11_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i50_51_LC_17_11_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i50_51_LC_17_11_5  (
            .in0(N__93924),
            .in1(N__76616),
            .in2(N__64186),
            .in3(N__82935),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93392),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i146_147_LC_17_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i146_147_LC_17_11_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i146_147_LC_17_11_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i146_147_LC_17_11_6  (
            .in0(N__76612),
            .in1(N__93925),
            .in2(N__64174),
            .in3(N__80266),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93392),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10865_3_lut_LC_17_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10865_3_lut_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10865_3_lut_LC_17_11_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10865_3_lut_LC_17_11_7  (
            .in0(N__64185),
            .in1(N__88341),
            .in2(_gnd_net_),
            .in3(N__64173),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.state_FSM_i3_LC_17_12_0 .C_ON=1'b0;
    defparam \usb3_if_inst.state_FSM_i3_LC_17_12_0 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.state_FSM_i3_LC_17_12_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \usb3_if_inst.state_FSM_i3_LC_17_12_0  (
            .in0(N__64068),
            .in1(N__64162),
            .in2(N__64150),
            .in3(N__64363),
            .lcout(\usb3_if_inst.n553 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.state_FSM_i3C_net ),
            .ce(),
            .sr(N__73685));
    defparam \bluejay_data_inst.i1_2_lut_3_lut_4_lut_LC_17_13_0 .C_ON=1'b0;
    defparam \bluejay_data_inst.i1_2_lut_3_lut_4_lut_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i1_2_lut_3_lut_4_lut_LC_17_13_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \bluejay_data_inst.i1_2_lut_3_lut_4_lut_LC_17_13_0  (
            .in0(N__64416),
            .in1(N__64481),
            .in2(N__64462),
            .in3(N__64439),
            .lcout(\bluejay_data_inst.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.state_FSM_i4_LC_17_13_1 .C_ON=1'b0;
    defparam \bluejay_data_inst.state_FSM_i4_LC_17_13_1 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.state_FSM_i4_LC_17_13_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \bluejay_data_inst.state_FSM_i4_LC_17_13_1  (
            .in0(N__78096),
            .in1(N__64420),
            .in2(N__64368),
            .in3(N__64395),
            .lcout(\bluejay_data_inst.bluejay_data_out_31__N_701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97376),
            .ce(),
            .sr(N__73556));
    defparam \bluejay_data_inst.i1_2_lut_adj_65_LC_17_13_2 .C_ON=1'b0;
    defparam \bluejay_data_inst.i1_2_lut_adj_65_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i1_2_lut_adj_65_LC_17_13_2 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \bluejay_data_inst.i1_2_lut_adj_65_LC_17_13_2  (
            .in0(N__64461),
            .in1(N__64483),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\bluejay_data_inst.n8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.state_FSM_i3_LC_17_13_3 .C_ON=1'b0;
    defparam \bluejay_data_inst.state_FSM_i3_LC_17_13_3 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.state_FSM_i3_LC_17_13_3 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \bluejay_data_inst.state_FSM_i3_LC_17_13_3  (
            .in0(N__64440),
            .in1(N__64489),
            .in2(N__64492),
            .in3(N__64698),
            .lcout(\bluejay_data_inst.n717 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97376),
            .ce(),
            .sr(N__73556));
    defparam \bluejay_data_inst.i1_4_lut_adj_61_LC_17_13_4 .C_ON=1'b0;
    defparam \bluejay_data_inst.i1_4_lut_adj_61_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i1_4_lut_adj_61_LC_17_13_4 .LUT_INIT=16'b0101000001010100;
    LogicCell40 \bluejay_data_inst.i1_4_lut_adj_61_LC_17_13_4  (
            .in0(N__64417),
            .in1(N__78094),
            .in2(N__68785),
            .in3(N__64354),
            .lcout(\bluejay_data_inst.n12_adj_1179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i1_2_lut_3_lut_LC_17_13_5 .C_ON=1'b0;
    defparam \bluejay_data_inst.i1_2_lut_3_lut_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i1_2_lut_3_lut_LC_17_13_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \bluejay_data_inst.i1_2_lut_3_lut_LC_17_13_5  (
            .in0(N__64482),
            .in1(N__64460),
            .in2(_gnd_net_),
            .in3(N__64441),
            .lcout(n7),
            .ltout(n7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.state_FSM_i2_LC_17_13_6 .C_ON=1'b0;
    defparam \bluejay_data_inst.state_FSM_i2_LC_17_13_6 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.state_FSM_i2_LC_17_13_6 .LUT_INIT=16'b1111111111001000;
    LogicCell40 \bluejay_data_inst.state_FSM_i2_LC_17_13_6  (
            .in0(N__64419),
            .in1(N__78095),
            .in2(N__64423),
            .in3(N__68604),
            .lcout(n718),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97376),
            .ce(),
            .sr(N__73556));
    defparam \bluejay_data_inst.i2_3_lut_4_lut_LC_17_13_7 .C_ON=1'b0;
    defparam \bluejay_data_inst.i2_3_lut_4_lut_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i2_3_lut_4_lut_LC_17_13_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \bluejay_data_inst.i2_3_lut_4_lut_LC_17_13_7  (
            .in0(N__78129),
            .in1(N__64418),
            .in2(N__64396),
            .in3(N__68635),
            .lcout(\bluejay_data_inst.n10745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.state_FSM_i7_LC_17_14_0 .C_ON=1'b0;
    defparam \bluejay_data_inst.state_FSM_i7_LC_17_14_0 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.state_FSM_i7_LC_17_14_0 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \bluejay_data_inst.state_FSM_i7_LC_17_14_0  (
            .in0(N__68528),
            .in1(N__78069),
            .in2(N__64367),
            .in3(N__64713),
            .lcout(\bluejay_data_inst.bluejay_data_out_31__N_702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97383),
            .ce(),
            .sr(N__73559));
    defparam \bluejay_data_inst.state_FSM_i6_LC_17_14_1 .C_ON=1'b0;
    defparam \bluejay_data_inst.state_FSM_i6_LC_17_14_1 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.state_FSM_i6_LC_17_14_1 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \bluejay_data_inst.state_FSM_i6_LC_17_14_1  (
            .in0(N__68602),
            .in1(N__64381),
            .in2(N__64714),
            .in3(N__64349),
            .lcout(\bluejay_data_inst.n714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97383),
            .ce(),
            .sr(N__73559));
    defparam \bluejay_data_inst.state_FSM_i5_LC_17_14_2 .C_ON=1'b0;
    defparam \bluejay_data_inst.state_FSM_i5_LC_17_14_2 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.state_FSM_i5_LC_17_14_2 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \bluejay_data_inst.state_FSM_i5_LC_17_14_2  (
            .in0(N__68527),
            .in1(N__68601),
            .in2(N__69096),
            .in3(N__78068),
            .lcout(\bluejay_data_inst.n715 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97383),
            .ce(),
            .sr(N__73559));
    defparam \bluejay_data_inst.state_FSM_i8_LC_17_14_3 .C_ON=1'b0;
    defparam \bluejay_data_inst.state_FSM_i8_LC_17_14_3 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.state_FSM_i8_LC_17_14_3 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \bluejay_data_inst.state_FSM_i8_LC_17_14_3  (
            .in0(N__68603),
            .in1(N__69060),
            .in2(N__64729),
            .in3(N__68864),
            .lcout(bluejay_data_out_31__N_703),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97383),
            .ce(),
            .sr(N__73559));
    defparam \bluejay_data_inst.state_FSM_i9_LC_17_14_4 .C_ON=1'b0;
    defparam \bluejay_data_inst.state_FSM_i9_LC_17_14_4 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.state_FSM_i9_LC_17_14_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \bluejay_data_inst.state_FSM_i9_LC_17_14_4  (
            .in0(N__68865),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64728),
            .lcout(bluejay_data_out_31__N_704),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97383),
            .ce(),
            .sr(N__73559));
    defparam \bluejay_data_inst.i2_3_lut_LC_17_14_5 .C_ON=1'b0;
    defparam \bluejay_data_inst.i2_3_lut_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i2_3_lut_LC_17_14_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \bluejay_data_inst.i2_3_lut_LC_17_14_5  (
            .in0(N__64709),
            .in1(N__68863),
            .in2(_gnd_net_),
            .in3(N__64699),
            .lcout(\bluejay_data_inst.n108 ),
            .ltout(\bluejay_data_inst.n108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i11119_3_lut_LC_17_14_6 .C_ON=1'b0;
    defparam \bluejay_data_inst.i11119_3_lut_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i11119_3_lut_LC_17_14_6 .LUT_INIT=16'b0101010100000101;
    LogicCell40 \bluejay_data_inst.i11119_3_lut_LC_17_14_6  (
            .in0(N__73560),
            .in1(_gnd_net_),
            .in2(N__64687),
            .in3(N__68599),
            .lcout(\bluejay_data_inst.n4062 ),
            .ltout(\bluejay_data_inst.n4062_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i1_3_lut_4_lut_LC_17_14_7 .C_ON=1'b0;
    defparam \bluejay_data_inst.i1_3_lut_4_lut_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i1_3_lut_4_lut_LC_17_14_7 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \bluejay_data_inst.i1_3_lut_4_lut_LC_17_14_7  (
            .in0(N__68600),
            .in1(N__69059),
            .in2(N__64684),
            .in3(N__64674),
            .lcout(\bluejay_data_inst.n4519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i7_LC_17_15_0 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i7_LC_17_15_0 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i7_LC_17_15_0 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i7_LC_17_15_0  (
            .in0(N__78791),
            .in1(N__64639),
            .in2(N__64801),
            .in3(N__64768),
            .lcout(mem_LUT_data_raw_r_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97390),
            .ce(N__78655),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_12338_LC_17_15_1 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_12338_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_12338_LC_17_15_1 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_12338_LC_17_15_1  (
            .in0(N__79014),
            .in1(N__64755),
            .in2(N__64786),
            .in3(N__78793),
            .lcout(\tx_fifo.lscc_fifo_inst.n13952 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i9_4_lut_LC_17_15_2 .C_ON=1'b0;
    defparam \usb3_if_inst.i9_4_lut_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i9_4_lut_LC_17_15_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \usb3_if_inst.i9_4_lut_LC_17_15_2  (
            .in0(N__64633),
            .in1(N__64615),
            .in2(N__64594),
            .in3(N__64573),
            .lcout(),
            .ltout(\usb3_if_inst.n20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i10_4_lut_LC_17_15_3 .C_ON=1'b0;
    defparam \usb3_if_inst.i10_4_lut_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i10_4_lut_LC_17_15_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \usb3_if_inst.i10_4_lut_LC_17_15_3  (
            .in0(N__64561),
            .in1(N__64543),
            .in2(N__64522),
            .in3(N__64807),
            .lcout(\usb3_if_inst.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.i5_2_lut_LC_17_15_4 .C_ON=1'b0;
    defparam \usb3_if_inst.i5_2_lut_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \usb3_if_inst.i5_2_lut_LC_17_15_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \usb3_if_inst.i5_2_lut_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__64843),
            .in2(_gnd_net_),
            .in3(N__64825),
            .lcout(\usb3_if_inst.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i8_LC_17_15_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i8_LC_17_15_5 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i8_LC_17_15_5 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i8_LC_17_15_5  (
            .in0(N__78910),
            .in1(N__64909),
            .in2(N__64927),
            .in3(N__78792),
            .lcout(mem_LUT_data_raw_r_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97390),
            .ce(N__78655),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i152_153_LC_17_16_0 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i152_153_LC_17_16_0 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i152_153_LC_17_16_0 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i152_153_LC_17_16_0  (
            .in0(N__74529),
            .in1(N__69621),
            .in2(N__64869),
            .in3(N__64797),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97399),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i248_249_LC_17_16_1 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i248_249_LC_17_16_1 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i248_249_LC_17_16_1 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i248_249_LC_17_16_1  (
            .in0(N__64779),
            .in1(N__74530),
            .in2(N__73992),
            .in3(N__64864),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97399),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i56_57_LC_17_16_2 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i56_57_LC_17_16_2 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i56_57_LC_17_16_2 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i56_57_LC_17_16_2  (
            .in0(N__74532),
            .in1(N__73986),
            .in2(N__64870),
            .in3(N__64767),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97399),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i344_345_LC_17_16_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i344_345_LC_17_16_3 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i344_345_LC_17_16_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i344_345_LC_17_16_3  (
            .in0(N__69622),
            .in1(N__74531),
            .in2(N__64756),
            .in3(N__64865),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97399),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.Rx_Recv_Byte_i5_LC_17_16_4 .C_ON=1'b0;
    defparam \spi0.Rx_Recv_Byte_i5_LC_17_16_4 .SEQ_MODE=4'b1000;
    defparam \spi0.Rx_Recv_Byte_i5_LC_17_16_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.Rx_Recv_Byte_i5_LC_17_16_4  (
            .in0(N__69255),
            .in1(N__64739),
            .in2(_gnd_net_),
            .in3(N__65160),
            .lcout(rx_buf_byte_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97399),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.rx_shift_reg_i5_LC_17_16_5 .C_ON=1'b0;
    defparam \spi0.rx_shift_reg_i5_LC_17_16_5 .SEQ_MODE=4'b1000;
    defparam \spi0.rx_shift_reg_i5_LC_17_16_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \spi0.rx_shift_reg_i5_LC_17_16_5  (
            .in0(N__64740),
            .in1(N__64941),
            .in2(_gnd_net_),
            .in3(N__65225),
            .lcout(rx_shift_reg_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97399),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.rx_shift_reg_i6_LC_17_16_6 .C_ON=1'b0;
    defparam \spi0.rx_shift_reg_i6_LC_17_16_6 .SEQ_MODE=4'b1000;
    defparam \spi0.rx_shift_reg_i6_LC_17_16_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi0.rx_shift_reg_i6_LC_17_16_6  (
            .in0(N__65226),
            .in1(N__64883),
            .in2(_gnd_net_),
            .in3(N__64741),
            .lcout(rx_shift_reg_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97399),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.rx_shift_reg_i4_LC_17_16_7 .C_ON=1'b0;
    defparam \spi0.rx_shift_reg_i4_LC_17_16_7 .SEQ_MODE=4'b1000;
    defparam \spi0.rx_shift_reg_i4_LC_17_16_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.rx_shift_reg_i4_LC_17_16_7  (
            .in0(N__65113),
            .in1(N__64940),
            .in2(_gnd_net_),
            .in3(N__65224),
            .lcout(rx_shift_reg_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97399),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i59_60_LC_17_17_0 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i59_60_LC_17_17_0 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i59_60_LC_17_17_0 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i59_60_LC_17_17_0  (
            .in0(N__69468),
            .in1(N__74471),
            .in2(N__73982),
            .in3(N__64920),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97407),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i347_348_LC_17_17_1 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i347_348_LC_17_17_1 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i347_348_LC_17_17_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i347_348_LC_17_17_1  (
            .in0(N__69605),
            .in1(N__79062),
            .in2(N__74528),
            .in3(N__69467),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97407),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i341_342_LC_17_17_2 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i341_342_LC_17_17_2 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i341_342_LC_17_17_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i341_342_LC_17_17_2  (
            .in0(N__69228),
            .in1(N__74467),
            .in2(N__69271),
            .in3(N__69604),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97407),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i155_156_LC_17_17_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i155_156_LC_17_17_3 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i155_156_LC_17_17_3 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i155_156_LC_17_17_3  (
            .in0(N__74466),
            .in1(N__64905),
            .in2(N__69620),
            .in3(N__69466),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97407),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.Rx_Recv_Byte_i7_LC_17_17_4 .C_ON=1'b0;
    defparam \spi0.Rx_Recv_Byte_i7_LC_17_17_4 .SEQ_MODE=4'b1000;
    defparam \spi0.Rx_Recv_Byte_i7_LC_17_17_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.Rx_Recv_Byte_i7_LC_17_17_4  (
            .in0(N__69465),
            .in1(N__64893),
            .in2(_gnd_net_),
            .in3(N__65159),
            .lcout(rx_buf_byte_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97407),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.rx_shift_reg_i7_LC_17_17_5 .C_ON=1'b0;
    defparam \spi0.rx_shift_reg_i7_LC_17_17_5 .SEQ_MODE=4'b1000;
    defparam \spi0.rx_shift_reg_i7_LC_17_17_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \spi0.rx_shift_reg_i7_LC_17_17_5  (
            .in0(N__64894),
            .in1(N__65223),
            .in2(_gnd_net_),
            .in3(N__64885),
            .lcout(rx_shift_reg_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97407),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.Rx_Recv_Byte_i2_LC_17_17_6 .C_ON=1'b0;
    defparam \spi0.Rx_Recv_Byte_i2_LC_17_17_6 .SEQ_MODE=4'b1000;
    defparam \spi0.Rx_Recv_Byte_i2_LC_17_17_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.Rx_Recv_Byte_i2_LC_17_17_6  (
            .in0(N__74196),
            .in1(N__65248),
            .in2(_gnd_net_),
            .in3(N__65157),
            .lcout(rx_buf_byte_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97407),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.Rx_Recv_Byte_i6_LC_17_17_7 .C_ON=1'b0;
    defparam \spi0.Rx_Recv_Byte_i6_LC_17_17_7 .SEQ_MODE=4'b1000;
    defparam \spi0.Rx_Recv_Byte_i6_LC_17_17_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi0.Rx_Recv_Byte_i6_LC_17_17_7  (
            .in0(N__65158),
            .in1(N__64884),
            .in2(_gnd_net_),
            .in3(N__64860),
            .lcout(rx_buf_byte_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97407),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.Rx_Recv_Byte_i0_LC_17_18_0 .C_ON=1'b0;
    defparam \spi0.Rx_Recv_Byte_i0_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \spi0.Rx_Recv_Byte_i0_LC_17_18_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi0.Rx_Recv_Byte_i0_LC_17_18_0  (
            .in0(N__65154),
            .in1(N__65283),
            .in2(_gnd_net_),
            .in3(N__69543),
            .lcout(rx_buf_byte_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97419),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.rx_shift_reg_i1_LC_17_18_1 .C_ON=1'b0;
    defparam \spi0.rx_shift_reg_i1_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \spi0.rx_shift_reg_i1_LC_17_18_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \spi0.rx_shift_reg_i1_LC_17_18_1  (
            .in0(N__65284),
            .in1(N__65220),
            .in2(_gnd_net_),
            .in3(N__65259),
            .lcout(rx_shift_reg_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97419),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.rx_shift_reg_i2_LC_17_18_2 .C_ON=1'b0;
    defparam \spi0.rx_shift_reg_i2_LC_17_18_2 .SEQ_MODE=4'b1000;
    defparam \spi0.rx_shift_reg_i2_LC_17_18_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \spi0.rx_shift_reg_i2_LC_17_18_2  (
            .in0(N__65260),
            .in1(N__65221),
            .in2(_gnd_net_),
            .in3(N__65246),
            .lcout(rx_shift_reg_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97419),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.Rx_Recv_Byte_i1_LC_17_18_3 .C_ON=1'b0;
    defparam \spi0.Rx_Recv_Byte_i1_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \spi0.Rx_Recv_Byte_i1_LC_17_18_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi0.Rx_Recv_Byte_i1_LC_17_18_3  (
            .in0(N__73873),
            .in1(N__65258),
            .in2(_gnd_net_),
            .in3(N__65155),
            .lcout(rx_buf_byte_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97419),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.rx_shift_reg_i3_LC_17_18_4 .C_ON=1'b0;
    defparam \spi0.rx_shift_reg_i3_LC_17_18_4 .SEQ_MODE=4'b1000;
    defparam \spi0.rx_shift_reg_i3_LC_17_18_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \spi0.rx_shift_reg_i3_LC_17_18_4  (
            .in0(N__65247),
            .in1(N__65222),
            .in2(_gnd_net_),
            .in3(N__65109),
            .lcout(rx_shift_reg_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97419),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i6_LC_17_18_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i6_LC_17_18_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i6_LC_17_18_5 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_buffer__i6_LC_17_18_5  (
            .in0(N__78562),
            .in1(N__80861),
            .in2(N__73476),
            .in3(N__65328),
            .lcout(fifo_data_out_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97419),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.Rx_Recv_Byte_i3_LC_17_18_6 .C_ON=1'b0;
    defparam \spi0.Rx_Recv_Byte_i3_LC_17_18_6 .SEQ_MODE=4'b1000;
    defparam \spi0.Rx_Recv_Byte_i3_LC_17_18_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi0.Rx_Recv_Byte_i3_LC_17_18_6  (
            .in0(N__65156),
            .in1(N__65108),
            .in2(_gnd_net_),
            .in3(N__74014),
            .lcout(rx_buf_byte_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97419),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i9_LC_17_19_0 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i9_LC_17_19_0 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i9_LC_17_19_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i9_LC_17_19_0  (
            .in0(N__68914),
            .in1(N__65095),
            .in2(_gnd_net_),
            .in3(N__69016),
            .lcout(DATA8_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i9C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i8_LC_17_19_1 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i8_LC_17_19_1 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i8_LC_17_19_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i8_LC_17_19_1  (
            .in0(N__69015),
            .in1(N__65050),
            .in2(_gnd_net_),
            .in3(N__68913),
            .lcout(DATA7_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i9C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i5_LC_17_19_2 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i5_LC_17_19_2 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i5_LC_17_19_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i5_LC_17_19_2  (
            .in0(N__68910),
            .in1(N__64996),
            .in2(_gnd_net_),
            .in3(N__69012),
            .lcout(DATA20_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i9C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i4_LC_17_19_3 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i4_LC_17_19_3 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i4_LC_17_19_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i4_LC_17_19_3  (
            .in0(N__69011),
            .in1(N__65536),
            .in2(_gnd_net_),
            .in3(N__68909),
            .lcout(DATA19_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i9C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i3_LC_17_19_4 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i3_LC_17_19_4 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i3_LC_17_19_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i3_LC_17_19_4  (
            .in0(N__68908),
            .in1(N__65482),
            .in2(_gnd_net_),
            .in3(N__69010),
            .lcout(DATA18_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i9C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i2_LC_17_19_5 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i2_LC_17_19_5 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i2_LC_17_19_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i2_LC_17_19_5  (
            .in0(N__69009),
            .in1(N__65428),
            .in2(_gnd_net_),
            .in3(N__68907),
            .lcout(DATA17_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i9C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i6_LC_17_19_6 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i6_LC_17_19_6 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i6_LC_17_19_6 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i6_LC_17_19_6  (
            .in0(N__68911),
            .in1(N__65380),
            .in2(_gnd_net_),
            .in3(N__69013),
            .lcout(DATA5_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i9C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i7_LC_17_19_7 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i7_LC_17_19_7 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i7_LC_17_19_7 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i7_LC_17_19_7  (
            .in0(N__69014),
            .in1(N__65329),
            .in2(_gnd_net_),
            .in3(N__68912),
            .lcout(DATA6_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i9C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i1311_3_lut_LC_17_20_2 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i1311_3_lut_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.i1311_3_lut_LC_17_20_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i1311_3_lut_LC_17_20_2  (
            .in0(N__74274),
            .in1(N__69889),
            .in2(_gnd_net_),
            .in3(N__74426),
            .lcout(),
            .ltout(wr_addr_p1_w_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_r__i2_LC_17_20_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_r__i2_LC_17_20_3 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_r__i2_LC_17_20_3 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.wr_addr_r__i2_LC_17_20_3  (
            .in0(N__69890),
            .in1(N__74350),
            .in2(N__65287),
            .in3(N__69938),
            .lcout(wr_addr_r_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97433),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_r__i1_LC_17_20_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_r__i1_LC_17_20_5 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_r__i1_LC_17_20_5 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.wr_addr_r__i1_LC_17_20_5  (
            .in0(N__74427),
            .in1(N__74275),
            .in2(N__78387),
            .in3(N__74349),
            .lcout(wr_addr_r_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97433),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.usb3_data_in_latched__i9_LC_18_1_0 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i9_LC_18_1_0 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i9_LC_18_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i9_LC_18_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65764),
            .lcout(\usb3_if_inst.usb3_data_in_latched_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93455),
            .ce(),
            .sr(N__73710));
    defparam \usb3_if_inst.usb3_data_in_latched__i3_LC_18_1_5 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i3_LC_18_1_5 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i3_LC_18_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i3_LC_18_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65752),
            .lcout(\usb3_if_inst.usb3_data_in_latched_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93455),
            .ce(),
            .sr(N__73710));
    defparam \usb3_if_inst.usb3_data_in_latched__i2_LC_18_1_7 .C_ON=1'b0;
    defparam \usb3_if_inst.usb3_data_in_latched__i2_LC_18_1_7 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.usb3_data_in_latched__i2_LC_18_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.usb3_data_in_latched__i2_LC_18_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65731),
            .lcout(\usb3_if_inst.usb3_data_in_latched_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93455),
            .ce(),
            .sr(N__73710));
    defparam \usb3_if_inst.dc32_fifo_data_in_i9_LC_18_2_0 .C_ON=1'b0;
    defparam \usb3_if_inst.dc32_fifo_data_in_i9_LC_18_2_0 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.dc32_fifo_data_in_i9_LC_18_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.dc32_fifo_data_in_i9_LC_18_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65710),
            .lcout(dc32_fifo_data_in_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVusb3_if_inst.dc32_fifo_data_in_i9C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1688_1689_LC_18_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1688_1689_LC_18_4_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1688_1689_LC_18_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1688_1689_LC_18_4_0  (
            .in0(N__96353),
            .in1(N__65703),
            .in2(_gnd_net_),
            .in3(N__66589),
            .lcout(REG_mem_17_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93438),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11864_LC_18_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11864_LC_18_4_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11864_LC_18_4_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11864_LC_18_4_1  (
            .in0(N__65545),
            .in1(N__92442),
            .in2(N__66091),
            .in3(N__88877),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13658_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13658_bdd_4_lut_LC_18_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13658_bdd_4_lut_LC_18_4_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13658_bdd_4_lut_LC_18_4_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13658_bdd_4_lut_LC_18_4_2  (
            .in0(N__92441),
            .in1(N__65704),
            .in2(N__65695),
            .in3(N__65554),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13661 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1592_1593_LC_18_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1592_1593_LC_18_4_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1592_1593_LC_18_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1592_1593_LC_18_4_3  (
            .in0(N__65553),
            .in1(N__96357),
            .in2(_gnd_net_),
            .in3(N__65692),
            .lcout(REG_mem_16_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93438),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1784_1785_LC_18_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1784_1785_LC_18_4_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1784_1785_LC_18_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1784_1785_LC_18_4_4  (
            .in0(N__96354),
            .in1(N__65544),
            .in2(_gnd_net_),
            .in3(N__67511),
            .lcout(REG_mem_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93438),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1880_1881_LC_18_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1880_1881_LC_18_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1880_1881_LC_18_4_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1880_1881_LC_18_4_5  (
            .in0(N__66087),
            .in1(N__96358),
            .in2(_gnd_net_),
            .in3(N__72114),
            .lcout(REG_mem_19_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93438),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i920_921_LC_18_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i920_921_LC_18_4_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i920_921_LC_18_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i920_921_LC_18_4_6  (
            .in0(N__96355),
            .in1(N__70152),
            .in2(_gnd_net_),
            .in3(N__67198),
            .lcout(REG_mem_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93438),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1016_1017_LC_18_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1016_1017_LC_18_4_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1016_1017_LC_18_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1016_1017_LC_18_4_7  (
            .in0(N__66072),
            .in1(N__96356),
            .in2(_gnd_net_),
            .in3(N__66997),
            .lcout(REG_mem_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93438),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11978_LC_18_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11978_LC_18_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11978_LC_18_5_0 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11978_LC_18_5_0  (
            .in0(N__91862),
            .in1(N__88851),
            .in2(N__66079),
            .in3(N__66061),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13778 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5132_5133_LC_18_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5132_5133_LC_18_5_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5132_5133_LC_18_5_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5132_5133_LC_18_5_1  (
            .in0(N__75806),
            .in1(N__95333),
            .in2(N__66045),
            .in3(N__77036),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93433),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3992_3993_LC_18_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3992_3993_LC_18_5_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3992_3993_LC_18_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3992_3993_LC_18_5_2  (
            .in0(N__96152),
            .in1(N__74571),
            .in2(_gnd_net_),
            .in3(N__66028),
            .lcout(REG_mem_41_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93433),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3896_3897_LC_18_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3896_3897_LC_18_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3896_3897_LC_18_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3896_3897_LC_18_5_3  (
            .in0(N__75222),
            .in1(N__96154),
            .in2(_gnd_net_),
            .in3(N__65902),
            .lcout(REG_mem_40_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93433),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4088_4089_LC_18_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4088_4089_LC_18_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4088_4089_LC_18_5_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4088_4089_LC_18_5_4  (
            .in0(N__96153),
            .in1(N__74586),
            .in2(_gnd_net_),
            .in3(N__68092),
            .lcout(REG_mem_42_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93433),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4184_4185_LC_18_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4184_4185_LC_18_5_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4184_4185_LC_18_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4184_4185_LC_18_5_5  (
            .in0(N__74607),
            .in1(N__96155),
            .in2(_gnd_net_),
            .in3(N__68298),
            .lcout(REG_mem_43_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93433),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i446_447_LC_18_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i446_447_LC_18_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i446_447_LC_18_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i446_447_LC_18_5_6  (
            .in0(N__77607),
            .in1(N__89277),
            .in2(_gnd_net_),
            .in3(N__72729),
            .lcout(REG_mem_4_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93433),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i632_633_LC_18_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i632_633_LC_18_5_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i632_633_LC_18_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i632_633_LC_18_5_7  (
            .in0(N__79152),
            .in1(N__96156),
            .in2(_gnd_net_),
            .in3(N__66429),
            .lcout(REG_mem_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93433),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4568_4569_LC_18_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4568_4569_LC_18_6_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4568_4569_LC_18_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4568_4569_LC_18_6_0  (
            .in0(N__71919),
            .in1(N__96350),
            .in2(_gnd_net_),
            .in3(N__66274),
            .lcout(REG_mem_47_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6104_6105_LC_18_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6104_6105_LC_18_6_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6104_6105_LC_18_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6104_6105_LC_18_6_1  (
            .in0(N__96349),
            .in1(N__71022),
            .in2(_gnd_net_),
            .in3(N__67714),
            .lcout(REG_mem_63_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10032_3_lut_LC_18_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10032_3_lut_LC_18_6_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10032_3_lut_LC_18_6_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10032_3_lut_LC_18_6_2  (
            .in0(N__71617),
            .in1(N__88835),
            .in2(_gnd_net_),
            .in3(N__66130),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11681_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11610_LC_18_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11610_LC_18_6_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11610_LC_18_6_3 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11610_LC_18_6_3  (
            .in0(N__91861),
            .in1(N__85627),
            .in2(N__66109),
            .in3(N__71032),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2846_2847_LC_18_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2846_2847_LC_18_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2846_2847_LC_18_6_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2846_2847_LC_18_6_4  (
            .in0(N__95323),
            .in1(N__89326),
            .in2(N__90435),
            .in3(N__71005),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_29_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2057_2058_LC_18_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2057_2058_LC_18_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2057_2058_LC_18_6_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2057_2058_LC_18_6_5  (
            .in0(N__96772),
            .in1(N__95324),
            .in2(N__71062),
            .in3(N__77035),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i536_537_LC_18_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i536_537_LC_18_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i536_537_LC_18_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i536_537_LC_18_6_6  (
            .in0(N__71157),
            .in1(N__96351),
            .in2(_gnd_net_),
            .in3(N__67873),
            .lcout(REG_mem_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i542_543_LC_18_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i542_543_LC_18_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i542_543_LC_18_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i542_543_LC_18_6_7  (
            .in0(N__89325),
            .in1(N__77628),
            .in2(_gnd_net_),
            .in3(N__67874),
            .lcout(REG_mem_5_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93427),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10158_3_lut_LC_18_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10158_3_lut_LC_18_7_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10158_3_lut_LC_18_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10158_3_lut_LC_18_7_0  (
            .in0(N__88778),
            .in1(N__66667),
            .in2(_gnd_net_),
            .in3(N__66838),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11525_LC_18_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11525_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11525_LC_18_7_1 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11525_LC_18_7_1  (
            .in0(N__85262),
            .in1(N__72274),
            .in2(N__92628),
            .in3(N__67021),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13238_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13238_bdd_4_lut_LC_18_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13238_bdd_4_lut_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13238_bdd_4_lut_LC_18_7_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13238_bdd_4_lut_LC_18_7_2  (
            .in0(N__66625),
            .in1(N__85261),
            .in2(N__67012),
            .in3(N__67009),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1004_1005_LC_18_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1004_1005_LC_18_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1004_1005_LC_18_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1004_1005_LC_18_7_3  (
            .in0(N__66837),
            .in1(N__75921),
            .in2(_gnd_net_),
            .in3(N__66995),
            .lcout(REG_mem_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93421),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1100_1101_LC_18_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1100_1101_LC_18_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1100_1101_LC_18_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1100_1101_LC_18_7_4  (
            .in0(N__75920),
            .in1(N__66666),
            .in2(_gnd_net_),
            .in3(N__66826),
            .lcout(REG_mem_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93421),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10157_3_lut_LC_18_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10157_3_lut_LC_18_7_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10157_3_lut_LC_18_7_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10157_3_lut_LC_18_7_5  (
            .in0(N__66658),
            .in1(N__88777),
            .in2(_gnd_net_),
            .in3(N__66637),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4946_4947_LC_18_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4946_4947_LC_18_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4946_4947_LC_18_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4946_4947_LC_18_7_6  (
            .in0(N__66603),
            .in1(N__76639),
            .in2(_gnd_net_),
            .in3(N__72265),
            .lcout(REG_mem_51_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93421),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12443_LC_18_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12443_LC_18_7_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12443_LC_18_7_7 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12443_LC_18_7_7  (
            .in0(N__92495),
            .in1(N__88779),
            .in2(N__66619),
            .in3(N__66604),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1694_1695_LC_18_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1694_1695_LC_18_8_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1694_1695_LC_18_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1694_1695_LC_18_8_0  (
            .in0(N__67542),
            .in1(N__89301),
            .in2(_gnd_net_),
            .in3(N__66588),
            .lcout(REG_mem_17_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12243_LC_18_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12243_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12243_LC_18_8_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12243_LC_18_8_1  (
            .in0(N__91815),
            .in1(N__88595),
            .in2(N__71941),
            .in3(N__67354),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14108_bdd_4_lut_LC_18_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14108_bdd_4_lut_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14108_bdd_4_lut_LC_18_8_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14108_bdd_4_lut_LC_18_8_2  (
            .in0(N__67543),
            .in1(N__91814),
            .in2(N__67531),
            .in3(N__67528),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11691 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3128_3129_LC_18_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3128_3129_LC_18_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3128_3129_LC_18_8_3 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3128_3129_LC_18_8_3  (
            .in0(N__96312),
            .in1(N__94828),
            .in2(N__79182),
            .in3(N__82954),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1790_1791_LC_18_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1790_1791_LC_18_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1790_1791_LC_18_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1790_1791_LC_18_8_4  (
            .in0(N__67353),
            .in1(N__89302),
            .in2(_gnd_net_),
            .in3(N__67503),
            .lcout(REG_mem_18_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2174_2175_LC_18_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2174_2175_LC_18_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2174_2175_LC_18_8_5 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2174_2175_LC_18_8_5  (
            .in0(N__89300),
            .in1(N__76344),
            .in2(N__72351),
            .in3(N__94829),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i830_831_LC_18_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i830_831_LC_18_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i830_831_LC_18_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i830_831_LC_18_8_6  (
            .in0(N__82986),
            .in1(N__89303),
            .in2(_gnd_net_),
            .in3(N__67345),
            .lcout(REG_mem_8_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i926_927_LC_18_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i926_927_LC_18_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i926_927_LC_18_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i926_927_LC_18_8_7  (
            .in0(N__89299),
            .in1(N__83007),
            .in2(_gnd_net_),
            .in3(N__67193),
            .lcout(REG_mem_9_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93414),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i434_435_LC_18_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i434_435_LC_18_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i434_435_LC_18_9_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i434_435_LC_18_9_0  (
            .in0(N__68109),
            .in1(N__76636),
            .in2(_gnd_net_),
            .in3(N__72712),
            .lcout(REG_mem_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93405),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13808_bdd_4_lut_LC_18_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13808_bdd_4_lut_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13808_bdd_4_lut_LC_18_9_1 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13808_bdd_4_lut_LC_18_9_1  (
            .in0(N__67057),
            .in1(N__91809),
            .in2(N__67045),
            .in3(N__67036),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11784 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10866_3_lut_LC_18_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10866_3_lut_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10866_3_lut_LC_18_9_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10866_3_lut_LC_18_9_2  (
            .in0(N__67740),
            .in1(N__88742),
            .in2(_gnd_net_),
            .in3(N__67728),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11973_LC_18_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11973_LC_18_9_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11973_LC_18_9_3 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11973_LC_18_9_3  (
            .in0(N__85735),
            .in1(N__91810),
            .in2(N__67921),
            .in3(N__68098),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13784_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13784_bdd_4_lut_LC_18_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13784_bdd_4_lut_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13784_bdd_4_lut_LC_18_9_4 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13784_bdd_4_lut_LC_18_9_4  (
            .in0(N__67909),
            .in1(N__85734),
            .in2(N__67903),
            .in3(N__67900),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i530_531_LC_18_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i530_531_LC_18_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i530_531_LC_18_9_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i530_531_LC_18_9_5  (
            .in0(N__76635),
            .in1(N__68121),
            .in2(_gnd_net_),
            .in3(N__67879),
            .lcout(REG_mem_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93405),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i242_243_LC_18_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i242_243_LC_18_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i242_243_LC_18_9_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i242_243_LC_18_9_6  (
            .in0(N__76637),
            .in1(N__94827),
            .in2(N__67741),
            .in3(N__80607),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93405),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i338_339_LC_18_9_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i338_339_LC_18_9_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i338_339_LC_18_9_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i338_339_LC_18_9_7  (
            .in0(N__94826),
            .in1(N__76638),
            .in2(N__67729),
            .in3(N__83290),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93405),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6110_6111_LC_18_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6110_6111_LC_18_10_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6110_6111_LC_18_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6110_6111_LC_18_10_0  (
            .in0(N__89275),
            .in1(N__67572),
            .in2(_gnd_net_),
            .in3(N__67674),
            .lcout(REG_mem_63_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11635_LC_18_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11635_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11635_LC_18_10_1 .LUT_INIT=16'b1100101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11635_LC_18_10_1  (
            .in0(N__68133),
            .in1(N__67573),
            .in2(N__88850),
            .in3(N__91808),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13382_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13382_bdd_4_lut_LC_18_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13382_bdd_4_lut_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13382_bdd_4_lut_LC_18_10_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13382_bdd_4_lut_LC_18_10_2  (
            .in0(N__67561),
            .in1(N__91732),
            .in2(N__67546),
            .in3(N__68310),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11874 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5918_5919_LC_18_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5918_5919_LC_18_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5918_5919_LC_18_10_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5918_5919_LC_18_10_3  (
            .in0(N__89437),
            .in1(N__95102),
            .in2(N__68311),
            .in3(N__70991),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4178_4179_LC_18_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4178_4179_LC_18_10_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4178_4179_LC_18_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4178_4179_LC_18_10_4  (
            .in0(N__68145),
            .in1(N__76743),
            .in2(_gnd_net_),
            .in3(N__68296),
            .lcout(REG_mem_43_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6014_6015_LC_18_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6014_6015_LC_18_10_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6014_6015_LC_18_10_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6014_6015_LC_18_10_5  (
            .in0(N__89438),
            .in1(N__95103),
            .in2(N__68134),
            .in3(N__77923),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10871_3_lut_LC_18_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10871_3_lut_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10871_3_lut_LC_18_10_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10871_3_lut_LC_18_10_6  (
            .in0(N__68122),
            .in1(N__88738),
            .in2(_gnd_net_),
            .in3(N__68110),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12520 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4094_4095_LC_18_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4094_4095_LC_18_10_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4094_4095_LC_18_10_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4094_4095_LC_18_10_7  (
            .in0(N__85917),
            .in1(N__89276),
            .in2(_gnd_net_),
            .in3(N__68086),
            .lcout(REG_mem_42_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93379),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.v_counter_i0_LC_18_11_0 .C_ON=1'b1;
    defparam \bluejay_data_inst.v_counter_i0_LC_18_11_0 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.v_counter_i0_LC_18_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \bluejay_data_inst.v_counter_i0_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(N__68724),
            .in2(N__68542),
            .in3(N__67933),
            .lcout(\bluejay_data_inst.v_counter_0 ),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\bluejay_data_inst.n10643 ),
            .clk(N__97362),
            .ce(N__68626),
            .sr(N__73561));
    defparam \bluejay_data_inst.v_counter_i1_LC_18_11_1 .C_ON=1'b1;
    defparam \bluejay_data_inst.v_counter_i1_LC_18_11_1 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.v_counter_i1_LC_18_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \bluejay_data_inst.v_counter_i1_LC_18_11_1  (
            .in0(_gnd_net_),
            .in1(N__68322),
            .in2(N__86582),
            .in3(N__67930),
            .lcout(\bluejay_data_inst.v_counter_1 ),
            .ltout(),
            .carryin(\bluejay_data_inst.n10643 ),
            .carryout(\bluejay_data_inst.n10644 ),
            .clk(N__97362),
            .ce(N__68626),
            .sr(N__73561));
    defparam \bluejay_data_inst.v_counter_i2_LC_18_11_2 .C_ON=1'b1;
    defparam \bluejay_data_inst.v_counter_i2_LC_18_11_2 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.v_counter_i2_LC_18_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \bluejay_data_inst.v_counter_i2_LC_18_11_2  (
            .in0(_gnd_net_),
            .in1(N__86513),
            .in2(N__68775),
            .in3(N__67927),
            .lcout(\bluejay_data_inst.v_counter_2 ),
            .ltout(),
            .carryin(\bluejay_data_inst.n10644 ),
            .carryout(\bluejay_data_inst.n10645 ),
            .clk(N__97362),
            .ce(N__68626),
            .sr(N__73561));
    defparam \bluejay_data_inst.v_counter_i3_LC_18_11_3 .C_ON=1'b1;
    defparam \bluejay_data_inst.v_counter_i3_LC_18_11_3 .SEQ_MODE=4'b1001;
    defparam \bluejay_data_inst.v_counter_i3_LC_18_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \bluejay_data_inst.v_counter_i3_LC_18_11_3  (
            .in0(_gnd_net_),
            .in1(N__68672),
            .in2(N__86583),
            .in3(N__67924),
            .lcout(\bluejay_data_inst.v_counter_3 ),
            .ltout(),
            .carryin(\bluejay_data_inst.n10645 ),
            .carryout(\bluejay_data_inst.n10646 ),
            .clk(N__97362),
            .ce(N__68626),
            .sr(N__73561));
    defparam \bluejay_data_inst.v_counter_i4_LC_18_11_4 .C_ON=1'b1;
    defparam \bluejay_data_inst.v_counter_i4_LC_18_11_4 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.v_counter_i4_LC_18_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \bluejay_data_inst.v_counter_i4_LC_18_11_4  (
            .in0(_gnd_net_),
            .in1(N__86517),
            .in2(N__68757),
            .in3(N__68389),
            .lcout(\bluejay_data_inst.v_counter_4 ),
            .ltout(),
            .carryin(\bluejay_data_inst.n10646 ),
            .carryout(\bluejay_data_inst.n10647 ),
            .clk(N__97362),
            .ce(N__68626),
            .sr(N__73561));
    defparam \bluejay_data_inst.v_counter_i5_LC_18_11_5 .C_ON=1'b1;
    defparam \bluejay_data_inst.v_counter_i5_LC_18_11_5 .SEQ_MODE=4'b1001;
    defparam \bluejay_data_inst.v_counter_i5_LC_18_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \bluejay_data_inst.v_counter_i5_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__68691),
            .in2(N__86584),
            .in3(N__68386),
            .lcout(\bluejay_data_inst.v_counter_5 ),
            .ltout(),
            .carryin(\bluejay_data_inst.n10647 ),
            .carryout(\bluejay_data_inst.n10648 ),
            .clk(N__97362),
            .ce(N__68626),
            .sr(N__73561));
    defparam \bluejay_data_inst.v_counter_i6_LC_18_11_6 .C_ON=1'b1;
    defparam \bluejay_data_inst.v_counter_i6_LC_18_11_6 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.v_counter_i6_LC_18_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \bluejay_data_inst.v_counter_i6_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__86521),
            .in2(N__68654),
            .in3(N__68383),
            .lcout(\bluejay_data_inst.v_counter_6 ),
            .ltout(),
            .carryin(\bluejay_data_inst.n10648 ),
            .carryout(\bluejay_data_inst.n10649 ),
            .clk(N__97362),
            .ce(N__68626),
            .sr(N__73561));
    defparam \bluejay_data_inst.v_counter_i7_LC_18_11_7 .C_ON=1'b1;
    defparam \bluejay_data_inst.v_counter_i7_LC_18_11_7 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.v_counter_i7_LC_18_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \bluejay_data_inst.v_counter_i7_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(N__68337),
            .in2(N__86585),
            .in3(N__68380),
            .lcout(\bluejay_data_inst.v_counter_7 ),
            .ltout(),
            .carryin(\bluejay_data_inst.n10649 ),
            .carryout(\bluejay_data_inst.n10650 ),
            .clk(N__97362),
            .ce(N__68626),
            .sr(N__73561));
    defparam \bluejay_data_inst.v_counter_i8_LC_18_12_0 .C_ON=1'b1;
    defparam \bluejay_data_inst.v_counter_i8_LC_18_12_0 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.v_counter_i8_LC_18_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \bluejay_data_inst.v_counter_i8_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(N__68739),
            .in2(N__86426),
            .in3(N__68377),
            .lcout(\bluejay_data_inst.v_counter_8 ),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\bluejay_data_inst.n10651 ),
            .clk(N__97377),
            .ce(N__68622),
            .sr(N__73557));
    defparam \bluejay_data_inst.v_counter_i9_LC_18_12_1 .C_ON=1'b1;
    defparam \bluejay_data_inst.v_counter_i9_LC_18_12_1 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.v_counter_i9_LC_18_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \bluejay_data_inst.v_counter_i9_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__68355),
            .in2(N__86425),
            .in3(N__68374),
            .lcout(\bluejay_data_inst.v_counter_9 ),
            .ltout(),
            .carryin(\bluejay_data_inst.n10651 ),
            .carryout(\bluejay_data_inst.n10652 ),
            .clk(N__97377),
            .ce(N__68622),
            .sr(N__73557));
    defparam \bluejay_data_inst.v_counter_i10_LC_18_12_2 .C_ON=1'b0;
    defparam \bluejay_data_inst.v_counter_i10_LC_18_12_2 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.v_counter_i10_LC_18_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \bluejay_data_inst.v_counter_i10_LC_18_12_2  (
            .in0(N__68367),
            .in1(N__86295),
            .in2(_gnd_net_),
            .in3(N__68371),
            .lcout(\bluejay_data_inst.v_counter_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97377),
            .ce(N__68622),
            .sr(N__73557));
    defparam \bluejay_data_inst.i6_4_lut_LC_18_13_0 .C_ON=1'b0;
    defparam \bluejay_data_inst.i6_4_lut_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i6_4_lut_LC_18_13_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \bluejay_data_inst.i6_4_lut_LC_18_13_0  (
            .in0(N__68368),
            .in1(N__68356),
            .in2(N__68344),
            .in3(N__68326),
            .lcout(\bluejay_data_inst.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i9770_2_lut_LC_18_13_1 .C_ON=1'b0;
    defparam \bluejay_data_inst.i9770_2_lut_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i9770_2_lut_LC_18_13_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \bluejay_data_inst.i9770_2_lut_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(N__68656),
            .in2(_gnd_net_),
            .in3(N__68704),
            .lcout(),
            .ltout(\bluejay_data_inst.n11418_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i1_4_lut_adj_60_LC_18_13_2 .C_ON=1'b0;
    defparam \bluejay_data_inst.i1_4_lut_adj_60_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i1_4_lut_adj_60_LC_18_13_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \bluejay_data_inst.i1_4_lut_adj_60_LC_18_13_2  (
            .in0(N__78127),
            .in1(N__68697),
            .in2(N__68788),
            .in3(N__68679),
            .lcout(\bluejay_data_inst.n11330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i2_2_lut_LC_18_13_3 .C_ON=1'b0;
    defparam \bluejay_data_inst.i2_2_lut_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i2_2_lut_LC_18_13_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \bluejay_data_inst.i2_2_lut_LC_18_13_3  (
            .in0(N__68776),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68758),
            .lcout(),
            .ltout(\bluejay_data_inst.n10_adj_1180_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i7_4_lut_LC_18_13_4 .C_ON=1'b0;
    defparam \bluejay_data_inst.i7_4_lut_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i7_4_lut_LC_18_13_4 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \bluejay_data_inst.i7_4_lut_LC_18_13_4  (
            .in0(N__68740),
            .in1(N__68728),
            .in2(N__68713),
            .in3(N__68710),
            .lcout(\bluejay_data_inst.n10 ),
            .ltout(\bluejay_data_inst.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i3_4_lut_LC_18_13_5 .C_ON=1'b0;
    defparam \bluejay_data_inst.i3_4_lut_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i3_4_lut_LC_18_13_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \bluejay_data_inst.i3_4_lut_LC_18_13_5  (
            .in0(N__68698),
            .in1(N__68680),
            .in2(N__68659),
            .in3(N__68655),
            .lcout(\bluejay_data_inst.n10781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i1_2_lut_adj_59_LC_18_13_6 .C_ON=1'b0;
    defparam \bluejay_data_inst.i1_2_lut_adj_59_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i1_2_lut_adj_59_LC_18_13_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \bluejay_data_inst.i1_2_lut_adj_59_LC_18_13_6  (
            .in0(N__73537),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78126),
            .lcout(\bluejay_data_inst.n4162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.state_FSM_i10_LC_18_13_7 .C_ON=1'b0;
    defparam \bluejay_data_inst.state_FSM_i10_LC_18_13_7 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.state_FSM_i10_LC_18_13_7 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \bluejay_data_inst.state_FSM_i10_LC_18_13_7  (
            .in0(N__68981),
            .in1(N__68605),
            .in2(N__68538),
            .in3(N__78128),
            .lcout(\bluejay_data_inst.n710 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97384),
            .ce(),
            .sr(N__73536));
    defparam \bluejay_data_inst.bluejay_data_out_i14_LC_18_14_0 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i14_LC_18_14_0 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i14_LC_18_14_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i14_LC_18_14_0  (
            .in0(N__68867),
            .in1(N__68506),
            .in2(_gnd_net_),
            .in3(N__68964),
            .lcout(DATA13_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i14C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i13_LC_18_14_1 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i13_LC_18_14_1 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i13_LC_18_14_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i13_LC_18_14_1  (
            .in0(N__68963),
            .in1(N__68440),
            .in2(_gnd_net_),
            .in3(N__68866),
            .lcout(DATA12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i14C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i11075_2_lut_LC_18_14_2 .C_ON=1'b0;
    defparam \bluejay_data_inst.i11075_2_lut_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i11075_2_lut_LC_18_14_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \bluejay_data_inst.i11075_2_lut_LC_18_14_2  (
            .in0(N__78046),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69153),
            .lcout(\bluejay_data_inst.n7424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i3240_2_lut_LC_18_14_3 .C_ON=1'b0;
    defparam \bluejay_data_inst.i3240_2_lut_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i3240_2_lut_LC_18_14_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \bluejay_data_inst.i3240_2_lut_LC_18_14_3  (
            .in0(N__69154),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69092),
            .lcout(\bluejay_data_inst.n4442 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.get_next_word_57_LC_18_14_4 .C_ON=1'b0;
    defparam \bluejay_data_inst.get_next_word_57_LC_18_14_4 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.get_next_word_57_LC_18_14_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \bluejay_data_inst.get_next_word_57_LC_18_14_4  (
            .in0(N__68869),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69061),
            .lcout(get_next_word),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i14C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i20_3_lut_LC_18_14_5 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i20_3_lut_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i20_3_lut_LC_18_14_5 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \timing_controller_inst.mux_855_i20_3_lut_LC_18_14_5  (
            .in0(N__84316),
            .in1(N__82291),
            .in2(_gnd_net_),
            .in3(N__82420),
            .lcout(\timing_controller_inst.n1735 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i21_3_lut_LC_18_14_6 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i21_3_lut_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i21_3_lut_LC_18_14_6 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \timing_controller_inst.mux_855_i21_3_lut_LC_18_14_6  (
            .in0(N__82292),
            .in1(_gnd_net_),
            .in2(N__82426),
            .in3(N__84796),
            .lcout(\timing_controller_inst.n1734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.bluejay_data_out_i15_LC_18_14_7 .C_ON=1'b0;
    defparam \bluejay_data_inst.bluejay_data_out_i15_LC_18_14_7 .SEQ_MODE=4'b1000;
    defparam \bluejay_data_inst.bluejay_data_out_i15_LC_18_14_7 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \bluejay_data_inst.bluejay_data_out_i15_LC_18_14_7  (
            .in0(N__68965),
            .in1(N__68938),
            .in2(_gnd_net_),
            .in3(N__68868),
            .lcout(DATA14_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVbluejay_data_inst.bluejay_data_out_i14C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11774_LC_18_15_1 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11774_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11774_LC_18_15_1 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11774_LC_18_15_1  (
            .in0(N__78771),
            .in1(N__69199),
            .in2(N__79024),
            .in3(N__69511),
            .lcout(),
            .ltout(\tx_fifo.lscc_fifo_inst.n13544_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i3_LC_18_15_2 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i3_LC_18_15_2 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i3_LC_18_15_2 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i3_LC_18_15_2  (
            .in0(N__74176),
            .in1(N__69213),
            .in2(N__68791),
            .in3(N__78768),
            .lcout(mem_LUT_data_raw_r_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97400),
            .ce(N__78654),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11949_LC_18_15_4 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11949_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11949_LC_18_15_4 .LUT_INIT=16'b1100101011110000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11949_LC_18_15_4  (
            .in0(N__69736),
            .in1(N__69652),
            .in2(N__79025),
            .in3(N__78772),
            .lcout(),
            .ltout(\tx_fifo.lscc_fifo_inst.n13694_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i5_LC_18_15_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i5_LC_18_15_5 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i5_LC_18_15_5 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i5_LC_18_15_5  (
            .in0(N__78769),
            .in1(N__69499),
            .in2(N__69235),
            .in3(N__69487),
            .lcout(mem_LUT_data_raw_r_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97400),
            .ce(N__78654),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_12103_LC_18_15_6 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_12103_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_12103_LC_18_15_6 .LUT_INIT=16'b1010110011110000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_12103_LC_18_15_6  (
            .in0(N__69232),
            .in1(N__69667),
            .in2(N__79026),
            .in3(N__78773),
            .lcout(),
            .ltout(\tx_fifo.lscc_fifo_inst.n13766_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i6_LC_18_15_7 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i6_LC_18_15_7 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i6_LC_18_15_7 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i6_LC_18_15_7  (
            .in0(N__78770),
            .in1(N__69301),
            .in2(N__69217),
            .in3(N__69286),
            .lcout(mem_LUT_data_raw_r_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97400),
            .ce(N__78654),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i137_138_LC_18_16_0 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i137_138_LC_18_16_0 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i137_138_LC_18_16_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i137_138_LC_18_16_0  (
            .in0(N__69613),
            .in1(N__74533),
            .in2(N__79107),
            .in3(N__73885),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97408),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i329_330_LC_18_16_1 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i329_330_LC_18_16_1 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i329_330_LC_18_16_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i329_330_LC_18_16_1  (
            .in0(N__74538),
            .in1(N__69617),
            .in2(N__73895),
            .in3(N__79134),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97408),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i140_141_LC_18_16_2 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i140_141_LC_18_16_2 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i140_141_LC_18_16_2 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i140_141_LC_18_16_2  (
            .in0(N__69614),
            .in1(N__74534),
            .in2(N__69214),
            .in3(N__74197),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97408),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i332_333_LC_18_16_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i332_333_LC_18_16_3 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i332_333_LC_18_16_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i332_333_LC_18_16_3  (
            .in0(N__74539),
            .in1(N__69618),
            .in2(N__74205),
            .in3(N__69198),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97408),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i143_144_LC_18_16_4 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i143_144_LC_18_16_4 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i143_144_LC_18_16_4 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i143_144_LC_18_16_4  (
            .in0(N__69615),
            .in1(N__74535),
            .in2(N__78891),
            .in3(N__74024),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97408),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i335_336_LC_18_16_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i335_336_LC_18_16_5 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i335_336_LC_18_16_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i335_336_LC_18_16_5  (
            .in0(N__74540),
            .in1(N__69619),
            .in2(N__74031),
            .in3(N__73854),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97408),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i236_237_LC_18_16_6 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i236_237_LC_18_16_6 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i236_237_LC_18_16_6 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i236_237_LC_18_16_6  (
            .in0(N__69510),
            .in1(N__74537),
            .in2(N__73987),
            .in3(N__74198),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97408),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i146_147_LC_18_16_7 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i146_147_LC_18_16_7 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i146_147_LC_18_16_7 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i146_147_LC_18_16_7  (
            .in0(N__74536),
            .in1(N__69498),
            .in2(N__69772),
            .in3(N__69616),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97408),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i38_39_LC_18_17_0 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i38_39_LC_18_17_0 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i38_39_LC_18_17_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i38_39_LC_18_17_0  (
            .in0(N__73945),
            .in1(N__74548),
            .in2(N__78849),
            .in3(N__69547),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97420),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i50_51_LC_18_17_1 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i50_51_LC_18_17_1 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i50_51_LC_18_17_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i50_51_LC_18_17_1  (
            .in0(N__74549),
            .in1(N__73946),
            .in2(N__69486),
            .in3(N__69773),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97420),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i239_240_LC_18_17_2 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i239_240_LC_18_17_2 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i239_240_LC_18_17_2 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i239_240_LC_18_17_2  (
            .in0(N__73839),
            .in1(N__74545),
            .in2(N__73970),
            .in3(N__74015),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97420),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i251_252_LC_18_17_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i251_252_LC_18_17_3 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i251_252_LC_18_17_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i251_252_LC_18_17_3  (
            .in0(N__74547),
            .in1(N__73944),
            .in2(N__79044),
            .in3(N__69469),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97420),
            .ce(),
            .sr(_gnd_net_));
    defparam tx_addr_byte_r_i0_i4_LC_18_17_4.C_ON=1'b0;
    defparam tx_addr_byte_r_i0_i4_LC_18_17_4.SEQ_MODE=4'b1000;
    defparam tx_addr_byte_r_i0_i4_LC_18_17_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 tx_addr_byte_r_i0_i4_LC_18_17_4 (
            .in0(N__69448),
            .in1(N__69412),
            .in2(_gnd_net_),
            .in3(N__69312),
            .lcout(tx_addr_byte_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97420),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i149_150_LC_18_17_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i149_150_LC_18_17_5 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i149_150_LC_18_17_5 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i149_150_LC_18_17_5  (
            .in0(N__74544),
            .in1(N__69585),
            .in2(N__69269),
            .in3(N__69297),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97420),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i53_54_LC_18_17_6 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i53_54_LC_18_17_6 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i53_54_LC_18_17_6 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i53_54_LC_18_17_6  (
            .in0(N__69282),
            .in1(N__74550),
            .in2(N__73971),
            .in3(N__69265),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97420),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i245_246_LC_18_17_7 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i245_246_LC_18_17_7 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i245_246_LC_18_17_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i245_246_LC_18_17_7  (
            .in0(N__74546),
            .in1(N__73943),
            .in2(N__69270),
            .in3(N__69663),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97420),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i338_339_LC_18_18_0 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i338_339_LC_18_18_0 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i338_339_LC_18_18_0 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i338_339_LC_18_18_0  (
            .in0(N__69774),
            .in1(N__74506),
            .in2(N__69612),
            .in3(N__69648),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97428),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i3_2_lut_3_lut_LC_18_18_1 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i3_2_lut_3_lut_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i3_2_lut_3_lut_LC_18_18_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i3_2_lut_3_lut_LC_18_18_1  (
            .in0(N__74259),
            .in1(N__69705),
            .in2(_gnd_net_),
            .in3(N__74378),
            .lcout(\tx_fifo.lscc_fifo_inst.n3_adj_1136 ),
            .ltout(\tx_fifo.lscc_fifo_inst.n3_adj_1136_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i134_135_LC_18_18_2 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i134_135_LC_18_18_2 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i134_135_LC_18_18_2 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i134_135_LC_18_18_2  (
            .in0(N__78810),
            .in1(N__74503),
            .in2(N__69637),
            .in3(N__69544),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97428),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i4_2_lut_3_lut_LC_18_18_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i4_2_lut_3_lut_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i4_2_lut_3_lut_LC_18_18_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i4_2_lut_3_lut_LC_18_18_3  (
            .in0(N__74260),
            .in1(N__69706),
            .in2(_gnd_net_),
            .in3(N__74379),
            .lcout(\tx_fifo.lscc_fifo_inst.n4 ),
            .ltout(\tx_fifo.lscc_fifo_inst.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i230_231_LC_18_18_4 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i230_231_LC_18_18_4 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i230_231_LC_18_18_4 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i230_231_LC_18_18_4  (
            .in0(N__69630),
            .in1(N__74504),
            .in2(N__69634),
            .in3(N__69545),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97428),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11759_LC_18_18_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11759_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11759_LC_18_18_5 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11759_LC_18_18_5  (
            .in0(N__78794),
            .in1(N__69523),
            .in2(N__79008),
            .in3(N__69631),
            .lcout(\tx_fifo.lscc_fifo_inst.n13496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i326_327_LC_18_18_6 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i326_327_LC_18_18_6 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i326_327_LC_18_18_6 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i326_327_LC_18_18_6  (
            .in0(N__69522),
            .in1(N__74505),
            .in2(N__69611),
            .in3(N__69546),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97428),
            .ce(),
            .sr(_gnd_net_));
    defparam i9776_4_lut_LC_18_19_0.C_ON=1'b0;
    defparam i9776_4_lut_LC_18_19_0.SEQ_MODE=4'b0000;
    defparam i9776_4_lut_LC_18_19_0.LUT_INIT=16'b1111101111111110;
    LogicCell40 i9776_4_lut_LC_18_19_0 (
            .in0(N__74321),
            .in1(N__74431),
            .in2(N__69919),
            .in3(N__78795),
            .lcout(),
            .ltout(n11424_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_LC_18_19_1.C_ON=1'b0;
    defparam i1_4_lut_4_lut_LC_18_19_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_LC_18_19_1.LUT_INIT=16'b0000111100000000;
    LogicCell40 i1_4_lut_4_lut_LC_18_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__69514),
            .in3(N__69703),
            .lcout(),
            .ltout(n15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.full_r_84_LC_18_19_2 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.full_r_84_LC_18_19_2 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.full_r_84_LC_18_19_2 .LUT_INIT=16'b0011001000110000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.full_r_84_LC_18_19_2  (
            .in0(N__69781),
            .in1(N__78414),
            .in2(N__69784),
            .in3(N__69898),
            .lcout(is_tx_fifo_full_flag),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97434),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_r_1__I_0_i1_2_lut_LC_18_19_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_r_1__I_0_i1_2_lut_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_r_1__I_0_i1_2_lut_LC_18_19_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.wr_addr_r_1__I_0_i1_2_lut_LC_18_19_3  (
            .in0(N__78961),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74258),
            .lcout(n1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1138_2_lut_3_lut_LC_18_19_4.C_ON=1'b0;
    defparam i1138_2_lut_3_lut_LC_18_19_4.SEQ_MODE=4'b0000;
    defparam i1138_2_lut_3_lut_LC_18_19_4.LUT_INIT=16'b1101110111001100;
    LogicCell40 i1138_2_lut_3_lut_LC_18_19_4 (
            .in0(N__69702),
            .in1(N__78413),
            .in2(_gnd_net_),
            .in3(N__74376),
            .lcout(n2207),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.wr_en_i_I_0_2_lut_LC_18_19_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.wr_en_i_I_0_2_lut_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.wr_en_i_I_0_2_lut_LC_18_19_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.wr_en_i_I_0_2_lut_LC_18_19_5  (
            .in0(N__74377),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69704),
            .lcout(full_nxt_r),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i242_243_LC_18_19_6 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i242_243_LC_18_19_6 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i242_243_LC_18_19_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i242_243_LC_18_19_6  (
            .in0(N__69775),
            .in1(N__74432),
            .in2(N__69735),
            .in3(N__73950),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97434),
            .ce(),
            .sr(_gnd_net_));
    defparam fifo_write_cmd_79_LC_18_19_7.C_ON=1'b0;
    defparam fifo_write_cmd_79_LC_18_19_7.SEQ_MODE=4'b1000;
    defparam fifo_write_cmd_79_LC_18_19_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 fifo_write_cmd_79_LC_18_19_7 (
            .in0(_gnd_net_),
            .in1(N__69718),
            .in2(_gnd_net_),
            .in3(N__69701),
            .lcout(fifo_write_cmd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97434),
            .ce(),
            .sr(_gnd_net_));
    defparam i9762_4_lut_LC_18_20_0.C_ON=1'b0;
    defparam i9762_4_lut_LC_18_20_0.SEQ_MODE=4'b0000;
    defparam i9762_4_lut_LC_18_20_0.LUT_INIT=16'b0111101111011110;
    LogicCell40 i9762_4_lut_LC_18_20_0 (
            .in0(N__69891),
            .in1(N__74428),
            .in2(N__69676),
            .in3(N__69682),
            .lcout(n11410),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i1326_2_lut_LC_18_20_1 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i1326_2_lut_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.i1326_2_lut_LC_18_20_1 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i1326_2_lut_LC_18_20_1  (
            .in0(N__78962),
            .in1(N__78796),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rd_addr_p1_w_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i1333_3_lut_LC_18_20_2 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i1333_3_lut_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.i1333_3_lut_LC_18_20_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i1333_3_lut_LC_18_20_2  (
            .in0(N__78797),
            .in1(N__69872),
            .in2(_gnd_net_),
            .in3(N__78963),
            .lcout(rd_addr_p1_w_2),
            .ltout(rd_addr_p1_w_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r__i2_LC_18_20_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r__i2_LC_18_20_3 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r__i2_LC_18_20_3 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_addr_r__i2_LC_18_20_3  (
            .in0(N__69873),
            .in1(N__74335),
            .in2(N__69964),
            .in3(N__69951),
            .lcout(rd_addr_r_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97440),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i1304_2_lut_LC_18_20_4 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i1304_2_lut_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.i1304_2_lut_LC_18_20_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i1304_2_lut_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__74261),
            .in2(_gnd_net_),
            .in3(N__74429),
            .lcout(),
            .ltout(\tx_fifo.lscc_fifo_inst.wr_addr_p1_w_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i2_4_lut_LC_18_20_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i2_4_lut_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.i2_4_lut_LC_18_20_5 .LUT_INIT=16'b1000001000000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i2_4_lut_LC_18_20_5  (
            .in0(N__69862),
            .in1(N__78798),
            .in2(N__69922),
            .in3(N__69918),
            .lcout(n10727),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_p1_w_2__I_0_i3_2_lut_4_lut_LC_18_20_6 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_p1_w_2__I_0_i3_2_lut_4_lut_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_p1_w_2__I_0_i3_2_lut_4_lut_LC_18_20_6 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.wr_addr_p1_w_2__I_0_i3_2_lut_4_lut_LC_18_20_6  (
            .in0(N__69892),
            .in1(N__74430),
            .in2(N__74268),
            .in3(N__69874),
            .lcout(\tx_fifo.lscc_fifo_inst.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11814_LC_19_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11814_LC_19_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11814_LC_19_4_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11814_LC_19_4_0  (
            .in0(N__92445),
            .in1(N__77656),
            .in2(N__70438),
            .in3(N__88843),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13598_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13598_bdd_4_lut_LC_19_4_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13598_bdd_4_lut_LC_19_4_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13598_bdd_4_lut_LC_19_4_1 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13598_bdd_4_lut_LC_19_4_1  (
            .in0(N__70456),
            .in1(N__92443),
            .in2(N__69856),
            .in3(N__69853),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11844_LC_19_4_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11844_LC_19_4_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11844_LC_19_4_2 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11844_LC_19_4_2  (
            .in0(N__92446),
            .in1(N__88844),
            .in2(N__70426),
            .in3(N__69829),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13634_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13634_bdd_4_lut_LC_19_4_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13634_bdd_4_lut_LC_19_4_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13634_bdd_4_lut_LC_19_4_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13634_bdd_4_lut_LC_19_4_3  (
            .in0(N__69811),
            .in1(N__92444),
            .in2(N__69796),
            .in3(N__96415),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13637_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12413_LC_19_4_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12413_LC_19_4_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12413_LC_19_4_4 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_12413_LC_19_4_4  (
            .in0(N__90348),
            .in1(N__85818),
            .in2(N__69793),
            .in3(N__69790),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13946 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3032_3033_LC_19_4_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3032_3033_LC_19_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3032_3033_LC_19_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3032_3033_LC_19_4_5  (
            .in0(N__96342),
            .in1(N__70434),
            .in2(_gnd_net_),
            .in3(N__72567),
            .lcout(REG_mem_31_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93448),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2552_2553_LC_19_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2552_2553_LC_19_4_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2552_2553_LC_19_4_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2552_2553_LC_19_4_6  (
            .in0(N__70422),
            .in1(N__96343),
            .in2(_gnd_net_),
            .in3(N__70336),
            .lcout(REG_mem_26_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93448),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3026_3027_LC_19_4_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3026_3027_LC_19_4_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3026_3027_LC_19_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3026_3027_LC_19_4_7  (
            .in0(N__70404),
            .in1(N__76588),
            .in2(_gnd_net_),
            .in3(N__72566),
            .lcout(REG_mem_31_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93448),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12183_LC_19_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12183_LC_19_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12183_LC_19_5_0 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12183_LC_19_5_0  (
            .in0(N__74784),
            .in1(N__92519),
            .in2(N__70198),
            .in3(N__88842),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14042 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2558_2559_LC_19_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2558_2559_LC_19_5_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2558_2559_LC_19_5_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2558_2559_LC_19_5_1  (
            .in0(N__70194),
            .in1(N__89389),
            .in2(_gnd_net_),
            .in3(N__70393),
            .lcout(REG_mem_26_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93439),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13778_bdd_4_lut_LC_19_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13778_bdd_4_lut_LC_19_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13778_bdd_4_lut_LC_19_5_2 .LUT_INIT=16'b1011101010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13778_bdd_4_lut_LC_19_5_2  (
            .in0(N__70183),
            .in1(N__92518),
            .in2(N__70177),
            .in3(N__70153),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1304_1305_LC_19_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1304_1305_LC_19_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1304_1305_LC_19_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1304_1305_LC_19_5_3  (
            .in0(N__74826),
            .in1(N__96352),
            .in2(_gnd_net_),
            .in3(N__70140),
            .lcout(REG_mem_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93439),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1961_1962_LC_19_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1961_1962_LC_19_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1961_1962_LC_19_5_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1961_1962_LC_19_5_4  (
            .in0(N__96728),
            .in1(N__95465),
            .in2(N__71047),
            .in3(N__77473),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93439),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2630_2631_LC_19_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2630_2631_LC_19_5_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2630_2631_LC_19_5_5 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2630_2631_LC_19_5_5  (
            .in0(N__71598),
            .in1(N__95464),
            .in2(N__69981),
            .in3(N__79755),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93439),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5702_5703_LC_19_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5702_5703_LC_19_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5702_5703_LC_19_5_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5702_5703_LC_19_5_6  (
            .in0(N__79754),
            .in1(N__71599),
            .in2(N__71092),
            .in3(N__95466),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93439),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10359_3_lut_LC_19_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10359_3_lut_LC_19_5_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10359_3_lut_LC_19_5_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10359_3_lut_LC_19_5_7  (
            .in0(N__88841),
            .in1(N__71091),
            .in2(_gnd_net_),
            .in3(N__71173),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12008 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10031_3_lut_LC_19_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10031_3_lut_LC_19_6_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10031_3_lut_LC_19_6_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10031_3_lut_LC_19_6_0  (
            .in0(N__71061),
            .in1(N__88837),
            .in2(_gnd_net_),
            .in3(N__71046),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12398_LC_19_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12398_LC_19_6_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12398_LC_19_6_1 .LUT_INIT=16'b1100101011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12398_LC_19_6_1  (
            .in0(N__70740),
            .in1(N__71023),
            .in2(N__88886),
            .in3(N__92517),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14294_bdd_4_lut_LC_19_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14294_bdd_4_lut_LC_19_6_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14294_bdd_4_lut_LC_19_6_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14294_bdd_4_lut_LC_19_6_2  (
            .in0(N__70752),
            .in1(N__92108),
            .in2(N__71011),
            .in3(N__70764),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5912_5913_LC_19_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5912_5913_LC_19_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5912_5913_LC_19_6_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5912_5913_LC_19_6_3  (
            .in0(N__96225),
            .in1(N__94666),
            .in2(N__70765),
            .in3(N__71006),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_61_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93434),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5816_5817_LC_19_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5816_5817_LC_19_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5816_5817_LC_19_6_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5816_5817_LC_19_6_4  (
            .in0(N__94665),
            .in1(N__70682),
            .in2(N__70753),
            .in3(N__96228),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_60_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93434),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6008_6009_LC_19_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6008_6009_LC_19_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6008_6009_LC_19_6_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6008_6009_LC_19_6_5  (
            .in0(N__96226),
            .in1(N__94667),
            .in2(N__70741),
            .in3(N__77969),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93434),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2744_2745_LC_19_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2744_2745_LC_19_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2744_2745_LC_19_6_6 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2744_2745_LC_19_6_6  (
            .in0(N__94664),
            .in1(N__70681),
            .in2(N__70455),
            .in3(N__96227),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_28_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93434),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2249_2250_LC_19_6_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2249_2250_LC_19_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2249_2250_LC_19_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2249_2250_LC_19_6_7  (
            .in0(N__71613),
            .in1(N__96727),
            .in2(_gnd_net_),
            .in3(N__75066),
            .lcout(REG_mem_23_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93434),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4856_4857_LC_19_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4856_4857_LC_19_7_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4856_4857_LC_19_7_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4856_4857_LC_19_7_2  (
            .in0(N__96209),
            .in1(N__75189),
            .in2(_gnd_net_),
            .in3(N__73051),
            .lcout(REG_mem_50_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93428),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5606_5607_LC_19_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5606_5607_LC_19_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5606_5607_LC_19_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5606_5607_LC_19_7_3  (
            .in0(N__71169),
            .in1(N__71597),
            .in2(_gnd_net_),
            .in3(N__79990),
            .lcout(REG_mem_58_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93428),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4286_4287_LC_19_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4286_4287_LC_19_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4286_4287_LC_19_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4286_4287_LC_19_7_5  (
            .in0(N__89715),
            .in1(N__89462),
            .in2(_gnd_net_),
            .in3(N__71741),
            .lcout(REG_mem_44_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93428),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i254_255_LC_19_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i254_255_LC_19_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i254_255_LC_19_7_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i254_255_LC_19_7_6  (
            .in0(N__89461),
            .in1(N__95155),
            .in2(N__83121),
            .in3(N__80604),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93428),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10139_3_lut_LC_19_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10139_3_lut_LC_19_7_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10139_3_lut_LC_19_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10139_3_lut_LC_19_7_7  (
            .in0(N__72583),
            .in1(N__88836),
            .in2(_gnd_net_),
            .in3(N__71158),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11788 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12458_LC_19_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12458_LC_19_8_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12458_LC_19_8_0 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12458_LC_19_8_0  (
            .in0(N__92272),
            .in1(N__71146),
            .in2(N__71125),
            .in3(N__88744),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5624_5625_LC_19_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5624_5625_LC_19_8_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5624_5625_LC_19_8_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5624_5625_LC_19_8_1  (
            .in0(_gnd_net_),
            .in1(N__71121),
            .in2(N__96341),
            .in3(N__79974),
            .lcout(REG_mem_58_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93422),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2444_2445_LC_19_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2444_2445_LC_19_8_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2444_2445_LC_19_8_2 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2444_2445_LC_19_8_2  (
            .in0(N__95152),
            .in1(N__75933),
            .in2(N__71109),
            .in3(N__97024),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93422),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10209_3_lut_LC_19_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10209_3_lut_LC_19_8_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10209_3_lut_LC_19_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10209_3_lut_LC_19_8_3  (
            .in0(N__88743),
            .in1(N__72307),
            .in2(_gnd_net_),
            .in3(N__72289),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11858 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2072_2073_LC_19_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2072_2073_LC_19_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2072_2073_LC_19_8_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2072_2073_LC_19_8_4  (
            .in0(N__95151),
            .in1(N__96269),
            .in2(N__75334),
            .in3(N__77015),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93422),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4952_4953_LC_19_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4952_4953_LC_19_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4952_4953_LC_19_8_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4952_4953_LC_19_8_5  (
            .in0(N__75201),
            .in1(_gnd_net_),
            .in2(N__96340),
            .in3(N__72233),
            .lcout(REG_mem_51_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93422),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5516_5517_LC_19_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5516_5517_LC_19_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5516_5517_LC_19_8_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5516_5517_LC_19_8_6  (
            .in0(N__95153),
            .in1(N__75934),
            .in2(N__75250),
            .in3(N__97025),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93422),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2462_2463_LC_19_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2462_2463_LC_19_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2462_2463_LC_19_8_7 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2462_2463_LC_19_8_7  (
            .in0(N__97023),
            .in1(N__89472),
            .in2(N__79473),
            .in3(N__95154),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93422),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1886_1887_LC_19_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1886_1887_LC_19_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1886_1887_LC_19_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1886_1887_LC_19_9_0  (
            .in0(N__89459),
            .in1(N__71937),
            .in2(_gnd_net_),
            .in3(N__72111),
            .lcout(REG_mem_19_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11640_LC_19_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11640_LC_19_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11640_LC_19_9_1 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11640_LC_19_9_1  (
            .in0(N__72739),
            .in1(N__92268),
            .in2(N__88772),
            .in3(N__71926),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4376_4377_LC_19_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4376_4377_LC_19_9_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4376_4377_LC_19_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4376_4377_LC_19_9_2  (
            .in0(N__96190),
            .in1(N__75387),
            .in2(_gnd_net_),
            .in3(N__71902),
            .lcout(REG_mem_45_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4280_4281_LC_19_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4280_4281_LC_19_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4280_4281_LC_19_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4280_4281_LC_19_9_3  (
            .in0(N__75408),
            .in1(N__96193),
            .in2(_gnd_net_),
            .in3(N__71736),
            .lcout(REG_mem_44_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4472_4473_LC_19_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4472_4473_LC_19_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4472_4473_LC_19_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4472_4473_LC_19_9_4  (
            .in0(N__96192),
            .in1(N__72738),
            .in2(_gnd_net_),
            .in3(N__89114),
            .lcout(REG_mem_46_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1982_1983_LC_19_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1982_1983_LC_19_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1982_1983_LC_19_9_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1982_1983_LC_19_9_5  (
            .in0(N__95156),
            .in1(N__89460),
            .in2(N__72334),
            .in3(N__77419),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i440_441_LC_19_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i440_441_LC_19_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i440_441_LC_19_9_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i440_441_LC_19_9_6  (
            .in0(N__96191),
            .in1(N__72711),
            .in2(_gnd_net_),
            .in3(N__72579),
            .lcout(REG_mem_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93415),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2942_2943_LC_19_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2942_2943_LC_19_10_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2942_2943_LC_19_10_0 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2942_2943_LC_19_10_0  (
            .in0(N__94603),
            .in1(N__72381),
            .in2(N__89516),
            .in3(N__77955),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3038_3039_LC_19_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3038_3039_LC_19_10_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3038_3039_LC_19_10_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3038_3039_LC_19_10_1  (
            .in0(N__72393),
            .in1(N__89463),
            .in2(_gnd_net_),
            .in3(N__72516),
            .lcout(REG_mem_31_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12158_LC_19_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12158_LC_19_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12158_LC_19_10_2 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12158_LC_19_10_2  (
            .in0(N__88590),
            .in1(N__91734),
            .in2(N__72397),
            .in3(N__72382),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12198_LC_19_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12198_LC_19_10_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12198_LC_19_10_3 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12198_LC_19_10_3  (
            .in0(N__91735),
            .in1(N__88591),
            .in2(N__72373),
            .in3(N__72352),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14060_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14060_bdd_4_lut_LC_19_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14060_bdd_4_lut_LC_19_10_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14060_bdd_4_lut_LC_19_10_4 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14060_bdd_4_lut_LC_19_10_4  (
            .in0(N__72333),
            .in1(N__91733),
            .in2(N__72319),
            .in3(N__72316),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11709 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2078_2079_LC_19_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2078_2079_LC_19_10_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2078_2079_LC_19_10_5 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2078_2079_LC_19_10_5  (
            .in0(N__72315),
            .in1(N__94604),
            .in2(N__89514),
            .in3(N__77020),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_21_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5330_5331_LC_19_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5330_5331_LC_19_10_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5330_5331_LC_19_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5330_5331_LC_19_10_6  (
            .in0(N__75376),
            .in1(N__76759),
            .in2(_gnd_net_),
            .in3(N__77244),
            .lcout(REG_mem_55_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4862_4863_LC_19_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4862_4863_LC_19_10_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4862_4863_LC_19_10_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4862_4863_LC_19_10_7  (
            .in0(N__72888),
            .in1(N__89464),
            .in2(_gnd_net_),
            .in3(N__73013),
            .lcout(REG_mem_50_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93393),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10533_3_lut_LC_19_11_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10533_3_lut_LC_19_11_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10533_3_lut_LC_19_11_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10533_3_lut_LC_19_11_1  (
            .in0(N__72877),
            .in1(N__85634),
            .in2(_gnd_net_),
            .in3(N__72862),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12182_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10534_3_lut_LC_19_11_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10534_3_lut_LC_19_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10534_3_lut_LC_19_11_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10534_3_lut_LC_19_11_2  (
            .in0(N__90211),
            .in1(_gnd_net_),
            .in2(N__72850),
            .in3(N__72847),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10513_3_lut_LC_19_11_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10513_3_lut_LC_19_11_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10513_3_lut_LC_19_11_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10513_3_lut_LC_19_11_3  (
            .in0(N__72838),
            .in1(N__90210),
            .in2(_gnd_net_),
            .in3(N__72829),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11829_LC_19_11_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11829_LC_19_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11829_LC_19_11_4 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11829_LC_19_11_4  (
            .in0(N__85635),
            .in1(N__72817),
            .in2(N__90290),
            .in3(N__72802),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13610_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13610_bdd_4_lut_LC_19_11_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13610_bdd_4_lut_LC_19_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13610_bdd_4_lut_LC_19_11_5 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13610_bdd_4_lut_LC_19_11_5  (
            .in0(N__72790),
            .in1(N__90212),
            .in2(N__72772),
            .in3(N__75358),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12246_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12188_LC_19_11_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12188_LC_19_11_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12188_LC_19_11_6 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_12188_LC_19_11_6  (
            .in0(N__81087),
            .in1(N__72769),
            .in2(N__72757),
            .in3(N__81273),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13442_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i5_LC_19_11_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i5_LC_19_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i5_LC_19_11_7 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i5_LC_19_11_7  (
            .in0(N__72754),
            .in1(N__81086),
            .in2(N__72748),
            .in3(N__72745),
            .lcout(REG_out_raw_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97370),
            .ce(N__80862),
            .sr(_gnd_net_));
    defparam i914_4_lut_4_lut_LC_19_12_0.C_ON=1'b0;
    defparam i914_4_lut_4_lut_LC_19_12_0.SEQ_MODE=4'b0000;
    defparam i914_4_lut_4_lut_LC_19_12_0.LUT_INIT=16'b0000100100000010;
    LogicCell40 i914_4_lut_4_lut_LC_19_12_0 (
            .in0(N__82175),
            .in1(N__81882),
            .in2(N__81754),
            .in3(N__83998),
            .lcout(n1876),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i1_2_lut_4_lut_adj_90_LC_19_12_1 .C_ON=1'b0;
    defparam \timing_controller_inst.i1_2_lut_4_lut_adj_90_LC_19_12_1 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i1_2_lut_4_lut_adj_90_LC_19_12_1 .LUT_INIT=16'b1111111100000001;
    LogicCell40 \timing_controller_inst.i1_2_lut_4_lut_adj_90_LC_19_12_1  (
            .in0(N__81884),
            .in1(N__82176),
            .in2(N__84017),
            .in3(N__73081),
            .lcout(\timing_controller_inst.n4200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i1_2_lut_3_lut_LC_19_12_2 .C_ON=1'b0;
    defparam \timing_controller_inst.i1_2_lut_3_lut_LC_19_12_2 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i1_2_lut_3_lut_LC_19_12_2 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \timing_controller_inst.i1_2_lut_3_lut_LC_19_12_2  (
            .in0(N__84004),
            .in1(_gnd_net_),
            .in2(N__81755),
            .in3(N__81883),
            .lcout(),
            .ltout(\timing_controller_inst.n11375_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_i1_LC_19_12_3 .C_ON=1'b0;
    defparam \timing_controller_inst.state_i1_LC_19_12_3 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_i1_LC_19_12_3 .LUT_INIT=16'b1101110100101110;
    LogicCell40 \timing_controller_inst.state_i1_LC_19_12_3  (
            .in0(N__84002),
            .in1(N__84074),
            .in2(N__73093),
            .in3(N__82177),
            .lcout(state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97385),
            .ce(N__73090),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_i2_LC_19_12_4 .C_ON=1'b0;
    defparam \timing_controller_inst.state_i2_LC_19_12_4 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_i2_LC_19_12_4 .LUT_INIT=16'b1001100011011100;
    LogicCell40 \timing_controller_inst.state_i2_LC_19_12_4  (
            .in0(N__84075),
            .in1(N__81886),
            .in2(N__82237),
            .in3(N__84003),
            .lcout(state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97385),
            .ce(N__73090),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i1_2_lut_adj_88_LC_19_12_5 .C_ON=1'b0;
    defparam \timing_controller_inst.i1_2_lut_adj_88_LC_19_12_5 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i1_2_lut_adj_88_LC_19_12_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \timing_controller_inst.i1_2_lut_adj_88_LC_19_12_5  (
            .in0(_gnd_net_),
            .in1(N__81738),
            .in2(_gnd_net_),
            .in3(N__84072),
            .lcout(n11376),
            .ltout(n11376_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11042_3_lut_4_lut_LC_19_12_6.C_ON=1'b0;
    defparam i11042_3_lut_4_lut_LC_19_12_6.SEQ_MODE=4'b0000;
    defparam i11042_3_lut_4_lut_LC_19_12_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 i11042_3_lut_4_lut_LC_19_12_6 (
            .in0(N__82174),
            .in1(N__81881),
            .in2(N__73075),
            .in3(N__83997),
            .lcout(n12601),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i2_3_lut_4_lut_LC_19_12_7 .C_ON=1'b0;
    defparam \timing_controller_inst.i2_3_lut_4_lut_LC_19_12_7 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i2_3_lut_4_lut_LC_19_12_7 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \timing_controller_inst.i2_3_lut_4_lut_LC_19_12_7  (
            .in0(N__81885),
            .in1(N__84073),
            .in2(N__82238),
            .in3(N__81739),
            .lcout(\timing_controller_inst.n11377 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_321_Mux_4_i15_4_lut_4_lut_LC_19_13_0 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_321_Mux_4_i15_4_lut_4_lut_LC_19_13_0 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_321_Mux_4_i15_4_lut_4_lut_LC_19_13_0 .LUT_INIT=16'b0100000001000010;
    LogicCell40 \timing_controller_inst.mux_321_Mux_4_i15_4_lut_4_lut_LC_19_13_0  (
            .in0(N__84089),
            .in1(N__82194),
            .in2(N__81908),
            .in3(N__84026),
            .lcout(\timing_controller_inst.invert_N_309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \usb3_if_inst.reset_per_frame_latched_82_LC_19_13_1 .C_ON=1'b0;
    defparam \usb3_if_inst.reset_per_frame_latched_82_LC_19_13_1 .SEQ_MODE=4'b1000;
    defparam \usb3_if_inst.reset_per_frame_latched_82_LC_19_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \usb3_if_inst.reset_per_frame_latched_82_LC_19_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73567),
            .lcout(\usb3_if_inst.reset_per_frame_latched ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97392),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.invert_55_i1_LC_19_13_2 .C_ON=1'b0;
    defparam \timing_controller_inst.invert_55_i1_LC_19_13_2 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.invert_55_i1_LC_19_13_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \timing_controller_inst.invert_55_i1_LC_19_13_2  (
            .in0(N__84087),
            .in1(N__82192),
            .in2(N__77998),
            .in3(N__84022),
            .lcout(reset_per_frame),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97392),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.invert_55_i2_LC_19_13_3 .C_ON=1'b0;
    defparam \timing_controller_inst.invert_55_i2_LC_19_13_3 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.invert_55_i2_LC_19_13_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \timing_controller_inst.invert_55_i2_LC_19_13_3  (
            .in0(N__82193),
            .in1(N__84088),
            .in2(N__84028),
            .in3(N__81892),
            .lcout(buffer_switch_done),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97392),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i13_3_lut_LC_19_13_4 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i13_3_lut_LC_19_13_4 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i13_3_lut_LC_19_13_4 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \timing_controller_inst.mux_855_i13_3_lut_LC_19_13_4  (
            .in0(N__82397),
            .in1(N__84526),
            .in2(_gnd_net_),
            .in3(N__82195),
            .lcout(\timing_controller_inst.n1742 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.invert_55_i0_LC_19_13_5 .C_ON=1'b0;
    defparam \timing_controller_inst.invert_55_i0_LC_19_13_5 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.invert_55_i0_LC_19_13_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \timing_controller_inst.invert_55_i0_LC_19_13_5  (
            .in0(N__82191),
            .in1(N__84086),
            .in2(N__84027),
            .in3(N__81891),
            .lcout(reset_all),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97392),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i6388_3_lut_LC_19_13_6 .C_ON=1'b0;
    defparam \timing_controller_inst.i6388_3_lut_LC_19_13_6 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i6388_3_lut_LC_19_13_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \timing_controller_inst.i6388_3_lut_LC_19_13_6  (
            .in0(N__81890),
            .in1(N__82190),
            .in2(_gnd_net_),
            .in3(N__84018),
            .lcout(n7566),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i19_3_lut_LC_19_13_7 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i19_3_lut_LC_19_13_7 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i19_3_lut_LC_19_13_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \timing_controller_inst.mux_855_i19_3_lut_LC_19_13_7  (
            .in0(N__82196),
            .in1(N__84355),
            .in2(_gnd_net_),
            .in3(N__82398),
            .lcout(\timing_controller_inst.n1736 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i30_4_lut_LC_19_14_0 .C_ON=1'b0;
    defparam \timing_controller_inst.i30_4_lut_LC_19_14_0 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i30_4_lut_LC_19_14_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \timing_controller_inst.i30_4_lut_LC_19_14_0  (
            .in0(N__78259),
            .in1(N__78253),
            .in2(N__78247),
            .in3(N__81820),
            .lcout(\timing_controller_inst.n62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Tx_Data_i6_LC_19_14_1 .C_ON=1'b0;
    defparam \pc_tx.r_Tx_Data_i6_LC_19_14_1 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Tx_Data_i6_LC_19_14_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pc_tx.r_Tx_Data_i6_LC_19_14_1  (
            .in0(N__81677),
            .in1(N__78153),
            .in2(_gnd_net_),
            .in3(N__73785),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97401),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Bit_Index_i0_LC_19_14_2 .C_ON=1'b0;
    defparam \pc_tx.r_Bit_Index_i0_LC_19_14_2 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Bit_Index_i0_LC_19_14_2 .LUT_INIT=16'b0011000000111000;
    LogicCell40 \pc_tx.r_Bit_Index_i0_LC_19_14_2  (
            .in0(N__83617),
            .in1(N__82693),
            .in2(N__83428),
            .in3(N__83404),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97401),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i4_LC_19_14_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i4_LC_19_14_3 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i4_LC_19_14_3 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i4_LC_19_14_3  (
            .in0(N__73828),
            .in1(N__78447),
            .in2(N__78331),
            .in3(N__73822),
            .lcout(fifo_temp_output_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97401),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Tx_Data_i4_LC_19_14_4 .C_ON=1'b0;
    defparam \pc_tx.r_Tx_Data_i4_LC_19_14_4 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Tx_Data_i4_LC_19_14_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \pc_tx.r_Tx_Data_i4_LC_19_14_4  (
            .in0(N__73821),
            .in1(N__77523),
            .in2(_gnd_net_),
            .in3(N__81675),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97401),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i5_LC_19_14_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i5_LC_19_14_5 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i5_LC_19_14_5 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i5_LC_19_14_5  (
            .in0(N__73813),
            .in1(N__78448),
            .in2(N__78332),
            .in3(N__73807),
            .lcout(fifo_temp_output_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97401),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Tx_Data_i5_LC_19_14_6 .C_ON=1'b0;
    defparam \pc_tx.r_Tx_Data_i5_LC_19_14_6 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Tx_Data_i5_LC_19_14_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \pc_tx.r_Tx_Data_i5_LC_19_14_6  (
            .in0(N__73806),
            .in1(N__77538),
            .in2(_gnd_net_),
            .in3(N__81676),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97401),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i6_LC_19_14_7 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i6_LC_19_14_7 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i6_LC_19_14_7 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i6_LC_19_14_7  (
            .in0(N__73798),
            .in1(N__78449),
            .in2(N__78333),
            .in3(N__73786),
            .lcout(fifo_temp_output_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97401),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i7_LC_19_15_0 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i7_LC_19_15_0 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i7_LC_19_15_0 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i7_LC_19_15_0  (
            .in0(N__73777),
            .in1(N__78435),
            .in2(N__78318),
            .in3(N__73768),
            .lcout(fifo_temp_output_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97409),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Tx_Data_i7_LC_19_15_1 .C_ON=1'b0;
    defparam \pc_tx.r_Tx_Data_i7_LC_19_15_1 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Tx_Data_i7_LC_19_15_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pc_tx.r_Tx_Data_i7_LC_19_15_1  (
            .in0(N__81679),
            .in1(N__73767),
            .in2(_gnd_net_),
            .in3(N__78168),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97409),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Tx_Data_i3_LC_19_15_3 .C_ON=1'b0;
    defparam \pc_tx.r_Tx_Data_i3_LC_19_15_3 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Tx_Data_i3_LC_19_15_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pc_tx.r_Tx_Data_i3_LC_19_15_3  (
            .in0(N__81678),
            .in1(N__77562),
            .in2(_gnd_net_),
            .in3(N__78271),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97409),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i17_4_lut_LC_19_15_4 .C_ON=1'b0;
    defparam \timing_controller_inst.i17_4_lut_LC_19_15_4 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i17_4_lut_LC_19_15_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \timing_controller_inst.i17_4_lut_LC_19_15_4  (
            .in0(N__86743),
            .in1(N__84372),
            .in2(N__83767),
            .in3(N__83848),
            .lcout(\timing_controller_inst.n49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i233_234_LC_19_15_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i233_234_LC_19_15_5 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i233_234_LC_19_15_5 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i233_234_LC_19_15_5  (
            .in0(N__73896),
            .in1(N__74556),
            .in2(N__73993),
            .in3(N__79122),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97409),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i44_45_LC_19_15_6 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i44_45_LC_19_15_6 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i44_45_LC_19_15_6 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i44_45_LC_19_15_6  (
            .in0(N__74557),
            .in1(N__73991),
            .in2(N__74212),
            .in3(N__74172),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97409),
            .ce(),
            .sr(_gnd_net_));
    defparam start_tx_81_LC_19_15_7.C_ON=1'b0;
    defparam start_tx_81_LC_19_15_7.SEQ_MODE=4'b1000;
    defparam start_tx_81_LC_19_15_7.LUT_INIT=16'b1111111000010000;
    LogicCell40 start_tx_81_LC_19_15_7 (
            .in0(N__80661),
            .in1(N__74899),
            .in2(N__81618),
            .in3(N__74329),
            .lcout(r_SM_Main_2_N_811_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97409),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi0.i6_4_lut_adj_30_LC_19_16_0 .C_ON=1'b0;
    defparam \spi0.i6_4_lut_adj_30_LC_19_16_0 .SEQ_MODE=4'b0000;
    defparam \spi0.i6_4_lut_adj_30_LC_19_16_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \spi0.i6_4_lut_adj_30_LC_19_16_0  (
            .in0(N__74161),
            .in1(N__74140),
            .in2(N__74116),
            .in3(N__74092),
            .lcout(\spi0.n14_adj_1140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i31_4_lut_LC_19_16_2 .C_ON=1'b0;
    defparam \timing_controller_inst.i31_4_lut_LC_19_16_2 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i31_4_lut_LC_19_16_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \timing_controller_inst.i31_4_lut_LC_19_16_2  (
            .in0(N__81931),
            .in1(N__74053),
            .in2(N__74044),
            .in3(N__81601),
            .lcout(n63),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i47_48_LC_19_16_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i47_48_LC_19_16_3 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i47_48_LC_19_16_3 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i47_48_LC_19_16_3  (
            .in0(N__74542),
            .in1(N__73976),
            .in2(N__74035),
            .in3(N__78873),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97421),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i41_42_LC_19_16_4 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i41_42_LC_19_16_4 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.i41_42_LC_19_16_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i41_42_LC_19_16_4  (
            .in0(N__73975),
            .in1(N__74541),
            .in2(N__73900),
            .in3(N__79086),
            .lcout(\tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97421),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11889_LC_19_16_6 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11889_LC_19_16_6 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11889_LC_19_16_6 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11889_LC_19_16_6  (
            .in0(N__78774),
            .in1(N__73855),
            .in2(N__73843),
            .in3(N__78988),
            .lcout(\tx_fifo.lscc_fifo_inst.n13556 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_en_i_I_0_2_lut_LC_19_17_0 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_en_i_I_0_2_lut_LC_19_17_0 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.rd_en_i_I_0_2_lut_LC_19_17_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_en_i_I_0_2_lut_LC_19_17_0  (
            .in0(_gnd_net_),
            .in1(N__74315),
            .in2(_gnd_net_),
            .in3(N__74898),
            .lcout(rd_fifo_en_w),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_19_18_1.C_ON=1'b0;
    defparam i1_4_lut_LC_19_18_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_19_18_1.LUT_INIT=16'b1000001001000001;
    LogicCell40 i1_4_lut_LC_19_18_1 (
            .in0(N__78960),
            .in1(N__74543),
            .in2(N__78799),
            .in3(N__74257),
            .lcout(),
            .ltout(n32_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_19_18_2.C_ON=1'b0;
    defparam i1_3_lut_LC_19_18_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_19_18_2.LUT_INIT=16'b0000000010100000;
    LogicCell40 i1_3_lut_LC_19_18_2 (
            .in0(N__74892),
            .in1(_gnd_net_),
            .in2(N__74383),
            .in3(N__74380),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r_86_LC_19_18_4 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r_86_LC_19_18_4 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r_86_LC_19_18_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r_86_LC_19_18_4  (
            .in0(N__74894),
            .in1(N__74311),
            .in2(_gnd_net_),
            .in3(N__78427),
            .lcout(\tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97435),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.i1_2_lut_3_lut_4_lut_LC_19_18_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i1_2_lut_3_lut_4_lut_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.i1_2_lut_3_lut_4_lut_LC_19_18_5 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i1_2_lut_3_lut_4_lut_LC_19_18_5  (
            .in0(N__78426),
            .in1(N__74356),
            .in2(N__74325),
            .in3(N__74893),
            .lcout(n4249),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam fifo_read_cmd_80_LC_19_18_7.C_ON=1'b0;
    defparam fifo_read_cmd_80_LC_19_18_7.SEQ_MODE=4'b1000;
    defparam fifo_read_cmd_80_LC_19_18_7.LUT_INIT=16'b0000000001010101;
    LogicCell40 fifo_read_cmd_80_LC_19_18_7 (
            .in0(N__80665),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74891),
            .lcout(fifo_read_cmd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97435),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r__i0_LC_19_19_0 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r__i0_LC_19_19_0 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r__i0_LC_19_19_0 .LUT_INIT=16'b0110011000110110;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_addr_r__i0_LC_19_19_0  (
            .in0(N__78425),
            .in1(N__78956),
            .in2(N__74326),
            .in3(N__74875),
            .lcout(rd_addr_r_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97441),
            .ce(),
            .sr(N__78424));
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_r__i0_LC_19_19_7 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_r__i0_LC_19_19_7 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.wr_addr_r__i0_LC_19_19_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.wr_addr_r__i0_LC_19_19_7  (
            .in0(N__74255),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74348),
            .lcout(wr_addr_r_0_adj_1181),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97441),
            .ce(),
            .sr(N__78424));
    defparam \tx_fifo.lscc_fifo_inst.i3110_2_lut_3_lut_LC_19_20_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.i3110_2_lut_3_lut_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.i3110_2_lut_3_lut_LC_19_20_3 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \tx_fifo.lscc_fifo_inst.i3110_2_lut_3_lut_LC_19_20_3  (
            .in0(N__74874),
            .in1(N__78389),
            .in2(_gnd_net_),
            .in3(N__74328),
            .lcout(empty_o_N_1116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_102_LC_19_20_6.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_102_LC_19_20_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_102_LC_19_20_6.LUT_INIT=16'b0000000000101000;
    LogicCell40 i1_2_lut_4_lut_adj_102_LC_19_20_6 (
            .in0(N__74327),
            .in1(N__74256),
            .in2(N__78984),
            .in3(N__74873),
            .lcout(),
            .ltout(n4_adj_1186_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.empty_r_85_LC_19_20_7 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.empty_r_85_LC_19_20_7 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.empty_r_85_LC_19_20_7 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \tx_fifo.lscc_fifo_inst.empty_r_85_LC_19_20_7  (
            .in0(N__74920),
            .in1(N__78388),
            .in2(N__74911),
            .in3(N__74908),
            .lcout(is_fifo_empty_flag),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97444),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13772_bdd_4_lut_LC_20_4_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13772_bdd_4_lut_LC_20_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13772_bdd_4_lut_LC_20_4_0 .LUT_INIT=16'b1010101011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13772_bdd_4_lut_LC_20_4_0  (
            .in0(N__74791),
            .in1(N__74848),
            .in2(N__74830),
            .in3(N__92447),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i56_57_LC_20_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i56_57_LC_20_5_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i56_57_LC_20_5_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i56_57_LC_20_5_0  (
            .in0(N__94222),
            .in1(N__96314),
            .in2(N__79206),
            .in3(N__82951),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93449),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11959_LC_20_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11959_LC_20_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11959_LC_20_5_1 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11959_LC_20_5_1  (
            .in0(N__88755),
            .in1(N__92635),
            .in2(N__74815),
            .in3(N__74623),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13772 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2654_2655_LC_20_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2654_2655_LC_20_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2654_2655_LC_20_5_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2654_2655_LC_20_5_3  (
            .in0(N__89388),
            .in1(N__94223),
            .in2(N__74785),
            .in3(N__79760),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_27_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93449),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1400_1401_LC_20_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1400_1401_LC_20_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1400_1401_LC_20_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1400_1401_LC_20_5_4  (
            .in0(N__74622),
            .in1(N__96313),
            .in2(_gnd_net_),
            .in3(N__74770),
            .lcout(REG_mem_14_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93449),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13004_bdd_4_lut_LC_20_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13004_bdd_4_lut_LC_20_5_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13004_bdd_4_lut_LC_20_5_5 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13004_bdd_4_lut_LC_20_5_5  (
            .in0(N__90353),
            .in1(N__75082),
            .in2(N__75097),
            .in3(N__75151),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13007 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11754_LC_20_5_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11754_LC_20_5_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11754_LC_20_5_6 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11754_LC_20_5_6  (
            .in0(N__92634),
            .in1(N__88754),
            .in2(N__74614),
            .in3(N__74596),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13520_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13520_bdd_4_lut_LC_20_5_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13520_bdd_4_lut_LC_20_5_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13520_bdd_4_lut_LC_20_5_7 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13520_bdd_4_lut_LC_20_5_7  (
            .in0(N__74575),
            .in1(N__92633),
            .in2(N__74560),
            .in3(N__75223),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11844 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11139_LC_20_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11139_LC_20_6_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11139_LC_20_6_0 .LUT_INIT=16'b1011110010110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11139_LC_20_6_0  (
            .in0(N__75205),
            .in1(N__92111),
            .in2(N__88852),
            .in3(N__75190),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12782_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12782_bdd_4_lut_LC_20_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12782_bdd_4_lut_LC_20_6_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12782_bdd_4_lut_LC_20_6_1 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12782_bdd_4_lut_LC_20_6_1  (
            .in0(N__75424),
            .in1(N__92109),
            .in2(N__75178),
            .in3(N__75175),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6002_6003_LC_20_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6002_6003_LC_20_6_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6002_6003_LC_20_6_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i6002_6003_LC_20_6_2  (
            .in0(N__76622),
            .in1(N__95150),
            .in2(N__75141),
            .in3(N__77974),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_62_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93440),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12473_LC_20_6_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12473_LC_20_6_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12473_LC_20_6_3 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12473_LC_20_6_3  (
            .in0(N__92112),
            .in1(N__88753),
            .in2(N__75124),
            .in3(N__75076),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14390_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14390_bdd_4_lut_LC_20_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14390_bdd_4_lut_LC_20_6_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14390_bdd_4_lut_LC_20_6_4 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14390_bdd_4_lut_LC_20_6_4  (
            .in0(N__75291),
            .in1(N__92110),
            .in2(N__75100),
            .in3(N__75276),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11340_LC_20_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11340_LC_20_6_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11340_LC_20_6_5 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11340_LC_20_6_5  (
            .in0(N__75088),
            .in1(N__76039),
            .in2(N__90400),
            .in3(N__85279),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13004 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5336_5337_LC_20_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5336_5337_LC_20_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5336_5337_LC_20_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5336_5337_LC_20_6_6  (
            .in0(N__75075),
            .in1(N__96251),
            .in2(_gnd_net_),
            .in3(N__77246),
            .lcout(REG_mem_55_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93440),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2264_2265_LC_20_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2264_2265_LC_20_7_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2264_2265_LC_20_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2264_2265_LC_20_7_0  (
            .in0(N__96243),
            .in1(N__75348),
            .in2(_gnd_net_),
            .in3(N__75067),
            .lcout(REG_mem_23_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93435),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11854_LC_20_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11854_LC_20_7_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11854_LC_20_7_1 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11854_LC_20_7_1  (
            .in0(N__75303),
            .in1(N__75349),
            .in2(N__92672),
            .in3(N__88857),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13646_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13646_bdd_4_lut_LC_20_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13646_bdd_4_lut_LC_20_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13646_bdd_4_lut_LC_20_7_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13646_bdd_4_lut_LC_20_7_2  (
            .in0(N__75315),
            .in1(N__92629),
            .in2(N__75337),
            .in3(N__75330),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13649 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1976_1977_LC_20_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1976_1977_LC_20_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1976_1977_LC_20_7_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1976_1977_LC_20_7_4  (
            .in0(N__96244),
            .in1(N__95148),
            .in2(N__75316),
            .in3(N__77471),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93435),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2168_2169_LC_20_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2168_2169_LC_20_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2168_2169_LC_20_7_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2168_2169_LC_20_7_5  (
            .in0(N__95146),
            .in1(N__96246),
            .in2(N__75304),
            .in3(N__76353),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_22_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93435),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5048_5049_LC_20_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5048_5049_LC_20_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5048_5049_LC_20_7_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5048_5049_LC_20_7_6  (
            .in0(N__96245),
            .in1(N__95149),
            .in2(N__75292),
            .in3(N__77472),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93435),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5144_5145_LC_20_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5144_5145_LC_20_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5144_5145_LC_20_7_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5144_5145_LC_20_7_7  (
            .in0(N__95147),
            .in1(N__96247),
            .in2(N__75277),
            .in3(N__77040),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93435),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5612_5613_LC_20_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5612_5613_LC_20_8_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5612_5613_LC_20_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5612_5613_LC_20_8_0  (
            .in0(N__75261),
            .in1(N__75936),
            .in2(_gnd_net_),
            .in3(N__79982),
            .lcout(REG_mem_58_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93429),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11924_LC_20_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11924_LC_20_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11924_LC_20_8_1 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11924_LC_20_8_1  (
            .in0(N__91820),
            .in1(N__75262),
            .in2(N__76018),
            .in3(N__88575),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13730_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13730_bdd_4_lut_LC_20_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13730_bdd_4_lut_LC_20_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13730_bdd_4_lut_LC_20_8_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13730_bdd_4_lut_LC_20_8_2  (
            .in0(N__76029),
            .in1(N__91816),
            .in2(N__75253),
            .in3(N__75249),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13733 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14372_bdd_4_lut_LC_20_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14372_bdd_4_lut_LC_20_8_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14372_bdd_4_lut_LC_20_8_3 .LUT_INIT=16'b1010111010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14372_bdd_4_lut_LC_20_8_3  (
            .in0(N__76069),
            .in1(N__93481),
            .in2(N__92169),
            .in3(N__76063),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5420_5421_LC_20_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5420_5421_LC_20_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5420_5421_LC_20_8_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5420_5421_LC_20_8_4  (
            .in0(N__95502),
            .in1(N__75938),
            .in2(N__76030),
            .in3(N__95985),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93429),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5708_5709_LC_20_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5708_5709_LC_20_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5708_5709_LC_20_8_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5708_5709_LC_20_8_5  (
            .in0(N__75935),
            .in1(N__95503),
            .in2(N__76017),
            .in3(N__79787),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93429),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2348_2349_LC_20_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2348_2349_LC_20_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2348_2349_LC_20_8_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2348_2349_LC_20_8_6  (
            .in0(N__95501),
            .in1(N__75937),
            .in2(N__75606),
            .in3(N__95984),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93429),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4664_4665_LC_20_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4664_4665_LC_20_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4664_4665_LC_20_8_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4664_4665_LC_20_8_7  (
            .in0(N__75420),
            .in1(_gnd_net_),
            .in2(N__96321),
            .in3(N__75588),
            .lcout(REG_mem_48_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93429),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13388_bdd_4_lut_LC_20_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13388_bdd_4_lut_LC_20_9_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13388_bdd_4_lut_LC_20_9_0 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13388_bdd_4_lut_LC_20_9_0  (
            .in0(N__92269),
            .in1(N__75409),
            .in2(N__75397),
            .in3(N__75388),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12328_LC_20_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12328_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12328_LC_20_9_1 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12328_LC_20_9_1  (
            .in0(N__77490),
            .in1(N__92270),
            .in2(N__88749),
            .in3(N__75375),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14216_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14216_bdd_4_lut_LC_20_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14216_bdd_4_lut_LC_20_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14216_bdd_4_lut_LC_20_9_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14216_bdd_4_lut_LC_20_9_2  (
            .in0(N__77502),
            .in1(N__92271),
            .in2(N__75361),
            .in3(N__76368),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12054 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5054_5055_LC_20_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5054_5055_LC_20_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5054_5055_LC_20_9_3 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5054_5055_LC_20_9_3  (
            .in0(N__77449),
            .in1(N__77067),
            .in2(N__95687),
            .in3(N__89474),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93423),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5042_5043_LC_20_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5042_5043_LC_20_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5042_5043_LC_20_9_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5042_5043_LC_20_9_4  (
            .in0(N__76705),
            .in1(N__95497),
            .in2(N__77503),
            .in3(N__77451),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_52_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93423),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5234_5235_LC_20_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5234_5235_LC_20_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5234_5235_LC_20_9_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5234_5235_LC_20_9_5  (
            .in0(N__95495),
            .in1(N__76706),
            .in2(N__77491),
            .in3(N__76352),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93423),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1970_1971_LC_20_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1970_1971_LC_20_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1970_1971_LC_20_9_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i1970_1971_LC_20_9_6  (
            .in0(N__76704),
            .in1(N__95496),
            .in2(N__77265),
            .in3(N__77450),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_20_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93423),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5342_5343_LC_20_10_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5342_5343_LC_20_10_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5342_5343_LC_20_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5342_5343_LC_20_10_0  (
            .in0(N__77079),
            .in1(N__89468),
            .in2(_gnd_net_),
            .in3(N__77245),
            .lcout(REG_mem_55_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11705_LC_20_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11705_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11705_LC_20_10_1 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11705_LC_20_10_1  (
            .in0(N__91738),
            .in1(N__88546),
            .in2(N__76084),
            .in3(N__77080),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13460_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13460_bdd_4_lut_LC_20_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13460_bdd_4_lut_LC_20_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13460_bdd_4_lut_LC_20_10_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13460_bdd_4_lut_LC_20_10_2  (
            .in0(N__77056),
            .in1(N__91737),
            .in2(N__77071),
            .in3(N__77068),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11853 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5150_5151_LC_20_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5150_5151_LC_20_10_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5150_5151_LC_20_10_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5150_5151_LC_20_10_3  (
            .in0(N__94660),
            .in1(N__77055),
            .in2(N__89517),
            .in3(N__77022),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5138_5139_LC_20_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5138_5139_LC_20_10_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5138_5139_LC_20_10_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5138_5139_LC_20_10_4  (
            .in0(N__77021),
            .in1(N__76758),
            .in2(N__76369),
            .in3(N__94663),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_53_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5246_5247_LC_20_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5246_5247_LC_20_10_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5246_5247_LC_20_10_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5246_5247_LC_20_10_5  (
            .in0(N__94661),
            .in1(N__89473),
            .in2(N__76083),
            .in3(N__76308),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_54_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2936_2937_LC_20_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2936_2937_LC_20_10_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2936_2937_LC_20_10_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2936_2937_LC_20_10_6  (
            .in0(N__96324),
            .in1(N__94662),
            .in2(N__77652),
            .in3(N__77956),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_30_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93406),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12824_bdd_4_lut_LC_20_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12824_bdd_4_lut_LC_20_10_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12824_bdd_4_lut_LC_20_10_7 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12824_bdd_4_lut_LC_20_10_7  (
            .in0(N__91736),
            .in1(N__77635),
            .in2(N__83050),
            .in3(N__77617),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12827 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.i10484_3_lut_LC_20_11_0 .C_ON=1'b0;
    defparam \pc_tx.i10484_3_lut_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i10484_3_lut_LC_20_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \pc_tx.i10484_3_lut_LC_20_11_0  (
            .in0(N__78508),
            .in1(N__78535),
            .in2(_gnd_net_),
            .in3(N__83446),
            .lcout(),
            .ltout(\pc_tx.n12133_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.n13790_bdd_4_lut_LC_20_11_1 .C_ON=1'b0;
    defparam \pc_tx.n13790_bdd_4_lut_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \pc_tx.n13790_bdd_4_lut_LC_20_11_1 .LUT_INIT=16'b1011101010011000;
    LogicCell40 \pc_tx.n13790_bdd_4_lut_LC_20_11_1  (
            .in0(N__77509),
            .in1(N__83490),
            .in2(N__77596),
            .in3(N__77551),
            .lcout(),
            .ltout(\pc_tx.o_Tx_Serial_N_840_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.o_Tx_Serial_44_LC_20_11_2 .C_ON=1'b0;
    defparam \pc_tx.o_Tx_Serial_44_LC_20_11_2 .SEQ_MODE=4'b1000;
    defparam \pc_tx.o_Tx_Serial_44_LC_20_11_2 .LUT_INIT=16'b1111101001010101;
    LogicCell40 \pc_tx.o_Tx_Serial_44_LC_20_11_2  (
            .in0(N__83674),
            .in1(_gnd_net_),
            .in2(N__77593),
            .in3(N__83613),
            .lcout(UART_TX_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97378),
            .ce(N__97117),
            .sr(_gnd_net_));
    defparam \pc_tx.i10485_3_lut_LC_20_11_3 .C_ON=1'b0;
    defparam \pc_tx.i10485_3_lut_LC_20_11_3 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i10485_3_lut_LC_20_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pc_tx.i10485_3_lut_LC_20_11_3  (
            .in0(N__83447),
            .in1(N__77569),
            .in2(_gnd_net_),
            .in3(N__78469),
            .lcout(\pc_tx.n12134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.i10490_3_lut_LC_20_11_4 .C_ON=1'b0;
    defparam \pc_tx.i10490_3_lut_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i10490_3_lut_LC_20_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \pc_tx.i10490_3_lut_LC_20_11_4  (
            .in0(N__77545),
            .in1(N__77527),
            .in2(_gnd_net_),
            .in3(N__83448),
            .lcout(),
            .ltout(\pc_tx.n12139_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Bit_Index_1__bdd_4_lut_LC_20_11_5 .C_ON=1'b0;
    defparam \pc_tx.r_Bit_Index_1__bdd_4_lut_LC_20_11_5 .SEQ_MODE=4'b0000;
    defparam \pc_tx.r_Bit_Index_1__bdd_4_lut_LC_20_11_5 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \pc_tx.r_Bit_Index_1__bdd_4_lut_LC_20_11_5  (
            .in0(N__83524),
            .in1(N__83491),
            .in2(N__77512),
            .in3(N__78142),
            .lcout(\pc_tx.n13790 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.i10491_3_lut_LC_20_11_6 .C_ON=1'b0;
    defparam \pc_tx.i10491_3_lut_LC_20_11_6 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i10491_3_lut_LC_20_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \pc_tx.i10491_3_lut_LC_20_11_6  (
            .in0(N__78178),
            .in1(N__78157),
            .in2(_gnd_net_),
            .in3(N__83449),
            .lcout(\pc_tx.n12140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \bluejay_data_inst.i2_3_lut_adj_68_LC_20_11_7 .C_ON=1'b0;
    defparam \bluejay_data_inst.i2_3_lut_adj_68_LC_20_11_7 .SEQ_MODE=4'b0000;
    defparam \bluejay_data_inst.i2_3_lut_adj_68_LC_20_11_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \bluejay_data_inst.i2_3_lut_adj_68_LC_20_11_7  (
            .in0(N__78136),
            .in1(N__78103),
            .in2(_gnd_net_),
            .in3(N__78079),
            .lcout(\bluejay_data_inst.n1137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i11069_2_lut_3_lut_4_lut_LC_20_12_0 .C_ON=1'b0;
    defparam \timing_controller_inst.i11069_2_lut_3_lut_4_lut_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i11069_2_lut_3_lut_4_lut_LC_20_12_0 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \timing_controller_inst.i11069_2_lut_3_lut_4_lut_LC_20_12_0  (
            .in0(N__84070),
            .in1(N__81887),
            .in2(N__84016),
            .in3(N__82184),
            .lcout(\timing_controller_inst.n4301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i2319_2_lut_LC_20_12_1 .C_ON=1'b0;
    defparam \timing_controller_inst.i2319_2_lut_LC_20_12_1 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i2319_2_lut_LC_20_12_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \timing_controller_inst.i2319_2_lut_LC_20_12_1  (
            .in0(N__82185),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83995),
            .lcout(n3514),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i1_2_lut_LC_20_12_2 .C_ON=1'b0;
    defparam \timing_controller_inst.i1_2_lut_LC_20_12_2 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i1_2_lut_LC_20_12_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \timing_controller_inst.i1_2_lut_LC_20_12_2  (
            .in0(_gnd_net_),
            .in1(N__81888),
            .in2(_gnd_net_),
            .in3(N__81756),
            .lcout(n4_adj_1182),
            .ltout(n4_adj_1182_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_i3_LC_20_12_3 .C_ON=1'b0;
    defparam \timing_controller_inst.state_i3_LC_20_12_3 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_i3_LC_20_12_3 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \timing_controller_inst.state_i3_LC_20_12_3  (
            .in0(N__77989),
            .in1(N__84071),
            .in2(N__77983),
            .in3(N__77980),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97393),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i15_3_lut_LC_20_12_4 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i15_3_lut_LC_20_12_4 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i15_3_lut_LC_20_12_4 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \timing_controller_inst.mux_855_i15_3_lut_LC_20_12_4  (
            .in0(N__84469),
            .in1(N__82186),
            .in2(_gnd_net_),
            .in3(N__82413),
            .lcout(\timing_controller_inst.n1740 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i16_3_lut_LC_20_12_5 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i16_3_lut_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i16_3_lut_LC_20_12_5 .LUT_INIT=16'b0101110001011100;
    LogicCell40 \timing_controller_inst.mux_855_i16_3_lut_LC_20_12_5  (
            .in0(N__82187),
            .in1(N__84430),
            .in2(N__82424),
            .in3(_gnd_net_),
            .lcout(\timing_controller_inst.n1739 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_3__I_0_59_Mux_0_i7_4_lut_LC_20_12_6 .C_ON=1'b0;
    defparam \timing_controller_inst.state_3__I_0_59_Mux_0_i7_4_lut_LC_20_12_6 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.state_3__I_0_59_Mux_0_i7_4_lut_LC_20_12_6 .LUT_INIT=16'b1000010010110111;
    LogicCell40 \timing_controller_inst.state_3__I_0_59_Mux_0_i7_4_lut_LC_20_12_6  (
            .in0(N__83996),
            .in1(N__81889),
            .in2(N__81773),
            .in3(N__82189),
            .lcout(\timing_controller_inst.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i1_3_lut_LC_20_12_7 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i1_3_lut_LC_20_12_7 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i1_3_lut_LC_20_12_7 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \timing_controller_inst.mux_855_i1_3_lut_LC_20_12_7  (
            .in0(N__82188),
            .in1(_gnd_net_),
            .in2(N__82425),
            .in3(N__83830),
            .lcout(\timing_controller_inst.n1754 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i21_4_lut_LC_20_13_0 .C_ON=1'b0;
    defparam \timing_controller_inst.i21_4_lut_LC_20_13_0 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i21_4_lut_LC_20_13_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \timing_controller_inst.i21_4_lut_LC_20_13_0  (
            .in0(N__84565),
            .in1(N__84229),
            .in2(N__86695),
            .in3(N__84480),
            .lcout(\timing_controller_inst.n53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i14_LC_20_13_1 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i14_LC_20_13_1 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i14_LC_20_13_1 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i14_LC_20_13_1  (
            .in0(N__81999),
            .in1(N__82083),
            .in2(N__82240),
            .in3(N__78238),
            .lcout(\timing_controller_inst.state_timeout_counter_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97402),
            .ce(N__86037),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i12_LC_20_13_2 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i12_LC_20_13_2 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i12_LC_20_13_2 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i12_LC_20_13_2  (
            .in0(N__82082),
            .in1(N__78232),
            .in2(N__82242),
            .in3(N__81998),
            .lcout(\timing_controller_inst.state_timeout_counter_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97402),
            .ce(N__86037),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i15_LC_20_13_3 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i15_LC_20_13_3 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i15_LC_20_13_3 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i15_LC_20_13_3  (
            .in0(N__82000),
            .in1(N__82084),
            .in2(N__82241),
            .in3(N__78226),
            .lcout(\timing_controller_inst.state_timeout_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97402),
            .ce(N__86037),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i18_LC_20_13_4 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i18_LC_20_13_4 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i18_LC_20_13_4 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i18_LC_20_13_4  (
            .in0(N__82085),
            .in1(N__78220),
            .in2(N__82243),
            .in3(N__82001),
            .lcout(\timing_controller_inst.state_timeout_counter_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97402),
            .ce(N__86037),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i0_LC_20_13_5 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i0_LC_20_13_5 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i0_LC_20_13_5 .LUT_INIT=16'b0011011100000100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i0_LC_20_13_5  (
            .in0(N__81997),
            .in1(N__82081),
            .in2(N__82239),
            .in3(N__78214),
            .lcout(\timing_controller_inst.state_timeout_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97402),
            .ce(N__86037),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i19_LC_20_13_6 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i19_LC_20_13_6 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i19_LC_20_13_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i19_LC_20_13_6  (
            .in0(N__82086),
            .in1(N__82206),
            .in2(N__78208),
            .in3(N__82002),
            .lcout(\timing_controller_inst.state_timeout_counter_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97402),
            .ce(N__86037),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i20_LC_20_13_7 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i20_LC_20_13_7 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i20_LC_20_13_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i20_LC_20_13_7  (
            .in0(N__82003),
            .in1(N__82087),
            .in2(N__78193),
            .in3(N__82213),
            .lcout(\timing_controller_inst.state_timeout_counter_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97402),
            .ce(N__86037),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r__i1_LC_20_14_0 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r__i1_LC_20_14_0 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r__i1_LC_20_14_0 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_addr_r__i1_LC_20_14_0  (
            .in0(N__78454),
            .in1(N__78657),
            .in2(N__79027),
            .in3(N__78704),
            .lcout(rd_addr_r_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97410),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i0_LC_20_14_1 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i0_LC_20_14_1 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i0_LC_20_14_1 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i0_LC_20_14_1  (
            .in0(N__78544),
            .in1(N__78450),
            .in2(N__78334),
            .in3(N__78667),
            .lcout(fifo_temp_output_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97410),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Tx_Data_i0_LC_20_14_2 .C_ON=1'b0;
    defparam \pc_tx.r_Tx_Data_i0_LC_20_14_2 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Tx_Data_i0_LC_20_14_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pc_tx.r_Tx_Data_i0_LC_20_14_2  (
            .in0(N__81672),
            .in1(N__78531),
            .in2(_gnd_net_),
            .in3(N__78543),
            .lcout(r_Tx_Data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97410),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i1_LC_20_14_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i1_LC_20_14_3 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i1_LC_20_14_3 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i1_LC_20_14_3  (
            .in0(N__79075),
            .in1(N__78451),
            .in2(N__78335),
            .in3(N__78520),
            .lcout(fifo_temp_output_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97410),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Tx_Data_i1_LC_20_14_4 .C_ON=1'b0;
    defparam \pc_tx.r_Tx_Data_i1_LC_20_14_4 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Tx_Data_i1_LC_20_14_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pc_tx.r_Tx_Data_i1_LC_20_14_4  (
            .in0(N__81673),
            .in1(N__78519),
            .in2(_gnd_net_),
            .in3(N__78504),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97410),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i2_LC_20_14_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i2_LC_20_14_5 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i2_LC_20_14_5 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i2_LC_20_14_5  (
            .in0(N__78493),
            .in1(N__78452),
            .in2(N__78336),
            .in3(N__78481),
            .lcout(fifo_temp_output_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97410),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Tx_Data_i2_LC_20_14_6 .C_ON=1'b0;
    defparam \pc_tx.r_Tx_Data_i2_LC_20_14_6 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Tx_Data_i2_LC_20_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pc_tx.r_Tx_Data_i2_LC_20_14_6  (
            .in0(N__81674),
            .in1(N__78480),
            .in2(_gnd_net_),
            .in3(N__78465),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97410),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i3_LC_20_14_7 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i3_LC_20_14_7 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i3_LC_20_14_7 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i3_LC_20_14_7  (
            .in0(N__78862),
            .in1(N__78453),
            .in2(N__78337),
            .in3(N__78270),
            .lcout(fifo_temp_output_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97410),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i23_4_lut_LC_20_15_0 .C_ON=1'b0;
    defparam \timing_controller_inst.i23_4_lut_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i23_4_lut_LC_20_15_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \timing_controller_inst.i23_4_lut_LC_20_15_0  (
            .in0(N__84739),
            .in1(N__84813),
            .in2(N__84453),
            .in3(N__84169),
            .lcout(\timing_controller_inst.n55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i24_4_lut_LC_20_15_1 .C_ON=1'b0;
    defparam \timing_controller_inst.i24_4_lut_LC_20_15_1 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i24_4_lut_LC_20_15_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \timing_controller_inst.i24_4_lut_LC_20_15_1  (
            .in0(N__86074),
            .in1(N__83737),
            .in2(N__84511),
            .in3(N__86716),
            .lcout(\timing_controller_inst.n56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11764_LC_20_15_2 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11764_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11764_LC_20_15_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_11764_LC_20_15_2  (
            .in0(N__79009),
            .in1(N__79141),
            .in2(N__78731),
            .in3(N__79123),
            .lcout(),
            .ltout(\tx_fifo.lscc_fifo_inst.n13538_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i2_LC_20_15_3 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i2_LC_20_15_3 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i2_LC_20_15_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i2_LC_20_15_3  (
            .in0(N__79111),
            .in1(N__78705),
            .in2(N__79090),
            .in3(N__79087),
            .lcout(mem_LUT_data_raw_r_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97422),
            .ce(N__78656),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_LC_20_15_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_LC_20_15_5 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_LC_20_15_5  (
            .in0(N__79069),
            .in1(N__78709),
            .in2(N__79051),
            .in3(N__79010),
            .lcout(\tx_fifo.lscc_fifo_inst.n14234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i4_LC_20_16_5 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i4_LC_20_16_5 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i4_LC_20_16_5 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i4_LC_20_16_5  (
            .in0(N__78732),
            .in1(N__78901),
            .in2(N__78895),
            .in3(N__78874),
            .lcout(mem_LUT_data_raw_r_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97429),
            .ce(N__78658),
            .sr(_gnd_net_));
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i1_LC_20_17_1 .C_ON=1'b0;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i1_LC_20_17_1 .SEQ_MODE=4'b1000;
    defparam \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i1_LC_20_17_1 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i1_LC_20_17_1  (
            .in0(N__78850),
            .in1(N__78832),
            .in2(N__78820),
            .in3(N__78733),
            .lcout(mem_LUT_data_raw_r_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97436),
            .ce(N__78635),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13946_bdd_4_lut_LC_22_4_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13946_bdd_4_lut_LC_22_4_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13946_bdd_4_lut_LC_22_4_6 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13946_bdd_4_lut_LC_22_4_6  (
            .in0(N__78601),
            .in1(N__90349),
            .in2(N__78589),
            .in3(N__78577),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13949 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i7_LC_22_5_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i7_LC_22_5_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i7_LC_22_5_0 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i7_LC_22_5_0  (
            .in0(N__81099),
            .in1(N__79297),
            .in2(N__79219),
            .in3(N__78568),
            .lcout(REG_out_raw_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97445),
            .ce(N__80871),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_LC_22_5_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_LC_22_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_LC_22_5_1 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_LC_22_5_1  (
            .in0(N__81481),
            .in1(N__81100),
            .in2(N__79252),
            .in3(N__79306),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11700_LC_22_5_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11700_LC_22_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11700_LC_22_5_2 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11700_LC_22_5_2  (
            .in0(N__79291),
            .in1(N__85503),
            .in2(N__90385),
            .in3(N__79279),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13370_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13370_bdd_4_lut_LC_22_5_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13370_bdd_4_lut_LC_22_5_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13370_bdd_4_lut_LC_22_5_3 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13370_bdd_4_lut_LC_22_5_3  (
            .in0(N__79270),
            .in1(N__90355),
            .in2(N__79255),
            .in3(N__79165),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10353_3_lut_LC_22_5_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10353_3_lut_LC_22_5_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10353_3_lut_LC_22_5_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10353_3_lut_LC_22_5_4  (
            .in0(N__79243),
            .in1(N__85502),
            .in2(_gnd_net_),
            .in3(N__79231),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12002_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10354_3_lut_LC_22_5_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10354_3_lut_LC_22_5_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10354_3_lut_LC_22_5_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10354_3_lut_LC_22_5_5  (
            .in0(N__79339),
            .in1(_gnd_net_),
            .in2(N__79222),
            .in3(N__90354),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12003 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10136_3_lut_LC_22_6_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10136_3_lut_LC_22_6_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10136_3_lut_LC_22_6_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10136_3_lut_LC_22_6_0  (
            .in0(N__79413),
            .in1(N__88906),
            .in2(_gnd_net_),
            .in3(N__79210),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11789_LC_22_6_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11789_LC_22_6_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11789_LC_22_6_1 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11789_LC_22_6_1  (
            .in0(N__92174),
            .in1(N__79401),
            .in2(N__88912),
            .in3(N__79428),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13568_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13568_bdd_4_lut_LC_22_6_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13568_bdd_4_lut_LC_22_6_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13568_bdd_4_lut_LC_22_6_2 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13568_bdd_4_lut_LC_22_6_2  (
            .in0(N__79371),
            .in1(N__92173),
            .in2(N__79189),
            .in3(N__79186),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11835 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10140_3_lut_LC_22_6_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10140_3_lut_LC_22_6_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10140_3_lut_LC_22_6_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10140_3_lut_LC_22_6_4  (
            .in0(N__79330),
            .in1(N__88907),
            .in2(_gnd_net_),
            .in3(N__79159),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3416_3417_LC_22_6_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3416_3417_LC_22_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3416_3417_LC_22_6_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3416_3417_LC_22_6_5  (
            .in0(N__95618),
            .in1(N__96345),
            .in2(N__79429),
            .in3(N__83377),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93453),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i152_153_LC_22_6_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i152_153_LC_22_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i152_153_LC_22_6_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i152_153_LC_22_6_6  (
            .in0(N__96344),
            .in1(N__95619),
            .in2(N__79414),
            .in3(N__80318),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93453),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3320_3321_LC_22_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3320_3321_LC_22_7_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3320_3321_LC_22_7_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3320_3321_LC_22_7_0  (
            .in0(N__96388),
            .in1(N__95623),
            .in2(N__79402),
            .in3(N__80606),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93450),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11779_LC_22_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11779_LC_22_7_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11779_LC_22_7_1 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_1__bdd_4_lut_11779_LC_22_7_1  (
            .in0(N__79387),
            .in1(N__92636),
            .in2(N__85381),
            .in3(N__79381),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13526 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3224_3225_LC_22_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3224_3225_LC_22_7_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3224_3225_LC_22_7_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3224_3225_LC_22_7_2  (
            .in0(N__96387),
            .in1(N__95622),
            .in2(N__79372),
            .in3(N__80312),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93450),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10137_3_lut_LC_22_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10137_3_lut_LC_22_7_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10137_3_lut_LC_22_7_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10137_3_lut_LC_22_7_3  (
            .in0(N__80007),
            .in1(N__88878),
            .in2(_gnd_net_),
            .in3(N__79317),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11786_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13526_bdd_4_lut_LC_22_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13526_bdd_4_lut_LC_22_7_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13526_bdd_4_lut_LC_22_7_4 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13526_bdd_4_lut_LC_22_7_4  (
            .in0(N__79357),
            .in1(N__79348),
            .in2(N__79342),
            .in3(N__85269),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13529 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i728_729_LC_22_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i728_729_LC_22_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i728_729_LC_22_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i728_729_LC_22_7_5  (
            .in0(N__79329),
            .in1(N__96389),
            .in2(_gnd_net_),
            .in3(N__89661),
            .lcout(REG_mem_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93450),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i248_249_LC_22_7_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i248_249_LC_22_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i248_249_LC_22_7_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i248_249_LC_22_7_6  (
            .in0(N__96386),
            .in1(N__95621),
            .in2(N__79318),
            .in3(N__80605),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93450),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i344_345_LC_22_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i344_345_LC_22_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i344_345_LC_22_7_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i344_345_LC_22_7_7  (
            .in0(N__95620),
            .in1(N__96390),
            .in2(N__80008),
            .in3(N__83376),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93450),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5630_5631_LC_22_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5630_5631_LC_22_8_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5630_5631_LC_22_8_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5630_5631_LC_22_8_0  (
            .in0(N__79833),
            .in1(_gnd_net_),
            .in2(N__89520),
            .in3(N__79981),
            .lcout(REG_mem_58_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93441),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11690_LC_22_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11690_LC_22_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11690_LC_22_8_1 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11690_LC_22_8_1  (
            .in0(N__92172),
            .in1(N__79834),
            .in2(N__79489),
            .in3(N__88900),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13448_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13448_bdd_4_lut_LC_22_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13448_bdd_4_lut_LC_22_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13448_bdd_4_lut_LC_22_8_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13448_bdd_4_lut_LC_22_8_2  (
            .in0(N__79809),
            .in1(N__92170),
            .in2(N__79825),
            .in3(N__79821),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11862 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5534_5535_LC_22_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5534_5535_LC_22_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5534_5535_LC_22_8_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5534_5535_LC_22_8_3  (
            .in0(N__95314),
            .in1(N__89487),
            .in2(N__79822),
            .in3(N__97055),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93441),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5438_5439_LC_22_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5438_5439_LC_22_8_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5438_5439_LC_22_8_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5438_5439_LC_22_8_4  (
            .in0(N__89483),
            .in1(N__95317),
            .in2(N__79810),
            .in3(N__95979),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93441),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5726_5727_LC_22_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5726_5727_LC_22_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5726_5727_LC_22_8_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5726_5727_LC_22_8_5  (
            .in0(N__95315),
            .in1(N__89488),
            .in2(N__79488),
            .in3(N__79788),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_59_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93441),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2366_2367_LC_22_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2366_2367_LC_22_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2366_2367_LC_22_8_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2366_2367_LC_22_8_6  (
            .in0(N__89482),
            .in1(N__95316),
            .in2(N__79441),
            .in3(N__95978),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93441),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14042_bdd_4_lut_LC_22_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14042_bdd_4_lut_LC_22_8_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14042_bdd_4_lut_LC_22_8_7 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14042_bdd_4_lut_LC_22_8_7  (
            .in0(N__92171),
            .in1(N__79474),
            .in2(N__79456),
            .in3(N__79440),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3230_3231_LC_22_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3230_3231_LC_22_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3230_3231_LC_22_9_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3230_3231_LC_22_9_0  (
            .in0(N__89490),
            .in1(N__95321),
            .in2(N__80638),
            .in3(N__80311),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_33_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93436),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12093_LC_22_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12093_LC_22_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12093_LC_22_9_1 .LUT_INIT=16'b1011110010110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_12093_LC_22_9_1  (
            .in0(N__80334),
            .in1(N__91223),
            .in2(N__88905),
            .in3(N__80346),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13928_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13928_bdd_4_lut_LC_22_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13928_bdd_4_lut_LC_22_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13928_bdd_4_lut_LC_22_9_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13928_bdd_4_lut_LC_22_9_2  (
            .in0(N__91222),
            .in1(N__80637),
            .in2(N__80623),
            .in3(N__80619),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11760 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3134_3135_LC_22_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3134_3135_LC_22_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3134_3135_LC_22_9_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3134_3135_LC_22_9_3  (
            .in0(N__95318),
            .in1(N__89492),
            .in2(N__80620),
            .in3(N__82925),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_32_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93436),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3326_3327_LC_22_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3326_3327_LC_22_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3326_3327_LC_22_9_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3326_3327_LC_22_9_4  (
            .in0(N__89491),
            .in1(N__95322),
            .in2(N__80347),
            .in3(N__80575),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_34_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93436),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3422_3423_LC_22_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3422_3423_LC_22_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3422_3423_LC_22_9_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i3422_3423_LC_22_9_5  (
            .in0(N__95319),
            .in1(N__89493),
            .in2(N__80335),
            .in3(N__83335),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_35_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93436),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i158_159_LC_22_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i158_159_LC_22_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i158_159_LC_22_9_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i158_159_LC_22_9_6  (
            .in0(N__89489),
            .in1(N__95320),
            .in2(N__83104),
            .in3(N__80310),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93436),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11440_LC_22_10_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11440_LC_22_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11440_LC_22_10_1 .LUT_INIT=16'b1010110011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11440_LC_22_10_1  (
            .in0(N__90418),
            .in1(N__80041),
            .in2(N__85820),
            .in3(N__90083),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13136_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13136_bdd_4_lut_LC_22_10_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13136_bdd_4_lut_LC_22_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13136_bdd_4_lut_LC_22_10_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13136_bdd_4_lut_LC_22_10_2  (
            .in0(N__90081),
            .in1(N__80032),
            .in2(N__80023),
            .in3(N__80020),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11898 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11390_LC_22_10_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11390_LC_22_10_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11390_LC_22_10_3 .LUT_INIT=16'b1010110011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11390_LC_22_10_3  (
            .in0(N__81562),
            .in1(N__81553),
            .in2(N__85819),
            .in3(N__90082),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13082_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13082_bdd_4_lut_LC_22_10_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13082_bdd_4_lut_LC_22_10_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13082_bdd_4_lut_LC_22_10_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13082_bdd_4_lut_LC_22_10_4  (
            .in0(N__90080),
            .in1(N__81544),
            .in2(N__81535),
            .in3(N__81532),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11913_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_11550_LC_22_10_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_11550_LC_22_10_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_11550_LC_22_10_5 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_4__bdd_4_lut_11550_LC_22_10_5  (
            .in0(N__81092),
            .in1(N__92707),
            .in2(N__81517),
            .in3(N__81450),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13058_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i9_LC_22_10_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i9_LC_22_10_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i9_LC_22_10_6 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_out_raw__i9_LC_22_10_6  (
            .in0(N__81106),
            .in1(N__81091),
            .in2(N__80905),
            .in3(N__89758),
            .lcout(REG_out_raw_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97411),
            .ce(N__80876),
            .sr(_gnd_net_));
    defparam \pc_tx.i11046_4_lut_4_lut_LC_22_11_0 .C_ON=1'b0;
    defparam \pc_tx.i11046_4_lut_4_lut_LC_22_11_0 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i11046_4_lut_4_lut_LC_22_11_0 .LUT_INIT=16'b1010000001000100;
    LogicCell40 \pc_tx.i11046_4_lut_4_lut_LC_22_11_0  (
            .in0(N__83599),
            .in1(N__81629),
            .in2(N__83563),
            .in3(N__83653),
            .lcout(),
            .ltout(n11339_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Tx_Active_46_LC_22_11_1 .C_ON=1'b0;
    defparam \pc_tx.r_Tx_Active_46_LC_22_11_1 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Tx_Active_46_LC_22_11_1 .LUT_INIT=16'b1000110011011100;
    LogicCell40 \pc_tx.r_Tx_Active_46_LC_22_11_1  (
            .in0(N__83909),
            .in1(N__80649),
            .in2(N__80668),
            .in3(N__83605),
            .lcout(tx_uart_active_flag),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97394),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_SM_Main_i2_LC_22_11_2 .C_ON=1'b0;
    defparam \pc_tx.r_SM_Main_i2_LC_22_11_2 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_SM_Main_i2_LC_22_11_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pc_tx.r_SM_Main_i2_LC_22_11_2  (
            .in0(N__83562),
            .in1(N__83606),
            .in2(N__83673),
            .in3(N__83908),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97394),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.i1_3_lut_4_lut_adj_22_LC_22_11_3 .C_ON=1'b0;
    defparam \pc_tx.i1_3_lut_4_lut_adj_22_LC_22_11_3 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i1_3_lut_4_lut_adj_22_LC_22_11_3 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \pc_tx.i1_3_lut_4_lut_adj_22_LC_22_11_3  (
            .in0(N__83906),
            .in1(N__83561),
            .in2(N__83671),
            .in3(N__83603),
            .lcout(n4133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.i2_3_lut_4_lut_LC_22_11_4 .C_ON=1'b0;
    defparam \pc_tx.i2_3_lut_4_lut_LC_22_11_4 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i2_3_lut_4_lut_LC_22_11_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \pc_tx.i2_3_lut_4_lut_LC_22_11_4  (
            .in0(N__83604),
            .in1(N__81631),
            .in2(N__83672),
            .in3(N__83907),
            .lcout(n3710),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.i11085_4_lut_LC_22_11_5 .C_ON=1'b0;
    defparam \pc_tx.i11085_4_lut_LC_22_11_5 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i11085_4_lut_LC_22_11_5 .LUT_INIT=16'b0100010001000101;
    LogicCell40 \pc_tx.i11085_4_lut_LC_22_11_5  (
            .in0(N__83904),
            .in1(N__83560),
            .in2(N__83670),
            .in3(N__83600),
            .lcout(\pc_tx.n4577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.i1_3_lut_4_lut_LC_22_11_6 .C_ON=1'b0;
    defparam \pc_tx.i1_3_lut_4_lut_LC_22_11_6 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i1_3_lut_4_lut_LC_22_11_6 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \pc_tx.i1_3_lut_4_lut_LC_22_11_6  (
            .in0(N__83602),
            .in1(N__83905),
            .in2(N__83536),
            .in3(N__83657),
            .lcout(\pc_tx.n4468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.i1627_3_lut_LC_22_11_7 .C_ON=1'b0;
    defparam \pc_tx.i1627_3_lut_LC_22_11_7 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i1627_3_lut_LC_22_11_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pc_tx.i1627_3_lut_LC_22_11_7  (
            .in0(N__81630),
            .in1(N__83601),
            .in2(_gnd_net_),
            .in3(N__83532),
            .lcout(\pc_tx.n2813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i18_4_lut_LC_22_12_0 .C_ON=1'b0;
    defparam \timing_controller_inst.i18_4_lut_LC_22_12_0 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i18_4_lut_LC_22_12_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \timing_controller_inst.i18_4_lut_LC_22_12_0  (
            .in0(N__84778),
            .in1(N__84208),
            .in2(N__84415),
            .in3(N__84145),
            .lcout(\timing_controller_inst.n50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i1_2_lut_3_lut_4_lut_LC_22_12_1 .C_ON=1'b0;
    defparam \timing_controller_inst.i1_2_lut_3_lut_4_lut_LC_22_12_1 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i1_2_lut_3_lut_4_lut_LC_22_12_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \timing_controller_inst.i1_2_lut_3_lut_4_lut_LC_22_12_1  (
            .in0(N__81910),
            .in1(N__81776),
            .in2(N__83991),
            .in3(N__84094),
            .lcout(\timing_controller_inst.n11368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i11088_2_lut_LC_22_12_2 .C_ON=1'b0;
    defparam \timing_controller_inst.i11088_2_lut_LC_22_12_2 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i11088_2_lut_LC_22_12_2 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \timing_controller_inst.i11088_2_lut_LC_22_12_2  (
            .in0(N__84093),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81909),
            .lcout(\timing_controller_inst.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.invert_55_i3_LC_22_12_3 .C_ON=1'b0;
    defparam \timing_controller_inst.invert_55_i3_LC_22_12_3 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.invert_55_i3_LC_22_12_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \timing_controller_inst.invert_55_i3_LC_22_12_3  (
            .in0(N__83965),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82247),
            .lcout(UPDATE_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97412),
            .ce(),
            .sr(N__81574));
    defparam i6317_2_lut_3_lut_LC_22_12_4.C_ON=1'b0;
    defparam i6317_2_lut_3_lut_LC_22_12_4.SEQ_MODE=4'b0000;
    defparam i6317_2_lut_3_lut_LC_22_12_4.LUT_INIT=16'b1110111010101010;
    LogicCell40 i6317_2_lut_3_lut_LC_22_12_4 (
            .in0(N__81775),
            .in1(N__82244),
            .in2(_gnd_net_),
            .in3(N__83960),
            .lcout(),
            .ltout(n7495_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i924_4_lut_LC_22_12_5 .C_ON=1'b0;
    defparam \timing_controller_inst.i924_4_lut_LC_22_12_5 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i924_4_lut_LC_22_12_5 .LUT_INIT=16'b0000000001001110;
    LogicCell40 \timing_controller_inst.i924_4_lut_LC_22_12_5  (
            .in0(N__81912),
            .in1(N__81796),
            .in2(N__81565),
            .in3(N__84095),
            .lcout(\timing_controller_inst.n1793 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i913_2_lut_3_lut_LC_22_12_6 .C_ON=1'b0;
    defparam \timing_controller_inst.i913_2_lut_3_lut_LC_22_12_6 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i913_2_lut_3_lut_LC_22_12_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \timing_controller_inst.i913_2_lut_3_lut_LC_22_12_6  (
            .in0(N__81778),
            .in1(N__82245),
            .in2(_gnd_net_),
            .in3(N__83964),
            .lcout(\timing_controller_inst.n1875 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i6413_3_lut_LC_22_12_7 .C_ON=1'b0;
    defparam \timing_controller_inst.i6413_3_lut_LC_22_12_7 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i6413_3_lut_LC_22_12_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \timing_controller_inst.i6413_3_lut_LC_22_12_7  (
            .in0(N__81911),
            .in1(N__81777),
            .in2(_gnd_net_),
            .in3(N__82246),
            .lcout(\timing_controller_inst.n7592 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3114_4_lut_LC_22_13_0.C_ON=1'b0;
    defparam i3114_4_lut_LC_22_13_0.SEQ_MODE=4'b0000;
    defparam i3114_4_lut_LC_22_13_0.LUT_INIT=16'b0111010000000000;
    LogicCell40 i3114_4_lut_LC_22_13_0 (
            .in0(N__81789),
            .in1(N__84112),
            .in2(N__81837),
            .in3(N__81760),
            .lcout(n1616),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i919_4_lut_LC_22_13_1.C_ON=1'b0;
    defparam i919_4_lut_LC_22_13_1.SEQ_MODE=4'b0000;
    defparam i919_4_lut_LC_22_13_1.LUT_INIT=16'b0101011100000010;
    LogicCell40 i919_4_lut_LC_22_13_1 (
            .in0(N__84113),
            .in1(N__81790),
            .in2(N__81774),
            .in3(N__81697),
            .lcout(n1721),
            .ltout(n1721_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i1_2_lut_adj_86_LC_22_13_2 .C_ON=1'b0;
    defparam \timing_controller_inst.i1_2_lut_adj_86_LC_22_13_2 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i1_2_lut_adj_86_LC_22_13_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \timing_controller_inst.i1_2_lut_adj_86_LC_22_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__81685),
            .in3(N__84667),
            .lcout(\timing_controller_inst.n11347 ),
            .ltout(\timing_controller_inst.n11347_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i11121_3_lut_4_lut_LC_22_13_3 .C_ON=1'b0;
    defparam \timing_controller_inst.i11121_3_lut_4_lut_LC_22_13_3 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i11121_3_lut_4_lut_LC_22_13_3 .LUT_INIT=16'b0100010111001111;
    LogicCell40 \timing_controller_inst.i11121_3_lut_4_lut_LC_22_13_3  (
            .in0(N__84114),
            .in1(N__82031),
            .in2(N__81682),
            .in3(N__81833),
            .lcout(\timing_controller_inst.n4589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i3384_2_lut_3_lut_LC_22_13_4 .C_ON=1'b0;
    defparam \timing_controller_inst.i3384_2_lut_3_lut_LC_22_13_4 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i3384_2_lut_3_lut_LC_22_13_4 .LUT_INIT=16'b0000101010101010;
    LogicCell40 \timing_controller_inst.i3384_2_lut_3_lut_LC_22_13_4  (
            .in0(N__82032),
            .in1(_gnd_net_),
            .in2(N__81838),
            .in3(N__84115),
            .lcout(\timing_controller_inst.n4586 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i1_LC_22_13_5 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i1_LC_22_13_5 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i1_LC_22_13_5 .LUT_INIT=16'b0100111001001110;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i1_LC_22_13_5  (
            .in0(N__82364),
            .in1(N__83794),
            .in2(N__82320),
            .in3(_gnd_net_),
            .lcout(\timing_controller_inst.state_timeout_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97423),
            .ce(N__86038),
            .sr(N__81922));
    defparam \timing_controller_inst.state_timeout_counter_i0_i2_LC_22_13_6 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i2_LC_22_13_6 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i2_LC_22_13_6 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i2_LC_22_13_6  (
            .in0(N__82365),
            .in1(N__83746),
            .in2(_gnd_net_),
            .in3(N__82297),
            .lcout(\timing_controller_inst.state_timeout_counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97423),
            .ce(N__86038),
            .sr(N__81922));
    defparam \timing_controller_inst.i1_2_lut_3_lut_adj_89_LC_22_13_7 .C_ON=1'b0;
    defparam \timing_controller_inst.i1_2_lut_3_lut_adj_89_LC_22_13_7 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i1_2_lut_3_lut_adj_89_LC_22_13_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \timing_controller_inst.i1_2_lut_3_lut_adj_89_LC_22_13_7  (
            .in0(N__82293),
            .in1(N__83966),
            .in2(_gnd_net_),
            .in3(N__81916),
            .lcout(n3929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i22_4_lut_LC_22_14_0 .C_ON=1'b0;
    defparam \timing_controller_inst.i22_4_lut_LC_22_14_0 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i22_4_lut_LC_22_14_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \timing_controller_inst.i22_4_lut_LC_22_14_0  (
            .in0(N__84244),
            .in1(N__84264),
            .in2(N__84339),
            .in3(N__84759),
            .lcout(\timing_controller_inst.n54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i5_LC_22_14_1 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i5_LC_22_14_1 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i5_LC_22_14_1 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i5_LC_22_14_1  (
            .in0(N__82058),
            .in1(N__84253),
            .in2(N__82324),
            .in3(_gnd_net_),
            .lcout(\timing_controller_inst.state_timeout_counter_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97430),
            .ce(N__86039),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i24_3_lut_LC_22_14_2 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i24_3_lut_LC_22_14_2 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i24_3_lut_LC_22_14_2 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \timing_controller_inst.mux_855_i24_3_lut_LC_22_14_2  (
            .in0(N__82310),
            .in1(N__82367),
            .in2(_gnd_net_),
            .in3(N__84721),
            .lcout(\timing_controller_inst.n1731 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i4_3_lut_LC_22_14_3 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i4_3_lut_LC_22_14_3 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i4_3_lut_LC_22_14_3 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \timing_controller_inst.mux_855_i4_3_lut_LC_22_14_3  (
            .in0(N__82368),
            .in1(N__83716),
            .in2(N__82322),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\timing_controller_inst.n1751_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i3_LC_22_14_4 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i3_LC_22_14_4 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i3_LC_22_14_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i3_LC_22_14_4  (
            .in0(N__82312),
            .in1(N__82057),
            .in2(N__81811),
            .in3(N__81977),
            .lcout(\timing_controller_inst.state_timeout_counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97430),
            .ce(N__86039),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i23_3_lut_LC_22_14_5 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i23_3_lut_LC_22_14_5 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i23_3_lut_LC_22_14_5 .LUT_INIT=16'b0100111001001110;
    LogicCell40 \timing_controller_inst.mux_855_i23_3_lut_LC_22_14_5  (
            .in0(N__82366),
            .in1(N__84748),
            .in2(N__82321),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\timing_controller_inst.n1732_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i22_LC_22_14_6 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i22_LC_22_14_6 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i22_LC_22_14_6 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i22_LC_22_14_6  (
            .in0(N__82311),
            .in1(N__82055),
            .in2(N__81808),
            .in3(N__81976),
            .lcout(\timing_controller_inst.state_timeout_counter_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97430),
            .ce(N__86039),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i23_LC_22_14_7 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i23_LC_22_14_7 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i23_LC_22_14_7 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i23_LC_22_14_7  (
            .in0(N__82056),
            .in1(N__81805),
            .in2(N__82323),
            .in3(N__81978),
            .lcout(\timing_controller_inst.state_timeout_counter_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97430),
            .ce(N__86039),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i25_3_lut_LC_22_15_0 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i25_3_lut_LC_22_15_0 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i25_3_lut_LC_22_15_0 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \timing_controller_inst.mux_855_i25_3_lut_LC_22_15_0  (
            .in0(N__82315),
            .in1(_gnd_net_),
            .in2(N__82411),
            .in3(N__84607),
            .lcout(),
            .ltout(\timing_controller_inst.n1730_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i24_LC_22_15_1 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i24_LC_22_15_1 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i24_LC_22_15_1 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i24_LC_22_15_1  (
            .in0(N__81980),
            .in1(N__82062),
            .in2(N__82432),
            .in3(N__82317),
            .lcout(\timing_controller_inst.state_timeout_counter_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97437),
            .ce(N__86056),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i4_LC_22_15_2 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i4_LC_22_15_2 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i4_LC_22_15_2 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i4_LC_22_15_2  (
            .in0(N__82318),
            .in1(N__82060),
            .in2(N__82412),
            .in3(N__84286),
            .lcout(\timing_controller_inst.state_timeout_counter_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97437),
            .ce(N__86056),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i10_3_lut_LC_22_15_3 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i10_3_lut_LC_22_15_3 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i10_3_lut_LC_22_15_3 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \timing_controller_inst.mux_855_i10_3_lut_LC_22_15_3  (
            .in0(N__84178),
            .in1(N__82313),
            .in2(_gnd_net_),
            .in3(N__82389),
            .lcout(),
            .ltout(\timing_controller_inst.n1745_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i9_LC_22_15_4 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i9_LC_22_15_4 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i9_LC_22_15_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i9_LC_22_15_4  (
            .in0(N__82319),
            .in1(N__82061),
            .in2(N__82429),
            .in3(N__81981),
            .lcout(\timing_controller_inst.state_timeout_counter_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97437),
            .ce(N__86056),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.mux_855_i11_3_lut_LC_22_15_5 .C_ON=1'b0;
    defparam \timing_controller_inst.mux_855_i11_3_lut_LC_22_15_5 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.mux_855_i11_3_lut_LC_22_15_5 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \timing_controller_inst.mux_855_i11_3_lut_LC_22_15_5  (
            .in0(N__84154),
            .in1(N__82314),
            .in2(_gnd_net_),
            .in3(N__82390),
            .lcout(),
            .ltout(\timing_controller_inst.n1744_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i10_LC_22_15_6 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i10_LC_22_15_6 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i10_LC_22_15_6 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i10_LC_22_15_6  (
            .in0(N__82316),
            .in1(N__82059),
            .in2(N__82006),
            .in3(N__81979),
            .lcout(\timing_controller_inst.state_timeout_counter_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97437),
            .ce(N__86056),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i20_4_lut_LC_22_15_7 .C_ON=1'b0;
    defparam \timing_controller_inst.i20_4_lut_LC_22_15_7 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i20_4_lut_LC_22_15_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \timing_controller_inst.i20_4_lut_LC_22_15_7  (
            .in0(N__84391),
            .in1(N__84297),
            .in2(N__83815),
            .in3(N__84618),
            .lcout(\timing_controller_inst.n52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i6_2_lut_LC_22_16_5 .C_ON=1'b0;
    defparam \timing_controller_inst.i6_2_lut_LC_22_16_5 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i6_2_lut_LC_22_16_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \timing_controller_inst.i6_2_lut_LC_22_16_5  (
            .in0(N__84544),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84189),
            .lcout(),
            .ltout(\timing_controller_inst.n38_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.i26_4_lut_LC_22_16_6 .C_ON=1'b0;
    defparam \timing_controller_inst.i26_4_lut_LC_22_16_6 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.i26_4_lut_LC_22_16_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \timing_controller_inst.i26_4_lut_LC_22_16_6  (
            .in0(N__81940),
            .in1(N__84582),
            .in2(N__81934),
            .in3(N__84598),
            .lcout(\timing_controller_inst.n58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i0_LC_23_5_0.C_ON=1'b1;
    defparam led_counter_1106_1179__i0_LC_23_5_0.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i0_LC_23_5_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i0_LC_23_5_0 (
            .in0(_gnd_net_),
            .in1(N__82504),
            .in2(_gnd_net_),
            .in3(N__82498),
            .lcout(n25_adj_1187),
            .ltout(),
            .carryin(bfn_23_5_0_),
            .carryout(n10670),
            .clk(N__97449),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i1_LC_23_5_1.C_ON=1'b1;
    defparam led_counter_1106_1179__i1_LC_23_5_1.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i1_LC_23_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i1_LC_23_5_1 (
            .in0(_gnd_net_),
            .in1(N__82495),
            .in2(_gnd_net_),
            .in3(N__82489),
            .lcout(n24_adj_1188),
            .ltout(),
            .carryin(n10670),
            .carryout(n10671),
            .clk(N__97449),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i2_LC_23_5_2.C_ON=1'b1;
    defparam led_counter_1106_1179__i2_LC_23_5_2.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i2_LC_23_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i2_LC_23_5_2 (
            .in0(_gnd_net_),
            .in1(N__82486),
            .in2(_gnd_net_),
            .in3(N__82480),
            .lcout(n23_adj_1189),
            .ltout(),
            .carryin(n10671),
            .carryout(n10672),
            .clk(N__97449),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i3_LC_23_5_3.C_ON=1'b1;
    defparam led_counter_1106_1179__i3_LC_23_5_3.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i3_LC_23_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i3_LC_23_5_3 (
            .in0(_gnd_net_),
            .in1(N__82477),
            .in2(_gnd_net_),
            .in3(N__82471),
            .lcout(n22_adj_1190),
            .ltout(),
            .carryin(n10672),
            .carryout(n10673),
            .clk(N__97449),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i4_LC_23_5_4.C_ON=1'b1;
    defparam led_counter_1106_1179__i4_LC_23_5_4.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i4_LC_23_5_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i4_LC_23_5_4 (
            .in0(_gnd_net_),
            .in1(N__82468),
            .in2(_gnd_net_),
            .in3(N__82462),
            .lcout(n21_adj_1191),
            .ltout(),
            .carryin(n10673),
            .carryout(n10674),
            .clk(N__97449),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i5_LC_23_5_5.C_ON=1'b1;
    defparam led_counter_1106_1179__i5_LC_23_5_5.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i5_LC_23_5_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i5_LC_23_5_5 (
            .in0(_gnd_net_),
            .in1(N__82459),
            .in2(_gnd_net_),
            .in3(N__82453),
            .lcout(n20_adj_1192),
            .ltout(),
            .carryin(n10674),
            .carryout(n10675),
            .clk(N__97449),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i6_LC_23_5_6.C_ON=1'b1;
    defparam led_counter_1106_1179__i6_LC_23_5_6.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i6_LC_23_5_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i6_LC_23_5_6 (
            .in0(_gnd_net_),
            .in1(N__82450),
            .in2(_gnd_net_),
            .in3(N__82444),
            .lcout(n19_adj_1193),
            .ltout(),
            .carryin(n10675),
            .carryout(n10676),
            .clk(N__97449),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i7_LC_23_5_7.C_ON=1'b1;
    defparam led_counter_1106_1179__i7_LC_23_5_7.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i7_LC_23_5_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i7_LC_23_5_7 (
            .in0(_gnd_net_),
            .in1(N__82441),
            .in2(_gnd_net_),
            .in3(N__82435),
            .lcout(n18_adj_1194),
            .ltout(),
            .carryin(n10676),
            .carryout(n10677),
            .clk(N__97449),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i8_LC_23_6_0.C_ON=1'b1;
    defparam led_counter_1106_1179__i8_LC_23_6_0.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i8_LC_23_6_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i8_LC_23_6_0 (
            .in0(_gnd_net_),
            .in1(N__82585),
            .in2(_gnd_net_),
            .in3(N__82579),
            .lcout(n17_adj_1195),
            .ltout(),
            .carryin(bfn_23_6_0_),
            .carryout(n10678),
            .clk(N__97446),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i9_LC_23_6_1.C_ON=1'b1;
    defparam led_counter_1106_1179__i9_LC_23_6_1.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i9_LC_23_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i9_LC_23_6_1 (
            .in0(_gnd_net_),
            .in1(N__82576),
            .in2(_gnd_net_),
            .in3(N__82570),
            .lcout(n16_adj_1196),
            .ltout(),
            .carryin(n10678),
            .carryout(n10679),
            .clk(N__97446),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i10_LC_23_6_2.C_ON=1'b1;
    defparam led_counter_1106_1179__i10_LC_23_6_2.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i10_LC_23_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i10_LC_23_6_2 (
            .in0(_gnd_net_),
            .in1(N__82567),
            .in2(_gnd_net_),
            .in3(N__82561),
            .lcout(n15_adj_1197),
            .ltout(),
            .carryin(n10679),
            .carryout(n10680),
            .clk(N__97446),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i11_LC_23_6_3.C_ON=1'b1;
    defparam led_counter_1106_1179__i11_LC_23_6_3.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i11_LC_23_6_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i11_LC_23_6_3 (
            .in0(_gnd_net_),
            .in1(N__82558),
            .in2(_gnd_net_),
            .in3(N__82552),
            .lcout(n14_adj_1198),
            .ltout(),
            .carryin(n10680),
            .carryout(n10681),
            .clk(N__97446),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i12_LC_23_6_4.C_ON=1'b1;
    defparam led_counter_1106_1179__i12_LC_23_6_4.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i12_LC_23_6_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i12_LC_23_6_4 (
            .in0(_gnd_net_),
            .in1(N__82549),
            .in2(_gnd_net_),
            .in3(N__82543),
            .lcout(n13),
            .ltout(),
            .carryin(n10681),
            .carryout(n10682),
            .clk(N__97446),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i13_LC_23_6_5.C_ON=1'b1;
    defparam led_counter_1106_1179__i13_LC_23_6_5.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i13_LC_23_6_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i13_LC_23_6_5 (
            .in0(_gnd_net_),
            .in1(N__82540),
            .in2(_gnd_net_),
            .in3(N__82534),
            .lcout(n12),
            .ltout(),
            .carryin(n10682),
            .carryout(n10683),
            .clk(N__97446),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i14_LC_23_6_6.C_ON=1'b1;
    defparam led_counter_1106_1179__i14_LC_23_6_6.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i14_LC_23_6_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i14_LC_23_6_6 (
            .in0(_gnd_net_),
            .in1(N__82531),
            .in2(_gnd_net_),
            .in3(N__82525),
            .lcout(n11),
            .ltout(),
            .carryin(n10683),
            .carryout(n10684),
            .clk(N__97446),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i15_LC_23_6_7.C_ON=1'b1;
    defparam led_counter_1106_1179__i15_LC_23_6_7.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i15_LC_23_6_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i15_LC_23_6_7 (
            .in0(_gnd_net_),
            .in1(N__82522),
            .in2(_gnd_net_),
            .in3(N__82516),
            .lcout(n10_adj_1199),
            .ltout(),
            .carryin(n10684),
            .carryout(n10685),
            .clk(N__97446),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i16_LC_23_7_0.C_ON=1'b1;
    defparam led_counter_1106_1179__i16_LC_23_7_0.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i16_LC_23_7_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i16_LC_23_7_0 (
            .in0(_gnd_net_),
            .in1(N__82513),
            .in2(_gnd_net_),
            .in3(N__82507),
            .lcout(n9),
            .ltout(),
            .carryin(bfn_23_7_0_),
            .carryout(n10686),
            .clk(N__97442),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i17_LC_23_7_1.C_ON=1'b1;
    defparam led_counter_1106_1179__i17_LC_23_7_1.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i17_LC_23_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i17_LC_23_7_1 (
            .in0(_gnd_net_),
            .in1(N__82675),
            .in2(_gnd_net_),
            .in3(N__82669),
            .lcout(n8),
            .ltout(),
            .carryin(n10686),
            .carryout(n10687),
            .clk(N__97442),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i18_LC_23_7_2.C_ON=1'b1;
    defparam led_counter_1106_1179__i18_LC_23_7_2.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i18_LC_23_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i18_LC_23_7_2 (
            .in0(_gnd_net_),
            .in1(N__82666),
            .in2(_gnd_net_),
            .in3(N__82660),
            .lcout(n7_adj_1200),
            .ltout(),
            .carryin(n10687),
            .carryout(n10688),
            .clk(N__97442),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i19_LC_23_7_3.C_ON=1'b1;
    defparam led_counter_1106_1179__i19_LC_23_7_3.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i19_LC_23_7_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i19_LC_23_7_3 (
            .in0(_gnd_net_),
            .in1(N__82657),
            .in2(_gnd_net_),
            .in3(N__82651),
            .lcout(n6),
            .ltout(),
            .carryin(n10688),
            .carryout(n10689),
            .clk(N__97442),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i20_LC_23_7_4.C_ON=1'b1;
    defparam led_counter_1106_1179__i20_LC_23_7_4.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i20_LC_23_7_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i20_LC_23_7_4 (
            .in0(_gnd_net_),
            .in1(N__82648),
            .in2(_gnd_net_),
            .in3(N__82642),
            .lcout(n5_adj_1201),
            .ltout(),
            .carryin(n10689),
            .carryout(n10690),
            .clk(N__97442),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i21_LC_23_7_5.C_ON=1'b1;
    defparam led_counter_1106_1179__i21_LC_23_7_5.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i21_LC_23_7_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i21_LC_23_7_5 (
            .in0(_gnd_net_),
            .in1(N__82639),
            .in2(_gnd_net_),
            .in3(N__82633),
            .lcout(n4_adj_1202),
            .ltout(),
            .carryin(n10690),
            .carryout(n10691),
            .clk(N__97442),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i22_LC_23_7_6.C_ON=1'b1;
    defparam led_counter_1106_1179__i22_LC_23_7_6.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i22_LC_23_7_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i22_LC_23_7_6 (
            .in0(_gnd_net_),
            .in1(N__82630),
            .in2(_gnd_net_),
            .in3(N__82624),
            .lcout(n3),
            .ltout(),
            .carryin(n10691),
            .carryout(n10692),
            .clk(N__97442),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i23_LC_23_7_7.C_ON=1'b1;
    defparam led_counter_1106_1179__i23_LC_23_7_7.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i23_LC_23_7_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i23_LC_23_7_7 (
            .in0(_gnd_net_),
            .in1(N__82621),
            .in2(_gnd_net_),
            .in3(N__82615),
            .lcout(n2_adj_1203),
            .ltout(),
            .carryin(n10692),
            .carryout(n10693),
            .clk(N__97442),
            .ce(),
            .sr(_gnd_net_));
    defparam led_counter_1106_1179__i24_LC_23_8_0.C_ON=1'b0;
    defparam led_counter_1106_1179__i24_LC_23_8_0.SEQ_MODE=4'b1000;
    defparam led_counter_1106_1179__i24_LC_23_8_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 led_counter_1106_1179__i24_LC_23_8_0 (
            .in0(_gnd_net_),
            .in1(N__82596),
            .in2(_gnd_net_),
            .in3(N__82612),
            .lcout(DEBUG_0_c_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97438),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i350_351_LC_23_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i350_351_LC_23_9_0 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i350_351_LC_23_9_0 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i350_351_LC_23_9_0  (
            .in0(N__83136),
            .in1(N__95104),
            .in2(N__89528),
            .in3(N__83342),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_3_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93442),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11385_LC_23_9_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11385_LC_23_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11385_LC_23_9_1 .LUT_INIT=16'b1101110110100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11385_LC_23_9_1  (
            .in0(N__91227),
            .in1(N__83137),
            .in2(N__83128),
            .in3(N__88899),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13070_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13070_bdd_4_lut_LC_23_9_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13070_bdd_4_lut_LC_23_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13070_bdd_4_lut_LC_23_9_2 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13070_bdd_4_lut_LC_23_9_2  (
            .in0(N__83103),
            .in1(N__82705),
            .in2(N__83089),
            .in3(N__91224),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13073 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11171_LC_23_9_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11171_LC_23_9_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11171_LC_23_9_3 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11171_LC_23_9_3  (
            .in0(N__91226),
            .in1(N__88898),
            .in2(N__83086),
            .in3(N__83065),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n12824 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14246_bdd_4_lut_LC_23_9_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14246_bdd_4_lut_LC_23_9_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14246_bdd_4_lut_LC_23_9_4 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14246_bdd_4_lut_LC_23_9_4  (
            .in0(N__83035),
            .in1(N__91225),
            .in2(N__83020),
            .in3(N__82996),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11646_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11575_LC_23_9_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11575_LC_23_9_5 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11575_LC_23_9_5 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11575_LC_23_9_5  (
            .in0(N__90302),
            .in1(N__85821),
            .in2(N__82975),
            .in3(N__82972),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i62_63_LC_23_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i62_63_LC_23_9_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i62_63_LC_23_9_6 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i62_63_LC_23_9_6  (
            .in0(N__82704),
            .in1(N__95105),
            .in2(N__89529),
            .in3(N__82926),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93442),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Bit_Index_i2_LC_23_10_0 .C_ON=1'b0;
    defparam \pc_tx.r_Bit_Index_i2_LC_23_10_0 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Bit_Index_i2_LC_23_10_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \pc_tx.r_Bit_Index_i2_LC_23_10_0  (
            .in0(N__83458),
            .in1(N__83476),
            .in2(_gnd_net_),
            .in3(N__83515),
            .lcout(\pc_tx.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97424),
            .ce(N__82686),
            .sr(N__83710));
    defparam \pc_tx.r_Bit_Index_i1_LC_23_10_1 .C_ON=1'b0;
    defparam \pc_tx.r_Bit_Index_i1_LC_23_10_1 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Bit_Index_i1_LC_23_10_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pc_tx.r_Bit_Index_i1_LC_23_10_1  (
            .in0(N__83514),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83457),
            .lcout(\pc_tx.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97424),
            .ce(N__82686),
            .sr(N__83710));
    defparam \pc_tx.i2_2_lut_LC_23_11_0 .C_ON=1'b0;
    defparam \pc_tx.i2_2_lut_LC_23_11_0 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i2_2_lut_LC_23_11_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pc_tx.i2_2_lut_LC_23_11_0  (
            .in0(_gnd_net_),
            .in1(N__97468),
            .in2(_gnd_net_),
            .in3(N__97486),
            .lcout(\pc_tx.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.i1_3_lut_LC_23_11_1 .C_ON=1'b0;
    defparam \pc_tx.i1_3_lut_LC_23_11_1 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i1_3_lut_LC_23_11_1 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \pc_tx.i1_3_lut_LC_23_11_1  (
            .in0(N__97579),
            .in1(N__89734),
            .in2(_gnd_net_),
            .in3(N__89749),
            .lcout(),
            .ltout(\pc_tx.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.i1_4_lut_LC_23_11_2 .C_ON=1'b0;
    defparam \pc_tx.i1_4_lut_LC_23_11_2 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i1_4_lut_LC_23_11_2 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \pc_tx.i1_4_lut_LC_23_11_2  (
            .in0(N__97564),
            .in1(N__97516),
            .in2(N__83698),
            .in3(N__97549),
            .lcout(\pc_tx.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.i5_4_lut_LC_23_11_3 .C_ON=1'b0;
    defparam \pc_tx.i5_4_lut_LC_23_11_3 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i5_4_lut_LC_23_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pc_tx.i5_4_lut_LC_23_11_3  (
            .in0(N__83695),
            .in1(N__97501),
            .in2(N__97534),
            .in3(N__83689),
            .lcout(r_SM_Main_2_N_808_1),
            .ltout(r_SM_Main_2_N_808_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_SM_Main_i0_LC_23_11_4 .C_ON=1'b0;
    defparam \pc_tx.r_SM_Main_i0_LC_23_11_4 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_SM_Main_i0_LC_23_11_4 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \pc_tx.r_SM_Main_i0_LC_23_11_4  (
            .in0(N__83683),
            .in1(_gnd_net_),
            .in2(N__83677),
            .in3(N__83651),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97403),
            .ce(),
            .sr(N__83914));
    defparam \pc_tx.r_SM_Main_i1_LC_23_11_5 .C_ON=1'b0;
    defparam \pc_tx.r_SM_Main_i1_LC_23_11_5 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_SM_Main_i1_LC_23_11_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \pc_tx.r_SM_Main_i1_LC_23_11_5  (
            .in0(N__83556),
            .in1(N__83652),
            .in2(_gnd_net_),
            .in3(N__83598),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97403),
            .ce(),
            .sr(N__83914));
    defparam \pc_tx.i6427_2_lut_4_lut_LC_23_11_6 .C_ON=1'b0;
    defparam \pc_tx.i6427_2_lut_4_lut_LC_23_11_6 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i6427_2_lut_4_lut_LC_23_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pc_tx.i6427_2_lut_4_lut_LC_23_11_6  (
            .in0(N__83456),
            .in1(N__83517),
            .in2(N__83484),
            .in3(N__83555),
            .lcout(\pc_tx.r_SM_Main_2_N_805_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.i2_2_lut_3_lut_LC_23_11_7 .C_ON=1'b0;
    defparam \pc_tx.i2_2_lut_3_lut_LC_23_11_7 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i2_2_lut_3_lut_LC_23_11_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pc_tx.i2_2_lut_3_lut_LC_23_11_7  (
            .in0(N__83516),
            .in1(N__83477),
            .in2(_gnd_net_),
            .in3(N__83455),
            .lcout(n11319),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_i0_LC_23_12_0 .C_ON=1'b0;
    defparam \timing_controller_inst.state_i0_LC_23_12_0 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_i0_LC_23_12_0 .LUT_INIT=16'b1111110001011100;
    LogicCell40 \timing_controller_inst.state_i0_LC_23_12_0  (
            .in0(N__84130),
            .in1(N__84124),
            .in2(N__84111),
            .in3(N__83959),
            .lcout(state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97425),
            .ce(N__83926),
            .sr(_gnd_net_));
    defparam \pc_tx.i1_1_lut_LC_23_12_1 .C_ON=1'b0;
    defparam \pc_tx.i1_1_lut_LC_23_12_1 .SEQ_MODE=4'b0000;
    defparam \pc_tx.i1_1_lut_LC_23_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pc_tx.i1_1_lut_LC_23_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83913),
            .lcout(\pc_tx.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_DEBUG_6_c_c_THRU_LUT4_0_LC_23_12_3.C_ON=1'b0;
    defparam GB_BUFFER_DEBUG_6_c_c_THRU_LUT4_0_LC_23_12_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_DEBUG_6_c_c_THRU_LUT4_0_LC_23_12_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_DEBUG_6_c_c_THRU_LUT4_0_LC_23_12_3 (
            .in0(N__93460),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_DEBUG_6_c_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_SLM_CLK_c_THRU_LUT4_0_LC_23_12_4.C_ON=1'b0;
    defparam GB_BUFFER_SLM_CLK_c_THRU_LUT4_0_LC_23_12_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_SLM_CLK_c_THRU_LUT4_0_LC_23_12_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_SLM_CLK_c_THRU_LUT4_0_LC_23_12_4 (
            .in0(N__97456),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_SLM_CLK_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_23_12_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_23_12_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_23_12_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_23_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.sub_31_add_2_2_lut_LC_23_13_0 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_2_lut_LC_23_13_0 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_2_lut_LC_23_13_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \timing_controller_inst.sub_31_add_2_2_lut_LC_23_13_0  (
            .in0(N__83784),
            .in1(N__83847),
            .in2(_gnd_net_),
            .in3(N__83818),
            .lcout(\timing_controller_inst.n12532 ),
            .ltout(),
            .carryin(bfn_23_13_0_),
            .carryout(\timing_controller_inst.n10588 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.sub_31_add_2_3_lut_LC_23_13_1 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_3_lut_LC_23_13_1 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_3_lut_LC_23_13_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_3_lut_LC_23_13_1  (
            .in0(N__84668),
            .in1(N__86215),
            .in2(N__83811),
            .in3(N__83788),
            .lcout(\timing_controller_inst.n12554 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10588 ),
            .carryout(\timing_controller_inst.n10589 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.sub_31_add_2_4_lut_LC_23_13_2 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_4_lut_LC_23_13_2 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_4_lut_LC_23_13_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \timing_controller_inst.sub_31_add_2_4_lut_LC_23_13_2  (
            .in0(N__83785),
            .in1(N__83757),
            .in2(N__86361),
            .in3(N__83740),
            .lcout(\timing_controller_inst.n12553 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10589 ),
            .carryout(\timing_controller_inst.n10590 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.sub_31_add_2_5_lut_LC_23_13_3 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_5_lut_LC_23_13_3 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_5_lut_LC_23_13_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_5_lut_LC_23_13_3  (
            .in0(N__84669),
            .in1(N__86219),
            .in2(N__83733),
            .in3(N__84304),
            .lcout(\timing_controller_inst.n12552 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10590 ),
            .carryout(\timing_controller_inst.n10591 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.sub_31_add_2_6_lut_LC_23_13_4 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_6_lut_LC_23_13_4 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_6_lut_LC_23_13_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_6_lut_LC_23_13_4  (
            .in0(N__84670),
            .in1(N__84301),
            .in2(N__86362),
            .in3(N__84277),
            .lcout(\timing_controller_inst.n12604 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10591 ),
            .carryout(\timing_controller_inst.n10592 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.sub_31_add_2_7_lut_LC_23_13_5 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_7_lut_LC_23_13_5 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_7_lut_LC_23_13_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_7_lut_LC_23_13_5  (
            .in0(N__84274),
            .in1(N__86223),
            .in2(N__84268),
            .in3(N__84247),
            .lcout(\timing_controller_inst.n12555 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10592 ),
            .carryout(\timing_controller_inst.n10593 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i6_LC_23_13_6 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i6_LC_23_13_6 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i6_LC_23_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i6_LC_23_13_6  (
            .in0(_gnd_net_),
            .in1(N__84243),
            .in2(N__86360),
            .in3(N__84232),
            .lcout(\timing_controller_inst.state_timeout_counter_6 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10593 ),
            .carryout(\timing_controller_inst.n10594 ),
            .clk(N__97431),
            .ce(N__86054),
            .sr(N__85981));
    defparam \timing_controller_inst.state_timeout_counter_i0_i7_LC_23_13_7 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i7_LC_23_13_7 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i7_LC_23_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i7_LC_23_13_7  (
            .in0(_gnd_net_),
            .in1(N__86214),
            .in2(N__84228),
            .in3(N__84211),
            .lcout(\timing_controller_inst.state_timeout_counter_7 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10594 ),
            .carryout(\timing_controller_inst.n10595 ),
            .clk(N__97431),
            .ce(N__86054),
            .sr(N__85981));
    defparam \timing_controller_inst.state_timeout_counter_i0_i8_LC_23_14_0 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i8_LC_23_14_0 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i8_LC_23_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i8_LC_23_14_0  (
            .in0(_gnd_net_),
            .in1(N__84204),
            .in2(N__86367),
            .in3(N__84193),
            .lcout(\timing_controller_inst.state_timeout_counter_8 ),
            .ltout(),
            .carryin(bfn_23_14_0_),
            .carryout(\timing_controller_inst.n10596 ),
            .clk(N__97439),
            .ce(N__86043),
            .sr(N__85982));
    defparam \timing_controller_inst.sub_31_add_2_11_lut_LC_23_14_1 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_11_lut_LC_23_14_1 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_11_lut_LC_23_14_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_11_lut_LC_23_14_1  (
            .in0(N__84671),
            .in1(N__84190),
            .in2(N__86365),
            .in3(N__84172),
            .lcout(\timing_controller_inst.n12551 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10596 ),
            .carryout(\timing_controller_inst.n10597 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.sub_31_add_2_12_lut_LC_23_14_2 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_12_lut_LC_23_14_2 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_12_lut_LC_23_14_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_12_lut_LC_23_14_2  (
            .in0(N__84673),
            .in1(N__84168),
            .in2(N__86368),
            .in3(N__84148),
            .lcout(\timing_controller_inst.n12550 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10597 ),
            .carryout(\timing_controller_inst.n10598 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i11_LC_23_14_3 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i11_LC_23_14_3 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i11_LC_23_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i11_LC_23_14_3  (
            .in0(_gnd_net_),
            .in1(N__84141),
            .in2(N__86363),
            .in3(N__84547),
            .lcout(\timing_controller_inst.state_timeout_counter_11 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10598 ),
            .carryout(\timing_controller_inst.n10599 ),
            .clk(N__97439),
            .ce(N__86043),
            .sr(N__85982));
    defparam \timing_controller_inst.sub_31_add_2_14_lut_LC_23_14_4 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_14_lut_LC_23_14_4 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_14_lut_LC_23_14_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_14_lut_LC_23_14_4  (
            .in0(N__84674),
            .in1(N__84543),
            .in2(N__86369),
            .in3(N__84514),
            .lcout(\timing_controller_inst.n12549 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10599 ),
            .carryout(\timing_controller_inst.n10600 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i13_LC_23_14_5 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i13_LC_23_14_5 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i13_LC_23_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i13_LC_23_14_5  (
            .in0(_gnd_net_),
            .in1(N__84501),
            .in2(N__86364),
            .in3(N__84490),
            .lcout(\timing_controller_inst.state_timeout_counter_13 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10600 ),
            .carryout(\timing_controller_inst.n10601 ),
            .clk(N__97439),
            .ce(N__86043),
            .sr(N__85982));
    defparam \timing_controller_inst.sub_31_add_2_16_lut_LC_23_14_6 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_16_lut_LC_23_14_6 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_16_lut_LC_23_14_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_16_lut_LC_23_14_6  (
            .in0(N__84675),
            .in1(N__84487),
            .in2(N__86370),
            .in3(N__84457),
            .lcout(\timing_controller_inst.n12548 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10601 ),
            .carryout(\timing_controller_inst.n10602 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.sub_31_add_2_17_lut_LC_23_14_7 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_17_lut_LC_23_14_7 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_17_lut_LC_23_14_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_17_lut_LC_23_14_7  (
            .in0(N__84672),
            .in1(N__84454),
            .in2(N__86366),
            .in3(N__84418),
            .lcout(\timing_controller_inst.n12547 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10602 ),
            .carryout(\timing_controller_inst.n10603 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i16_LC_23_15_0 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i16_LC_23_15_0 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i16_LC_23_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i16_LC_23_15_0  (
            .in0(_gnd_net_),
            .in1(N__84405),
            .in2(N__86371),
            .in3(N__84394),
            .lcout(\timing_controller_inst.state_timeout_counter_16 ),
            .ltout(),
            .carryin(bfn_23_15_0_),
            .carryout(\timing_controller_inst.n10604 ),
            .clk(N__97443),
            .ce(N__86055),
            .sr(N__85984));
    defparam \timing_controller_inst.state_timeout_counter_i0_i17_LC_23_15_1 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i17_LC_23_15_1 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i17_LC_23_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i17_LC_23_15_1  (
            .in0(_gnd_net_),
            .in1(N__84390),
            .in2(N__86375),
            .in3(N__84379),
            .lcout(\timing_controller_inst.state_timeout_counter_17 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10604 ),
            .carryout(\timing_controller_inst.n10605 ),
            .clk(N__97443),
            .ce(N__86055),
            .sr(N__85984));
    defparam \timing_controller_inst.sub_31_add_2_20_lut_LC_23_15_2 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_20_lut_LC_23_15_2 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_20_lut_LC_23_15_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_20_lut_LC_23_15_2  (
            .in0(N__84694),
            .in1(N__84376),
            .in2(N__86372),
            .in3(N__84343),
            .lcout(\timing_controller_inst.n12545 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10605 ),
            .carryout(\timing_controller_inst.n10606 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.sub_31_add_2_21_lut_LC_23_15_3 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_21_lut_LC_23_15_3 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_21_lut_LC_23_15_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_21_lut_LC_23_15_3  (
            .in0(N__84697),
            .in1(N__86254),
            .in2(N__84340),
            .in3(N__84820),
            .lcout(\timing_controller_inst.n12544 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10606 ),
            .carryout(\timing_controller_inst.n10607 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.sub_31_add_2_22_lut_LC_23_15_4 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_22_lut_LC_23_15_4 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_22_lut_LC_23_15_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_22_lut_LC_23_15_4  (
            .in0(N__84695),
            .in1(N__84817),
            .in2(N__86373),
            .in3(N__84781),
            .lcout(\timing_controller_inst.n12542 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10607 ),
            .carryout(\timing_controller_inst.n10608 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i21_LC_23_15_5 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i21_LC_23_15_5 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i21_LC_23_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i21_LC_23_15_5  (
            .in0(_gnd_net_),
            .in1(N__84774),
            .in2(N__86376),
            .in3(N__84763),
            .lcout(\timing_controller_inst.state_timeout_counter_21 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10608 ),
            .carryout(\timing_controller_inst.n10609 ),
            .clk(N__97443),
            .ce(N__86055),
            .sr(N__85984));
    defparam \timing_controller_inst.sub_31_add_2_24_lut_LC_23_15_6 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_24_lut_LC_23_15_6 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_24_lut_LC_23_15_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_24_lut_LC_23_15_6  (
            .in0(N__84696),
            .in1(N__84760),
            .in2(N__86374),
            .in3(N__84742),
            .lcout(\timing_controller_inst.n12541 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10609 ),
            .carryout(\timing_controller_inst.n10610 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.sub_31_add_2_25_lut_LC_23_15_7 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_25_lut_LC_23_15_7 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_25_lut_LC_23_15_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_25_lut_LC_23_15_7  (
            .in0(N__84698),
            .in1(N__84732),
            .in2(N__86377),
            .in3(N__84715),
            .lcout(\timing_controller_inst.n12540 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10610 ),
            .carryout(\timing_controller_inst.n10611 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.sub_31_add_2_26_lut_LC_23_16_0 .C_ON=1'b1;
    defparam \timing_controller_inst.sub_31_add_2_26_lut_LC_23_16_0 .SEQ_MODE=4'b0000;
    defparam \timing_controller_inst.sub_31_add_2_26_lut_LC_23_16_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \timing_controller_inst.sub_31_add_2_26_lut_LC_23_16_0  (
            .in0(N__84705),
            .in1(N__84619),
            .in2(N__86509),
            .in3(N__84601),
            .lcout(\timing_controller_inst.n12539 ),
            .ltout(),
            .carryin(bfn_23_16_0_),
            .carryout(\timing_controller_inst.n10612 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \timing_controller_inst.state_timeout_counter_i0_i25_LC_23_16_1 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i25_LC_23_16_1 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i25_LC_23_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i25_LC_23_16_1  (
            .in0(_gnd_net_),
            .in1(N__84597),
            .in2(N__86506),
            .in3(N__84586),
            .lcout(\timing_controller_inst.state_timeout_counter_25 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10612 ),
            .carryout(\timing_controller_inst.n10613 ),
            .clk(N__97447),
            .ce(N__86044),
            .sr(N__85983));
    defparam \timing_controller_inst.state_timeout_counter_i0_i26_LC_23_16_2 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i26_LC_23_16_2 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i26_LC_23_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i26_LC_23_16_2  (
            .in0(_gnd_net_),
            .in1(N__86381),
            .in2(N__84583),
            .in3(N__84568),
            .lcout(\timing_controller_inst.state_timeout_counter_26 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10613 ),
            .carryout(\timing_controller_inst.n10614 ),
            .clk(N__97447),
            .ce(N__86044),
            .sr(N__85983));
    defparam \timing_controller_inst.state_timeout_counter_i0_i27_LC_23_16_3 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i27_LC_23_16_3 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i27_LC_23_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i27_LC_23_16_3  (
            .in0(_gnd_net_),
            .in1(N__84558),
            .in2(N__86507),
            .in3(N__86746),
            .lcout(\timing_controller_inst.state_timeout_counter_27 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10614 ),
            .carryout(\timing_controller_inst.n10615 ),
            .clk(N__97447),
            .ce(N__86044),
            .sr(N__85983));
    defparam \timing_controller_inst.state_timeout_counter_i0_i28_LC_23_16_4 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i28_LC_23_16_4 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i28_LC_23_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i28_LC_23_16_4  (
            .in0(_gnd_net_),
            .in1(N__86385),
            .in2(N__86736),
            .in3(N__86719),
            .lcout(\timing_controller_inst.state_timeout_counter_28 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10615 ),
            .carryout(\timing_controller_inst.n10616 ),
            .clk(N__97447),
            .ce(N__86044),
            .sr(N__85983));
    defparam \timing_controller_inst.state_timeout_counter_i0_i29_LC_23_16_5 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i29_LC_23_16_5 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i29_LC_23_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i29_LC_23_16_5  (
            .in0(_gnd_net_),
            .in1(N__86709),
            .in2(N__86508),
            .in3(N__86698),
            .lcout(\timing_controller_inst.state_timeout_counter_29 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10616 ),
            .carryout(\timing_controller_inst.n10617 ),
            .clk(N__97447),
            .ce(N__86044),
            .sr(N__85983));
    defparam \timing_controller_inst.state_timeout_counter_i0_i30_LC_23_16_6 .C_ON=1'b1;
    defparam \timing_controller_inst.state_timeout_counter_i0_i30_LC_23_16_6 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i30_LC_23_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i30_LC_23_16_6  (
            .in0(_gnd_net_),
            .in1(N__86389),
            .in2(N__86688),
            .in3(N__86671),
            .lcout(\timing_controller_inst.state_timeout_counter_30 ),
            .ltout(),
            .carryin(\timing_controller_inst.n10617 ),
            .carryout(\timing_controller_inst.n10618 ),
            .clk(N__97447),
            .ce(N__86044),
            .sr(N__85983));
    defparam \timing_controller_inst.state_timeout_counter_i0_i31_LC_23_16_7 .C_ON=1'b0;
    defparam \timing_controller_inst.state_timeout_counter_i0_i31_LC_23_16_7 .SEQ_MODE=4'b1000;
    defparam \timing_controller_inst.state_timeout_counter_i0_i31_LC_23_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \timing_controller_inst.state_timeout_counter_i0_i31_LC_23_16_7  (
            .in0(N__86067),
            .in1(N__86390),
            .in2(_gnd_net_),
            .in3(N__86077),
            .lcout(\timing_controller_inst.state_timeout_counter_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97447),
            .ce(N__86044),
            .sr(N__85983));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11919_LC_24_7_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11919_LC_24_7_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11919_LC_24_7_0 .LUT_INIT=16'b1011110010110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11919_LC_24_7_0  (
            .in0(N__85942),
            .in1(N__92676),
            .in2(N__88911),
            .in3(N__85924),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13724_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13724_bdd_4_lut_LC_24_7_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13724_bdd_4_lut_LC_24_7_1 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13724_bdd_4_lut_LC_24_7_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13724_bdd_4_lut_LC_24_7_1  (
            .in0(N__92674),
            .in1(N__85903),
            .in2(N__85882),
            .in3(N__85879),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11811_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11425_LC_24_7_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11425_LC_24_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11425_LC_24_7_2 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_2__bdd_4_lut_11425_LC_24_7_2  (
            .in0(N__90352),
            .in1(N__85387),
            .in2(N__84847),
            .in3(N__89677),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11849_LC_24_7_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11849_LC_24_7_3 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11849_LC_24_7_3 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.rd_addr_r_0__bdd_4_lut_11849_LC_24_7_3  (
            .in0(N__92675),
            .in1(N__88901),
            .in2(N__88981),
            .in3(N__84844),
            .lcout(),
            .ltout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13640_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13640_bdd_4_lut_LC_24_7_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13640_bdd_4_lut_LC_24_7_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13640_bdd_4_lut_LC_24_7_4 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13640_bdd_4_lut_LC_24_7_4  (
            .in0(N__89719),
            .in1(N__92673),
            .in2(N__89704),
            .in3(N__89701),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11820 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i713_714_LC_24_7_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i713_714_LC_24_7_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i713_714_LC_24_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i713_714_LC_24_7_5  (
            .in0(N__89541),
            .in1(N__96734),
            .in2(_gnd_net_),
            .in3(N__89662),
            .lcout(REG_mem_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93456),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4478_4479_LC_24_7_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4478_4479_LC_24_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4478_4479_LC_24_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i4478_4479_LC_24_7_7  (
            .in0(N__88977),
            .in1(N__89504),
            .in2(_gnd_net_),
            .in3(N__89128),
            .lcout(REG_mem_46_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93456),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10034_3_lut_LC_24_8_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10034_3_lut_LC_24_8_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10034_3_lut_LC_24_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10034_3_lut_LC_24_8_0  (
            .in0(N__88935),
            .in1(N__88947),
            .in2(_gnd_net_),
            .in3(N__88770),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11683 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2345_2346_LC_24_8_1 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2345_2346_LC_24_8_1 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2345_2346_LC_24_8_1 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2345_2346_LC_24_8_1  (
            .in0(N__96735),
            .in1(N__95980),
            .in2(N__88948),
            .in3(N__95460),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93454),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2441_2442_LC_24_8_2 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2441_2442_LC_24_8_2 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2441_2442_LC_24_8_2 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2441_2442_LC_24_8_2  (
            .in0(N__95459),
            .in1(N__96736),
            .in2(N__88936),
            .in3(N__97054),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_25_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93454),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5417_5418_LC_24_8_3 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5417_5418_LC_24_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5417_5418_LC_24_8_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5417_5418_LC_24_8_3  (
            .in0(N__96737),
            .in1(N__95981),
            .in2(N__88924),
            .in3(N__95461),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93454),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10076_3_lut_LC_24_8_4 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10076_3_lut_LC_24_8_4 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10076_3_lut_LC_24_8_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i10076_3_lut_LC_24_8_4  (
            .in0(N__96429),
            .in1(N__88923),
            .in2(_gnd_net_),
            .in3(N__88771),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11725 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5513_5514_LC_24_8_5 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5513_5514_LC_24_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5513_5514_LC_24_8_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5513_5514_LC_24_8_5  (
            .in0(N__97053),
            .in1(N__96738),
            .in2(N__96430),
            .in3(N__95463),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_57_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93454),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2360_2361_LC_24_8_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2360_2361_LC_24_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2360_2361_LC_24_8_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i2360_2361_LC_24_8_6  (
            .in0(N__95458),
            .in1(N__96323),
            .in2(N__96408),
            .in3(N__95983),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_24_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93454),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5432_5433_LC_24_8_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5432_5433_LC_24_8_7 .SEQ_MODE=4'b1000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5432_5433_LC_24_8_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.i5432_5433_LC_24_8_7  (
            .in0(N__96322),
            .in1(N__95982),
            .in2(N__93477),
            .in3(N__95462),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.REG_mem_56_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__93454),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13130_bdd_4_lut_LC_24_9_0 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13130_bdd_4_lut_LC_24_9_0 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13130_bdd_4_lut_LC_24_9_0 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13130_bdd_4_lut_LC_24_9_0  (
            .in0(N__90351),
            .in1(N__92740),
            .in2(N__92728),
            .in3(N__92716),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11901 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14012_bdd_4_lut_LC_24_9_6 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14012_bdd_4_lut_LC_24_9_6 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14012_bdd_4_lut_LC_24_9_6 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n14012_bdd_4_lut_LC_24_9_6  (
            .in0(N__92695),
            .in1(N__91228),
            .in2(N__90460),
            .in3(N__90442),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11736 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13304_bdd_4_lut_LC_24_10_7 .C_ON=1'b0;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13304_bdd_4_lut_LC_24_10_7 .SEQ_MODE=4'b0000;
    defparam \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13304_bdd_4_lut_LC_24_10_7 .LUT_INIT=16'b1011101010011000;
    LogicCell40 \fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n13304_bdd_4_lut_LC_24_10_7  (
            .in0(N__90406),
            .in1(N__90398),
            .in2(N__89776),
            .in3(N__89767),
            .lcout(\fifo_dc_32_lut_gen_inst.lscc_fifo_dc_inst.n11880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc_tx.r_Clock_Count_1113__i0_LC_24_11_0 .C_ON=1'b1;
    defparam \pc_tx.r_Clock_Count_1113__i0_LC_24_11_0 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Clock_Count_1113__i0_LC_24_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_tx.r_Clock_Count_1113__i0_LC_24_11_0  (
            .in0(_gnd_net_),
            .in1(N__89748),
            .in2(_gnd_net_),
            .in3(N__89737),
            .lcout(\pc_tx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(bfn_24_11_0_),
            .carryout(\pc_tx.n10712 ),
            .clk(N__97413),
            .ce(N__97110),
            .sr(N__97077));
    defparam \pc_tx.r_Clock_Count_1113__i1_LC_24_11_1 .C_ON=1'b1;
    defparam \pc_tx.r_Clock_Count_1113__i1_LC_24_11_1 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Clock_Count_1113__i1_LC_24_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_tx.r_Clock_Count_1113__i1_LC_24_11_1  (
            .in0(_gnd_net_),
            .in1(N__89733),
            .in2(_gnd_net_),
            .in3(N__89722),
            .lcout(\pc_tx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\pc_tx.n10712 ),
            .carryout(\pc_tx.n10713 ),
            .clk(N__97413),
            .ce(N__97110),
            .sr(N__97077));
    defparam \pc_tx.r_Clock_Count_1113__i2_LC_24_11_2 .C_ON=1'b1;
    defparam \pc_tx.r_Clock_Count_1113__i2_LC_24_11_2 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Clock_Count_1113__i2_LC_24_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_tx.r_Clock_Count_1113__i2_LC_24_11_2  (
            .in0(_gnd_net_),
            .in1(N__97578),
            .in2(_gnd_net_),
            .in3(N__97567),
            .lcout(\pc_tx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\pc_tx.n10713 ),
            .carryout(\pc_tx.n10714 ),
            .clk(N__97413),
            .ce(N__97110),
            .sr(N__97077));
    defparam \pc_tx.r_Clock_Count_1113__i3_LC_24_11_3 .C_ON=1'b1;
    defparam \pc_tx.r_Clock_Count_1113__i3_LC_24_11_3 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Clock_Count_1113__i3_LC_24_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_tx.r_Clock_Count_1113__i3_LC_24_11_3  (
            .in0(_gnd_net_),
            .in1(N__97563),
            .in2(_gnd_net_),
            .in3(N__97552),
            .lcout(\pc_tx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\pc_tx.n10714 ),
            .carryout(\pc_tx.n10715 ),
            .clk(N__97413),
            .ce(N__97110),
            .sr(N__97077));
    defparam \pc_tx.r_Clock_Count_1113__i4_LC_24_11_4 .C_ON=1'b1;
    defparam \pc_tx.r_Clock_Count_1113__i4_LC_24_11_4 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Clock_Count_1113__i4_LC_24_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_tx.r_Clock_Count_1113__i4_LC_24_11_4  (
            .in0(_gnd_net_),
            .in1(N__97548),
            .in2(_gnd_net_),
            .in3(N__97537),
            .lcout(\pc_tx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\pc_tx.n10715 ),
            .carryout(\pc_tx.n10716 ),
            .clk(N__97413),
            .ce(N__97110),
            .sr(N__97077));
    defparam \pc_tx.r_Clock_Count_1113__i5_LC_24_11_5 .C_ON=1'b1;
    defparam \pc_tx.r_Clock_Count_1113__i5_LC_24_11_5 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Clock_Count_1113__i5_LC_24_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_tx.r_Clock_Count_1113__i5_LC_24_11_5  (
            .in0(_gnd_net_),
            .in1(N__97530),
            .in2(_gnd_net_),
            .in3(N__97519),
            .lcout(\pc_tx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\pc_tx.n10716 ),
            .carryout(\pc_tx.n10717 ),
            .clk(N__97413),
            .ce(N__97110),
            .sr(N__97077));
    defparam \pc_tx.r_Clock_Count_1113__i6_LC_24_11_6 .C_ON=1'b1;
    defparam \pc_tx.r_Clock_Count_1113__i6_LC_24_11_6 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Clock_Count_1113__i6_LC_24_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_tx.r_Clock_Count_1113__i6_LC_24_11_6  (
            .in0(_gnd_net_),
            .in1(N__97515),
            .in2(_gnd_net_),
            .in3(N__97504),
            .lcout(\pc_tx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\pc_tx.n10717 ),
            .carryout(\pc_tx.n10718 ),
            .clk(N__97413),
            .ce(N__97110),
            .sr(N__97077));
    defparam \pc_tx.r_Clock_Count_1113__i7_LC_24_11_7 .C_ON=1'b1;
    defparam \pc_tx.r_Clock_Count_1113__i7_LC_24_11_7 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Clock_Count_1113__i7_LC_24_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_tx.r_Clock_Count_1113__i7_LC_24_11_7  (
            .in0(_gnd_net_),
            .in1(N__97500),
            .in2(_gnd_net_),
            .in3(N__97489),
            .lcout(\pc_tx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(\pc_tx.n10718 ),
            .carryout(\pc_tx.n10719 ),
            .clk(N__97413),
            .ce(N__97110),
            .sr(N__97077));
    defparam \pc_tx.r_Clock_Count_1113__i8_LC_24_12_0 .C_ON=1'b1;
    defparam \pc_tx.r_Clock_Count_1113__i8_LC_24_12_0 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Clock_Count_1113__i8_LC_24_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pc_tx.r_Clock_Count_1113__i8_LC_24_12_0  (
            .in0(_gnd_net_),
            .in1(N__97485),
            .in2(_gnd_net_),
            .in3(N__97474),
            .lcout(\pc_tx.r_Clock_Count_8 ),
            .ltout(),
            .carryin(bfn_24_12_0_),
            .carryout(\pc_tx.n10720 ),
            .clk(N__97432),
            .ce(N__97098),
            .sr(N__97084));
    defparam \pc_tx.r_Clock_Count_1113__i9_LC_24_12_1 .C_ON=1'b0;
    defparam \pc_tx.r_Clock_Count_1113__i9_LC_24_12_1 .SEQ_MODE=4'b1000;
    defparam \pc_tx.r_Clock_Count_1113__i9_LC_24_12_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pc_tx.r_Clock_Count_1113__i9_LC_24_12_1  (
            .in0(N__97467),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__97471),
            .lcout(\pc_tx.r_Clock_Count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97432),
            .ce(N__97098),
            .sr(N__97084));
endmodule // top

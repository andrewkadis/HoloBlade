
module unsaved (
	clk_clk,
	reset_reset_n,
	rs232_0_clk_clk);	

	input		clk_clk;
	input		reset_reset_n;
	input		rs232_0_clk_clk;
endmodule

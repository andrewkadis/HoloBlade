// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Mon Jun 15 23:03:04 2020
//
// Verilog Description of module top
//

module top (ICE_SYSCLK, DCD, DSR, DTR, CTS, RST, UART_RX, UART_TX, 
            SEN, SCK, SOUT, SDAT, UPDATE, RESET, SLM_CLK, INVERT, 
            SYNC, VALID, DATA31, DATA0, DATA30, DATA29, DATA1, 
            DATA28, DATA27, DATA2, DATA26, DATA25, DATA3, DATA24, 
            DATA23, DATA4, DATA22, DATA21, DATA5, DATA20, DATA19, 
            DATA6, DATA18, DATA17, DATA7, DATA16, DATA15, DATA8, 
            DATA14, DATA13, DATA12, DATA11, DATA9, DATA10, FT_OE, 
            FT_RD, FT_WR, FT_SIWU, FR_RXF, FT_TXE, FIFO_BE3, FIFO_BE2, 
            FIFO_BE1, FIFO_BE0, FIFO_D31, FIFO_D30, FIFO_D29, FIFO_D28, 
            FIFO_D27, FIFO_CLK, FIFO_D26, FIFO_D25, FIFO_D24, FIFO_D23, 
            FIFO_D22, FIFO_D21, FIFO_D20, FIFO_D19, FIFO_D18, FIFO_D17, 
            FIFO_D16, FIFO_D15, FIFO_D14, FIFO_D13, FIFO_D12, FIFO_D11, 
            FIFO_D10, FIFO_D9, FIFO_D8, FIFO_D7, FIFO_D6, FIFO_D5, 
            FIFO_D4, FIFO_D3, FIFO_D2, FIFO_D1, FIFO_D0, DEBUG_0, 
            DEBUG_1, DEBUG_2, DEBUG_3, DEBUG_5, DEBUG_6, DEBUG_8, 
            DEBUG_9, ICE_CLK, ICE_CDONE, ICE_CREST) /* synthesis syn_module_defined=1 */ ;   // src/top.v(5[8:11])
    input ICE_SYSCLK;   // src/top.v(8[11:21])
    output DCD;   // src/top.v(11[12:15])
    output DSR;   // src/top.v(12[12:15])
    output DTR;   // src/top.v(13[12:15])
    output CTS;   // src/top.v(14[12:15])
    output RST;   // src/top.v(15[12:15])
    input UART_RX;   // src/top.v(16[12:19])
    output UART_TX;   // src/top.v(17[12:19])
    output SEN;   // src/top.v(20[12:15])
    output SCK;   // src/top.v(21[12:15])
    input SOUT;   // src/top.v(22[12:16])
    output SDAT;   // src/top.v(23[12:16])
    output UPDATE;   // src/top.v(27[12:18])
    output RESET;   // src/top.v(28[12:17])
    output SLM_CLK;   // src/top.v(29[12:19])
    output INVERT;   // src/top.v(30[12:18])
    output SYNC;   // src/top.v(31[12:16])
    output VALID;   // src/top.v(32[12:17])
    output DATA31;   // src/top.v(34[12:18])
    output DATA0;   // src/top.v(35[12:17])
    output DATA30;   // src/top.v(36[12:18])
    output DATA29;   // src/top.v(37[12:18])
    output DATA1;   // src/top.v(38[12:17])
    output DATA28;   // src/top.v(39[12:18])
    output DATA27;   // src/top.v(40[12:18])
    output DATA2;   // src/top.v(41[12:17])
    output DATA26;   // src/top.v(42[12:18])
    output DATA25;   // src/top.v(43[12:18])
    output DATA3;   // src/top.v(44[12:17])
    output DATA24;   // src/top.v(45[12:18])
    output DATA23;   // src/top.v(46[12:18])
    output DATA4;   // src/top.v(47[12:17])
    output DATA22;   // src/top.v(48[12:18])
    output DATA21;   // src/top.v(49[12:18])
    output DATA5;   // src/top.v(50[12:17])
    output DATA20;   // src/top.v(51[12:18])
    output DATA19;   // src/top.v(52[12:18])
    output DATA6;   // src/top.v(53[12:17])
    output DATA18;   // src/top.v(54[12:18])
    output DATA17;   // src/top.v(55[12:18])
    output DATA7;   // src/top.v(56[12:17])
    output DATA16;   // src/top.v(57[12:18])
    output DATA15;   // src/top.v(58[12:18])
    output DATA8;   // src/top.v(59[12:17])
    output DATA14;   // src/top.v(60[12:18])
    output DATA13;   // src/top.v(61[12:18])
    output DATA12;   // src/top.v(62[12:18])
    output DATA11;   // src/top.v(63[12:18])
    output DATA9;   // src/top.v(64[12:17])
    output DATA10;   // src/top.v(65[12:18])
    output FT_OE;   // src/top.v(69[12:17])
    output FT_RD;   // src/top.v(70[12:17])
    output FT_WR;   // src/top.v(71[12:17])
    output FT_SIWU;   // src/top.v(72[12:19])
    input FR_RXF;   // src/top.v(73[12:18])
    input FT_TXE;   // src/top.v(74[12:18])
    input FIFO_BE3;   // src/top.v(75[12:20])
    input FIFO_BE2;   // src/top.v(76[12:20])
    input FIFO_BE1;   // src/top.v(77[12:20])
    input FIFO_BE0;   // src/top.v(78[12:20])
    input FIFO_D31;   // src/top.v(79[12:20])
    input FIFO_D30;   // src/top.v(80[12:20])
    input FIFO_D29;   // src/top.v(81[12:20])
    input FIFO_D28;   // src/top.v(82[12:20])
    input FIFO_D27;   // src/top.v(83[12:20])
    input FIFO_CLK;   // src/top.v(84[12:20])
    input FIFO_D26;   // src/top.v(85[12:20])
    input FIFO_D25;   // src/top.v(86[12:20])
    input FIFO_D24;   // src/top.v(87[12:20])
    input FIFO_D23;   // src/top.v(88[12:20])
    input FIFO_D22;   // src/top.v(89[12:20])
    input FIFO_D21;   // src/top.v(90[12:20])
    input FIFO_D20;   // src/top.v(91[12:20])
    input FIFO_D19;   // src/top.v(92[12:20])
    input FIFO_D18;   // src/top.v(93[12:20])
    input FIFO_D17;   // src/top.v(94[12:20])
    input FIFO_D16;   // src/top.v(95[12:20])
    input FIFO_D15;   // src/top.v(97[11:19])
    input FIFO_D14;   // src/top.v(98[11:19])
    input FIFO_D13;   // src/top.v(99[11:19])
    input FIFO_D12;   // src/top.v(100[11:19])
    input FIFO_D11;   // src/top.v(101[11:19])
    input FIFO_D10;   // src/top.v(102[11:19])
    input FIFO_D9;   // src/top.v(103[11:18])
    input FIFO_D8;   // src/top.v(104[11:18])
    input FIFO_D7;   // src/top.v(105[11:18])
    input FIFO_D6;   // src/top.v(106[11:18])
    input FIFO_D5;   // src/top.v(107[11:18])
    input FIFO_D4;   // src/top.v(108[11:18])
    input FIFO_D3;   // src/top.v(109[11:18])
    input FIFO_D2;   // src/top.v(110[11:18])
    input FIFO_D1;   // src/top.v(111[11:18])
    input FIFO_D0;   // src/top.v(112[11:18])
    output DEBUG_0;   // src/top.v(115[12:19])
    output DEBUG_1;   // src/top.v(116[12:19])
    output DEBUG_2;   // src/top.v(117[12:19])
    output DEBUG_3;   // src/top.v(118[12:19])
    output DEBUG_5;   // src/top.v(119[12:19])
    output DEBUG_6;   // src/top.v(120[12:19])
    output DEBUG_8;   // src/top.v(121[12:19])
    output DEBUG_9;   // src/top.v(122[12:19])
    output ICE_CLK;   // src/top.v(125[12:19])
    output ICE_CDONE;   // src/top.v(126[12:21])
    output ICE_CREST;   // src/top.v(127[12:21])
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire DEBUG_6_c_c /* synthesis is_clock=1, SET_AS_NETWORK=DEBUG_6_c_c */ ;   // src/top.v(84[12:20])
    
    wire GND_net, VCC_net, ICE_SYSCLK_c, UART_RX_c, UART_TX_c, SEN_c_1, 
        SCK_c_0, SOUT_c, SDAT_c_15, UPDATE_c_3, RESET_c, INVERT_c_4, 
        SYNC_c, VALID_c, DATA15_c, DATA16_c, DATA14_c, DATA13_c, 
        DATA17_c, DATA12_c, DATA11_c, DATA18_c, DATA10_c, DATA9_c, 
        DATA19_c, DATA8_c, DATA7_c, DATA20_c, DATA6_c, DATA5_c, 
        FT_OE_c, DEBUG_3_c, DEBUG_2_c_c, FIFO_D15_c_15, FIFO_D14_c_14, 
        FIFO_D13_c_13, FIFO_D12_c_12, FIFO_D11_c_11, FIFO_D10_c_10, 
        FIFO_D9_c_9, FIFO_D8_c_8, FIFO_D7_c_7, FIFO_D6_c_6, FIFO_D5_c_5, 
        FIFO_D4_c_4, FIFO_D3_c_3, FIFO_D2_c_2, FIFO_D1_c_1, DEBUG_1_c_0_c, 
        DEBUG_0_c_24, DEBUG_5_c, DEBUG_9_c, debug_led3, reset_all_w;
    wire [3:0]reset_clk_counter;   // src/top.v(242[10:27])
    
    wire reset_all, reset_per_frame, buffer_switch_done, \REG.mem_14_1 , 
        \REG.mem_14_0 , \REG.mem_11_0 , n11424, \REG.mem_12_15 , \REG.mem_12_14 , 
        \REG.mem_12_13 , \REG.mem_12_12 , \REG.mem_12_11 , \REG.mem_12_10 , 
        \REG.mem_12_9 ;
    wire [31:0]dc32_fifo_data_in;   // src/top.v(500[13:30])
    
    wire dc32_fifo_almost_empty, get_next_word, \REG.mem_9_3 , \REG.mem_9_2 , 
        \REG.mem_9_1 , \REG.mem_9_0 ;
    wire [31:0]fifo_data_out;   // src/top.v(535[12:25])
    wire [7:0]pc_data_rx;   // src/top.v(675[11:21])
    
    wire tx_uart_active_flag, spi_start_transfer_r, multi_byte_spi_trans_flag_r;
    wire [7:0]tx_addr_byte;   // src/top.v(797[11:23])
    wire [7:0]tx_data_byte;   // src/top.v(799[11:23])
    wire [7:0]rx_buf_byte;   // src/top.v(806[11:22])
    
    wire is_tx_fifo_full_flag, fifo_write_cmd, spi_rx_byte_ready, fifo_read_cmd, 
        is_fifo_empty_flag;
    wire [31:0]fifo_temp_output;   // src/top.v(896[12:28])
    
    wire even_byte_flag, uart_rx_complete_rising_edge, uart_rx_complete_prev;
    wire [3:0]state;   // src/timing_controller.v(48[11:16])
    
    wire reset_all_w_N_61, start_tx_N_64, pll_clk_unbuf, n718, multi_byte_spi_trans_flag_r_N_72, 
        \REG.mem_8_15 , \REG.mem_8_14 , \REG.mem_8_13 , \REG.mem_8_12 , 
        \REG.mem_8_11 , \REG.mem_8_10 , \REG.mem_8_9 , \REG.mem_8_8 , 
        \REG.mem_8_7 , \REG.mem_8_6 , \REG.mem_8_5 , \REG.mem_8_4 , 
        n11376, \REG.mem_18_15 , \REG.mem_18_14 , \REG.mem_18_13 , \REG.mem_18_12 , 
        \REG.mem_18_11 , \REG.mem_18_10 , \REG.mem_18_9 , \REG.mem_18_8 , 
        \REG.mem_18_7 , \REG.mem_18_6 , \REG.mem_18_5 , \REG.mem_18_4 , 
        \REG.mem_18_3 , \REG.mem_18_2 , \REG.mem_18_1 , \REG.mem_18_0 , 
        \REG.mem_17_15 , \REG.mem_17_14 , \REG.mem_17_13 , \REG.mem_17_12 , 
        \REG.mem_17_11 , \REG.mem_17_10 , \REG.mem_17_9 , \REG.mem_17_8 , 
        \REG.mem_17_7 , \REG.mem_17_6 , \REG.mem_17_5 , \REG.mem_17_4 , 
        \REG.mem_17_3 , \REG.mem_17_2 , \REG.mem_17_1 , \REG.mem_17_0 , 
        n7383, \REG.mem_16_15 , \REG.mem_16_14 , \REG.mem_16_13 , \REG.mem_16_12 , 
        \REG.mem_16_11 , \REG.mem_16_10 , \REG.mem_16_9 , \REG.mem_16_8 , 
        \REG.mem_16_7 , \REG.mem_16_6 , \REG.mem_16_5 , \REG.mem_16_4 , 
        \REG.mem_16_3 , \REG.mem_16_2 , \REG.mem_16_1 , \REG.mem_16_0 , 
        \REG.mem_15_15 , \REG.mem_15_14 , \REG.mem_15_13 , \REG.mem_15_12 , 
        \REG.mem_15_11 , \REG.mem_15_10 , \REG.mem_15_9 , \REG.mem_15_8 , 
        \REG.mem_15_7 , \REG.mem_15_6 , \REG.mem_15_5 , \REG.mem_15_4 , 
        \REG.mem_15_3 , \REG.mem_15_2 , \REG.mem_15_1 , \REG.mem_15_0 , 
        \REG.mem_14_15 , \REG.mem_14_14 , \REG.mem_14_13 , \REG.mem_14_12 , 
        \REG.mem_14_11 , \REG.mem_14_10 , \REG.mem_14_9 , \REG.mem_14_8 , 
        \REG.mem_14_7 , \REG.mem_14_6 , \REG.mem_14_5 , \REG.mem_14_4 , 
        \REG.mem_8_3 , \REG.mem_8_2 , \REG.mem_8_1 , \REG.mem_8_0 , 
        \REG.mem_7_15 , \REG.mem_7_14 , \REG.mem_7_13 , \REG.mem_7_12 , 
        \REG.mem_7_11 , \REG.mem_7_10 , \REG.mem_7_9 , \REG.mem_7_8 , 
        \REG.mem_7_7 , \REG.mem_7_6 , \REG.mem_7_5 , \REG.mem_7_4 , 
        \REG.mem_14_3 , n1876, buffer_switch_done_latched, \REG.mem_11_15 , 
        \REG.mem_11_14 , \REG.mem_14_2 , n4002, \REG.mem_10_1 , \REG.mem_11_2 , 
        \REG.mem_11_1 , n4724, \REG.mem_7_3 , \REG.mem_7_2 , \REG.mem_7_1 , 
        \REG.mem_7_0 , \REG.mem_10_0 ;
    wire [7:0]state_timeout_counter_adj_1218;   // src/bluejay_data.v(52[11:32])
    
    wire n11089, \REG.mem_12_7 , \REG.mem_12_8 , \REG.mem_11_7 , \REG.mem_11_6 , 
        \REG.mem_11_5 , \REG.mem_11_4 , \REG.mem_11_3 , \REG.mem_12_5 , 
        n4703, n4700, n4697, bluejay_data_out_31__N_703, bluejay_data_out_31__N_704, 
        n11412, r_Rx_Data, \REG.mem_10_9 , \REG.mem_10_8 , \REG.mem_10_7 , 
        \REG.mem_10_6 , \REG.mem_10_5 , \REG.mem_10_4 , n4686, \REG.mem_12_6 , 
        \REG.mem_12_4 , \REG.mem_12_3 , n4679;
    wire [2:0]r_SM_Main_adj_1225;   // src/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_1227;   // src/uart_tx.v(33[16:27])
    wire [7:0]r_Tx_Data;   // src/uart_tx.v(34[16:25])
    wire [2:0]r_SM_Main_2__N_811;
    
    wire n11410;
    wire [2:0]r_SM_Main_2__N_808;
    
    wire \REG.mem_13_15 , n7596, \REG.mem_12_2 , \REG.mem_12_1 , \REG.mem_13_14 , 
        \REG.mem_9_15 , n4443, \REG.mem_9_14 , \REG.mem_9_13 , \REG.mem_9_12 ;
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    wire [15:0]rx_shift_reg;   // src/spi.v(72[12:24])
    
    wire \REG.mem_13_13 , \REG.mem_13_12 , \REG.mem_9_11 , \REG.mem_9_10 , 
        \REG.mem_9_9 , \REG.mem_9_8 , \REG.mem_9_7 , \REG.mem_9_6 , 
        \REG.mem_9_5 , \REG.mem_9_4 , n2207, \REG.mem_11_11 , \REG.mem_11_10 , 
        \REG.mem_11_9 , \REG.mem_11_8 , \REG.mem_13_11 , \REG.mem_10_3 , 
        \REG.mem_10_2 , n4674, n4670, \REG.mem_6_15 , \REG.mem_6_14 , 
        \REG.mem_6_13 , \REG.mem_6_12 , \REG.mem_6_11 , \REG.mem_6_10 , 
        \REG.mem_6_9 , \REG.mem_6_8 , n4249, \REG.mem_12_0 , \REG.mem_11_12 , 
        \REG.mem_11_13 , \REG.mem_6_7 , \REG.mem_6_6 , \REG.mem_6_5 , 
        \REG.mem_6_4 , \REG.mem_6_3 , \REG.mem_6_2 , \REG.mem_6_1 , 
        \REG.mem_6_0 ;
    wire [6:0]wr_addr_r;   // src/fifo_dc_32_lut_gen.v(196[29:38])
    wire [6:0]wr_addr_nxt_c;   // src/fifo_dc_32_lut_gen.v(198[29:42])
    wire [6:0]wr_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(200[30:42])
    wire [6:0]rp_sync1_r;   // src/fifo_dc_32_lut_gen.v(201[37:47])
    wire [6:0]wr_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(204[37:51])
    wire [6:0]rd_addr_r;   // src/fifo_dc_32_lut_gen.v(217[29:38])
    wire [6:0]wp_sync1_r;   // src/fifo_dc_32_lut_gen.v(222[37:47])
    wire [6:0]rd_grey_sync_r;   // src/fifo_dc_32_lut_gen.v(225[37:51])
    wire [6:0]rd_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(233[30:44])
    
    wire \aempty_flag_impl.ae_flag_nxt_w , t_rd_fifo_en_w;
    wire [31:0]\REG.out_raw ;   // src/fifo_dc_32_lut_gen.v(879[47:54])
    wire [6:0]\afull_flag_impl.af_flag_p_w_N_603 ;
    wire [6:0]rd_addr_nxt_c_6__N_465;
    
    wire n4, n4667, \REG.mem_13_10 , \REG.mem_5_15 , \REG.mem_5_14 , 
        \REG.mem_5_13 , \REG.mem_5_12 , \REG.mem_5_11 , \REG.mem_5_10 , 
        \REG.mem_5_9 , \REG.mem_5_8 , \REG.mem_5_7 , \REG.mem_5_6 , 
        \REG.mem_5_5 , \REG.mem_5_4 , \REG.mem_5_3 , \REG.mem_5_2 , 
        \REG.mem_5_1 , \REG.mem_5_0 , n7566, n11319, \REG.mem_4_15 , 
        \REG.mem_4_14 , \REG.mem_4_13 , \REG.mem_4_12 , \REG.mem_4_11 , 
        \REG.mem_4_10 , \REG.mem_4_9 , \REG.mem_4_8 , \REG.mem_4_7 , 
        \REG.mem_4_6 , \REG.mem_4_5 , \REG.mem_4_4 , \REG.mem_4_3 , 
        \REG.mem_4_2 , \REG.mem_4_1 , \REG.mem_4_0 , rd_fifo_en_w;
    wire [2:0]wr_addr_r_adj_1249;   // src/fifo_quad_word_mod.v(65[31:40])
    wire [2:0]wr_addr_p1_w_adj_1251;   // src/fifo_quad_word_mod.v(67[32:44])
    wire [2:0]rd_addr_r_adj_1252;   // src/fifo_quad_word_mod.v(69[31:40])
    wire [2:0]rd_addr_p1_w_adj_1254;   // src/fifo_quad_word_mod.v(71[32:44])
    
    wire full_nxt_r, n7495;
    wire [31:0]\mem_LUT.data_raw_r ;   // src/fifo_quad_word_mod.v(449[42:52])
    
    wire empty_o_N_1116, n7455, n2679, n2766, n4654, n5905, n5902, 
        n5899, n4646, \REG.mem_10_10 , \REG.mem_10_11 , \REG.mem_10_12 , 
        n5896, n5893, n5890, n5887, n5884, n1928, n4644, n5881, 
        \REG.mem_19_15 , \REG.mem_13_9 , \REG.mem_13_8 , \REG.mem_13_7 , 
        \REG.mem_13_6 , \REG.mem_13_5 , \REG.mem_13_4 , \REG.mem_13_3 , 
        \REG.mem_13_2 , \REG.mem_13_1 , \REG.mem_13_0 , \REG.mem_10_15 , 
        \REG.mem_10_14 , \REG.mem_10_13 , \REG.mem_19_14 , \REG.mem_19_13 , 
        \REG.mem_19_12 , n1721, n1616, \REG.mem_19_11 , \REG.mem_19_10 , 
        \REG.mem_19_9 , \REG.mem_19_8 , \REG.mem_19_7 , \REG.mem_19_6 , 
        \REG.mem_19_5 , \REG.mem_19_4 , \REG.mem_19_3 , \REG.mem_19_2 , 
        \REG.mem_19_1 , \REG.mem_19_0 , \REG.mem_23_0 , \REG.mem_23_1 , 
        \REG.mem_23_2 , \REG.mem_23_3 , \REG.mem_23_4 , \REG.mem_23_5 , 
        \REG.mem_23_6 , \REG.mem_23_7 , \REG.mem_23_8 , \REG.mem_23_9 , 
        \REG.mem_23_10 , \REG.mem_23_11 , \REG.mem_23_12 , \REG.mem_23_13 , 
        \REG.mem_23_14 , \REG.mem_23_15 , n10681, n10680, \REG.mem_26_0 , 
        \REG.mem_26_1 , \REG.mem_26_2 , \REG.mem_26_3 , \REG.mem_26_4 , 
        \REG.mem_26_5 , \REG.mem_26_6 , \REG.mem_26_7 , \REG.mem_26_8 , 
        \REG.mem_26_9 , \REG.mem_26_10 , \REG.mem_26_11 , \REG.mem_26_12 , 
        \REG.mem_26_13 , \REG.mem_26_14 , \REG.mem_26_15 , n15, n11015, 
        n32, \REG.mem_31_0 , \REG.mem_31_1 , \REG.mem_31_2 , \REG.mem_31_3 , 
        \REG.mem_31_4 , \REG.mem_31_5 , \REG.mem_31_6 , \REG.mem_31_7 , 
        \REG.mem_31_8 , \REG.mem_31_9 , \REG.mem_31_10 , \REG.mem_31_11 , 
        \REG.mem_31_12 , \REG.mem_31_13 , \REG.mem_31_14 , \REG.mem_31_15 , 
        n11141, n24, n3929, \REG.mem_36_0 , \REG.mem_36_1 , \REG.mem_36_2 , 
        \REG.mem_36_3 , \REG.mem_36_4 , \REG.mem_36_5 , \REG.mem_36_6 , 
        \REG.mem_36_7 , \REG.mem_36_8 , \REG.mem_36_9 , \REG.mem_36_10 , 
        \REG.mem_36_11 , \REG.mem_36_12 , \REG.mem_36_13 , \REG.mem_36_14 , 
        \REG.mem_36_15 , n5870, \REG.mem_37_0 , \REG.mem_37_1 , \REG.mem_37_2 , 
        \REG.mem_37_3 , \REG.mem_37_4 , \REG.mem_37_5 , \REG.mem_37_6 , 
        \REG.mem_37_7 , \REG.mem_37_8 , \REG.mem_37_9 , \REG.mem_37_10 , 
        \REG.mem_37_11 , \REG.mem_37_12 , \REG.mem_37_13 , \REG.mem_37_14 , 
        \REG.mem_37_15 , n5869, n10679, \REG.mem_38_0 , \REG.mem_38_1 , 
        \REG.mem_38_2 , \REG.mem_38_3 , \REG.mem_38_4 , \REG.mem_38_5 , 
        \REG.mem_38_6 , \REG.mem_38_7 , \REG.mem_38_8 , \REG.mem_38_9 , 
        \REG.mem_38_10 , \REG.mem_38_11 , \REG.mem_38_12 , \REG.mem_38_13 , 
        \REG.mem_38_14 , \REG.mem_38_15 , \REG.mem_39_0 , \REG.mem_39_1 , 
        \REG.mem_39_2 , \REG.mem_39_3 , \REG.mem_39_4 , \REG.mem_39_5 , 
        \REG.mem_39_6 , \REG.mem_39_7 , \REG.mem_39_8 , \REG.mem_39_9 , 
        \REG.mem_39_10 , \REG.mem_39_11 , \REG.mem_39_12 , \REG.mem_39_13 , 
        \REG.mem_39_14 , \REG.mem_39_15 , \REG.mem_40_0 , \REG.mem_40_1 , 
        \REG.mem_40_2 , \REG.mem_40_3 , \REG.mem_40_4 , \REG.mem_40_5 , 
        \REG.mem_40_6 , \REG.mem_40_7 , \REG.mem_40_8 , \REG.mem_40_9 , 
        \REG.mem_40_10 , \REG.mem_40_11 , \REG.mem_40_12 , \REG.mem_40_13 , 
        \REG.mem_40_14 , \REG.mem_40_15 , \REG.mem_41_0 , \REG.mem_41_1 , 
        \REG.mem_41_2 , \REG.mem_41_3 , \REG.mem_41_4 , \REG.mem_41_5 , 
        \REG.mem_41_6 , \REG.mem_41_7 , \REG.mem_41_8 , \REG.mem_41_9 , 
        \REG.mem_41_10 , \REG.mem_41_11 , \REG.mem_41_12 , \REG.mem_41_13 , 
        \REG.mem_41_14 , \REG.mem_41_15 , \REG.mem_42_0 , \REG.mem_42_1 , 
        \REG.mem_42_2 , \REG.mem_42_3 , \REG.mem_42_4 , \REG.mem_42_5 , 
        \REG.mem_42_6 , \REG.mem_42_7 , \REG.mem_42_8 , \REG.mem_42_9 , 
        \REG.mem_42_10 , \REG.mem_42_11 , \REG.mem_42_12 , \REG.mem_42_13 , 
        \REG.mem_42_14 , \REG.mem_42_15 , n3204, \REG.mem_43_0 , \REG.mem_43_1 , 
        \REG.mem_43_2 , \REG.mem_43_3 , \REG.mem_43_4 , \REG.mem_43_5 , 
        \REG.mem_43_6 , \REG.mem_43_7 , \REG.mem_43_8 , \REG.mem_43_9 , 
        \REG.mem_43_10 , \REG.mem_43_11 , \REG.mem_43_12 , \REG.mem_43_13 , 
        \REG.mem_43_14 , \REG.mem_43_15 , \REG.mem_44_0 , \REG.mem_44_1 , 
        \REG.mem_44_2 , \REG.mem_44_3 , \REG.mem_44_4 , \REG.mem_44_5 , 
        \REG.mem_44_6 , \REG.mem_44_7 , \REG.mem_44_8 , \REG.mem_44_9 , 
        \REG.mem_44_10 , \REG.mem_44_11 , \REG.mem_44_12 , \REG.mem_44_13 , 
        \REG.mem_44_14 , \REG.mem_44_15 , \REG.mem_45_0 , \REG.mem_45_1 , 
        \REG.mem_45_2 , \REG.mem_45_3 , \REG.mem_45_4 , \REG.mem_45_5 , 
        \REG.mem_45_6 , \REG.mem_45_7 , \REG.mem_45_8 , \REG.mem_45_9 , 
        \REG.mem_45_10 , \REG.mem_45_11 , \REG.mem_45_12 , \REG.mem_45_13 , 
        \REG.mem_45_14 , \REG.mem_45_15 , \REG.mem_46_0 , \REG.mem_46_1 , 
        \REG.mem_46_2 , \REG.mem_46_3 , \REG.mem_46_4 , \REG.mem_46_5 , 
        \REG.mem_46_6 , \REG.mem_46_7 , \REG.mem_46_8 , \REG.mem_46_9 , 
        \REG.mem_46_10 , \REG.mem_46_11 , \REG.mem_46_12 , \REG.mem_46_13 , 
        \REG.mem_46_14 , \REG.mem_46_15 , n5861, \REG.mem_47_0 , \REG.mem_47_1 , 
        \REG.mem_47_2 , \REG.mem_47_3 , \REG.mem_47_4 , \REG.mem_47_5 , 
        \REG.mem_47_6 , \REG.mem_47_7 , \REG.mem_47_8 , \REG.mem_47_9 , 
        \REG.mem_47_10 , \REG.mem_47_11 , \REG.mem_47_12 , \REG.mem_47_13 , 
        \REG.mem_47_14 , \REG.mem_47_15 , \REG.mem_48_0 , \REG.mem_48_1 , 
        \REG.mem_48_2 , \REG.mem_48_3 , \REG.mem_48_4 , \REG.mem_48_5 , 
        \REG.mem_48_6 , \REG.mem_48_7 , \REG.mem_48_8 , \REG.mem_48_9 , 
        \REG.mem_48_10 , \REG.mem_48_11 , \REG.mem_48_12 , \REG.mem_48_13 , 
        \REG.mem_48_14 , \REG.mem_48_15 , n5858, \REG.mem_49_0 , \REG.mem_49_1 , 
        \REG.mem_49_2 , \REG.mem_49_3 , \REG.mem_49_4 , \REG.mem_49_5 , 
        \REG.mem_49_6 , \REG.mem_49_7 , \REG.mem_49_8 , \REG.mem_49_9 , 
        \REG.mem_49_10 , \REG.mem_49_11 , \REG.mem_49_12 , \REG.mem_49_13 , 
        \REG.mem_49_14 , \REG.mem_49_15 , n5857, n10921, \REG.mem_50_0 , 
        \REG.mem_50_1 , \REG.mem_50_2 , \REG.mem_50_3 , \REG.mem_50_4 , 
        \REG.mem_50_5 , \REG.mem_50_6 , \REG.mem_50_7 , \REG.mem_50_8 , 
        \REG.mem_50_9 , \REG.mem_50_10 , \REG.mem_50_11 , \REG.mem_50_12 , 
        \REG.mem_50_13 , \REG.mem_50_14 , \REG.mem_50_15 , n10678, n5854, 
        \REG.mem_51_0 , \REG.mem_51_1 , \REG.mem_51_2 , \REG.mem_51_3 , 
        \REG.mem_51_4 , \REG.mem_51_5 , \REG.mem_51_6 , \REG.mem_51_7 , 
        \REG.mem_51_8 , \REG.mem_51_9 , \REG.mem_51_10 , \REG.mem_51_11 , 
        \REG.mem_51_12 , \REG.mem_51_13 , \REG.mem_51_14 , \REG.mem_51_15 , 
        n4_adj_1182, n10677, n10676, \REG.mem_55_0 , \REG.mem_55_1 , 
        \REG.mem_55_2 , \REG.mem_55_3 , \REG.mem_55_4 , \REG.mem_55_5 , 
        \REG.mem_55_6 , \REG.mem_55_7 , \REG.mem_55_8 , \REG.mem_55_9 , 
        \REG.mem_55_10 , \REG.mem_55_11 , \REG.mem_55_12 , \REG.mem_55_13 , 
        \REG.mem_55_14 , \REG.mem_55_15 , \REG.mem_58_0 , \REG.mem_58_1 , 
        \REG.mem_58_2 , \REG.mem_58_3 , \REG.mem_58_4 , \REG.mem_58_5 , 
        \REG.mem_58_6 , \REG.mem_58_7 , \REG.mem_58_8 , \REG.mem_58_9 , 
        \REG.mem_58_10 , \REG.mem_58_11 , \REG.mem_58_12 , \REG.mem_58_13 , 
        \REG.mem_58_14 , \REG.mem_58_15 , n11324, n10727, n10847, 
        \REG.mem_63_0 , \REG.mem_63_1 , \REG.mem_63_2 , \REG.mem_63_3 , 
        \REG.mem_63_4 , \REG.mem_63_5 , \REG.mem_63_6 , \REG.mem_63_7 , 
        \REG.mem_63_8 , \REG.mem_63_9 , \REG.mem_63_10 , \REG.mem_63_11 , 
        \REG.mem_63_12 , \REG.mem_63_13 , \REG.mem_63_14 , \REG.mem_63_15 , 
        n7, n2, n7_adj_1183, n10, n14, n15_adj_1184, n16, n17, 
        n18, n19, n20, n21, n22, n23, n24_adj_1185, n25, n26, 
        n27, n28, n29, n34, n39, n42, n46, n47, n48, n49, 
        n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
        n60, n61, n11097, n11143, n11137, n5844, n5843, n5842, 
        n5841, n5840, n5839, n5838, n63, n5827, n5826, n5789, 
        n5788, n5787, n5786, n4_adj_1186, n5785, n5784, n5783, 
        n5782, n5781, n5780, n5779, n5778, n5777, n5776, n5775, 
        n11135, n5773, n5756, n5755, n5754, n5753, n5752, n5751, 
        n5750, n5733, n5732, n5731, n5730, n5729, n5728, n5727, 
        n11139, n5709, n5708, n5707, n5706, n3997, n5705, n5704, 
        n5686, n5685, n5684, n5683, n5682, n5681, n5680, n5679, 
        n5678, n5677, n5676, n5675, n5674, n5, n5673, n5672, 
        n5671, n5670, n5669, n5668, n5667, n5666, n5665, n5664, 
        n5662, n5660, n3514, n5626, n12601, n5625, n5624, n5623, 
        n5622, n5621, n5620, n5619, n5618, n5617, n5616, n5615, 
        n5614, n5613, n5612, n5610, n11007, n5609, n5608, n5607, 
        n5606, n5605, n5604, n5603, n5586, n5585, n5584, n5583, 
        n5582, n11073, n10675, n10674, n10673, n10672, n10671, 
        n5548, n5547, n5546, n10670, n10562, n5545, n5544, n5543, 
        n5542, n5541, n5540, n5539, n5538, n5537, n5536, n5535, 
        n5534, n5533, n5532, n5531, n5530, n4133, n5529, n5528, 
        n5527, n5526, n5525, n5524, n5523, n5522, n5521, n5520, 
        n5519, n5518, n5517, n5516, n5515, n5514, n5513, n5512, 
        n5511, n5510, n5509, n5508, n5507, n5506, n5505, n5504, 
        n5503, n5502, n5501, n5500, n5499, n5498, n5497, n5496, 
        n5495, n5494, n5492, n5491, n5490, n5489, n5488, n5487, 
        n5486, n5485, n5484, n5483, n5482, n5481, n5480, n5479, 
        n5478, n5477, n5476, n5474, n5472, n5471, n5470, n5469, 
        n5468, n5467, n5466, n5465, n5464, n5463, n5462, n5461, 
        n5460, n5459, n5458, n5457, n5456, n5455, n5454, n5453, 
        n5452, n5451, n5450, n5449, n5448, n5447, n5446, n5445, 
        n5444, n5443, n5442, n5441, n5440, n5439, n5438, n5437, 
        n5436, n5435, n5434, n5433, n5432, n5431, n5430, n5429, 
        n5428, n5427, n5426, n5425, n5424, n5423, n5422, n5421, 
        n5420, n5419, n5418, n5417, n5416, n5415, n5414, n5413, 
        n5412, n5411, n5410, n5409, n5408, n5407, n5406, n5405, 
        n5404, n5403, n5402, n5401, n5400, n5399, n5398, n5397, 
        n5396, n5395, n5394, n5393, n5392, n11071, n5390, n5389, 
        n5388, n5387, n5386, n5385, n5384, n5383, n5382, n5381, 
        n5380, n5379, n5378, n5377, n5376, n5375, n5374, n5373, 
        n5372, n5371, n5370, n10693, n5369, n5368, n5367, n5366, 
        n5365, n5364, n5363, n5362, n5361, n5360, n5358, n5357, 
        n5356, n5355, n5354, n10692, n5353, n5352, n5351, n5350, 
        n5349, n5348, n5347, n5346, n5345, n5344, n5343, n5342, 
        n5341, n5340, n5339, n5338, n10691, n5337, n5336, n5335, 
        n5334, n5333, n5332, n5331, n5330, n5329, n5328, n5327, 
        n5326, n5325, n5324, n5323, n5322, n10690, n5321, n5320, 
        n5319, n5318, n5317, n5316, n5315, n5314, n5313, n5312, 
        n5311, n5310, n5309, n5308, n5307, n5306, n5305, n5304, 
        n5303, n5302, n5301, n5300, n5299, n5298, n5297, n5296, 
        n5295, n5294, n5293, n5292, n5291, n5290, n5289, n5288, 
        n5286, n5285, n5284, n5283, n5282, n5281, n5280, n5279, 
        n5278, n5277, n5276, n5275, n5274, n5273, n5272, n5271, 
        n5270, n11069, n4639, n130, n129, n128, n127, n126, 
        n125, n124, n123, n122, n121, n120, n119, n118, n117, 
        n116, n115, n114, n113, n112, n111, n110, n109, n108, 
        n107, n106, n5202, n5201, n5200, n5199, n5198, n5197, 
        n5196, n5195, n5194, n10689, n5193, n5192, n5191, n5190, 
        n5189, n5188, n5187, n10688, n10687, n10686, n25_adj_1187, 
        n24_adj_1188, n23_adj_1189, n22_adj_1190, n21_adj_1191, n5121, 
        n5120, n5119, n5118, n5117, n5116, n5115, n5114, n5113, 
        n20_adj_1192, n19_adj_1193, n18_adj_1194, n17_adj_1195, n16_adj_1196, 
        n15_adj_1197, n14_adj_1198, n13, n12, n11, n10_adj_1199, 
        n9, n8, n7_adj_1200, n6, n5_adj_1201, n5112, n5111, n5110, 
        n5109, n5108, n5107, n5106, n4_adj_1202, n3, n2_adj_1203, 
        n25_adj_1204, n5073, n5072, n5071, n5070, n5069, n5068, 
        n5067, n5066, n5065, n5064, n5063, n5062, n5061, n5060, 
        n5059, n5058, n4638, n4637, n4632, n4631, n10685, n5006, 
        n5005, n5004, n5003, n5002, n5001, n5000, n4999, n4998, 
        n4997, n4996, n4995, n4994, n4993, n4992, n4991, n4990, 
        n4989, n4988, n4987, n4986, n4985, n4984, n4983, n4982, 
        n4981, n4980, n4979, n4978, n4977, n4976, n4975, n4974, 
        n4973, n4972, n4971, n4970, n4969, n4968, n4967, n4966, 
        n4965, n4964, n4963, n4962, n4961, n4960, n4958, n4957, 
        n4956, n4955, n4954, n4953, n4952, n4951, n4950, n4949, 
        n10684, n4948, n4947, n4946, n4945, n4944, n4943, n4942, 
        n4941, n4940, n4939, n4938, n4937, n4936, n4935, n4934, 
        n4933, n4932, n4931, n4930, n4929, n4928, n4927, n4926, 
        n4925, n4924, n4923, n4922, n4921, n4920, n4919, n4918, 
        n4917, n4916, n4915, n4914, n4913, n4912, n4911, n4910, 
        n4909, n4908, n4907, n10683, n4612, n4609, n4906, n4905, 
        n4904, n4903, n4902, n4901, n4900, n4899, n4898, n4897, 
        n4896, n4895, n4894, n4893, n4892, n4891, n10682, n4890, 
        n4889, n4888, n4887, n4886, n4885, n4884, n4883, n4882, 
        n4881, n4880, n4879, n4878, n4877, n4876, n4875, n4874, 
        n4873, n4872, n4871, n4870, n4869, n4868, n4867, n4866, 
        n4865, n4864, n4863, n4862, n4861, n4860, n4859, n4858, 
        n4857, n4856, n4855, n4854, n4853, n4852, n4851, n4850, 
        n4849, n4848, n4847, n4846, n4845, n4844, n4843, n4842, 
        n4841, n4840, n4839, n4838, n4837, n4836, n4835, n4834, 
        n4833, n4832, n4831, n4830, n4829, n4828, n4827, n4826, 
        n4825, n4824, n4823, n4822, n4821, n4820, n4819, n4818, 
        n4817, n4816, n4815, n4814, n4813, n4812, n4811, n4810, 
        n4809, n4808, n4807, n4806, n4805, n4804, n4803, n4802, 
        n4801, n4800, n4799, n4798, n4797, n4796, n4795, n4794, 
        n4793, n4792, n4791, n14424, n11133, n4790, n4789, n4788, 
        n4787, n4786, n4785, n4784, n4783, n11339, n4779, n4778, 
        n4777, n4776, n4775, n4774, n4773, n4772, n4771, n4093, 
        n4770, n4769, n4768, n4767, n4766, n4765, n4764, n4763, 
        n11119, n4762, n4761, n4760, n4759, n4758, n4757, n4756, 
        n4755, n11342, n4754, n4753, n4752, n4070, n4751, n4750, 
        n4749, n11471, n4748, n4_adj_1205, n4747, n4746, n4745, 
        n4744, n4743, n4742, n4740, n4_adj_1206, n10802, n10800, 
        n10798, n1, n3710, n14415, n11095;
    
    VCC i2 (.Y(VCC_net));
    timing_controller timing_controller_inst (.state({state}), .SLM_CLK_c(SLM_CLK_c), 
            .n1721(n1721), .GND_net(GND_net), .VCC_net(VCC_net), .n63(n63), 
            .n4(n4_adj_1182), .n11342(n11342), .reset_per_frame(reset_per_frame), 
            .n1616(n1616), .n7383(n7383), .INVERT_c_4(INVERT_c_4), .reset_all(reset_all), 
            .n7495(n7495), .buffer_switch_done(buffer_switch_done), .n11015(n11015), 
            .n3514(n3514), .n7566(n7566), .n11376(n11376), .UPDATE_c_3(UPDATE_c_3), 
            .n3929(n3929)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(442[19] 454[2])
    SB_LUT4 i4580_3_lut (.I0(\REG.mem_63_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n2), .I3(GND_net), .O(n5782));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4580_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF fifo_read_cmd_80 (.Q(fifo_read_cmd), .C(SLM_CLK_c), .D(start_tx_N_64));   // src/top.v(900[8] 918[4])
    SB_LUT4 i4581_3_lut (.I0(\REG.mem_63_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n2), .I3(GND_net), .O(n5783));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4581_3_lut.LUT_INIT = 16'hcaca;
    bluejay_data bluejay_data_inst (.VCC_net(VCC_net), .VALID_c(VALID_c), 
            .SLM_CLK_c(SLM_CLK_c), .\state_timeout_counter[3] (state_timeout_counter_adj_1218[3]), 
            .buffer_switch_done_latched(buffer_switch_done_latched), .bluejay_data_out_31__N_704(bluejay_data_out_31__N_704), 
            .n5870(n5870), .DATA16_c(DATA16_c), .DATA15_c(DATA15_c), .DATA14_c(DATA14_c), 
            .DATA13_c(DATA13_c), .DATA12_c(DATA12_c), .DATA11_c(DATA11_c), 
            .DATA10_c(DATA10_c), .DATA9_c(DATA9_c), .DATA8_c(DATA8_c), 
            .DATA7_c(DATA7_c), .n5827(n5827), .DATA6_c(DATA6_c), .n5826(n5826), 
            .DATA5_c(DATA5_c), .DATA20_c(DATA20_c), .DATA19_c(DATA19_c), 
            .DATA18_c(DATA18_c), .DATA17_c(DATA17_c), .GND_net(GND_net), 
            .SYNC_c(SYNC_c), .buffer_switch_done(buffer_switch_done), .bluejay_data_out_31__N_703(bluejay_data_out_31__N_703), 
            .n14424(n14424), .n718(n718), .n7(n7), .n5(n5), .\rd_sig_diff0_w[0] (rd_sig_diff0_w[0]), 
            .\rd_sig_diff0_w[1] (rd_sig_diff0_w[1]), .get_next_word(get_next_word), 
            .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .DEBUG_9_c(DEBUG_9_c), .dc32_fifo_almost_empty(dc32_fifo_almost_empty), 
            .DEBUG_5_c(DEBUG_5_c), .reset_all(reset_all), .n4667(n4667), 
            .\fifo_data_out[15] (fifo_data_out[15]), .\fifo_data_out[14] (fifo_data_out[14]), 
            .\fifo_data_out[13] (fifo_data_out[13]), .\fifo_data_out[12] (fifo_data_out[12]), 
            .\fifo_data_out[11] (fifo_data_out[11]), .\fifo_data_out[10] (fifo_data_out[10]), 
            .\fifo_data_out[9] (fifo_data_out[9]), .\fifo_data_out[8] (fifo_data_out[8]), 
            .\fifo_data_out[7] (fifo_data_out[7]), .\fifo_data_out[4] (fifo_data_out[4]), 
            .\fifo_data_out[3] (fifo_data_out[3]), .\fifo_data_out[2] (fifo_data_out[2]), 
            .\fifo_data_out[1] (fifo_data_out[1])) /* synthesis syn_module_defined=1 */ ;   // src/top.v(616[14] 629[2])
    SB_LUT4 i1_2_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_1204));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_GB clk_gb (.GLOBAL_BUFFER_OUTPUT(SLM_CLK_c), .USER_SIGNAL_TO_GLOBAL_BUFFER(pll_clk_unbuf)) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/clock.v(82[7:96])
    SB_DFF uart_rx_complete_prev_83 (.Q(uart_rx_complete_prev), .C(SLM_CLK_c), 
           .D(debug_led3));   // src/top.v(1055[8] 1061[4])
    SB_IO UART_TX_pad (.PACKAGE_PIN(UART_TX), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UART_TX_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_TX_pad.PIN_TYPE = 6'b011001;
    defparam UART_TX_pad.PULLUP = 1'b0;
    defparam UART_TX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_TX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4582_3_lut (.I0(\REG.mem_63_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n2), .I3(GND_net), .O(n5784));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4265_3_lut (.I0(\REG.mem_47_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n18), .I3(GND_net), .O(n5467));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4266_3_lut (.I0(\REG.mem_47_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n18), .I3(GND_net), .O(n5468));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4583_3_lut (.I0(\REG.mem_63_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n2), .I3(GND_net), .O(n5785));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4267_3_lut (.I0(\REG.mem_47_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n18), .I3(GND_net), .O(n5469));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4268_3_lut (.I0(\REG.mem_47_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n18), .I3(GND_net), .O(n5470));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4269_3_lut (.I0(\REG.mem_47_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n18), .I3(GND_net), .O(n5471));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3985_3_lut (.I0(\REG.mem_31_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n34), .I3(GND_net), .O(n5187));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4584_3_lut (.I0(\REG.mem_63_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n2), .I3(GND_net), .O(n5786));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3986_3_lut (.I0(\REG.mem_31_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n34), .I3(GND_net), .O(n5188));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3987_3_lut (.I0(\REG.mem_31_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n34), .I3(GND_net), .O(n5189));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4585_3_lut (.I0(\REG.mem_63_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n2), .I3(GND_net), .O(n5787));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4586_3_lut (.I0(\REG.mem_63_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n2), .I3(GND_net), .O(n5788));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3988_3_lut (.I0(\REG.mem_31_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n34), .I3(GND_net), .O(n5190));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4270_3_lut (.I0(\REG.mem_47_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n18), .I3(GND_net), .O(n5472));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3989_3_lut (.I0(\REG.mem_31_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n34), .I3(GND_net), .O(n5191));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3990_3_lut (.I0(\REG.mem_31_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n34), .I3(GND_net), .O(n5192));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3991_3_lut (.I0(\REG.mem_31_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n34), .I3(GND_net), .O(n5193));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3992_3_lut (.I0(\REG.mem_31_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n34), .I3(GND_net), .O(n5194));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3993_3_lut (.I0(\REG.mem_31_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n34), .I3(GND_net), .O(n5195));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3993_3_lut.LUT_INIT = 16'hcaca;
    SB_IO RST_pad (.PACKAGE_PIN(RST), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RST_pad.PIN_TYPE = 6'b011001;
    defparam RST_pad.PULLUP = 1'b0;
    defparam RST_pad.NEG_TRIGGER = 1'b0;
    defparam RST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i3994_3_lut (.I0(\REG.mem_31_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n34), .I3(GND_net), .O(n5196));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3995_3_lut (.I0(\REG.mem_31_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n34), .I3(GND_net), .O(n5197));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3996_3_lut (.I0(\REG.mem_31_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n34), .I3(GND_net), .O(n5198));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3997_3_lut (.I0(\REG.mem_31_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n34), .I3(GND_net), .O(n5199));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3998_3_lut (.I0(\REG.mem_31_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n34), .I3(GND_net), .O(n5200));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3999_3_lut (.I0(\REG.mem_31_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n34), .I3(GND_net), .O(n5201));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4000_3_lut (.I0(\REG.mem_31_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n34), .I3(GND_net), .O(n5202));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19_4_lut (.I0(n3514), .I1(n12601), .I2(state[3]), .I3(n4_adj_1182), 
            .O(n11015));   // src/timing_controller.v(53[8] 129[4])
    defparam i19_4_lut.LUT_INIT = 16'hfcac;
    SB_DFF reset_all_r_77 (.Q(reset_all_w), .C(SLM_CLK_c), .D(reset_all_w_N_61));   // src/top.v(246[8] 264[4])
    SB_LUT4 i4587_3_lut (.I0(\REG.mem_63_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n2), .I3(GND_net), .O(n5789));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4272_2_lut (.I0(reset_all), .I1(wr_addr_nxt_c[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5474));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4272_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4274_3_lut (.I0(\REG.mem_48_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n17), .I3(GND_net), .O(n5476));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4275_3_lut (.I0(\REG.mem_48_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n17), .I3(GND_net), .O(n5477));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4276_3_lut (.I0(\REG.mem_48_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n17), .I3(GND_net), .O(n5478));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4277_3_lut (.I0(\REG.mem_48_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n17), .I3(GND_net), .O(n5479));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4278_3_lut (.I0(\REG.mem_48_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n17), .I3(GND_net), .O(n5480));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4279_3_lut (.I0(\REG.mem_48_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n17), .I3(GND_net), .O(n5481));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4280_3_lut (.I0(\REG.mem_48_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n17), .I3(GND_net), .O(n5482));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4068_3_lut (.I0(\REG.mem_36_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n29), .I3(GND_net), .O(n5270));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4069_3_lut (.I0(\REG.mem_36_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n29), .I3(GND_net), .O(n5271));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4070_3_lut (.I0(\REG.mem_36_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n29), .I3(GND_net), .O(n5272));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4071_3_lut (.I0(\REG.mem_36_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n29), .I3(GND_net), .O(n5273));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4072_3_lut (.I0(\REG.mem_36_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n29), .I3(GND_net), .O(n5274));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4073_3_lut (.I0(\REG.mem_36_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n29), .I3(GND_net), .O(n5275));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4074_3_lut (.I0(\REG.mem_36_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n29), .I3(GND_net), .O(n5276));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4075_3_lut (.I0(\REG.mem_36_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n29), .I3(GND_net), .O(n5277));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4076_3_lut (.I0(\REG.mem_36_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n29), .I3(GND_net), .O(n5278));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4077_3_lut (.I0(\REG.mem_36_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n29), .I3(GND_net), .O(n5279));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4281_3_lut (.I0(\REG.mem_48_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n17), .I3(GND_net), .O(n5483));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4078_3_lut (.I0(\REG.mem_36_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n29), .I3(GND_net), .O(n5280));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4079_3_lut (.I0(\REG.mem_36_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n29), .I3(GND_net), .O(n5281));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4282_3_lut (.I0(\REG.mem_48_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n17), .I3(GND_net), .O(n5484));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4283_3_lut (.I0(\REG.mem_48_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n17), .I3(GND_net), .O(n5485));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4283_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_LUT4 i4284_3_lut (.I0(\REG.mem_48_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n17), .I3(GND_net), .O(n5486));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4285_3_lut (.I0(\REG.mem_48_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n17), .I3(GND_net), .O(n5487));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4080_3_lut (.I0(\REG.mem_36_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n29), .I3(GND_net), .O(n5282));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4286_3_lut (.I0(\REG.mem_48_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n17), .I3(GND_net), .O(n5488));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4081_3_lut (.I0(\REG.mem_36_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n29), .I3(GND_net), .O(n5283));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4287_3_lut (.I0(\REG.mem_48_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n17), .I3(GND_net), .O(n5489));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4288_3_lut (.I0(\REG.mem_48_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n17), .I3(GND_net), .O(n5490));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4082_3_lut (.I0(\REG.mem_36_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n29), .I3(GND_net), .O(n5284));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4289_2_lut (.I0(reset_all), .I1(wr_addr_nxt_c[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5491));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i4289_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4083_3_lut (.I0(\REG.mem_36_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n29), .I3(GND_net), .O(n5285));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4083_3_lut.LUT_INIT = 16'hcaca;
    SB_IO CTS_pad (.PACKAGE_PIN(CTS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CTS_pad.PIN_TYPE = 6'b011001;
    defparam CTS_pad.PULLUP = 1'b0;
    defparam CTS_pad.NEG_TRIGGER = 1'b0;
    defparam CTS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DTR_pad (.PACKAGE_PIN(DTR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DTR_pad.PIN_TYPE = 6'b011001;
    defparam DTR_pad.PULLUP = 1'b0;
    defparam DTR_pad.NEG_TRIGGER = 1'b0;
    defparam DTR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DSR_pad (.PACKAGE_PIN(DSR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DSR_pad.PIN_TYPE = 6'b011001;
    defparam DSR_pad.PULLUP = 1'b0;
    defparam DSR_pad.NEG_TRIGGER = 1'b0;
    defparam DSR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4084_3_lut (.I0(\REG.mem_37_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n28), .I3(GND_net), .O(n5286));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3472_4_lut (.I0(RESET_c), .I1(rd_addr_r_adj_1252[2]), .I2(rd_addr_p1_w_adj_1254[2]), 
            .I3(empty_o_N_1116), .O(n4674));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i3472_4_lut.LUT_INIT = 16'ha088;
    SB_IO DCD_pad (.PACKAGE_PIN(DCD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DCD_pad.PIN_TYPE = 6'b011001;
    defparam DCD_pad.PULLUP = 1'b0;
    defparam DCD_pad.NEG_TRIGGER = 1'b0;
    defparam DCD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4086_3_lut (.I0(\REG.mem_37_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n28), .I3(GND_net), .O(n5288));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4087_3_lut (.I0(\REG.mem_37_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n28), .I3(GND_net), .O(n5289));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4088_3_lut (.I0(\REG.mem_37_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n28), .I3(GND_net), .O(n5290));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4089_3_lut (.I0(\REG.mem_37_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n28), .I3(GND_net), .O(n5291));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4290_3_lut (.I0(\REG.mem_48_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n17), .I3(GND_net), .O(n5492));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4090_3_lut (.I0(\REG.mem_37_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n28), .I3(GND_net), .O(n5292));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4091_3_lut (.I0(\REG.mem_37_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n28), .I3(GND_net), .O(n5293));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4091_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DEBUG_1_c_0_pad (.PACKAGE_PIN(FIFO_D0), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(DEBUG_1_c_0_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_1_c_0_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_1_c_0_pad.PULLUP = 1'b0;
    defparam DEBUG_1_c_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_1_c_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4092_3_lut (.I0(\REG.mem_37_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n28), .I3(GND_net), .O(n5294));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4093_3_lut (.I0(\REG.mem_37_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n28), .I3(GND_net), .O(n5295));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4292_3_lut (.I0(tx_data_byte[7]), .I1(pc_data_rx[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5494));   // src/top.v(1064[8] 1131[4])
    defparam i4292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4293_3_lut (.I0(tx_data_byte[6]), .I1(pc_data_rx[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5495));   // src/top.v(1064[8] 1131[4])
    defparam i4293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4094_3_lut (.I0(\REG.mem_37_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n28), .I3(GND_net), .O(n5296));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4294_3_lut (.I0(tx_data_byte[5]), .I1(pc_data_rx[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5496));   // src/top.v(1064[8] 1131[4])
    defparam i4294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4095_3_lut (.I0(\REG.mem_37_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n28), .I3(GND_net), .O(n5297));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4096_3_lut (.I0(\REG.mem_37_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n28), .I3(GND_net), .O(n5298));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4295_3_lut (.I0(tx_data_byte[4]), .I1(pc_data_rx[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5497));   // src/top.v(1064[8] 1131[4])
    defparam i4295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4097_3_lut (.I0(\REG.mem_37_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n28), .I3(GND_net), .O(n5299));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4098_3_lut (.I0(\REG.mem_37_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n28), .I3(GND_net), .O(n5300));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4296_3_lut (.I0(tx_data_byte[3]), .I1(pc_data_rx[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5498));   // src/top.v(1064[8] 1131[4])
    defparam i4296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4099_3_lut (.I0(\REG.mem_37_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n28), .I3(GND_net), .O(n5301));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4100_3_lut (.I0(\REG.mem_37_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n28), .I3(GND_net), .O(n5302));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4101_3_lut (.I0(tx_addr_byte[7]), .I1(tx_data_byte[7]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5303));   // src/top.v(1064[8] 1131[4])
    defparam i4101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4297_3_lut (.I0(tx_data_byte[2]), .I1(pc_data_rx[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5499));   // src/top.v(1064[8] 1131[4])
    defparam i4297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4102_3_lut (.I0(tx_addr_byte[6]), .I1(tx_data_byte[6]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5304));   // src/top.v(1064[8] 1131[4])
    defparam i4102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4103_3_lut (.I0(tx_addr_byte[5]), .I1(tx_data_byte[5]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5305));   // src/top.v(1064[8] 1131[4])
    defparam i4103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4104_3_lut (.I0(tx_addr_byte[4]), .I1(tx_data_byte[4]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5306));   // src/top.v(1064[8] 1131[4])
    defparam i4104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4298_3_lut (.I0(tx_data_byte[1]), .I1(pc_data_rx[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5500));   // src/top.v(1064[8] 1131[4])
    defparam i4298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4105_3_lut (.I0(tx_addr_byte[3]), .I1(tx_data_byte[3]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5307));   // src/top.v(1064[8] 1131[4])
    defparam i4105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4299_3_lut (.I0(\REG.mem_49_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n16), .I3(GND_net), .O(n5501));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4106_3_lut (.I0(\REG.mem_38_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n27), .I3(GND_net), .O(n5308));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4300_3_lut (.I0(\REG.mem_49_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n16), .I3(GND_net), .O(n5502));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4107_3_lut (.I0(\REG.mem_38_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n27), .I3(GND_net), .O(n5309));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4301_3_lut (.I0(\REG.mem_49_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n16), .I3(GND_net), .O(n5503));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4301_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_1107__i3 (.Q(reset_clk_counter[3]), .C(SLM_CLK_c), 
           .D(n10802));   // src/top.v(259[27:51])
    SB_LUT4 i4302_3_lut (.I0(\REG.mem_49_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n16), .I3(GND_net), .O(n5504));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4303_3_lut (.I0(\REG.mem_49_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n16), .I3(GND_net), .O(n5505));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4304_3_lut (.I0(\REG.mem_49_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n16), .I3(GND_net), .O(n5506));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4305_3_lut (.I0(\REG.mem_49_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n16), .I3(GND_net), .O(n5507));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4108_3_lut (.I0(\REG.mem_38_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n27), .I3(GND_net), .O(n5310));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4109_3_lut (.I0(\REG.mem_38_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n27), .I3(GND_net), .O(n5311));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4109_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1106_1179__i0 (.Q(n25_adj_1187), .C(SLM_CLK_c), .D(n130));   // src/top.v(203[20:35])
    SB_DFF reset_clk_counter_i3_1107__i2 (.Q(reset_clk_counter[2]), .C(SLM_CLK_c), 
           .D(n10800));   // src/top.v(259[27:51])
    SB_LUT4 i4306_3_lut (.I0(\REG.mem_49_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n16), .I3(GND_net), .O(n5508));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4307_3_lut (.I0(\REG.mem_49_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n16), .I3(GND_net), .O(n5509));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4307_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_1107__i1 (.Q(reset_clk_counter[1]), .C(SLM_CLK_c), 
           .D(n10798));   // src/top.v(259[27:51])
    SB_DFF led_counter_1106_1179__i24 (.Q(DEBUG_0_c_24), .C(SLM_CLK_c), 
           .D(n106));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i23 (.Q(n2_adj_1203), .C(SLM_CLK_c), .D(n107));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i22 (.Q(n3), .C(SLM_CLK_c), .D(n108));   // src/top.v(203[20:35])
    SB_LUT4 i4308_3_lut (.I0(\REG.mem_49_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n16), .I3(GND_net), .O(n5510));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4308_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1106_1179__i21 (.Q(n4_adj_1202), .C(SLM_CLK_c), .D(n109));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i20 (.Q(n5_adj_1201), .C(SLM_CLK_c), .D(n110));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i19 (.Q(n6), .C(SLM_CLK_c), .D(n111));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i18 (.Q(n7_adj_1200), .C(SLM_CLK_c), .D(n112));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i17 (.Q(n8), .C(SLM_CLK_c), .D(n113));   // src/top.v(203[20:35])
    SB_LUT4 i4110_3_lut (.I0(\REG.mem_38_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n27), .I3(GND_net), .O(n5312));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4309_3_lut (.I0(\REG.mem_49_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n16), .I3(GND_net), .O(n5511));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4111_3_lut (.I0(\REG.mem_38_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n27), .I3(GND_net), .O(n5313));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4310_3_lut (.I0(\REG.mem_49_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n16), .I3(GND_net), .O(n5512));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4311_3_lut (.I0(\REG.mem_49_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n16), .I3(GND_net), .O(n5513));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4312_3_lut (.I0(\REG.mem_49_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n16), .I3(GND_net), .O(n5514));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 reset_all_w_I_0_1_lut (.I0(reset_all_w), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(RESET_c));   // src/top.v(295[16:28])
    defparam reset_all_w_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4313_3_lut (.I0(\REG.mem_49_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n16), .I3(GND_net), .O(n5515));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4313_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1106_1179__i16 (.Q(n9), .C(SLM_CLK_c), .D(n114));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i15 (.Q(n10_adj_1199), .C(SLM_CLK_c), 
           .D(n115));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i14 (.Q(n11), .C(SLM_CLK_c), .D(n116));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i13 (.Q(n12), .C(SLM_CLK_c), .D(n117));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i12 (.Q(n13), .C(SLM_CLK_c), .D(n118));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i11 (.Q(n14_adj_1198), .C(SLM_CLK_c), 
           .D(n119));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i10 (.Q(n15_adj_1197), .C(SLM_CLK_c), 
           .D(n120));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i9 (.Q(n16_adj_1196), .C(SLM_CLK_c), .D(n121));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i8 (.Q(n17_adj_1195), .C(SLM_CLK_c), .D(n122));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i7 (.Q(n18_adj_1194), .C(SLM_CLK_c), .D(n123));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i6 (.Q(n19_adj_1193), .C(SLM_CLK_c), .D(n124));   // src/top.v(203[20:35])
    SB_LUT4 i4112_3_lut (.I0(\REG.mem_38_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n27), .I3(GND_net), .O(n5314));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4112_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF led_counter_1106_1179__i5 (.Q(n20_adj_1192), .C(SLM_CLK_c), .D(n125));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i4 (.Q(n21_adj_1191), .C(SLM_CLK_c), .D(n126));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i3 (.Q(n22_adj_1190), .C(SLM_CLK_c), .D(n127));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i2 (.Q(n23_adj_1189), .C(SLM_CLK_c), .D(n128));   // src/top.v(203[20:35])
    SB_DFF led_counter_1106_1179__i1 (.Q(n24_adj_1188), .C(SLM_CLK_c), .D(n129));   // src/top.v(203[20:35])
    SB_LUT4 i4314_3_lut (.I0(\REG.mem_49_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n16), .I3(GND_net), .O(n5516));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4113_3_lut (.I0(\REG.mem_38_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n27), .I3(GND_net), .O(n5315));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4315_3_lut (.I0(\REG.mem_50_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5517));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4114_3_lut (.I0(\REG.mem_38_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n27), .I3(GND_net), .O(n5316));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4316_3_lut (.I0(\REG.mem_50_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5518));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4115_3_lut (.I0(\REG.mem_38_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n27), .I3(GND_net), .O(n5317));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4116_3_lut (.I0(\REG.mem_38_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n27), .I3(GND_net), .O(n5318));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4317_3_lut (.I0(\REG.mem_50_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5519));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4318_3_lut (.I0(\REG.mem_50_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5520));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4117_3_lut (.I0(\REG.mem_38_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n27), .I3(GND_net), .O(n5319));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4319_3_lut (.I0(\REG.mem_50_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5521));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4118_3_lut (.I0(\REG.mem_38_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n27), .I3(GND_net), .O(n5320));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4320_3_lut (.I0(\REG.mem_50_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5522));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4119_3_lut (.I0(\REG.mem_38_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n27), .I3(GND_net), .O(n5321));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4119_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF fifo_write_cmd_79 (.Q(fifo_write_cmd), .C(SLM_CLK_c), .D(n4703));   // src/top.v(879[8] 888[4])
    SB_LUT4 i4321_3_lut (.I0(\REG.mem_50_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5523));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4322_3_lut (.I0(\REG.mem_50_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5524));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4323_3_lut (.I0(\REG.mem_50_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5525));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4324_3_lut (.I0(\REG.mem_50_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5526));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4120_3_lut (.I0(\REG.mem_38_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n27), .I3(GND_net), .O(n5322));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4325_3_lut (.I0(\REG.mem_50_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5527));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4326_3_lut (.I0(\REG.mem_50_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5528));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4327_3_lut (.I0(\REG.mem_50_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5529));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4328_3_lut (.I0(\REG.mem_50_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5530));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4329_3_lut (.I0(\REG.mem_50_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5531));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4636_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[1]), .I2(n4_adj_1206), 
            .I3(n4002), .O(n5838));   // src/uart_rx.v(49[10] 144[8])
    defparam i4636_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4121_3_lut (.I0(\REG.mem_38_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n27), .I3(GND_net), .O(n5323));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4637_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[2]), .I2(n4), 
            .I3(n3997), .O(n5839));   // src/uart_rx.v(49[10] 144[8])
    defparam i4637_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4638_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[3]), .I2(n4), 
            .I3(n4002), .O(n5840));   // src/uart_rx.v(49[10] 144[8])
    defparam i4638_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4122_3_lut (.I0(tx_addr_byte[2]), .I1(tx_data_byte[2]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5324));   // src/top.v(1064[8] 1131[4])
    defparam i4122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4330_3_lut (.I0(\REG.mem_50_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n15_adj_1184), .I3(GND_net), .O(n5532));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4123_3_lut (.I0(tx_addr_byte[1]), .I1(tx_data_byte[1]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n5325));   // src/top.v(1064[8] 1131[4])
    defparam i4123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4331_3_lut (.I0(\REG.mem_51_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n14), .I3(GND_net), .O(n5533));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4124_3_lut (.I0(\REG.mem_39_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n26), .I3(GND_net), .O(n5326));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4332_3_lut (.I0(\REG.mem_51_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n14), .I3(GND_net), .O(n5534));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4639_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[4]), .I2(n4_adj_1205), 
            .I3(n3997), .O(n5841));   // src/uart_rx.v(49[10] 144[8])
    defparam i4639_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4125_3_lut (.I0(\REG.mem_39_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n26), .I3(GND_net), .O(n5327));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4640_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[5]), .I2(n4_adj_1205), 
            .I3(n4002), .O(n5842));   // src/uart_rx.v(49[10] 144[8])
    defparam i4640_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4333_3_lut (.I0(\REG.mem_51_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n14), .I3(GND_net), .O(n5535));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4126_3_lut (.I0(\REG.mem_39_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n26), .I3(GND_net), .O(n5328));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4641_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[6]), .I2(n7455), 
            .I3(n3997), .O(n5843));   // src/uart_rx.v(49[10] 144[8])
    defparam i4641_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i4334_3_lut (.I0(\REG.mem_51_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n14), .I3(GND_net), .O(n5536));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4642_4_lut (.I0(r_Rx_Data), .I1(pc_data_rx[7]), .I2(n7455), 
            .I3(n4002), .O(n5844));   // src/uart_rx.v(49[10] 144[8])
    defparam i4642_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1582_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n2766));   // src/top.v(1064[8] 1131[4])
    defparam i1582_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4335_3_lut (.I0(\REG.mem_51_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n14), .I3(GND_net), .O(n5537));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4127_3_lut (.I0(\REG.mem_39_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n26), .I3(GND_net), .O(n5329));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4336_3_lut (.I0(\REG.mem_51_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n14), .I3(GND_net), .O(n5538));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4128_3_lut (.I0(\REG.mem_39_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n26), .I3(GND_net), .O(n5330));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4337_3_lut (.I0(\REG.mem_51_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n14), .I3(GND_net), .O(n5539));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4338_3_lut (.I0(\REG.mem_51_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n14), .I3(GND_net), .O(n5540));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4129_3_lut (.I0(\REG.mem_39_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n26), .I3(GND_net), .O(n5331));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4339_3_lut (.I0(\REG.mem_51_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n14), .I3(GND_net), .O(n5541));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4130_3_lut (.I0(\REG.mem_39_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n26), .I3(GND_net), .O(n5332));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4131_3_lut (.I0(\REG.mem_39_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n26), .I3(GND_net), .O(n5333));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4132_3_lut (.I0(\REG.mem_39_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n26), .I3(GND_net), .O(n5334));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4340_3_lut (.I0(\REG.mem_51_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n14), .I3(GND_net), .O(n5542));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4341_3_lut (.I0(\REG.mem_51_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n14), .I3(GND_net), .O(n5543));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4133_3_lut (.I0(\REG.mem_39_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n26), .I3(GND_net), .O(n5335));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4342_3_lut (.I0(\REG.mem_51_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n14), .I3(GND_net), .O(n5544));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4343_3_lut (.I0(\REG.mem_51_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n14), .I3(GND_net), .O(n5545));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4134_3_lut (.I0(\REG.mem_39_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n26), .I3(GND_net), .O(n5336));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4135_3_lut (.I0(\REG.mem_39_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n26), .I3(GND_net), .O(n5337));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4344_3_lut (.I0(\REG.mem_51_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n14), .I3(GND_net), .O(n5546));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4345_3_lut (.I0(\REG.mem_51_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n14), .I3(GND_net), .O(n5547));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4136_3_lut (.I0(\REG.mem_39_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n26), .I3(GND_net), .O(n5338));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4655_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[0]), .I2(\mem_LUT.data_raw_r [0]), 
            .I3(n4249), .O(n5857));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4655_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4346_3_lut (.I0(\REG.mem_51_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n14), .I3(GND_net), .O(n5548));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(rd_addr_r_adj_1252[1]), .I1(rd_addr_r_adj_1252[0]), 
            .I2(wr_addr_r_adj_1249[1]), .I3(wr_addr_r_adj_1249[0]), .O(n32));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 i1_3_lut (.I0(is_fifo_empty_flag), .I1(fifo_write_cmd), .I2(n32), 
            .I3(GND_net), .O(n24));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i4659_4_lut (.I0(n4133), .I1(r_Bit_Index_adj_1227[0]), .I2(n11319), 
            .I3(r_SM_Main_adj_1225[1]), .O(n5861));   // src/uart_tx.v(38[10] 141[8])
    defparam i4659_4_lut.LUT_INIT = 16'h4644;
    SB_LUT4 i9762_4_lut (.I0(rd_addr_p1_w_adj_1254[2]), .I1(rd_addr_p1_w_adj_1254[1]), 
            .I2(wr_addr_r_adj_1249[2]), .I3(wr_addr_r_adj_1249[1]), .O(n11410));
    defparam i9762_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_91 (.I0(reset_all_w), .I1(n11410), .I2(n24), 
            .I3(n4_adj_1186), .O(n11324));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_91.LUT_INIT = 16'hfbfa;
    SB_LUT4 i4137_3_lut (.I0(\REG.mem_39_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n26), .I3(GND_net), .O(n5339));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4138_3_lut (.I0(\REG.mem_39_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n26), .I3(GND_net), .O(n5340));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4667_3_lut (.I0(pc_data_rx[0]), .I1(r_Rx_Data), .I2(n10847), 
            .I3(GND_net), .O(n5869));   // src/uart_rx.v(49[10] 144[8])
    defparam i4667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut (.I0(tx_shift_reg[0]), .I1(n1928), .I2(n4070), .I3(tx_data_byte[0]), 
            .O(n11007));   // src/spi.v(76[8] 221[4])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i4139_3_lut (.I0(\REG.mem_39_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n26), .I3(GND_net), .O(n5341));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4140_3_lut (.I0(\REG.mem_40_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n25), .I3(GND_net), .O(n5342));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4141_3_lut (.I0(\REG.mem_40_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n25), .I3(GND_net), .O(n5343));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4142_3_lut (.I0(\REG.mem_40_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n25), .I3(GND_net), .O(n5344));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4143_3_lut (.I0(\REG.mem_40_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n25), .I3(GND_net), .O(n5345));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4144_3_lut (.I0(\REG.mem_40_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n25), .I3(GND_net), .O(n5346));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4145_3_lut (.I0(\REG.mem_40_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n25), .I3(GND_net), .O(n5347));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4146_3_lut (.I0(\REG.mem_40_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n25), .I3(GND_net), .O(n5348));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4146_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF start_tx_81 (.Q(r_SM_Main_2__N_811[0]), .C(SLM_CLK_c), .D(n5858));   // src/top.v(900[8] 918[4])
    SB_LUT4 i4147_3_lut (.I0(\REG.mem_40_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n25), .I3(GND_net), .O(n5349));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4148_3_lut (.I0(\REG.mem_40_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n25), .I3(GND_net), .O(n5350));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4149_3_lut (.I0(\REG.mem_40_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n25), .I3(GND_net), .O(n5351));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4150_3_lut (.I0(\REG.mem_40_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n25), .I3(GND_net), .O(n5352));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4151_3_lut (.I0(\REG.mem_40_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n25), .I3(GND_net), .O(n5353));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4152_3_lut (.I0(\REG.mem_40_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n25), .I3(GND_net), .O(n5354));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4152_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF spi_start_transfer_r_84 (.Q(spi_start_transfer_r), .C(SLM_CLK_c), 
           .D(n2766));   // src/top.v(1064[8] 1131[4])
    SB_LUT4 i4153_3_lut (.I0(\REG.mem_40_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n25), .I3(GND_net), .O(n5355));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4154_3_lut (.I0(\REG.mem_40_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n25), .I3(GND_net), .O(n5356));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4155_3_lut (.I0(\REG.mem_40_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n25), .I3(GND_net), .O(n5357));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9776_4_lut (.I0(n1), .I1(fifo_read_cmd), .I2(wr_addr_r_adj_1249[1]), 
            .I3(rd_addr_r_adj_1252[1]), .O(n11424));
    defparam i9776_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i4156_3_lut (.I0(\REG.mem_41_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5358));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_92 (.I0(reset_all_w), .I1(n15), .I2(full_nxt_r), 
            .I3(n10727), .O(n10921));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_adj_92.LUT_INIT = 16'h5444;
    SB_LUT4 i4158_3_lut (.I0(\REG.mem_41_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5360));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4679_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[1]), .I2(\mem_LUT.data_raw_r [1]), 
            .I3(n4249), .O(n5881));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4679_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4159_3_lut (.I0(\REG.mem_41_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5361));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4160_3_lut (.I0(\REG.mem_41_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5362));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4682_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[2]), .I2(\mem_LUT.data_raw_r [2]), 
            .I3(n4249), .O(n5884));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4682_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4380_2_lut (.I0(reset_all), .I1(wp_sync1_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n5582));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4380_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4685_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[3]), .I2(\mem_LUT.data_raw_r [3]), 
            .I3(n4249), .O(n5887));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4685_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4161_3_lut (.I0(\REG.mem_41_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5363));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4162_3_lut (.I0(\REG.mem_41_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5364));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4163_3_lut (.I0(\REG.mem_41_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5365));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4164_3_lut (.I0(\REG.mem_41_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5366));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4688_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[4]), .I2(\mem_LUT.data_raw_r [4]), 
            .I3(n4249), .O(n5890));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4688_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i4381_2_lut (.I0(reset_all), .I1(wp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5583));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4381_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4382_2_lut (.I0(reset_all), .I1(wp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5584));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4382_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4165_3_lut (.I0(\REG.mem_41_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5367));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1106_1179_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(DEBUG_0_c_24), .I3(n10693), .O(n106)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4166_3_lut (.I0(\REG.mem_41_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5368));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4697_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[5]), .I2(\mem_LUT.data_raw_r [5]), 
            .I3(n4249), .O(n5899));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4697_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 led_counter_1106_1179_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n2_adj_1203), .I3(n10692), .O(n107)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1106_1179_add_4_25 (.CI(n10692), .I0(GND_net), 
            .I1(n2_adj_1203), .CO(n10693));
    SB_LUT4 led_counter_1106_1179_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3), .I3(n10691), .O(n108)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1106_1179_add_4_24 (.CI(n10691), .I0(GND_net), 
            .I1(n3), .CO(n10692));
    SB_LUT4 led_counter_1106_1179_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_1202), .I3(n10690), .O(n109)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4383_2_lut (.I0(reset_all), .I1(wp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5585));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4383_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY led_counter_1106_1179_add_4_23 (.CI(n10690), .I0(GND_net), 
            .I1(n4_adj_1202), .CO(n10691));
    SB_LUT4 i4167_3_lut (.I0(\REG.mem_41_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5369));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4168_3_lut (.I0(\REG.mem_41_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5370));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1106_1179_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_1201), .I3(n10689), .O(n110)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4384_2_lut (.I0(reset_all), .I1(wp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5586));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4384_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4700_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[6]), .I2(\mem_LUT.data_raw_r [6]), 
            .I3(n4249), .O(n5902));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4700_4_lut.LUT_INIT = 16'h5044;
    SB_CARRY led_counter_1106_1179_add_4_22 (.CI(n10689), .I0(GND_net), 
            .I1(n5_adj_1201), .CO(n10690));
    SB_LUT4 led_counter_1106_1179_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6), .I3(n10688), .O(n111)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11042_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(n11376), .O(n12601));
    defparam i11042_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY led_counter_1106_1179_add_4_21 (.CI(n10688), .I0(GND_net), 
            .I1(n6), .CO(n10689));
    SB_LUT4 led_counter_1106_1179_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_1200), .I3(n10687), .O(n112)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4703_4_lut (.I0(reset_all_w), .I1(fifo_temp_output[7]), .I2(\mem_LUT.data_raw_r [7]), 
            .I3(n4249), .O(n5905));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    defparam i4703_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i3501_2_lut (.I0(is_tx_fifo_full_flag), .I1(spi_rx_byte_ready), 
            .I2(GND_net), .I3(GND_net), .O(n4703));   // src/top.v(879[8] 888[4])
    defparam i3501_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY led_counter_1106_1179_add_4_20 (.CI(n10687), .I0(GND_net), 
            .I1(n7_adj_1200), .CO(n10688));
    SB_LUT4 i4169_3_lut (.I0(\REG.mem_41_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5371));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1106_1179_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8), .I3(n10686), .O(n113)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1106_1179_add_4_19 (.CI(n10686), .I0(GND_net), 
            .I1(n8), .CO(n10687));
    SB_LUT4 i4170_3_lut (.I0(\REG.mem_41_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5372));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4171_3_lut (.I0(\REG.mem_41_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5373));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4172_3_lut (.I0(\REG.mem_41_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n24_adj_1185), .I3(GND_net), .O(n5374));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4173_3_lut (.I0(\REG.mem_42_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n23), .I3(GND_net), .O(n5375));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4174_3_lut (.I0(\REG.mem_42_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n23), .I3(GND_net), .O(n5376));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4175_3_lut (.I0(\REG.mem_42_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n23), .I3(GND_net), .O(n5377));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4176_3_lut (.I0(\REG.mem_42_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n23), .I3(GND_net), .O(n5378));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1106_1179_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9), .I3(n10685), .O(n114)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4177_3_lut (.I0(\REG.mem_42_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n23), .I3(GND_net), .O(n5379));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4178_3_lut (.I0(\REG.mem_42_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n23), .I3(GND_net), .O(n5380));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4179_3_lut (.I0(\REG.mem_42_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n23), .I3(GND_net), .O(n5381));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4180_3_lut (.I0(\REG.mem_42_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n23), .I3(GND_net), .O(n5382));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4181_3_lut (.I0(\REG.mem_42_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n23), .I3(GND_net), .O(n5383));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_93 (.I0(reset_clk_counter[3]), .I1(reset_clk_counter[2]), 
            .I2(n10562), .I3(GND_net), .O(n10802));
    defparam i1_3_lut_adj_93.LUT_INIT = 16'ha9a9;
    SB_LUT4 i4182_3_lut (.I0(\REG.mem_42_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n23), .I3(GND_net), .O(n5384));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4183_3_lut (.I0(\REG.mem_42_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n23), .I3(GND_net), .O(n5385));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4183_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1106_1179_add_4_18 (.CI(n10685), .I0(GND_net), 
            .I1(n9), .CO(n10686));
    SB_IO FIFO_D1_pad (.PACKAGE_PIN(FIFO_D1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D1_c_1));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D1_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D1_pad.PULLUP = 1'b0;
    defparam FIFO_D1_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D2_pad (.PACKAGE_PIN(FIFO_D2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D2_c_2));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D2_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D2_pad.PULLUP = 1'b0;
    defparam FIFO_D2_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 led_counter_1106_1179_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_1199), .I3(n10684), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_IO FIFO_D3_pad (.PACKAGE_PIN(FIFO_D3), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D3_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D3_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D3_pad.PULLUP = 1'b0;
    defparam FIFO_D3_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4184_3_lut (.I0(\REG.mem_42_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n23), .I3(GND_net), .O(n5386));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4184_3_lut.LUT_INIT = 16'hcaca;
    SB_IO FIFO_D4_pad (.PACKAGE_PIN(FIFO_D4), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D4_c_4));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D4_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D4_pad.PULLUP = 1'b0;
    defparam FIFO_D4_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D5_pad (.PACKAGE_PIN(FIFO_D5), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D5_c_5));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D5_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D5_pad.PULLUP = 1'b0;
    defparam FIFO_D5_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D6_pad (.PACKAGE_PIN(FIFO_D6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D6_c_6));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D6_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D6_pad.PULLUP = 1'b0;
    defparam FIFO_D6_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D7_pad (.PACKAGE_PIN(FIFO_D7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D7_c_7));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D7_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D7_pad.PULLUP = 1'b0;
    defparam FIFO_D7_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D8_pad (.PACKAGE_PIN(FIFO_D8), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D8_c_8));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D8_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D8_pad.PULLUP = 1'b0;
    defparam FIFO_D8_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D9_pad (.PACKAGE_PIN(FIFO_D9), .OUTPUT_ENABLE(VCC_net), .D_IN_0(FIFO_D9_c_9));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D9_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D9_pad.PULLUP = 1'b0;
    defparam FIFO_D9_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D10_pad (.PACKAGE_PIN(FIFO_D10), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D10_c_10));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D10_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D10_pad.PULLUP = 1'b0;
    defparam FIFO_D10_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4185_3_lut (.I0(\REG.mem_42_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n23), .I3(GND_net), .O(n5387));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4185_3_lut.LUT_INIT = 16'hcaca;
    SB_IO FIFO_D11_pad (.PACKAGE_PIN(FIFO_D11), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D11_c_11));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D11_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D11_pad.PULLUP = 1'b0;
    defparam FIFO_D11_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D12_pad (.PACKAGE_PIN(FIFO_D12), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D12_c_12));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D12_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D12_pad.PULLUP = 1'b0;
    defparam FIFO_D12_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4186_3_lut (.I0(\REG.mem_42_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n23), .I3(GND_net), .O(n5388));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4186_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1106_1179_add_4_17 (.CI(n10684), .I0(GND_net), 
            .I1(n10_adj_1199), .CO(n10685));
    SB_IO FIFO_D13_pad (.PACKAGE_PIN(FIFO_D13), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D13_c_13));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D13_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D13_pad.PULLUP = 1'b0;
    defparam FIFO_D13_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D14_pad (.PACKAGE_PIN(FIFO_D14), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D14_c_14));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D14_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D14_pad.PULLUP = 1'b0;
    defparam FIFO_D14_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FIFO_D15_pad (.PACKAGE_PIN(FIFO_D15), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(FIFO_D15_c_15));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FIFO_D15_pad.PIN_TYPE = 6'b000001;
    defparam FIFO_D15_pad.PULLUP = 1'b0;
    defparam FIFO_D15_pad.NEG_TRIGGER = 1'b0;
    defparam FIFO_D15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO DEBUG_6_c_pad (.PACKAGE_PIN(FIFO_CLK), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(DEBUG_6_c_c));   // src/top.v(84[12:20])
    defparam DEBUG_6_c_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_6_c_pad.PULLUP = 1'b0;
    defparam DEBUG_6_c_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_6_c_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4401_2_lut (.I0(reset_all), .I1(wp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5603));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4401_2_lut.LUT_INIT = 16'h4444;
    SB_IO DEBUG_2_c_pad (.PACKAGE_PIN(FR_RXF), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(DEBUG_2_c_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_2_c_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_2_c_pad.PULLUP = 1'b0;
    defparam DEBUG_2_c_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_2_c_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SOUT_pad (.PACKAGE_PIN(SOUT), .OUTPUT_ENABLE(VCC_net), .D_IN_0(SOUT_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SOUT_pad.PIN_TYPE = 6'b000001;
    defparam SOUT_pad.PULLUP = 1'b0;
    defparam SOUT_pad.NEG_TRIGGER = 1'b0;
    defparam SOUT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UART_RX_pad (.PACKAGE_PIN(UART_RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(UART_RX_c)) /* synthesis IO_FF_IN=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UART_RX_pad.PIN_TYPE = 6'b000001;
    defparam UART_RX_pad.PULLUP = 1'b0;
    defparam UART_RX_pad.NEG_TRIGGER = 1'b0;
    defparam UART_RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4187_3_lut (.I0(\REG.mem_42_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n23), .I3(GND_net), .O(n5389));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4187_3_lut.LUT_INIT = 16'hcaca;
    SB_IO ICE_SYSCLK_pad (.PACKAGE_PIN(ICE_SYSCLK), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ICE_SYSCLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_SYSCLK_pad.PIN_TYPE = 6'b000001;
    defparam ICE_SYSCLK_pad.PULLUP = 1'b0;
    defparam ICE_SYSCLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_SYSCLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CREST_pad (.PACKAGE_PIN(ICE_CREST), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CREST_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CREST_pad.PULLUP = 1'b0;
    defparam ICE_CREST_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CREST_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CDONE_pad (.PACKAGE_PIN(ICE_CDONE), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CDONE_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CDONE_pad.PULLUP = 1'b0;
    defparam ICE_CDONE_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CDONE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ICE_CLK_pad (.PACKAGE_PIN(ICE_CLK), .OUTPUT_ENABLE(GND_net), .D_OUT_0(GND_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ICE_CLK_pad.PIN_TYPE = 6'b101001;
    defparam ICE_CLK_pad.PULLUP = 1'b0;
    defparam ICE_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam ICE_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4402_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n5604));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4402_2_lut.LUT_INIT = 16'h4444;
    SB_IO DEBUG_9_pad (.PACKAGE_PIN(DEBUG_9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_9_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_9_pad.PULLUP = 1'b0;
    defparam DEBUG_9_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_8_pad (.PACKAGE_PIN(DEBUG_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(\afull_flag_impl.af_flag_p_w_N_603 [3]));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_8_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_8_pad.PULLUP = 1'b0;
    defparam DEBUG_8_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 led_counter_1106_1179_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11), .I3(n10683), .O(n116)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_IO DEBUG_6_pad (.PACKAGE_PIN(DEBUG_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_6_c_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_6_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_6_pad.PULLUP = 1'b0;
    defparam DEBUG_6_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_5_pad (.PACKAGE_PIN(DEBUG_5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_5_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_5_pad.PULLUP = 1'b0;
    defparam DEBUG_5_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_3_pad (.PACKAGE_PIN(DEBUG_3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_3_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_3_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_3_pad.PULLUP = 1'b0;
    defparam DEBUG_3_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_2_pad (.PACKAGE_PIN(DEBUG_2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_2_c_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_2_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_2_pad.PULLUP = 1'b0;
    defparam DEBUG_2_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_1_pad (.PACKAGE_PIN(DEBUG_1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_1_c_0_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_1_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_1_pad.PULLUP = 1'b0;
    defparam DEBUG_1_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_0_pad (.PACKAGE_PIN(DEBUG_0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_0_c_24));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_0_pad.PIN_TYPE = 6'b011001;
    defparam DEBUG_0_pad.PULLUP = 1'b0;
    defparam DEBUG_0_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_SIWU_pad (.PACKAGE_PIN(FT_SIWU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_SIWU_pad.PIN_TYPE = 6'b011001;
    defparam FT_SIWU_pad.PULLUP = 1'b0;
    defparam FT_SIWU_pad.NEG_TRIGGER = 1'b0;
    defparam FT_SIWU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_WR_pad (.PACKAGE_PIN(FT_WR), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_WR_pad.PIN_TYPE = 6'b011001;
    defparam FT_WR_pad.PULLUP = 1'b0;
    defparam FT_WR_pad.NEG_TRIGGER = 1'b0;
    defparam FT_WR_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4403_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5605));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4403_2_lut.LUT_INIT = 16'h4444;
    SB_IO FT_RD_pad (.PACKAGE_PIN(FT_RD), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DEBUG_3_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_RD_pad.PIN_TYPE = 6'b011001;
    defparam FT_RD_pad.PULLUP = 1'b0;
    defparam FT_RD_pad.NEG_TRIGGER = 1'b0;
    defparam FT_RD_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO FT_OE_pad (.PACKAGE_PIN(FT_OE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(FT_OE_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam FT_OE_pad.PIN_TYPE = 6'b011001;
    defparam FT_OE_pad.PULLUP = 1'b0;
    defparam FT_OE_pad.NEG_TRIGGER = 1'b0;
    defparam FT_OE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA10_pad (.PACKAGE_PIN(DATA10), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA10_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA10_pad.PIN_TYPE = 6'b011001;
    defparam DATA10_pad.PULLUP = 1'b0;
    defparam DATA10_pad.NEG_TRIGGER = 1'b0;
    defparam DATA10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA9_pad (.PACKAGE_PIN(DATA9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA9_pad.PIN_TYPE = 6'b011001;
    defparam DATA9_pad.PULLUP = 1'b0;
    defparam DATA9_pad.NEG_TRIGGER = 1'b0;
    defparam DATA9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA11_pad (.PACKAGE_PIN(DATA11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA11_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA11_pad.PIN_TYPE = 6'b011001;
    defparam DATA11_pad.PULLUP = 1'b0;
    defparam DATA11_pad.NEG_TRIGGER = 1'b0;
    defparam DATA11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA12_pad (.PACKAGE_PIN(DATA12), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA12_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA12_pad.PIN_TYPE = 6'b011001;
    defparam DATA12_pad.PULLUP = 1'b0;
    defparam DATA12_pad.NEG_TRIGGER = 1'b0;
    defparam DATA12_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY led_counter_1106_1179_add_4_16 (.CI(n10683), .I0(GND_net), 
            .I1(n11), .CO(n10684));
    SB_IO DATA13_pad (.PACKAGE_PIN(DATA13), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA13_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA13_pad.PIN_TYPE = 6'b011001;
    defparam DATA13_pad.PULLUP = 1'b0;
    defparam DATA13_pad.NEG_TRIGGER = 1'b0;
    defparam DATA13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA14_pad (.PACKAGE_PIN(DATA14), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA14_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA14_pad.PIN_TYPE = 6'b011001;
    defparam DATA14_pad.PULLUP = 1'b0;
    defparam DATA14_pad.NEG_TRIGGER = 1'b0;
    defparam DATA14_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA8_pad (.PACKAGE_PIN(DATA8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA8_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA8_pad.PIN_TYPE = 6'b011001;
    defparam DATA8_pad.PULLUP = 1'b0;
    defparam DATA8_pad.NEG_TRIGGER = 1'b0;
    defparam DATA8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA15_pad (.PACKAGE_PIN(DATA15), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA15_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA15_pad.PIN_TYPE = 6'b011001;
    defparam DATA15_pad.PULLUP = 1'b0;
    defparam DATA15_pad.NEG_TRIGGER = 1'b0;
    defparam DATA15_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4188_3_lut (.I0(\REG.mem_42_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n23), .I3(GND_net), .O(n5390));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4188_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DATA16_pad (.PACKAGE_PIN(DATA16), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA16_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA16_pad.PIN_TYPE = 6'b011001;
    defparam DATA16_pad.PULLUP = 1'b0;
    defparam DATA16_pad.NEG_TRIGGER = 1'b0;
    defparam DATA16_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA7_pad (.PACKAGE_PIN(DATA7), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA7_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA7_pad.PIN_TYPE = 6'b011001;
    defparam DATA7_pad.PULLUP = 1'b0;
    defparam DATA7_pad.NEG_TRIGGER = 1'b0;
    defparam DATA7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 led_counter_1106_1179_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12), .I3(n10682), .O(n117)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_IO DATA17_pad (.PACKAGE_PIN(DATA17), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA17_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA17_pad.PIN_TYPE = 6'b011001;
    defparam DATA17_pad.PULLUP = 1'b0;
    defparam DATA17_pad.NEG_TRIGGER = 1'b0;
    defparam DATA17_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA18_pad (.PACKAGE_PIN(DATA18), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA18_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA18_pad.PIN_TYPE = 6'b011001;
    defparam DATA18_pad.PULLUP = 1'b0;
    defparam DATA18_pad.NEG_TRIGGER = 1'b0;
    defparam DATA18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA6_pad (.PACKAGE_PIN(DATA6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA6_pad.PIN_TYPE = 6'b011001;
    defparam DATA6_pad.PULLUP = 1'b0;
    defparam DATA6_pad.NEG_TRIGGER = 1'b0;
    defparam DATA6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA19_pad (.PACKAGE_PIN(DATA19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA19_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA19_pad.PIN_TYPE = 6'b011001;
    defparam DATA19_pad.PULLUP = 1'b0;
    defparam DATA19_pad.NEG_TRIGGER = 1'b0;
    defparam DATA19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA20_pad (.PACKAGE_PIN(DATA20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA20_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA20_pad.PIN_TYPE = 6'b011001;
    defparam DATA20_pad.PULLUP = 1'b0;
    defparam DATA20_pad.NEG_TRIGGER = 1'b0;
    defparam DATA20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA5_pad (.PACKAGE_PIN(DATA5), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA5_pad.PIN_TYPE = 6'b011001;
    defparam DATA5_pad.PULLUP = 1'b0;
    defparam DATA5_pad.NEG_TRIGGER = 1'b0;
    defparam DATA5_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA21_pad (.PACKAGE_PIN(DATA21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA5_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA21_pad.PIN_TYPE = 6'b011001;
    defparam DATA21_pad.PULLUP = 1'b0;
    defparam DATA21_pad.NEG_TRIGGER = 1'b0;
    defparam DATA21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA22_pad (.PACKAGE_PIN(DATA22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA6_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA22_pad.PIN_TYPE = 6'b011001;
    defparam DATA22_pad.PULLUP = 1'b0;
    defparam DATA22_pad.NEG_TRIGGER = 1'b0;
    defparam DATA22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA4_pad (.PACKAGE_PIN(DATA4), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA20_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA4_pad.PIN_TYPE = 6'b011001;
    defparam DATA4_pad.PULLUP = 1'b0;
    defparam DATA4_pad.NEG_TRIGGER = 1'b0;
    defparam DATA4_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA23_pad (.PACKAGE_PIN(DATA23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA7_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA23_pad.PIN_TYPE = 6'b011001;
    defparam DATA23_pad.PULLUP = 1'b0;
    defparam DATA23_pad.NEG_TRIGGER = 1'b0;
    defparam DATA23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA24_pad (.PACKAGE_PIN(DATA24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA8_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA24_pad.PIN_TYPE = 6'b011001;
    defparam DATA24_pad.PULLUP = 1'b0;
    defparam DATA24_pad.NEG_TRIGGER = 1'b0;
    defparam DATA24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA3_pad (.PACKAGE_PIN(DATA3), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA19_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA3_pad.PIN_TYPE = 6'b011001;
    defparam DATA3_pad.PULLUP = 1'b0;
    defparam DATA3_pad.NEG_TRIGGER = 1'b0;
    defparam DATA3_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA25_pad (.PACKAGE_PIN(DATA25), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA9_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA25_pad.PIN_TYPE = 6'b011001;
    defparam DATA25_pad.PULLUP = 1'b0;
    defparam DATA25_pad.NEG_TRIGGER = 1'b0;
    defparam DATA25_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA26_pad (.PACKAGE_PIN(DATA26), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA10_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA26_pad.PIN_TYPE = 6'b011001;
    defparam DATA26_pad.PULLUP = 1'b0;
    defparam DATA26_pad.NEG_TRIGGER = 1'b0;
    defparam DATA26_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4404_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5606));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4404_2_lut.LUT_INIT = 16'h4444;
    SB_IO DATA2_pad (.PACKAGE_PIN(DATA2), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA18_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA2_pad.PIN_TYPE = 6'b011001;
    defparam DATA2_pad.PULLUP = 1'b0;
    defparam DATA2_pad.NEG_TRIGGER = 1'b0;
    defparam DATA2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA27_pad (.PACKAGE_PIN(DATA27), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA11_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA27_pad.PIN_TYPE = 6'b011001;
    defparam DATA27_pad.PULLUP = 1'b0;
    defparam DATA27_pad.NEG_TRIGGER = 1'b0;
    defparam DATA27_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA28_pad (.PACKAGE_PIN(DATA28), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA12_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA28_pad.PIN_TYPE = 6'b011001;
    defparam DATA28_pad.PULLUP = 1'b0;
    defparam DATA28_pad.NEG_TRIGGER = 1'b0;
    defparam DATA28_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA1_pad (.PACKAGE_PIN(DATA1), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA17_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA1_pad.PIN_TYPE = 6'b011001;
    defparam DATA1_pad.PULLUP = 1'b0;
    defparam DATA1_pad.NEG_TRIGGER = 1'b0;
    defparam DATA1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4405_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5607));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4405_2_lut.LUT_INIT = 16'h4444;
    SB_IO DATA29_pad (.PACKAGE_PIN(DATA29), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA13_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA29_pad.PIN_TYPE = 6'b011001;
    defparam DATA29_pad.PULLUP = 1'b0;
    defparam DATA29_pad.NEG_TRIGGER = 1'b0;
    defparam DATA29_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA30_pad (.PACKAGE_PIN(DATA30), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA14_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA30_pad.PIN_TYPE = 6'b011001;
    defparam DATA30_pad.PULLUP = 1'b0;
    defparam DATA30_pad.NEG_TRIGGER = 1'b0;
    defparam DATA30_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DATA0_pad (.PACKAGE_PIN(DATA0), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA16_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA0_pad.PIN_TYPE = 6'b011001;
    defparam DATA0_pad.PULLUP = 1'b0;
    defparam DATA0_pad.NEG_TRIGGER = 1'b0;
    defparam DATA0_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i6317_2_lut_3_lut (.I0(state[1]), .I1(state[0]), .I2(n63), 
            .I3(GND_net), .O(n7495));
    defparam i6317_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_IO DATA31_pad (.PACKAGE_PIN(DATA31), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DATA15_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DATA31_pad.PIN_TYPE = 6'b011001;
    defparam DATA31_pad.PULLUP = 1'b0;
    defparam DATA31_pad.NEG_TRIGGER = 1'b0;
    defparam DATA31_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO VALID_pad (.PACKAGE_PIN(VALID), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VALID_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam VALID_pad.PIN_TYPE = 6'b011001;
    defparam VALID_pad.PULLUP = 1'b0;
    defparam VALID_pad.NEG_TRIGGER = 1'b0;
    defparam VALID_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SYNC_pad (.PACKAGE_PIN(SYNC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SYNC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SYNC_pad.PIN_TYPE = 6'b011001;
    defparam SYNC_pad.PULLUP = 1'b0;
    defparam SYNC_pad.NEG_TRIGGER = 1'b0;
    defparam SYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4190_3_lut (.I0(\REG.mem_43_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n22), .I3(GND_net), .O(n5392));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4190_3_lut.LUT_INIT = 16'hcaca;
    SB_IO INVERT_pad (.PACKAGE_PIN(INVERT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INVERT_c_4)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INVERT_pad.PIN_TYPE = 6'b011001;
    defparam INVERT_pad.PULLUP = 1'b0;
    defparam INVERT_pad.NEG_TRIGGER = 1'b0;
    defparam INVERT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SLM_CLK_pad (.PACKAGE_PIN(SLM_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SLM_CLK_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SLM_CLK_pad.PIN_TYPE = 6'b011001;
    defparam SLM_CLK_pad.PULLUP = 1'b0;
    defparam SLM_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam SLM_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO RESET_pad (.PACKAGE_PIN(RESET), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(RESET_c));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RESET_pad.PIN_TYPE = 6'b011001;
    defparam RESET_pad.PULLUP = 1'b0;
    defparam RESET_pad.NEG_TRIGGER = 1'b0;
    defparam RESET_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO UPDATE_pad (.PACKAGE_PIN(UPDATE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(UPDATE_c_3));   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam UPDATE_pad.PIN_TYPE = 6'b011001;
    defparam UPDATE_pad.PULLUP = 1'b0;
    defparam UPDATE_pad.NEG_TRIGGER = 1'b0;
    defparam UPDATE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF tx_data_byte_r_i0_i1 (.Q(tx_data_byte[1]), .C(SLM_CLK_c), .D(n5500));   // src/top.v(1064[8] 1131[4])
    SB_DFF tx_data_byte_r_i0_i2 (.Q(tx_data_byte[2]), .C(SLM_CLK_c), .D(n5499));   // src/top.v(1064[8] 1131[4])
    SB_IO SDAT_pad (.PACKAGE_PIN(SDAT), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SDAT_c_15)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SDAT_pad.PIN_TYPE = 6'b011001;
    defparam SDAT_pad.PULLUP = 1'b0;
    defparam SDAT_pad.NEG_TRIGGER = 1'b0;
    defparam SDAT_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SCK_pad (.PACKAGE_PIN(SCK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SCK_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SCK_pad.PIN_TYPE = 6'b011001;
    defparam SCK_pad.PULLUP = 1'b0;
    defparam SCK_pad.NEG_TRIGGER = 1'b0;
    defparam SCK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SEN_pad (.PACKAGE_PIN(SEN), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(SEN_c_1)) /* synthesis IO_FF_OUT=TRUE */ ;   // D:/ProgramFiles/Lattice/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SEN_pad.PIN_TYPE = 6'b011001;
    defparam SEN_pad.PULLUP = 1'b0;
    defparam SEN_pad.NEG_TRIGGER = 1'b0;
    defparam SEN_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4191_3_lut (.I0(\REG.mem_43_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n22), .I3(GND_net), .O(n5393));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4192_3_lut (.I0(\REG.mem_43_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n22), .I3(GND_net), .O(n5394));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4406_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5608));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4406_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4193_3_lut (.I0(\REG.mem_43_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n22), .I3(GND_net), .O(n5395));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4194_3_lut (.I0(\REG.mem_43_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n22), .I3(GND_net), .O(n5396));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4194_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_data_byte_r_i0_i3 (.Q(tx_data_byte[3]), .C(SLM_CLK_c), .D(n5498));   // src/top.v(1064[8] 1131[4])
    SB_DFF tx_data_byte_r_i0_i4 (.Q(tx_data_byte[4]), .C(SLM_CLK_c), .D(n5497));   // src/top.v(1064[8] 1131[4])
    SB_DFF tx_data_byte_r_i0_i5 (.Q(tx_data_byte[5]), .C(SLM_CLK_c), .D(n5496));   // src/top.v(1064[8] 1131[4])
    SB_DFF tx_data_byte_r_i0_i6 (.Q(tx_data_byte[6]), .C(SLM_CLK_c), .D(n5495));   // src/top.v(1064[8] 1131[4])
    SB_DFF tx_data_byte_r_i0_i7 (.Q(tx_data_byte[7]), .C(SLM_CLK_c), .D(n5494));   // src/top.v(1064[8] 1131[4])
    SB_LUT4 i4195_3_lut (.I0(\REG.mem_43_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n22), .I3(GND_net), .O(n5397));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[3]), 
            .I3(n4_adj_1182), .O(n11342));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i4196_3_lut (.I0(\REG.mem_43_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n22), .I3(GND_net), .O(n5398));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4197_3_lut (.I0(\REG.mem_43_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n22), .I3(GND_net), .O(n5399));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4198_3_lut (.I0(\REG.mem_43_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n22), .I3(GND_net), .O(n5400));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4198_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF uart_rx_complete_rising_edge_82 (.Q(uart_rx_complete_rising_edge), 
           .C(SLM_CLK_c), .D(n4686));   // src/top.v(1055[8] 1061[4])
    SB_LUT4 i4199_3_lut (.I0(\REG.mem_43_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n22), .I3(GND_net), .O(n5401));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4200_3_lut (.I0(\REG.mem_43_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n22), .I3(GND_net), .O(n5402));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4407_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5609));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i4407_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4408_3_lut (.I0(\REG.mem_55_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n10), .I3(GND_net), .O(n5610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4201_3_lut (.I0(\REG.mem_43_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n22), .I3(GND_net), .O(n5403));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4202_3_lut (.I0(\REG.mem_43_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n22), .I3(GND_net), .O(n5404));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4203_3_lut (.I0(\REG.mem_43_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n22), .I3(GND_net), .O(n5405));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4410_3_lut (.I0(\REG.mem_55_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n10), .I3(GND_net), .O(n5612));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4204_3_lut (.I0(\REG.mem_43_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n22), .I3(GND_net), .O(n5406));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4411_3_lut (.I0(\REG.mem_55_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n10), .I3(GND_net), .O(n5613));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4411_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1106_1179_add_4_15 (.CI(n10682), .I0(GND_net), 
            .I1(n12), .CO(n10683));
    SB_LUT4 i4412_3_lut (.I0(\REG.mem_55_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n10), .I3(GND_net), .O(n5614));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4413_3_lut (.I0(\REG.mem_55_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n10), .I3(GND_net), .O(n5615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4205_3_lut (.I0(\REG.mem_43_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n22), .I3(GND_net), .O(n5407));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4414_3_lut (.I0(\REG.mem_55_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n10), .I3(GND_net), .O(n5616));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4415_3_lut (.I0(\REG.mem_55_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n10), .I3(GND_net), .O(n5617));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4416_3_lut (.I0(\REG.mem_55_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n10), .I3(GND_net), .O(n5618));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1106_1179_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13), .I3(n10681), .O(n118)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4417_3_lut (.I0(\REG.mem_55_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n10), .I3(GND_net), .O(n5619));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4417_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1106_1179_add_4_14 (.CI(n10681), .I0(GND_net), 
            .I1(n13), .CO(n10682));
    SB_LUT4 led_counter_1106_1179_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_1198), .I3(n10680), .O(n119)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4207_3_lut (.I0(\REG.mem_44_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n21), .I3(GND_net), .O(n5409));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4208_3_lut (.I0(\REG.mem_44_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n21), .I3(GND_net), .O(n5410));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4418_3_lut (.I0(\REG.mem_55_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n10), .I3(GND_net), .O(n5620));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4418_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1106_1179_add_4_13 (.CI(n10680), .I0(GND_net), 
            .I1(n14_adj_1198), .CO(n10681));
    SB_LUT4 led_counter_1106_1179_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_1197), .I3(n10679), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4209_3_lut (.I0(\REG.mem_44_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n21), .I3(GND_net), .O(n5411));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4209_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1106_1179_add_4_12 (.CI(n10679), .I0(GND_net), 
            .I1(n15_adj_1197), .CO(n10680));
    SB_LUT4 i4210_3_lut (.I0(\REG.mem_44_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n21), .I3(GND_net), .O(n5412));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4419_3_lut (.I0(\REG.mem_55_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n10), .I3(GND_net), .O(n5621));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4420_3_lut (.I0(\REG.mem_55_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n10), .I3(GND_net), .O(n5622));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4211_3_lut (.I0(\REG.mem_44_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n21), .I3(GND_net), .O(n5413));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4421_3_lut (.I0(\REG.mem_55_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n10), .I3(GND_net), .O(n5623));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1106_1179_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_1196), .I3(n10678), .O(n121)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4212_3_lut (.I0(\REG.mem_44_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n21), .I3(GND_net), .O(n5414));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4213_3_lut (.I0(\REG.mem_44_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n21), .I3(GND_net), .O(n5415));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4214_3_lut (.I0(\REG.mem_44_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n21), .I3(GND_net), .O(n5416));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4422_3_lut (.I0(\REG.mem_55_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n10), .I3(GND_net), .O(n5624));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4215_3_lut (.I0(\REG.mem_44_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n21), .I3(GND_net), .O(n5417));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4216_3_lut (.I0(\REG.mem_44_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n21), .I3(GND_net), .O(n5418));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4423_3_lut (.I0(\REG.mem_55_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n10), .I3(GND_net), .O(n5625));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4217_3_lut (.I0(\REG.mem_44_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n21), .I3(GND_net), .O(n5419));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4218_3_lut (.I0(\REG.mem_44_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n21), .I3(GND_net), .O(n5420));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4219_3_lut (.I0(\REG.mem_44_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n21), .I3(GND_net), .O(n5421));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4219_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF tx_addr_byte_r_i0_i1 (.Q(tx_addr_byte[1]), .C(SLM_CLK_c), .D(n5325));   // src/top.v(1064[8] 1131[4])
    SB_DFF tx_addr_byte_r_i0_i2 (.Q(tx_addr_byte[2]), .C(SLM_CLK_c), .D(n5324));   // src/top.v(1064[8] 1131[4])
    SB_DFF tx_addr_byte_r_i0_i3 (.Q(tx_addr_byte[3]), .C(SLM_CLK_c), .D(n5307));   // src/top.v(1064[8] 1131[4])
    SB_DFF tx_addr_byte_r_i0_i4 (.Q(tx_addr_byte[4]), .C(SLM_CLK_c), .D(n5306));   // src/top.v(1064[8] 1131[4])
    SB_DFF tx_addr_byte_r_i0_i5 (.Q(tx_addr_byte[5]), .C(SLM_CLK_c), .D(n5305));   // src/top.v(1064[8] 1131[4])
    SB_DFF tx_addr_byte_r_i0_i6 (.Q(tx_addr_byte[6]), .C(SLM_CLK_c), .D(n5304));   // src/top.v(1064[8] 1131[4])
    SB_DFF tx_addr_byte_r_i0_i7 (.Q(tx_addr_byte[7]), .C(SLM_CLK_c), .D(n5303));   // src/top.v(1064[8] 1131[4])
    SB_LUT4 i4220_3_lut (.I0(\REG.mem_44_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n21), .I3(GND_net), .O(n5422));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i919_4_lut (.I0(n1876), .I1(n7566), .I2(state[3]), .I3(n63), 
            .O(n1721));   // src/timing_controller.v(48[11:16])
    defparam i919_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i4221_3_lut (.I0(\REG.mem_44_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n21), .I3(GND_net), .O(n5423));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4222_3_lut (.I0(\REG.mem_44_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n21), .I3(GND_net), .O(n5424));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4223_3_lut (.I0(\REG.mem_45_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n20), .I3(GND_net), .O(n5425));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4224_3_lut (.I0(\REG.mem_45_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n20), .I3(GND_net), .O(n5426));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4224_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1106_1179_add_4_11 (.CI(n10678), .I0(GND_net), 
            .I1(n16_adj_1196), .CO(n10679));
    SB_LUT4 i4424_3_lut (.I0(\REG.mem_55_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n10), .I3(GND_net), .O(n5626));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4225_3_lut (.I0(\REG.mem_45_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n20), .I3(GND_net), .O(n5427));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4226_3_lut (.I0(\REG.mem_45_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n20), .I3(GND_net), .O(n5428));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4226_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF reset_clk_counter_i3_1107__i0 (.Q(reset_clk_counter[0]), .C(SLM_CLK_c), 
           .D(n25_adj_1204));   // src/top.v(259[27:51])
    SB_LUT4 i4227_3_lut (.I0(\REG.mem_45_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n20), .I3(GND_net), .O(n5429));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4228_3_lut (.I0(\REG.mem_45_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n20), .I3(GND_net), .O(n5430));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4229_3_lut (.I0(\REG.mem_45_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n20), .I3(GND_net), .O(n5431));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4230_3_lut (.I0(\REG.mem_45_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n20), .I3(GND_net), .O(n5432));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4231_3_lut (.I0(\REG.mem_45_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n20), .I3(GND_net), .O(n5433));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4232_3_lut (.I0(\REG.mem_45_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n20), .I3(GND_net), .O(n5434));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4233_3_lut (.I0(\REG.mem_45_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n20), .I3(GND_net), .O(n5435));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4234_3_lut (.I0(\REG.mem_45_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n20), .I3(GND_net), .O(n5436));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4235_3_lut (.I0(\REG.mem_45_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n20), .I3(GND_net), .O(n5437));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4236_3_lut (.I0(\REG.mem_45_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n20), .I3(GND_net), .O(n5438));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 led_counter_1106_1179_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_1195), .I3(n10677), .O(n122)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4237_3_lut (.I0(\REG.mem_45_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n20), .I3(GND_net), .O(n5439));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4238_3_lut (.I0(\REG.mem_45_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n20), .I3(GND_net), .O(n5440));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4239_3_lut (.I0(\REG.mem_46_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n19), .I3(GND_net), .O(n5441));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4240_3_lut (.I0(\REG.mem_46_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n19), .I3(GND_net), .O(n5442));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4241_3_lut (.I0(\REG.mem_46_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n19), .I3(GND_net), .O(n5443));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4242_3_lut (.I0(\REG.mem_46_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n19), .I3(GND_net), .O(n5444));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4243_3_lut (.I0(\REG.mem_46_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n19), .I3(GND_net), .O(n5445));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4244_3_lut (.I0(\REG.mem_46_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n19), .I3(GND_net), .O(n5446));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4245_3_lut (.I0(\REG.mem_46_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n19), .I3(GND_net), .O(n5447));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4246_3_lut (.I0(\REG.mem_46_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n19), .I3(GND_net), .O(n5448));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4247_3_lut (.I0(\REG.mem_46_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n19), .I3(GND_net), .O(n5449));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4248_3_lut (.I0(\REG.mem_46_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n19), .I3(GND_net), .O(n5450));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4248_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1106_1179_add_4_10 (.CI(n10677), .I0(GND_net), 
            .I1(n17_adj_1195), .CO(n10678));
    SB_LUT4 led_counter_1106_1179_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_1194), .I3(n10676), .O(n123)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF tx_addr_byte_r_i0_i0 (.Q(tx_addr_byte[0]), .C(SLM_CLK_c), .D(n4654));   // src/top.v(1064[8] 1131[4])
    SB_LUT4 i3484_2_lut (.I0(uart_rx_complete_prev), .I1(debug_led3), .I2(GND_net), 
            .I3(GND_net), .O(n4686));   // src/top.v(1055[8] 1061[4])
    defparam i3484_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4249_3_lut (.I0(\REG.mem_46_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n19), .I3(GND_net), .O(n5451));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4250_3_lut (.I0(\REG.mem_46_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n19), .I3(GND_net), .O(n5452));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4251_3_lut (.I0(\REG.mem_46_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n19), .I3(GND_net), .O(n5453));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4252_3_lut (.I0(\REG.mem_46_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n19), .I3(GND_net), .O(n5454));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4252_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF even_byte_flag_89 (.Q(even_byte_flag), .C(SLM_CLK_c), .D(n2679));   // src/top.v(1064[8] 1131[4])
    SB_LUT4 i4253_3_lut (.I0(\REG.mem_46_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n19), .I3(GND_net), .O(n5455));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4458_2_lut (.I0(reset_all), .I1(rd_addr_nxt_c_6__N_465[5]), 
            .I2(GND_net), .I3(GND_net), .O(n5660));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i4458_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4254_3_lut (.I0(\REG.mem_46_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n19), .I3(GND_net), .O(n5456));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4254_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1106_1179_add_4_9 (.CI(n10676), .I0(GND_net), .I1(n18_adj_1194), 
            .CO(n10677));
    SB_LUT4 i4255_3_lut (.I0(\REG.mem_47_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n18), .I3(GND_net), .O(n5457));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4460_2_lut (.I0(reset_all), .I1(rd_addr_nxt_c_6__N_465[3]), 
            .I2(GND_net), .I3(GND_net), .O(n5662));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i4460_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4256_3_lut (.I0(\REG.mem_47_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n18), .I3(GND_net), .O(n5458));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4257_3_lut (.I0(\REG.mem_47_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n18), .I3(GND_net), .O(n5459));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4258_3_lut (.I0(\REG.mem_47_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n18), .I3(GND_net), .O(n5460));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4259_3_lut (.I0(\REG.mem_47_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n18), .I3(GND_net), .O(n5461));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4260_3_lut (.I0(\REG.mem_47_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n18), .I3(GND_net), .O(n5462));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4261_3_lut (.I0(\REG.mem_47_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n18), .I3(GND_net), .O(n5463));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4462_2_lut (.I0(reset_all), .I1(rd_addr_nxt_c_6__N_465[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5664));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i4462_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4262_3_lut (.I0(\REG.mem_47_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n18), .I3(GND_net), .O(n5464));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4463_2_lut (.I0(reset_all), .I1(rp_sync1_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n5665));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4463_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4263_3_lut (.I0(\REG.mem_47_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n18), .I3(GND_net), .O(n5465));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4264_3_lut (.I0(\REG.mem_47_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n18), .I3(GND_net), .O(n5466));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4464_2_lut (.I0(reset_all), .I1(rp_sync1_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5666));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4464_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4465_3_lut (.I0(\REG.mem_58_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5667));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4466_3_lut (.I0(\REG.mem_58_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5668));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4467_3_lut (.I0(\REG.mem_58_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5669));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4468_3_lut (.I0(\REG.mem_58_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5670));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4469_3_lut (.I0(\REG.mem_58_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5671));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4470_3_lut (.I0(\REG.mem_58_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5672));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4471_3_lut (.I0(\REG.mem_58_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5673));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4472_3_lut (.I0(\REG.mem_58_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5674));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4473_3_lut (.I0(\REG.mem_58_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5675));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4474_3_lut (.I0(\REG.mem_58_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5676));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4475_3_lut (.I0(\REG.mem_58_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5677));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4476_3_lut (.I0(\REG.mem_58_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5678));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4477_3_lut (.I0(\REG.mem_58_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5679));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4478_3_lut (.I0(\REG.mem_58_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5680));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4479_3_lut (.I0(\REG.mem_58_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5681));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4480_3_lut (.I0(\REG.mem_58_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n7_adj_1183), .I3(GND_net), .O(n5682));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4481_2_lut (.I0(reset_all), .I1(rp_sync1_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5683));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4481_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3522_3_lut (.I0(r_Tx_Data[7]), .I1(fifo_temp_output[7]), .I2(n3710), 
            .I3(GND_net), .O(n4724));   // src/uart_tx.v(38[10] 141[8])
    defparam i3522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4482_2_lut (.I0(reset_all), .I1(rp_sync1_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5684));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4482_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4483_2_lut (.I0(reset_all), .I1(rp_sync1_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5685));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4483_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4484_2_lut (.I0(reset_all), .I1(rp_sync1_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5686));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4484_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4502_2_lut (.I0(reset_all), .I1(rd_addr_r[6]), .I2(GND_net), 
            .I3(GND_net), .O(n5704));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4502_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i6205_1_lut (.I0(n1616), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n7383));   // src/timing_controller.v(48[11:16])
    defparam i6205_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 led_counter_1106_1179_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_1193), .I3(n10675), .O(n124)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4503_2_lut (.I0(reset_all), .I1(rd_grey_sync_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5705));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4503_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4504_2_lut (.I0(reset_all), .I1(rd_grey_sync_r[4]), .I2(GND_net), 
            .I3(GND_net), .O(n5706));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4504_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4505_2_lut (.I0(reset_all), .I1(rd_grey_sync_r[3]), .I2(GND_net), 
            .I3(GND_net), .O(n5707));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4505_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4506_2_lut (.I0(reset_all), .I1(rd_grey_sync_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5708));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4506_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4507_2_lut (.I0(reset_all), .I1(rd_grey_sync_r[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5709));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i4507_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3_4_lut (.I0(reset_clk_counter[0]), .I1(reset_clk_counter[2]), 
            .I2(reset_clk_counter[3]), .I3(reset_clk_counter[1]), .O(reset_all_w_N_61));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3114_4_lut (.I0(n63), .I1(n3929), .I2(n7566), .I3(state[3]), 
            .O(n1616));   // src/timing_controller.v(48[11:16])
    defparam i3114_4_lut.LUT_INIT = 16'h0a88;
    SB_CARRY led_counter_1106_1179_add_4_8 (.CI(n10675), .I0(GND_net), .I1(n19_adj_1193), 
            .CO(n10676));
    SB_LUT4 i4525_3_lut (.I0(rx_buf_byte[7]), .I1(rx_shift_reg[7]), .I2(n3204), 
            .I3(GND_net), .O(n5727));   // src/spi.v(76[8] 221[4])
    defparam i4525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4526_3_lut (.I0(rx_buf_byte[6]), .I1(rx_shift_reg[6]), .I2(n3204), 
            .I3(GND_net), .O(n5728));   // src/spi.v(76[8] 221[4])
    defparam i4526_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4527_3_lut (.I0(rx_buf_byte[5]), .I1(rx_shift_reg[5]), .I2(n3204), 
            .I3(GND_net), .O(n5729));   // src/spi.v(76[8] 221[4])
    defparam i4527_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4528_3_lut (.I0(rx_buf_byte[4]), .I1(rx_shift_reg[4]), .I2(n3204), 
            .I3(GND_net), .O(n5730));   // src/spi.v(76[8] 221[4])
    defparam i4528_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4529_3_lut (.I0(rx_buf_byte[3]), .I1(rx_shift_reg[3]), .I2(n3204), 
            .I3(GND_net), .O(n5731));   // src/spi.v(76[8] 221[4])
    defparam i4529_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4530_3_lut (.I0(rx_buf_byte[2]), .I1(rx_shift_reg[2]), .I2(n3204), 
            .I3(GND_net), .O(n5732));   // src/spi.v(76[8] 221[4])
    defparam i4530_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4531_3_lut (.I0(rx_buf_byte[1]), .I1(rx_shift_reg[1]), .I2(n3204), 
            .I3(GND_net), .O(n5733));   // src/spi.v(76[8] 221[4])
    defparam i4531_3_lut.LUT_INIT = 16'hacac;
    SB_DFF tx_data_byte_r_i0_i0 (.Q(tx_data_byte[0]), .C(SLM_CLK_c), .D(n4609));   // src/top.v(1064[8] 1131[4])
    SB_LUT4 led_counter_1106_1179_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_1192), .I3(n10674), .O(n125)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1106_1179_add_4_7 (.CI(n10674), .I0(GND_net), .I1(n20_adj_1192), 
            .CO(n10675));
    SB_LUT4 led_counter_1106_1179_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_1191), .I3(n10673), .O(n126)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR multi_byte_spi_trans_flag_r_86 (.Q(multi_byte_spi_trans_flag_r), 
            .C(SLM_CLK_c), .D(multi_byte_spi_trans_flag_r_N_72), .R(n4443));   // src/top.v(1064[8] 1131[4])
    SB_CARRY led_counter_1106_1179_add_4_6 (.CI(n10673), .I0(GND_net), .I1(n21_adj_1191), 
            .CO(n10674));
    SB_LUT4 led_counter_1106_1179_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_1190), .I3(n10672), .O(n127)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1106_1179_add_4_5 (.CI(n10672), .I0(GND_net), .I1(n22_adj_1190), 
            .CO(n10673));
    SB_LUT4 led_counter_1106_1179_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_1189), .I3(n10671), .O(n128)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1106_1179_add_4_4 (.CI(n10671), .I0(GND_net), .I1(n23_adj_1189), 
            .CO(n10672));
    SB_LUT4 led_counter_1106_1179_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_1188), .I3(n10670), .O(n129)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY led_counter_1106_1179_add_4_3 (.CI(n10670), .I0(GND_net), .I1(n24_adj_1188), 
            .CO(n10671));
    SB_LUT4 led_counter_1106_1179_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_1187), .I3(VCC_net), .O(n130)) /* synthesis syn_instantiated=1 */ ;
    defparam led_counter_1106_1179_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4548_3_lut (.I0(rx_shift_reg[7]), .I1(rx_shift_reg[6]), .I2(n4093), 
            .I3(GND_net), .O(n5750));   // src/spi.v(76[8] 221[4])
    defparam i4548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4549_3_lut (.I0(rx_shift_reg[6]), .I1(rx_shift_reg[5]), .I2(n4093), 
            .I3(GND_net), .O(n5751));   // src/spi.v(76[8] 221[4])
    defparam i4549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4550_3_lut (.I0(rx_shift_reg[5]), .I1(rx_shift_reg[4]), .I2(n4093), 
            .I3(GND_net), .O(n5752));   // src/spi.v(76[8] 221[4])
    defparam i4550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4551_3_lut (.I0(rx_shift_reg[4]), .I1(rx_shift_reg[3]), .I2(n4093), 
            .I3(GND_net), .O(n5753));   // src/spi.v(76[8] 221[4])
    defparam i4551_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY led_counter_1106_1179_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(n25_adj_1187), .CO(n10670));
    SB_LUT4 i4552_3_lut (.I0(rx_shift_reg[3]), .I1(rx_shift_reg[2]), .I2(n4093), 
            .I3(GND_net), .O(n5754));   // src/spi.v(76[8] 221[4])
    defparam i4552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4553_3_lut (.I0(rx_shift_reg[2]), .I1(rx_shift_reg[1]), .I2(n4093), 
            .I3(GND_net), .O(n5755));   // src/spi.v(76[8] 221[4])
    defparam i4553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4554_3_lut (.I0(rx_shift_reg[1]), .I1(rx_shift_reg[0]), .I2(n4093), 
            .I3(GND_net), .O(n5756));   // src/spi.v(76[8] 221[4])
    defparam i4554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4571_3_lut (.I0(\REG.mem_63_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n2), .I3(GND_net), .O(n5773));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4573_3_lut (.I0(\REG.mem_63_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n2), .I3(GND_net), .O(n5775));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4574_3_lut (.I0(\REG.mem_63_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n2), .I3(GND_net), .O(n5776));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4575_3_lut (.I0(\REG.mem_63_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n2), .I3(GND_net), .O(n5777));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4576_3_lut (.I0(\REG.mem_63_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n2), .I3(GND_net), .O(n5778));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4577_3_lut (.I0(\REG.mem_63_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n2), .I3(GND_net), .O(n5779));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11062_2_lut (.I0(is_fifo_empty_flag), .I1(tx_uart_active_flag), 
            .I2(GND_net), .I3(GND_net), .O(start_tx_N_64));
    defparam i11062_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i4578_3_lut (.I0(\REG.mem_63_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n2), .I3(GND_net), .O(n5780));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4579_3_lut (.I0(\REG.mem_63_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n2), .I3(GND_net), .O(n5781));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i4579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3919_3_lut (.I0(\REG.mem_26_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n39), .I3(GND_net), .O(n5121));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3918_3_lut (.I0(\REG.mem_26_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n39), .I3(GND_net), .O(n5120));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3917_3_lut (.I0(\REG.mem_26_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n39), .I3(GND_net), .O(n5119));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3916_3_lut (.I0(\REG.mem_26_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n39), .I3(GND_net), .O(n5118));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3915_3_lut (.I0(\REG.mem_26_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n39), .I3(GND_net), .O(n5117));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3914_3_lut (.I0(\REG.mem_26_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n39), .I3(GND_net), .O(n5116));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3913_3_lut (.I0(\REG.mem_26_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n39), .I3(GND_net), .O(n5115));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3912_3_lut (.I0(\REG.mem_26_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n39), .I3(GND_net), .O(n5114));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3911_3_lut (.I0(\REG.mem_26_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n39), .I3(GND_net), .O(n5113));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3910_3_lut (.I0(\REG.mem_26_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n39), .I3(GND_net), .O(n5112));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3909_3_lut (.I0(\REG.mem_26_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n39), .I3(GND_net), .O(n5111));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3908_3_lut (.I0(\REG.mem_26_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n39), .I3(GND_net), .O(n5110));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3907_3_lut (.I0(\REG.mem_26_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n39), .I3(GND_net), .O(n5109));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3906_3_lut (.I0(\REG.mem_26_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n39), .I3(GND_net), .O(n5108));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3905_3_lut (.I0(\REG.mem_26_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n39), .I3(GND_net), .O(n5107));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3904_3_lut (.I0(\REG.mem_26_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n39), .I3(GND_net), .O(n5106));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3871_3_lut (.I0(\REG.mem_23_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n42), .I3(GND_net), .O(n5073));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3870_3_lut (.I0(\REG.mem_23_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n42), .I3(GND_net), .O(n5072));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3869_3_lut (.I0(\REG.mem_23_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n42), .I3(GND_net), .O(n5071));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3868_3_lut (.I0(\REG.mem_23_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n42), .I3(GND_net), .O(n5070));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3867_3_lut (.I0(\REG.mem_23_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n42), .I3(GND_net), .O(n5069));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3866_3_lut (.I0(\REG.mem_23_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n42), .I3(GND_net), .O(n5068));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3865_3_lut (.I0(\REG.mem_23_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n42), .I3(GND_net), .O(n5067));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3864_3_lut (.I0(\REG.mem_23_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n42), .I3(GND_net), .O(n5066));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3863_3_lut (.I0(\REG.mem_23_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n42), .I3(GND_net), .O(n5065));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3862_3_lut (.I0(\REG.mem_23_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n42), .I3(GND_net), .O(n5064));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3861_3_lut (.I0(\REG.mem_23_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n42), .I3(GND_net), .O(n5063));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3860_3_lut (.I0(\REG.mem_23_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n42), .I3(GND_net), .O(n5062));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3859_3_lut (.I0(\REG.mem_23_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n42), .I3(GND_net), .O(n5061));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3858_3_lut (.I0(\REG.mem_23_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n42), .I3(GND_net), .O(n5060));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3857_3_lut (.I0(\REG.mem_23_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n42), .I3(GND_net), .O(n5059));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3856_3_lut (.I0(\REG.mem_23_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n42), .I3(GND_net), .O(n5058));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3241_1_lut_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n4443));   // src/top.v(1064[8] 1131[4])
    defparam i3241_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i3410_2_lut_4_lut (.I0(reset_all), .I1(wr_addr_r[0]), .I2(wr_addr_p1_w[0]), 
            .I3(n7596), .O(n4612));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    defparam i3410_2_lut_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i3429_4_lut_4_lut (.I0(tx_uart_active_flag), .I1(r_SM_Main_adj_1225[1]), 
            .I2(r_SM_Main_adj_1225[2]), .I3(n11339), .O(n4631));   // src/uart_tx.v(38[10] 141[8])
    defparam i3429_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i3495_4_lut_4_lut (.I0(reset_all_w), .I1(wr_addr_r_adj_1249[1]), 
            .I2(wr_addr_r_adj_1249[0]), .I3(n2207), .O(n4697));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i3495_4_lut_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i3804_3_lut (.I0(\REG.mem_19_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n46), .I3(GND_net), .O(n5006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3803_3_lut (.I0(\REG.mem_19_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n46), .I3(GND_net), .O(n5005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3802_3_lut (.I0(\REG.mem_19_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n46), .I3(GND_net), .O(n5004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3801_3_lut (.I0(\REG.mem_19_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n46), .I3(GND_net), .O(n5003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3800_3_lut (.I0(\REG.mem_19_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n46), .I3(GND_net), .O(n5002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3799_3_lut (.I0(\REG.mem_19_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n46), .I3(GND_net), .O(n5001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3798_3_lut (.I0(\REG.mem_19_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n46), .I3(GND_net), .O(n5000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3797_3_lut (.I0(\REG.mem_19_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n46), .I3(GND_net), .O(n4999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3796_3_lut (.I0(\REG.mem_19_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n46), .I3(GND_net), .O(n4998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3795_3_lut (.I0(\REG.mem_19_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n46), .I3(GND_net), .O(n4997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3794_3_lut (.I0(\REG.mem_19_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n46), .I3(GND_net), .O(n4996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3793_3_lut (.I0(\REG.mem_19_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n46), .I3(GND_net), .O(n4995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3792_3_lut (.I0(\REG.mem_19_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n46), .I3(GND_net), .O(n4994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3791_3_lut (.I0(\REG.mem_19_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n46), .I3(GND_net), .O(n4993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3790_3_lut (.I0(\REG.mem_19_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n46), .I3(GND_net), .O(n4992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3789_3_lut (.I0(\REG.mem_19_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n46), .I3(GND_net), .O(n4991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3788_3_lut (.I0(\REG.mem_18_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n47), .I3(GND_net), .O(n4990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3787_3_lut (.I0(\REG.mem_18_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n47), .I3(GND_net), .O(n4989));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3786_3_lut (.I0(\REG.mem_18_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n47), .I3(GND_net), .O(n4988));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3785_3_lut (.I0(\REG.mem_18_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n47), .I3(GND_net), .O(n4987));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3784_3_lut (.I0(\REG.mem_18_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n47), .I3(GND_net), .O(n4986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3783_3_lut (.I0(\REG.mem_18_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n47), .I3(GND_net), .O(n4985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3782_3_lut (.I0(\REG.mem_18_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n47), .I3(GND_net), .O(n4984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3781_3_lut (.I0(\REG.mem_18_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n47), .I3(GND_net), .O(n4983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3780_3_lut (.I0(\REG.mem_18_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n47), .I3(GND_net), .O(n4982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3779_3_lut (.I0(\REG.mem_18_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n47), .I3(GND_net), .O(n4981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3778_3_lut (.I0(\REG.mem_18_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n47), .I3(GND_net), .O(n4980));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3777_3_lut (.I0(\REG.mem_18_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n47), .I3(GND_net), .O(n4979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3776_3_lut (.I0(\REG.mem_18_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n47), .I3(GND_net), .O(n4978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3775_3_lut (.I0(\REG.mem_18_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n47), .I3(GND_net), .O(n4977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3774_3_lut (.I0(\REG.mem_18_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n47), .I3(GND_net), .O(n4976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3452_3_lut (.I0(tx_addr_byte[0]), .I1(tx_data_byte[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4654));   // src/top.v(1064[8] 1131[4])
    defparam i3452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3773_3_lut (.I0(\REG.mem_18_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n47), .I3(GND_net), .O(n4975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3772_3_lut (.I0(\REG.mem_17_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n48), .I3(GND_net), .O(n4974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3771_3_lut (.I0(\REG.mem_17_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n48), .I3(GND_net), .O(n4973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3770_3_lut (.I0(\REG.mem_17_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n48), .I3(GND_net), .O(n4972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3769_3_lut (.I0(\REG.mem_17_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n48), .I3(GND_net), .O(n4971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3768_3_lut (.I0(\REG.mem_17_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n48), .I3(GND_net), .O(n4970));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3767_3_lut (.I0(\REG.mem_17_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n48), .I3(GND_net), .O(n4969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3766_3_lut (.I0(\REG.mem_17_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n48), .I3(GND_net), .O(n4968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3765_3_lut (.I0(\REG.mem_17_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n48), .I3(GND_net), .O(n4967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3764_3_lut (.I0(\REG.mem_17_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n48), .I3(GND_net), .O(n4966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3763_3_lut (.I0(\REG.mem_17_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n48), .I3(GND_net), .O(n4965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3762_3_lut (.I0(\REG.mem_17_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n48), .I3(GND_net), .O(n4964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3761_3_lut (.I0(\REG.mem_17_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n48), .I3(GND_net), .O(n4963));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3760_3_lut (.I0(\REG.mem_17_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n48), .I3(GND_net), .O(n4962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3759_3_lut (.I0(\REG.mem_17_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n48), .I3(GND_net), .O(n4961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3758_3_lut (.I0(\REG.mem_17_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n48), .I3(GND_net), .O(n4960));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3498_4_lut (.I0(RESET_c), .I1(wr_addr_r_adj_1249[2]), .I2(wr_addr_p1_w_adj_1251[2]), 
            .I3(n2207), .O(n4700));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i3498_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i3756_3_lut (.I0(\REG.mem_17_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n48), .I3(GND_net), .O(n4958));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3755_3_lut (.I0(\REG.mem_16_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n49), .I3(GND_net), .O(n4957));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3754_3_lut (.I0(\REG.mem_16_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n49), .I3(GND_net), .O(n4956));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3753_3_lut (.I0(\REG.mem_16_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n49), .I3(GND_net), .O(n4955));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3752_3_lut (.I0(\REG.mem_16_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n49), .I3(GND_net), .O(n4954));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3751_3_lut (.I0(\REG.mem_16_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n49), .I3(GND_net), .O(n4953));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3750_3_lut (.I0(\REG.mem_16_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n49), .I3(GND_net), .O(n4952));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3749_3_lut (.I0(\REG.mem_16_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n49), .I3(GND_net), .O(n4951));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3748_3_lut (.I0(\REG.mem_16_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n49), .I3(GND_net), .O(n4950));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1507_2_lut (.I0(even_byte_flag), .I1(uart_rx_complete_rising_edge), 
            .I2(GND_net), .I3(GND_net), .O(n2679));   // src/top.v(1064[8] 1131[4])
    defparam i1507_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3747_3_lut (.I0(\REG.mem_16_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n49), .I3(GND_net), .O(n4949));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3746_3_lut (.I0(\REG.mem_16_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n49), .I3(GND_net), .O(n4948));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3745_3_lut (.I0(\REG.mem_16_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n49), .I3(GND_net), .O(n4947));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9054_2_lut_3_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(reset_clk_counter[1]), .I3(GND_net), .O(n10562));   // src/top.v(259[27:51])
    defparam i9054_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i3744_3_lut (.I0(\REG.mem_16_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n49), .I3(GND_net), .O(n4946));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3743_3_lut (.I0(\REG.mem_16_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n49), .I3(GND_net), .O(n4945));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3742_3_lut (.I0(\REG.mem_16_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n49), .I3(GND_net), .O(n4944));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3741_3_lut (.I0(\REG.mem_16_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n49), .I3(GND_net), .O(n4943));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3740_3_lut (.I0(\REG.mem_16_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n49), .I3(GND_net), .O(n4942));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3739_3_lut (.I0(\REG.mem_15_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n50), .I3(GND_net), .O(n4941));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(reset_all_w_N_61), .I1(reset_clk_counter[0]), 
            .I2(reset_clk_counter[1]), .I3(GND_net), .O(n10798));   // src/top.v(259[27:51])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i3738_3_lut (.I0(\REG.mem_15_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n50), .I3(GND_net), .O(n4940));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3737_3_lut (.I0(\REG.mem_15_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n50), .I3(GND_net), .O(n4939));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3736_3_lut (.I0(\REG.mem_15_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n50), .I3(GND_net), .O(n4938));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3735_3_lut (.I0(\REG.mem_15_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n50), .I3(GND_net), .O(n4937));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3734_3_lut (.I0(\REG.mem_15_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n50), .I3(GND_net), .O(n4936));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3733_3_lut (.I0(\REG.mem_15_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n50), .I3(GND_net), .O(n4935));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3732_3_lut (.I0(\REG.mem_15_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n50), .I3(GND_net), .O(n4934));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3731_3_lut (.I0(\REG.mem_15_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n50), .I3(GND_net), .O(n4933));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3730_3_lut (.I0(\REG.mem_15_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n50), .I3(GND_net), .O(n4932));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3729_3_lut (.I0(\REG.mem_15_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n50), .I3(GND_net), .O(n4931));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3728_3_lut (.I0(\REG.mem_15_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n50), .I3(GND_net), .O(n4930));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3727_3_lut (.I0(\REG.mem_15_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n50), .I3(GND_net), .O(n4929));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3726_3_lut (.I0(\REG.mem_15_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n50), .I3(GND_net), .O(n4928));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3725_3_lut (.I0(\REG.mem_15_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n50), .I3(GND_net), .O(n4927));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3724_3_lut (.I0(\REG.mem_15_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n50), .I3(GND_net), .O(n4926));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3723_3_lut (.I0(\REG.mem_14_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n51), .I3(GND_net), .O(n4925));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3722_3_lut (.I0(\REG.mem_14_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n51), .I3(GND_net), .O(n4924));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3721_3_lut (.I0(\REG.mem_14_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n51), .I3(GND_net), .O(n4923));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3720_3_lut (.I0(\REG.mem_14_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n51), .I3(GND_net), .O(n4922));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3719_3_lut (.I0(\REG.mem_14_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n51), .I3(GND_net), .O(n4921));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3718_3_lut (.I0(\REG.mem_14_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n51), .I3(GND_net), .O(n4920));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3717_3_lut (.I0(\REG.mem_14_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n51), .I3(GND_net), .O(n4919));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3716_3_lut (.I0(\REG.mem_14_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n51), .I3(GND_net), .O(n4918));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3715_3_lut (.I0(\REG.mem_14_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n51), .I3(GND_net), .O(n4917));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3714_3_lut (.I0(\REG.mem_14_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n51), .I3(GND_net), .O(n4916));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3713_3_lut (.I0(\REG.mem_14_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n51), .I3(GND_net), .O(n4915));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3712_3_lut (.I0(\REG.mem_14_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n51), .I3(GND_net), .O(n4914));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3711_3_lut (.I0(\REG.mem_14_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n51), .I3(GND_net), .O(n4913));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3710_3_lut (.I0(\REG.mem_14_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n51), .I3(GND_net), .O(n4912));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3709_3_lut (.I0(\REG.mem_14_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n51), .I3(GND_net), .O(n4911));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3708_3_lut (.I0(\REG.mem_14_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n51), .I3(GND_net), .O(n4910));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3707_3_lut (.I0(\REG.mem_13_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n52), .I3(GND_net), .O(n4909));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3706_3_lut (.I0(\REG.mem_13_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n52), .I3(GND_net), .O(n4908));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3705_3_lut (.I0(\REG.mem_13_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n52), .I3(GND_net), .O(n4907));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3704_3_lut (.I0(\REG.mem_13_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n52), .I3(GND_net), .O(n4906));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3703_3_lut (.I0(\REG.mem_13_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n52), .I3(GND_net), .O(n4905));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3702_3_lut (.I0(\REG.mem_13_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n52), .I3(GND_net), .O(n4904));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3701_3_lut (.I0(\REG.mem_13_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n52), .I3(GND_net), .O(n4903));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3700_3_lut (.I0(\REG.mem_13_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n52), .I3(GND_net), .O(n4902));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3699_3_lut (.I0(\REG.mem_13_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n52), .I3(GND_net), .O(n4901));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3698_3_lut (.I0(\REG.mem_13_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n52), .I3(GND_net), .O(n4900));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3697_3_lut (.I0(\REG.mem_13_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n52), .I3(GND_net), .O(n4899));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3696_3_lut (.I0(\REG.mem_13_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n52), .I3(GND_net), .O(n4898));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3695_3_lut (.I0(\REG.mem_13_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n52), .I3(GND_net), .O(n4897));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3694_3_lut (.I0(\REG.mem_13_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n52), .I3(GND_net), .O(n4896));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3694_3_lut.LUT_INIT = 16'hcaca;
    fifo_dc_32_lut_gen2 fifo_dc_32_lut_gen_inst (.\REG.mem_58_4 (\REG.mem_58_4 ), 
            .GND_net(GND_net), .\REG.mem_14_8 (\REG.mem_14_8 ), .\REG.mem_15_8 (\REG.mem_15_8 ), 
            .\dc32_fifo_data_in[10] (dc32_fifo_data_in[10]), .\dc32_fifo_data_in[9] (dc32_fifo_data_in[9]), 
            .DEBUG_6_c_c(DEBUG_6_c_c), .\REG.mem_13_8 (\REG.mem_13_8 ), 
            .\REG.mem_12_8 (\REG.mem_12_8 ), .\dc32_fifo_data_in[8] (dc32_fifo_data_in[8]), 
            .\REG.mem_10_10 (\REG.mem_10_10 ), .\REG.mem_11_10 (\REG.mem_11_10 ), 
            .\REG.mem_9_10 (\REG.mem_9_10 ), .\REG.mem_8_10 (\REG.mem_8_10 ), 
            .t_rd_fifo_en_w(t_rd_fifo_en_w), .\REG.out_raw[0] (\REG.out_raw [0]), 
            .SLM_CLK_c(SLM_CLK_c), .\dc32_fifo_data_in[7] (dc32_fifo_data_in[7]), 
            .\REG.mem_10_13 (\REG.mem_10_13 ), .\REG.mem_11_13 (\REG.mem_11_13 ), 
            .\REG.mem_9_13 (\REG.mem_9_13 ), .\REG.mem_8_13 (\REG.mem_8_13 ), 
            .\dc32_fifo_data_in[6] (dc32_fifo_data_in[6]), .DEBUG_9_c(DEBUG_9_c), 
            .n7596(n7596), .\wr_addr_nxt_c[4] (wr_addr_nxt_c[4]), .\REG.mem_26_14 (\REG.mem_26_14 ), 
            .\dc32_fifo_data_in[5] (dc32_fifo_data_in[5]), .\REG.mem_42_2 (\REG.mem_42_2 ), 
            .\REG.mem_43_2 (\REG.mem_43_2 ), .\REG.mem_41_2 (\REG.mem_41_2 ), 
            .\REG.mem_40_2 (\REG.mem_40_2 ), .\REG.mem_14_10 (\REG.mem_14_10 ), 
            .\REG.mem_15_10 (\REG.mem_15_10 ), .reset_all(reset_all), .\REG.mem_55_8 (\REG.mem_55_8 ), 
            .\REG.mem_13_10 (\REG.mem_13_10 ), .\REG.mem_12_10 (\REG.mem_12_10 ), 
            .\dc32_fifo_data_in[4] (dc32_fifo_data_in[4]), .\REG.mem_42_3 (\REG.mem_42_3 ), 
            .\REG.mem_43_3 (\REG.mem_43_3 ), .\REG.mem_41_3 (\REG.mem_41_3 ), 
            .\REG.mem_40_3 (\REG.mem_40_3 ), .\rd_grey_sync_r[0] (rd_grey_sync_r[0]), 
            .\dc32_fifo_data_in[3] (dc32_fifo_data_in[3]), .\REG.mem_58_8 (\REG.mem_58_8 ), 
            .DEBUG_5_c(DEBUG_5_c), .wr_grey_sync_r({wr_grey_sync_r}), .\REG.mem_48_5 (\REG.mem_48_5 ), 
            .\REG.mem_49_5 (\REG.mem_49_5 ), .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .dc32_fifo_almost_empty(dc32_fifo_almost_empty), .\dc32_fifo_data_in[2] (dc32_fifo_data_in[2]), 
            .\REG.mem_55_11 (\REG.mem_55_11 ), .\REG.mem_50_5 (\REG.mem_50_5 ), 
            .\REG.mem_51_5 (\REG.mem_51_5 ), .\dc32_fifo_data_in[1] (dc32_fifo_data_in[1]), 
            .\REG.mem_55_5 (\REG.mem_55_5 ), .\REG.mem_63_4 (\REG.mem_63_4 ), 
            .\REG.mem_23_11 (\REG.mem_23_11 ), .\dc32_fifo_data_in[0] (dc32_fifo_data_in[0]), 
            .\REG.mem_10_12 (\REG.mem_10_12 ), .\REG.mem_11_12 (\REG.mem_11_12 ), 
            .\REG.mem_9_12 (\REG.mem_9_12 ), .\REG.mem_8_12 (\REG.mem_8_12 ), 
            .\REG.mem_38_11 (\REG.mem_38_11 ), .\REG.mem_39_11 (\REG.mem_39_11 ), 
            .\REG.mem_37_11 (\REG.mem_37_11 ), .\REG.mem_36_11 (\REG.mem_36_11 ), 
            .\REG.mem_14_12 (\REG.mem_14_12 ), .\REG.mem_15_12 (\REG.mem_15_12 ), 
            .\REG.mem_14_13 (\REG.mem_14_13 ), .\REG.mem_15_13 (\REG.mem_15_13 ), 
            .\REG.mem_6_12 (\REG.mem_6_12 ), .\REG.mem_7_12 (\REG.mem_7_12 ), 
            .\REG.mem_4_12 (\REG.mem_4_12 ), .\REG.mem_5_12 (\REG.mem_5_12 ), 
            .\REG.mem_13_13 (\REG.mem_13_13 ), .\REG.mem_12_13 (\REG.mem_12_13 ), 
            .\REG.mem_13_12 (\REG.mem_13_12 ), .\REG.mem_12_12 (\REG.mem_12_12 ), 
            .\REG.mem_23_15 (\REG.mem_23_15 ), .\REG.mem_18_12 (\REG.mem_18_12 ), 
            .\REG.mem_19_12 (\REG.mem_19_12 ), .\REG.mem_6_8 (\REG.mem_6_8 ), 
            .\REG.mem_7_8 (\REG.mem_7_8 ), .\REG.mem_17_12 (\REG.mem_17_12 ), 
            .\REG.mem_16_12 (\REG.mem_16_12 ), .\wr_addr_nxt_c[2] (wr_addr_nxt_c[2]), 
            .\REG.mem_26_0 (\REG.mem_26_0 ), .\REG.mem_42_10 (\REG.mem_42_10 ), 
            .\REG.mem_43_10 (\REG.mem_43_10 ), .\REG.mem_18_8 (\REG.mem_18_8 ), 
            .\REG.mem_19_8 (\REG.mem_19_8 ), .\REG.mem_14_15 (\REG.mem_14_15 ), 
            .\REG.mem_15_15 (\REG.mem_15_15 ), .\REG.mem_17_8 (\REG.mem_17_8 ), 
            .\REG.mem_16_8 (\REG.mem_16_8 ), .\REG.mem_41_10 (\REG.mem_41_10 ), 
            .\REG.mem_40_10 (\REG.mem_40_10 ), .n60(n60), .\REG.mem_18_13 (\REG.mem_18_13 ), 
            .\REG.mem_19_13 (\REG.mem_19_13 ), .\REG.mem_17_13 (\REG.mem_17_13 ), 
            .\REG.mem_16_13 (\REG.mem_16_13 ), .n28(n28), .\REG.mem_13_15 (\REG.mem_13_15 ), 
            .\REG.mem_12_15 (\REG.mem_12_15 ), .\REG.mem_26_3 (\REG.mem_26_3 ), 
            .\REG.mem_46_6 (\REG.mem_46_6 ), .\REG.mem_47_6 (\REG.mem_47_6 ), 
            .\REG.mem_45_6 (\REG.mem_45_6 ), .\REG.mem_44_6 (\REG.mem_44_6 ), 
            .\REG.mem_63_8 (\REG.mem_63_8 ), .\REG.mem_46_2 (\REG.mem_46_2 ), 
            .\REG.mem_47_2 (\REG.mem_47_2 ), .\REG.mem_45_2 (\REG.mem_45_2 ), 
            .\REG.mem_44_2 (\REG.mem_44_2 ), .\dc32_fifo_data_in[15] (dc32_fifo_data_in[15]), 
            .\dc32_fifo_data_in[14] (dc32_fifo_data_in[14]), .\REG.mem_6_7 (\REG.mem_6_7 ), 
            .\REG.mem_7_7 (\REG.mem_7_7 ), .\dc32_fifo_data_in[13] (dc32_fifo_data_in[13]), 
            .\REG.mem_46_11 (\REG.mem_46_11 ), .\REG.mem_47_11 (\REG.mem_47_11 ), 
            .\dc32_fifo_data_in[12] (dc32_fifo_data_in[12]), .\REG.mem_5_7 (\REG.mem_5_7 ), 
            .\REG.mem_4_7 (\REG.mem_4_7 ), .\dc32_fifo_data_in[11] (dc32_fifo_data_in[11]), 
            .\REG.mem_45_11 (\REG.mem_45_11 ), .\REG.mem_44_11 (\REG.mem_44_11 ), 
            .\REG.mem_23_13 (\REG.mem_23_13 ), .\REG.mem_58_5 (\REG.mem_58_5 ), 
            .\REG.mem_23_8 (\REG.mem_23_8 ), .\REG.mem_46_3 (\REG.mem_46_3 ), 
            .\REG.mem_47_3 (\REG.mem_47_3 ), .\REG.mem_10_7 (\REG.mem_10_7 ), 
            .\REG.mem_11_7 (\REG.mem_11_7 ), .\REG.mem_45_3 (\REG.mem_45_3 ), 
            .\REG.mem_44_3 (\REG.mem_44_3 ), .\REG.mem_8_2 (\REG.mem_8_2 ), 
            .\REG.mem_9_2 (\REG.mem_9_2 ), .\REG.mem_9_7 (\REG.mem_9_7 ), 
            .\REG.mem_8_7 (\REG.mem_8_7 ), .\REG.mem_31_14 (\REG.mem_31_14 ), 
            .\REG.mem_10_2 (\REG.mem_10_2 ), .\REG.mem_11_2 (\REG.mem_11_2 ), 
            .\REG.mem_58_13 (\REG.mem_58_13 ), .\REG.mem_26_8 (\REG.mem_26_8 ), 
            .\REG.mem_14_2 (\REG.mem_14_2 ), .\REG.mem_15_2 (\REG.mem_15_2 ), 
            .\REG.mem_12_2 (\REG.mem_12_2 ), .\REG.mem_13_2 (\REG.mem_13_2 ), 
            .\REG.mem_14_7 (\REG.mem_14_7 ), .\REG.mem_15_7 (\REG.mem_15_7 ), 
            .\REG.mem_13_7 (\REG.mem_13_7 ), .\REG.mem_12_7 (\REG.mem_12_7 ), 
            .\REG.mem_26_13 (\REG.mem_26_13 ), .\REG.mem_6_3 (\REG.mem_6_3 ), 
            .\REG.mem_7_3 (\REG.mem_7_3 ), .\REG.mem_5_3 (\REG.mem_5_3 ), 
            .\REG.mem_4_3 (\REG.mem_4_3 ), .\REG.mem_40_1 (\REG.mem_40_1 ), 
            .\REG.mem_41_1 (\REG.mem_41_1 ), .\REG.mem_14_5 (\REG.mem_14_5 ), 
            .\REG.mem_15_5 (\REG.mem_15_5 ), .\REG.mem_13_5 (\REG.mem_13_5 ), 
            .\REG.mem_12_5 (\REG.mem_12_5 ), .\REG.mem_42_1 (\REG.mem_42_1 ), 
            .\REG.mem_43_1 (\REG.mem_43_1 ), .\REG.mem_46_1 (\REG.mem_46_1 ), 
            .\REG.mem_47_1 (\REG.mem_47_1 ), .\REG.mem_44_1 (\REG.mem_44_1 ), 
            .\REG.mem_45_1 (\REG.mem_45_1 ), .\REG.mem_31_8 (\REG.mem_31_8 ), 
            .\REG.mem_26_10 (\REG.mem_26_10 ), .\REG.mem_18_2 (\REG.mem_18_2 ), 
            .\REG.mem_19_2 (\REG.mem_19_2 ), .\REG.mem_31_3 (\REG.mem_31_3 ), 
            .\REG.mem_17_2 (\REG.mem_17_2 ), .\REG.mem_16_2 (\REG.mem_16_2 ), 
            .n61(n61), .\REG.mem_63_13 (\REG.mem_63_13 ), .n34(n34), .n29(n29), 
            .\REG.mem_50_6 (\REG.mem_50_6 ), .\REG.mem_51_6 (\REG.mem_51_6 ), 
            .n58(n58), .\REG.mem_6_14 (\REG.mem_6_14 ), .\REG.mem_7_14 (\REG.mem_7_14 ), 
            .n26(n26), .\REG.mem_6_10 (\REG.mem_6_10 ), .\REG.mem_7_10 (\REG.mem_7_10 ), 
            .\REG.mem_4_10 (\REG.mem_4_10 ), .\REG.mem_5_10 (\REG.mem_5_10 ), 
            .\REG.mem_4_14 (\REG.mem_4_14 ), .\REG.mem_5_14 (\REG.mem_5_14 ), 
            .n5896(n5896), .VCC_net(VCC_net), .\fifo_data_out[6] (fifo_data_out[6]), 
            .n5893(n5893), .\fifo_data_out[5] (fifo_data_out[5]), .\REG.mem_16_10 (\REG.mem_16_10 ), 
            .\REG.mem_17_10 (\REG.mem_17_10 ), .\REG.mem_18_10 (\REG.mem_18_10 ), 
            .\REG.mem_19_10 (\REG.mem_19_10 ), .n11119(n11119), .\fifo_data_out[7] (fifo_data_out[7]), 
            .\REG.mem_18_7 (\REG.mem_18_7 ), .\REG.mem_19_7 (\REG.mem_19_7 ), 
            .n11139(n11139), .\fifo_data_out[3] (fifo_data_out[3]), .\REG.mem_17_7 (\REG.mem_17_7 ), 
            .\REG.mem_16_7 (\REG.mem_16_7 ), .\REG.mem_50_2 (\REG.mem_50_2 ), 
            .\REG.mem_51_2 (\REG.mem_51_2 ), .\REG.mem_46_0 (\REG.mem_46_0 ), 
            .\REG.mem_47_0 (\REG.mem_47_0 ), .\REG.mem_46_9 (\REG.mem_46_9 ), 
            .\REG.mem_47_9 (\REG.mem_47_9 ), .\REG.mem_45_9 (\REG.mem_45_9 ), 
            .\REG.mem_44_9 (\REG.mem_44_9 ), .\REG.mem_49_6 (\REG.mem_49_6 ), 
            .\REG.mem_48_6 (\REG.mem_48_6 ), .\REG.mem_49_2 (\REG.mem_49_2 ), 
            .\REG.mem_48_2 (\REG.mem_48_2 ), .n11097(n11097), .\fifo_data_out[8] (fifo_data_out[8]), 
            .n5854(n5854), .\fifo_data_out[0] (fifo_data_out[0]), .\REG.mem_5_8 (\REG.mem_5_8 ), 
            .\REG.mem_4_8 (\REG.mem_4_8 ), .\REG.mem_6_11 (\REG.mem_6_11 ), 
            .\REG.mem_7_11 (\REG.mem_7_11 ), .\REG.mem_58_1 (\REG.mem_58_1 ), 
            .\REG.mem_26_15 (\REG.mem_26_15 ), .n11095(n11095), .\fifo_data_out[9] (fifo_data_out[9]), 
            .\REG.mem_23_7 (\REG.mem_23_7 ), .n11143(n11143), .\fifo_data_out[1] (fifo_data_out[1]), 
            .n11141(n11141), .\fifo_data_out[2] (fifo_data_out[2]), .n11089(n11089), 
            .\fifo_data_out[10] (fifo_data_out[10]), .n11135(n11135), .\fifo_data_out[11] (fifo_data_out[11]), 
            .\REG.mem_50_3 (\REG.mem_50_3 ), .\REG.mem_51_3 (\REG.mem_51_3 ), 
            .\REG.mem_31_13 (\REG.mem_31_13 ), .\REG.mem_49_3 (\REG.mem_49_3 ), 
            .\REG.mem_48_3 (\REG.mem_48_3 ), .\REG.mem_10_9 (\REG.mem_10_9 ), 
            .\REG.mem_11_9 (\REG.mem_11_9 ), .\REG.mem_9_9 (\REG.mem_9_9 ), 
            .\REG.mem_8_9 (\REG.mem_8_9 ), .\REG.mem_23_10 (\REG.mem_23_10 ), 
            .\REG.mem_26_1 (\REG.mem_26_1 ), .n47(n47), .n5789(n5789), 
            .\REG.mem_63_15 (\REG.mem_63_15 ), .n5788(n5788), .\REG.mem_63_14 (\REG.mem_63_14 ), 
            .n5787(n5787), .\REG.mem_31_11 (\REG.mem_31_11 ), .\REG.mem_5_11 (\REG.mem_5_11 ), 
            .\REG.mem_4_11 (\REG.mem_4_11 ), .\REG.mem_31_1 (\REG.mem_31_1 ), 
            .\REG.mem_23_12 (\REG.mem_23_12 ), .n5786(n5786), .\REG.mem_63_12 (\REG.mem_63_12 ), 
            .n5785(n5785), .\REG.mem_63_11 (\REG.mem_63_11 ), .n5784(n5784), 
            .\REG.mem_63_10 (\REG.mem_63_10 ), .n5783(n5783), .\REG.mem_63_9 (\REG.mem_63_9 ), 
            .\REG.mem_14_9 (\REG.mem_14_9 ), .\REG.mem_15_9 (\REG.mem_15_9 ), 
            .n5782(n5782), .n5781(n5781), .\REG.mem_63_7 (\REG.mem_63_7 ), 
            .n5780(n5780), .\REG.mem_63_6 (\REG.mem_63_6 ), .n5779(n5779), 
            .\REG.mem_63_5 (\REG.mem_63_5 ), .n5778(n5778), .n5777(n5777), 
            .\REG.mem_63_3 (\REG.mem_63_3 ), .n5776(n5776), .\REG.mem_63_2 (\REG.mem_63_2 ), 
            .n5775(n5775), .\REG.mem_63_1 (\REG.mem_63_1 ), .n11133(n11133), 
            .\fifo_data_out[12] (fifo_data_out[12]), .n5773(n5773), .\REG.mem_63_0 (\REG.mem_63_0 ), 
            .\REG.mem_13_9 (\REG.mem_13_9 ), .\REG.mem_12_9 (\REG.mem_12_9 ), 
            .\REG.mem_38_10 (\REG.mem_38_10 ), .\REG.mem_39_10 (\REG.mem_39_10 ), 
            .n15(n15_adj_1184), .\REG.mem_36_10 (\REG.mem_36_10 ), .\REG.mem_37_10 (\REG.mem_37_10 ), 
            .\REG.mem_8_1 (\REG.mem_8_1 ), .\REG.mem_9_1 (\REG.mem_9_1 ), 
            .\REG.mem_10_1 (\REG.mem_10_1 ), .\REG.mem_11_1 (\REG.mem_11_1 ), 
            .n11137(n11137), .\fifo_data_out[4] (fifo_data_out[4]), .\REG.mem_14_1 (\REG.mem_14_1 ), 
            .\REG.mem_15_1 (\REG.mem_15_1 ), .\REG.mem_12_1 (\REG.mem_12_1 ), 
            .\REG.mem_13_1 (\REG.mem_13_1 ), .\REG.mem_38_12 (\REG.mem_38_12 ), 
            .\REG.mem_39_12 (\REG.mem_39_12 ), .\REG.mem_36_12 (\REG.mem_36_12 ), 
            .\REG.mem_37_12 (\REG.mem_37_12 ), .\REG.mem_38_5 (\REG.mem_38_5 ), 
            .\REG.mem_39_5 (\REG.mem_39_5 ), .n5709(n5709), .rp_sync1_r({rp_sync1_r}), 
            .n5708(n5708), .n5707(n5707), .n5706(n5706), .n5705(n5705), 
            .\REG.mem_36_5 (\REG.mem_36_5 ), .\REG.mem_37_5 (\REG.mem_37_5 ), 
            .\REG.mem_48_12 (\REG.mem_48_12 ), .\REG.mem_49_12 (\REG.mem_49_12 ), 
            .\wr_addr_r[0] (wr_addr_r[0]), .\REG.mem_50_12 (\REG.mem_50_12 ), 
            .\REG.mem_51_12 (\REG.mem_51_12 ), .\REG.mem_55_12 (\REG.mem_55_12 ), 
            .\wr_addr_p1_w[6] (wr_addr_p1_w[6]), .n5704(n5704), .\rd_sig_diff0_w[1] (rd_sig_diff0_w[1]), 
            .n5686(n5686), .n5685(n5685), .n5684(n5684), .n5683(n5683), 
            .n5682(n5682), .\REG.mem_58_15 (\REG.mem_58_15 ), .n5681(n5681), 
            .\REG.mem_58_14 (\REG.mem_58_14 ), .n5680(n5680), .n5679(n5679), 
            .\REG.mem_58_12 (\REG.mem_58_12 ), .n5678(n5678), .\REG.mem_58_11 (\REG.mem_58_11 ), 
            .n5677(n5677), .\REG.mem_58_10 (\REG.mem_58_10 ), .n5676(n5676), 
            .\REG.mem_58_9 (\REG.mem_58_9 ), .n5675(n5675), .n5674(n5674), 
            .\REG.mem_58_7 (\REG.mem_58_7 ), .n5673(n5673), .\REG.mem_58_6 (\REG.mem_58_6 ), 
            .\REG.mem_26_7 (\REG.mem_26_7 ), .\rd_sig_diff0_w[0] (rd_sig_diff0_w[0]), 
            .n5672(n5672), .n5671(n5671), .n5670(n5670), .\REG.mem_58_3 (\REG.mem_58_3 ), 
            .n5669(n5669), .\REG.mem_58_2 (\REG.mem_58_2 ), .n5668(n5668), 
            .n5667(n5667), .\REG.mem_58_0 (\REG.mem_58_0 ), .n5666(n5666), 
            .n5665(n5665), .n5664(n5664), .n5662(n5662), .n5660(n5660), 
            .\rd_addr_r[6] (rd_addr_r[6]), .\REG.out_raw[15] (\REG.out_raw [15]), 
            .\REG.out_raw[14] (\REG.out_raw [14]), .\REG.out_raw[13] (\REG.out_raw [13]), 
            .\REG.out_raw[12] (\REG.out_raw [12]), .\REG.out_raw[11] (\REG.out_raw [11]), 
            .\REG.out_raw[10] (\REG.out_raw [10]), .\REG.out_raw[9] (\REG.out_raw [9]), 
            .\REG.out_raw[8] (\REG.out_raw [8]), .\REG.out_raw[7] (\REG.out_raw [7]), 
            .\REG.out_raw[6] (\REG.out_raw [6]), .\REG.out_raw[5] (\REG.out_raw [5]), 
            .\REG.out_raw[4] (\REG.out_raw [4]), .\REG.out_raw[3] (\REG.out_raw [3]), 
            .\REG.out_raw[2] (\REG.out_raw [2]), .\REG.out_raw[1] (\REG.out_raw [1]), 
            .\REG.mem_31_7 (\REG.mem_31_7 ), .\REG.mem_42_11 (\REG.mem_42_11 ), 
            .\REG.mem_43_11 (\REG.mem_43_11 ), .\REG.mem_41_11 (\REG.mem_41_11 ), 
            .\REG.mem_40_11 (\REG.mem_40_11 ), .n2(n2), .\REG.mem_6_1 (\REG.mem_6_1 ), 
            .\REG.mem_7_1 (\REG.mem_7_1 ), .\REG.mem_4_1 (\REG.mem_4_1 ), 
            .\REG.mem_5_1 (\REG.mem_5_1 ), .\REG.mem_38_4 (\REG.mem_38_4 ), 
            .\REG.mem_39_4 (\REG.mem_39_4 ), .\REG.mem_16_1 (\REG.mem_16_1 ), 
            .\REG.mem_17_1 (\REG.mem_17_1 ), .\REG.mem_37_4 (\REG.mem_37_4 ), 
            .\REG.mem_36_4 (\REG.mem_36_4 ), .\REG.mem_55_2 (\REG.mem_55_2 ), 
            .\REG.mem_18_1 (\REG.mem_18_1 ), .\REG.mem_19_1 (\REG.mem_19_1 ), 
            .n5626(n5626), .\REG.mem_55_15 (\REG.mem_55_15 ), .\REG.mem_23_1 (\REG.mem_23_1 ), 
            .\REG.mem_31_10 (\REG.mem_31_10 ), .n5625(n5625), .\REG.mem_55_14 (\REG.mem_55_14 ), 
            .n5624(n5624), .\REG.mem_55_13 (\REG.mem_55_13 ), .n5623(n5623), 
            .n5622(n5622), .n5621(n5621), .\REG.mem_55_10 (\REG.mem_55_10 ), 
            .n5620(n5620), .\REG.mem_55_9 (\REG.mem_55_9 ), .n5619(n5619), 
            .n5618(n5618), .\REG.mem_55_7 (\REG.mem_55_7 ), .n5617(n5617), 
            .\REG.mem_55_6 (\REG.mem_55_6 ), .n5616(n5616), .n5615(n5615), 
            .\REG.mem_55_4 (\REG.mem_55_4 ), .n5614(n5614), .\REG.mem_55_3 (\REG.mem_55_3 ), 
            .n5613(n5613), .n5612(n5612), .\REG.mem_55_1 (\REG.mem_55_1 ), 
            .n11073(n11073), .\fifo_data_out[13] (fifo_data_out[13]), .n5610(n5610), 
            .\REG.mem_55_0 (\REG.mem_55_0 ), .n5609(n5609), .wp_sync1_r({wp_sync1_r}), 
            .n5608(n5608), .n5607(n5607), .n5606(n5606), .n5605(n5605), 
            .n5604(n5604), .n5603(n5603), .n5586(n5586), .n5585(n5585), 
            .n5584(n5584), .n5583(n5583), .n5582(n5582), .n11071(n11071), 
            .\fifo_data_out[14] (fifo_data_out[14]), .\REG.mem_38_1 (\REG.mem_38_1 ), 
            .\REG.mem_39_1 (\REG.mem_39_1 ), .\REG.mem_36_1 (\REG.mem_36_1 ), 
            .\REG.mem_37_1 (\REG.mem_37_1 ), .\REG.mem_6_2 (\REG.mem_6_2 ), 
            .\REG.mem_7_2 (\REG.mem_7_2 ), .\REG.mem_5_2 (\REG.mem_5_2 ), 
            .\REG.mem_4_2 (\REG.mem_4_2 ), .n5548(n5548), .\REG.mem_51_15 (\REG.mem_51_15 ), 
            .n5547(n5547), .\REG.mem_51_14 (\REG.mem_51_14 ), .n5546(n5546), 
            .\REG.mem_51_13 (\REG.mem_51_13 ), .n5545(n5545), .n5544(n5544), 
            .\REG.mem_51_11 (\REG.mem_51_11 ), .n5543(n5543), .\REG.mem_51_10 (\REG.mem_51_10 ), 
            .n5542(n5542), .\REG.mem_51_9 (\REG.mem_51_9 ), .n5541(n5541), 
            .\REG.mem_51_8 (\REG.mem_51_8 ), .n5540(n5540), .\REG.mem_51_7 (\REG.mem_51_7 ), 
            .n5539(n5539), .n5538(n5538), .n5537(n5537), .\REG.mem_51_4 (\REG.mem_51_4 ), 
            .n5536(n5536), .n5535(n5535), .n5534(n5534), .\REG.mem_51_1 (\REG.mem_51_1 ), 
            .n5533(n5533), .\REG.mem_51_0 (\REG.mem_51_0 ), .n5532(n5532), 
            .\REG.mem_50_15 (\REG.mem_50_15 ), .\REG.mem_48_1 (\REG.mem_48_1 ), 
            .\REG.mem_49_1 (\REG.mem_49_1 ), .n5531(n5531), .\REG.mem_50_14 (\REG.mem_50_14 ), 
            .n5530(n5530), .\REG.mem_50_13 (\REG.mem_50_13 ), .n5529(n5529), 
            .n5528(n5528), .\REG.mem_50_11 (\REG.mem_50_11 ), .n5527(n5527), 
            .\REG.mem_50_10 (\REG.mem_50_10 ), .n5526(n5526), .\REG.mem_50_9 (\REG.mem_50_9 ), 
            .n5525(n5525), .\REG.mem_50_8 (\REG.mem_50_8 ), .n5524(n5524), 
            .\REG.mem_50_7 (\REG.mem_50_7 ), .n5523(n5523), .n5522(n5522), 
            .n5521(n5521), .\REG.mem_50_4 (\REG.mem_50_4 ), .n5520(n5520), 
            .n5519(n5519), .n5518(n5518), .\REG.mem_50_1 (\REG.mem_50_1 ), 
            .n5517(n5517), .\REG.mem_50_0 (\REG.mem_50_0 ), .n5516(n5516), 
            .\REG.mem_49_15 (\REG.mem_49_15 ), .n5515(n5515), .\REG.mem_49_14 (\REG.mem_49_14 ), 
            .\REG.mem_31_12 (\REG.mem_31_12 ), .\REG.mem_26_11 (\REG.mem_26_11 ), 
            .n5514(n5514), .\REG.mem_49_13 (\REG.mem_49_13 ), .n5513(n5513), 
            .n5512(n5512), .\REG.mem_49_11 (\REG.mem_49_11 ), .n5511(n5511), 
            .\REG.mem_49_10 (\REG.mem_49_10 ), .n5510(n5510), .\REG.mem_49_9 (\REG.mem_49_9 ), 
            .n5509(n5509), .\REG.mem_49_8 (\REG.mem_49_8 ), .n5508(n5508), 
            .\REG.mem_49_7 (\REG.mem_49_7 ), .n5507(n5507), .n5506(n5506), 
            .n5505(n5505), .\REG.mem_49_4 (\REG.mem_49_4 ), .n5504(n5504), 
            .n5503(n5503), .n5502(n5502), .n5501(n5501), .\REG.mem_49_0 (\REG.mem_49_0 ), 
            .\REG.mem_31_0 (\REG.mem_31_0 ), .\REG.mem_26_4 (\REG.mem_26_4 ), 
            .n5492(n5492), .\REG.mem_48_15 (\REG.mem_48_15 ), .n5491(n5491), 
            .n5490(n5490), .\REG.mem_48_14 (\REG.mem_48_14 ), .n5489(n5489), 
            .\REG.mem_48_13 (\REG.mem_48_13 ), .n5488(n5488), .n5487(n5487), 
            .\REG.mem_48_11 (\REG.mem_48_11 ), .n5486(n5486), .\REG.mem_48_10 (\REG.mem_48_10 ), 
            .n5485(n5485), .\REG.mem_48_9 (\REG.mem_48_9 ), .n5484(n5484), 
            .\REG.mem_48_8 (\REG.mem_48_8 ), .n5483(n5483), .\REG.mem_48_7 (\REG.mem_48_7 ), 
            .\REG.mem_46_10 (\REG.mem_46_10 ), .\REG.mem_47_10 (\REG.mem_47_10 ), 
            .n5482(n5482), .n5481(n5481), .n5480(n5480), .\REG.mem_48_4 (\REG.mem_48_4 ), 
            .n5479(n5479), .n5478(n5478), .n5477(n5477), .n5476(n5476), 
            .\REG.mem_48_0 (\REG.mem_48_0 ), .n5474(n5474), .n5472(n5472), 
            .\REG.mem_47_15 (\REG.mem_47_15 ), .n5471(n5471), .\REG.mem_47_14 (\REG.mem_47_14 ), 
            .n5470(n5470), .\REG.mem_47_13 (\REG.mem_47_13 ), .n5469(n5469), 
            .\REG.mem_47_12 (\REG.mem_47_12 ), .n5468(n5468), .n5467(n5467), 
            .\REG.mem_45_0 (\REG.mem_45_0 ), .\REG.mem_44_0 (\REG.mem_44_0 ), 
            .\REG.mem_45_10 (\REG.mem_45_10 ), .\REG.mem_44_10 (\REG.mem_44_10 ), 
            .n5466(n5466), .n5465(n5465), .\REG.mem_47_8 (\REG.mem_47_8 ), 
            .n5464(n5464), .\REG.mem_47_7 (\REG.mem_47_7 ), .n5463(n5463), 
            .n5462(n5462), .\REG.mem_47_5 (\REG.mem_47_5 ), .n5461(n5461), 
            .\REG.mem_47_4 (\REG.mem_47_4 ), .n5460(n5460), .n5459(n5459), 
            .n5458(n5458), .n5457(n5457), .n5456(n5456), .\REG.mem_46_15 (\REG.mem_46_15 ), 
            .n5455(n5455), .\REG.mem_46_14 (\REG.mem_46_14 ), .n5454(n5454), 
            .\REG.mem_46_13 (\REG.mem_46_13 ), .n5453(n5453), .\REG.mem_46_12 (\REG.mem_46_12 ), 
            .n5452(n5452), .n5451(n5451), .n5450(n5450), .n5449(n5449), 
            .\REG.mem_46_8 (\REG.mem_46_8 ), .n5448(n5448), .\REG.mem_46_7 (\REG.mem_46_7 ), 
            .n5447(n5447), .n5446(n5446), .\REG.mem_46_5 (\REG.mem_46_5 ), 
            .n5445(n5445), .\REG.mem_46_4 (\REG.mem_46_4 ), .n5444(n5444), 
            .n5443(n5443), .n5442(n5442), .n5441(n5441), .n5440(n5440), 
            .\REG.mem_45_15 (\REG.mem_45_15 ), .n5439(n5439), .\REG.mem_45_14 (\REG.mem_45_14 ), 
            .n5438(n5438), .\REG.mem_45_13 (\REG.mem_45_13 ), .n5437(n5437), 
            .\REG.mem_45_12 (\REG.mem_45_12 ), .n5436(n5436), .n5435(n5435), 
            .n5434(n5434), .\REG.mem_38_7 (\REG.mem_38_7 ), .\REG.mem_39_7 (\REG.mem_39_7 ), 
            .\REG.mem_37_7 (\REG.mem_37_7 ), .\REG.mem_36_7 (\REG.mem_36_7 ), 
            .n5433(n5433), .\REG.mem_45_8 (\REG.mem_45_8 ), .n5432(n5432), 
            .\REG.mem_45_7 (\REG.mem_45_7 ), .n5431(n5431), .n5430(n5430), 
            .\REG.mem_45_5 (\REG.mem_45_5 ), .n5429(n5429), .\REG.mem_45_4 (\REG.mem_45_4 ), 
            .n5428(n5428), .n5427(n5427), .n5426(n5426), .n5425(n5425), 
            .n5424(n5424), .\REG.mem_44_15 (\REG.mem_44_15 ), .n5423(n5423), 
            .\REG.mem_44_14 (\REG.mem_44_14 ), .n5422(n5422), .\REG.mem_44_13 (\REG.mem_44_13 ), 
            .n5421(n5421), .\REG.mem_44_12 (\REG.mem_44_12 ), .n5420(n5420), 
            .n5419(n5419), .\REG.mem_10_0 (\REG.mem_10_0 ), .\REG.mem_11_0 (\REG.mem_11_0 ), 
            .n5418(n5418), .\REG.mem_9_0 (\REG.mem_9_0 ), .\REG.mem_8_0 (\REG.mem_8_0 ), 
            .n5417(n5417), .\REG.mem_44_8 (\REG.mem_44_8 ), .n5416(n5416), 
            .\REG.mem_44_7 (\REG.mem_44_7 ), .n5415(n5415), .n5414(n5414), 
            .\REG.mem_44_5 (\REG.mem_44_5 ), .n5413(n5413), .\REG.mem_44_4 (\REG.mem_44_4 ), 
            .n5412(n5412), .n5411(n5411), .n5410(n5410), .n5409(n5409), 
            .n5408(n5408), .n5407(n5407), .\REG.mem_43_15 (\REG.mem_43_15 ), 
            .n5406(n5406), .\REG.mem_43_14 (\REG.mem_43_14 ), .n5405(n5405), 
            .\REG.mem_43_13 (\REG.mem_43_13 ), .n5404(n5404), .\REG.mem_43_12 (\REG.mem_43_12 ), 
            .n5403(n5403), .n5402(n5402), .\REG.mem_10_5 (\REG.mem_10_5 ), 
            .\REG.mem_11_5 (\REG.mem_11_5 ), .\REG.mem_9_5 (\REG.mem_9_5 ), 
            .\REG.mem_8_5 (\REG.mem_8_5 ), .\wr_addr_p1_w[0] (wr_addr_p1_w[0]), 
            .n5401(n5401), .\REG.mem_43_9 (\REG.mem_43_9 ), .n5400(n5400), 
            .\REG.mem_43_8 (\REG.mem_43_8 ), .n5399(n5399), .\REG.mem_43_7 (\REG.mem_43_7 ), 
            .n5398(n5398), .\REG.mem_43_6 (\REG.mem_43_6 ), .n5397(n5397), 
            .\REG.mem_43_5 (\REG.mem_43_5 ), .n5396(n5396), .\REG.mem_43_4 (\REG.mem_43_4 ), 
            .n5395(n5395), .n5394(n5394), .n5393(n5393), .n5392(n5392), 
            .\REG.mem_43_0 (\REG.mem_43_0 ), .n11069(n11069), .\fifo_data_out[15] (fifo_data_out[15]), 
            .n5390(n5390), .\REG.mem_42_15 (\REG.mem_42_15 ), .n5389(n5389), 
            .\REG.mem_42_14 (\REG.mem_42_14 ), .n5388(n5388), .\REG.mem_42_13 (\REG.mem_42_13 ), 
            .n5387(n5387), .\REG.mem_42_12 (\REG.mem_42_12 ), .n5386(n5386), 
            .\REG.mem_42_4 (\REG.mem_42_4 ), .\REG.mem_41_4 (\REG.mem_41_4 ), 
            .\REG.mem_40_4 (\REG.mem_40_4 ), .n5385(n5385), .n5384(n5384), 
            .\REG.mem_42_9 (\REG.mem_42_9 ), .n5383(n5383), .\REG.mem_42_8 (\REG.mem_42_8 ), 
            .n5382(n5382), .\REG.mem_42_7 (\REG.mem_42_7 ), .n5381(n5381), 
            .\REG.mem_42_6 (\REG.mem_42_6 ), .n5380(n5380), .\REG.mem_42_5 (\REG.mem_42_5 ), 
            .n5379(n5379), .n5378(n5378), .n5377(n5377), .n5376(n5376), 
            .n5375(n5375), .\REG.mem_42_0 (\REG.mem_42_0 ), .n5374(n5374), 
            .\REG.mem_41_15 (\REG.mem_41_15 ), .n5373(n5373), .\REG.mem_41_14 (\REG.mem_41_14 ), 
            .n5372(n5372), .\REG.mem_41_13 (\REG.mem_41_13 ), .n5371(n5371), 
            .\REG.mem_41_12 (\REG.mem_41_12 ), .n4667(n4667), .n5370(n5370), 
            .n5369(n5369), .n5368(n5368), .\REG.mem_41_9 (\REG.mem_41_9 ), 
            .n5367(n5367), .\REG.mem_41_8 (\REG.mem_41_8 ), .n5366(n5366), 
            .\REG.mem_41_7 (\REG.mem_41_7 ), .n5365(n5365), .\REG.mem_41_6 (\REG.mem_41_6 ), 
            .n5364(n5364), .\REG.mem_41_5 (\REG.mem_41_5 ), .n5363(n5363), 
            .n5362(n5362), .n5361(n5361), .n5360(n5360), .n5358(n5358), 
            .\REG.mem_41_0 (\REG.mem_41_0 ), .n5357(n5357), .\REG.mem_40_15 (\REG.mem_40_15 ), 
            .n5356(n5356), .\REG.mem_40_14 (\REG.mem_40_14 ), .n5355(n5355), 
            .\REG.mem_40_13 (\REG.mem_40_13 ), .n5354(n5354), .\REG.mem_40_12 (\REG.mem_40_12 ), 
            .\REG.mem_38_13 (\REG.mem_38_13 ), .\REG.mem_39_13 (\REG.mem_39_13 ), 
            .\REG.mem_37_13 (\REG.mem_37_13 ), .\REG.mem_36_13 (\REG.mem_36_13 ), 
            .n5353(n5353), .n5352(n5352), .n5351(n5351), .\REG.mem_40_9 (\REG.mem_40_9 ), 
            .n5350(n5350), .\REG.mem_40_8 (\REG.mem_40_8 ), .n5349(n5349), 
            .\REG.mem_40_7 (\REG.mem_40_7 ), .n5348(n5348), .\REG.mem_40_6 (\REG.mem_40_6 ), 
            .n5347(n5347), .\REG.mem_40_5 (\REG.mem_40_5 ), .n5346(n5346), 
            .n5345(n5345), .n5344(n5344), .n5343(n5343), .n5342(n5342), 
            .\REG.mem_40_0 (\REG.mem_40_0 ), .n5341(n5341), .\REG.mem_39_15 (\REG.mem_39_15 ), 
            .n5340(n5340), .\REG.mem_39_14 (\REG.mem_39_14 ), .n5339(n5339), 
            .\REG.mem_23_5 (\REG.mem_23_5 ), .\REG.mem_14_0 (\REG.mem_14_0 ), 
            .\REG.mem_15_0 (\REG.mem_15_0 ), .\REG.mem_13_0 (\REG.mem_13_0 ), 
            .\REG.mem_12_0 (\REG.mem_12_0 ), .n5338(n5338), .n5337(n5337), 
            .n5336(n5336), .n5335(n5335), .\REG.mem_39_9 (\REG.mem_39_9 ), 
            .n5334(n5334), .\REG.mem_39_8 (\REG.mem_39_8 ), .n5333(n5333), 
            .n5332(n5332), .\REG.mem_39_6 (\REG.mem_39_6 ), .n5331(n5331), 
            .n5330(n5330), .n5329(n5329), .\REG.mem_39_3 (\REG.mem_39_3 ), 
            .n5328(n5328), .\REG.mem_39_2 (\REG.mem_39_2 ), .n5327(n5327), 
            .n5326(n5326), .\REG.mem_39_0 (\REG.mem_39_0 ), .n5323(n5323), 
            .\REG.mem_38_15 (\REG.mem_38_15 ), .n5322(n5322), .\REG.mem_38_14 (\REG.mem_38_14 ), 
            .n5321(n5321), .n5320(n5320), .n5319(n5319), .n5318(n5318), 
            .n5317(n5317), .\REG.mem_38_9 (\REG.mem_38_9 ), .n5316(n5316), 
            .\REG.mem_38_8 (\REG.mem_38_8 ), .n5315(n5315), .n5314(n5314), 
            .\REG.mem_38_6 (\REG.mem_38_6 ), .n5313(n5313), .n5312(n5312), 
            .n5311(n5311), .\REG.mem_38_3 (\REG.mem_38_3 ), .n5310(n5310), 
            .\REG.mem_38_2 (\REG.mem_38_2 ), .n5309(n5309), .n5308(n5308), 
            .\REG.mem_38_0 (\REG.mem_38_0 ), .n5302(n5302), .\REG.mem_37_15 (\REG.mem_37_15 ), 
            .n5301(n5301), .\REG.mem_37_14 (\REG.mem_37_14 ), .n5300(n5300), 
            .n5299(n5299), .n5298(n5298), .n5297(n5297), .n5296(n5296), 
            .\REG.mem_37_9 (\REG.mem_37_9 ), .n5295(n5295), .\REG.mem_37_8 (\REG.mem_37_8 ), 
            .n5294(n5294), .n5293(n5293), .\REG.mem_37_6 (\REG.mem_37_6 ), 
            .n5292(n5292), .n5291(n5291), .n5290(n5290), .\REG.mem_37_3 (\REG.mem_37_3 ), 
            .n5289(n5289), .\REG.mem_37_2 (\REG.mem_37_2 ), .n5288(n5288), 
            .n5286(n5286), .\REG.mem_37_0 (\REG.mem_37_0 ), .n5285(n5285), 
            .\REG.mem_36_15 (\REG.mem_36_15 ), .n5284(n5284), .\REG.mem_36_14 (\REG.mem_36_14 ), 
            .n5283(n5283), .n5282(n5282), .n5281(n5281), .n5280(n5280), 
            .n5279(n5279), .\REG.mem_36_9 (\REG.mem_36_9 ), .n5278(n5278), 
            .\REG.mem_36_8 (\REG.mem_36_8 ), .n5277(n5277), .n5276(n5276), 
            .\REG.mem_36_6 (\REG.mem_36_6 ), .n5275(n5275), .n5274(n5274), 
            .n5273(n5273), .\REG.mem_36_3 (\REG.mem_36_3 ), .n5272(n5272), 
            .\REG.mem_36_2 (\REG.mem_36_2 ), .n5271(n5271), .n5270(n5270), 
            .\REG.mem_36_0 (\REG.mem_36_0 ), .\REG.mem_26_12 (\REG.mem_26_12 ), 
            .\REG.mem_10_3 (\REG.mem_10_3 ), .\REG.mem_11_3 (\REG.mem_11_3 ), 
            .n5202(n5202), .\REG.mem_31_15 (\REG.mem_31_15 ), .n5201(n5201), 
            .n5200(n5200), .n5199(n5199), .n5198(n5198), .n5197(n5197), 
            .n5196(n5196), .\REG.mem_31_9 (\REG.mem_31_9 ), .n5195(n5195), 
            .n5194(n5194), .n5193(n5193), .\REG.mem_31_6 (\REG.mem_31_6 ), 
            .n5192(n5192), .\REG.mem_31_5 (\REG.mem_31_5 ), .n5191(n5191), 
            .\REG.mem_31_4 (\REG.mem_31_4 ), .n5190(n5190), .n5189(n5189), 
            .\REG.mem_31_2 (\REG.mem_31_2 ), .\REG.mem_9_3 (\REG.mem_9_3 ), 
            .\REG.mem_8_3 (\REG.mem_8_3 ), .n5188(n5188), .n5187(n5187), 
            .\REG.mem_10_14 (\REG.mem_10_14 ), .\REG.mem_11_14 (\REG.mem_11_14 ), 
            .\REG.mem_9_14 (\REG.mem_9_14 ), .\REG.mem_8_14 (\REG.mem_8_14 ), 
            .\REG.mem_23_2 (\REG.mem_23_2 ), .n5121(n5121), .n5120(n5120), 
            .n5119(n5119), .n5118(n5118), .n5117(n5117), .n5116(n5116), 
            .n5115(n5115), .\REG.mem_26_9 (\REG.mem_26_9 ), .n5114(n5114), 
            .n5113(n5113), .n5112(n5112), .\REG.mem_26_6 (\REG.mem_26_6 ), 
            .n5111(n5111), .\REG.mem_26_5 (\REG.mem_26_5 ), .n5110(n5110), 
            .n5109(n5109), .n5108(n5108), .\REG.mem_26_2 (\REG.mem_26_2 ), 
            .n5107(n5107), .n5106(n5106), .n5073(n5073), .n5072(n5072), 
            .\REG.mem_23_14 (\REG.mem_23_14 ), .n5071(n5071), .n5070(n5070), 
            .n5069(n5069), .n5068(n5068), .n5067(n5067), .\REG.mem_23_9 (\REG.mem_23_9 ), 
            .n5066(n5066), .\rd_grey_sync_r[5] (rd_grey_sync_r[5]), .\rd_grey_sync_r[4] (rd_grey_sync_r[4]), 
            .\REG.mem_10_6 (\REG.mem_10_6 ), .\REG.mem_11_6 (\REG.mem_11_6 ), 
            .\rd_grey_sync_r[3] (rd_grey_sync_r[3]), .\rd_grey_sync_r[2] (rd_grey_sync_r[2]), 
            .\rd_grey_sync_r[1] (rd_grey_sync_r[1]), .n5065(n5065), .n5064(n5064), 
            .\REG.mem_23_6 (\REG.mem_23_6 ), .n5063(n5063), .n5062(n5062), 
            .\REG.mem_23_4 (\REG.mem_23_4 ), .n5061(n5061), .\REG.mem_23_3 (\REG.mem_23_3 ), 
            .n5060(n5060), .n5059(n5059), .n5058(n5058), .\REG.mem_23_0 (\REG.mem_23_0 ), 
            .\REG.mem_9_6 (\REG.mem_9_6 ), .\REG.mem_8_6 (\REG.mem_8_6 ), 
            .n5(n5), .\REG.mem_14_6 (\REG.mem_14_6 ), .\REG.mem_15_6 (\REG.mem_15_6 ), 
            .\REG.mem_13_6 (\REG.mem_13_6 ), .\REG.mem_12_6 (\REG.mem_12_6 ), 
            .n5006(n5006), .\REG.mem_19_15 (\REG.mem_19_15 ), .n5005(n5005), 
            .\REG.mem_19_14 (\REG.mem_19_14 ), .n5004(n5004), .n5003(n5003), 
            .n5002(n5002), .\REG.mem_19_11 (\REG.mem_19_11 ), .n5001(n5001), 
            .n5000(n5000), .\REG.mem_19_9 (\REG.mem_19_9 ), .n4999(n4999), 
            .n4998(n4998), .n4997(n4997), .\REG.mem_19_6 (\REG.mem_19_6 ), 
            .n4996(n4996), .\REG.mem_19_5 (\REG.mem_19_5 ), .n4995(n4995), 
            .\REG.mem_19_4 (\REG.mem_19_4 ), .n4994(n4994), .\REG.mem_19_3 (\REG.mem_19_3 ), 
            .n4993(n4993), .n4992(n4992), .n4991(n4991), .\REG.mem_19_0 (\REG.mem_19_0 ), 
            .n4990(n4990), .\REG.mem_18_15 (\REG.mem_18_15 ), .n4989(n4989), 
            .\REG.mem_18_14 (\REG.mem_18_14 ), .n4988(n4988), .n4987(n4987), 
            .n4986(n4986), .\REG.mem_18_11 (\REG.mem_18_11 ), .n4985(n4985), 
            .n4984(n4984), .\REG.mem_18_9 (\REG.mem_18_9 ), .n4983(n4983), 
            .n4982(n4982), .n4981(n4981), .\REG.mem_18_6 (\REG.mem_18_6 ), 
            .n4980(n4980), .\REG.mem_18_5 (\REG.mem_18_5 ), .n4979(n4979), 
            .\REG.mem_18_4 (\REG.mem_18_4 ), .n4978(n4978), .\REG.mem_18_3 (\REG.mem_18_3 ), 
            .n4977(n4977), .n4976(n4976), .n4975(n4975), .\REG.mem_18_0 (\REG.mem_18_0 ), 
            .n4974(n4974), .\REG.mem_17_15 (\REG.mem_17_15 ), .n4973(n4973), 
            .\REG.mem_17_14 (\REG.mem_17_14 ), .n4972(n4972), .n4971(n4971), 
            .n4970(n4970), .\REG.mem_17_11 (\REG.mem_17_11 ), .n4969(n4969), 
            .n4968(n4968), .\REG.mem_17_9 (\REG.mem_17_9 ), .n4967(n4967), 
            .n4966(n4966), .n4965(n4965), .\REG.mem_17_6 (\REG.mem_17_6 ), 
            .n4964(n4964), .\REG.mem_17_5 (\REG.mem_17_5 ), .n4963(n4963), 
            .\REG.mem_17_4 (\REG.mem_17_4 ), .n4962(n4962), .\REG.mem_17_3 (\REG.mem_17_3 ), 
            .n4961(n4961), .n4960(n4960), .n4958(n4958), .\REG.mem_17_0 (\REG.mem_17_0 ), 
            .n4957(n4957), .\REG.mem_16_15 (\REG.mem_16_15 ), .n4956(n4956), 
            .\REG.mem_16_14 (\REG.mem_16_14 ), .n4955(n4955), .n4954(n4954), 
            .n4953(n4953), .\REG.mem_16_11 (\REG.mem_16_11 ), .n4952(n4952), 
            .n51(n51), .n4951(n4951), .\REG.mem_16_9 (\REG.mem_16_9 ), 
            .n4950(n4950), .n4949(n4949), .n4948(n4948), .\REG.mem_16_6 (\REG.mem_16_6 ), 
            .n4947(n4947), .\REG.mem_16_5 (\REG.mem_16_5 ), .n4946(n4946), 
            .\REG.mem_16_4 (\REG.mem_16_4 ), .n4945(n4945), .\REG.mem_16_3 (\REG.mem_16_3 ), 
            .n4944(n4944), .n4943(n4943), .n4942(n4942), .\REG.mem_16_0 (\REG.mem_16_0 ), 
            .n4941(n4941), .n4940(n4940), .\REG.mem_15_14 (\REG.mem_15_14 ), 
            .n4939(n4939), .n4938(n4938), .n4937(n4937), .\REG.mem_15_11 (\REG.mem_15_11 ), 
            .\rd_addr_nxt_c_6__N_465[5] (rd_addr_nxt_c_6__N_465[5]), .n19(n19), 
            .n4936(n4936), .n4935(n4935), .get_next_word(get_next_word), 
            .\rd_addr_nxt_c_6__N_465[3] (rd_addr_nxt_c_6__N_465[3]), .n4934(n4934), 
            .n4933(n4933), .n4932(n4932), .n4931(n4931), .n4930(n4930), 
            .\REG.mem_15_4 (\REG.mem_15_4 ), .n4929(n4929), .\REG.mem_15_3 (\REG.mem_15_3 ), 
            .n4928(n4928), .n4927(n4927), .n4926(n4926), .n4925(n4925), 
            .n4924(n4924), .\REG.mem_14_14 (\REG.mem_14_14 ), .n4923(n4923), 
            .n4922(n4922), .n4921(n4921), .\REG.mem_14_11 (\REG.mem_14_11 ), 
            .n4920(n4920), .n4919(n4919), .n4918(n4918), .\rd_addr_nxt_c_6__N_465[1] (rd_addr_nxt_c_6__N_465[1]), 
            .\state_timeout_counter[3] (state_timeout_counter_adj_1218[3]), 
            .n718(n718), .n7(n7), .n14424(n14424), .n4917(n4917), .n4916(n4916), 
            .n4915(n4915), .n4914(n4914), .\REG.mem_14_4 (\REG.mem_14_4 ), 
            .n4913(n4913), .\REG.mem_14_3 (\REG.mem_14_3 ), .n4912(n4912), 
            .n4911(n4911), .n4910(n4910), .\REG.mem_6_15 (\REG.mem_6_15 ), 
            .\REG.mem_7_15 (\REG.mem_7_15 ), .\REG.mem_5_15 (\REG.mem_5_15 ), 
            .\REG.mem_4_15 (\REG.mem_4_15 ), .\REG.mem_10_15 (\REG.mem_10_15 ), 
            .\REG.mem_11_15 (\REG.mem_11_15 ), .\REG.mem_9_15 (\REG.mem_9_15 ), 
            .\REG.mem_8_15 (\REG.mem_8_15 ), .n50(n50), .n52(n52), .n20(n20), 
            .n18(n18), .n4909(n4909), .n4908(n4908), .\REG.mem_13_14 (\REG.mem_13_14 ), 
            .n4907(n4907), .n4906(n4906), .n4905(n4905), .\REG.mem_13_11 (\REG.mem_13_11 ), 
            .n4904(n4904), .n4903(n4903), .n4902(n4902), .n4901(n4901), 
            .n46(n46), .n4900(n4900), .n4899(n4899), .n14(n14), .\REG.mem_10_11 (\REG.mem_10_11 ), 
            .\REG.mem_11_11 (\REG.mem_11_11 ), .n4898(n4898), .\REG.mem_13_4 (\REG.mem_13_4 ), 
            .n4897(n4897), .\REG.mem_13_3 (\REG.mem_13_3 ), .\REG.mem_9_11 (\REG.mem_9_11 ), 
            .\REG.mem_8_11 (\REG.mem_8_11 ), .\REG.mem_12_14 (\REG.mem_12_14 ), 
            .\REG.mem_12_11 (\REG.mem_12_11 ), .n4896(n4896), .n4895(n4895), 
            .n4894(n4894), .n4893(n4893), .n4892(n4892), .n53(n53), 
            .n4891(n4891), .n4890(n4890), .n21(n21), .n4889(n4889), 
            .n4888(n4888), .n4887(n4887), .n4886(n4886), .n4885(n4885), 
            .n4884(n4884), .n4883(n4883), .n4882(n4882), .\REG.mem_12_4 (\REG.mem_12_4 ), 
            .n4881(n4881), .\REG.mem_12_3 (\REG.mem_12_3 ), .n4880(n4880), 
            .n4879(n4879), .n4878(n4878), .n4646(n4646), .n4644(n4644), 
            .n4639(n4639), .n4877(n4877), .n4876(n4876), .n4875(n4875), 
            .n4874(n4874), .n4873(n4873), .n4872(n4872), .n4871(n4871), 
            .n4870(n4870), .\REG.mem_11_8 (\REG.mem_11_8 ), .n4869(n4869), 
            .n4638(n4638), .n4868(n4868), .n4867(n4867), .n4866(n4866), 
            .\REG.mem_11_4 (\REG.mem_11_4 ), .n4865(n4865), .n4864(n4864), 
            .n4863(n4863), .n4862(n4862), .n4861(n4861), .n4860(n4860), 
            .n4859(n4859), .n54(n54), .n22(n22), .n39(n39), .n7_adj_4(n7_adj_1183), 
            .n4858(n4858), .n4857(n4857), .n4856(n4856), .n4855(n4855), 
            .n4854(n4854), .\REG.mem_10_8 (\REG.mem_10_8 ), .n4853(n4853), 
            .n4852(n4852), .n4851(n4851), .n56(n56), .n24(n24_adj_1185), 
            .n4850(n4850), .\REG.mem_10_4 (\REG.mem_10_4 ), .n4849(n4849), 
            .n4848(n4848), .n4847(n4847), .n4846(n4846), .n4845(n4845), 
            .n4844(n4844), .n4843(n4843), .n4842(n4842), .n4841(n4841), 
            .n4840(n4840), .n4839(n4839), .\afull_flag_impl.af_flag_p_w_N_603[3] (\afull_flag_impl.af_flag_p_w_N_603 [3]), 
            .n4838(n4838), .\REG.mem_9_8 (\REG.mem_9_8 ), .n4837(n4837), 
            .n4836(n4836), .n4835(n4835), .n4834(n4834), .\REG.mem_9_4 (\REG.mem_9_4 ), 
            .n4833(n4833), .n4832(n4832), .n4831(n4831), .n4830(n4830), 
            .n4829(n4829), .n4828(n4828), .n4827(n4827), .n4826(n4826), 
            .n4825(n4825), .n4824(n4824), .n4823(n4823), .n4822(n4822), 
            .\REG.mem_8_8 (\REG.mem_8_8 ), .n4821(n4821), .n4820(n4820), 
            .n4819(n4819), .n4818(n4818), .\REG.mem_8_4 (\REG.mem_8_4 ), 
            .n4817(n4817), .n4816(n4816), .n4815(n4815), .n4814(n4814), 
            .n4813(n4813), .n4812(n4812), .n4811(n4811), .\REG.mem_7_13 (\REG.mem_7_13 ), 
            .n4810(n4810), .n4809(n4809), .n4808(n4808), .n4807(n4807), 
            .\REG.mem_7_9 (\REG.mem_7_9 ), .n4806(n4806), .n4805(n4805), 
            .n4804(n4804), .\REG.mem_7_6 (\REG.mem_7_6 ), .n4803(n4803), 
            .\REG.mem_7_5 (\REG.mem_7_5 ), .n4802(n4802), .\REG.mem_7_4 (\REG.mem_7_4 ), 
            .n4801(n4801), .n4800(n4800), .n4799(n4799), .n4798(n4798), 
            .\REG.mem_7_0 (\REG.mem_7_0 ), .n4797(n4797), .n4796(n4796), 
            .n4795(n4795), .\REG.mem_6_13 (\REG.mem_6_13 ), .n4794(n4794), 
            .n4793(n4793), .n4792(n4792), .n4791(n4791), .\REG.mem_6_9 (\REG.mem_6_9 ), 
            .n4790(n4790), .n4789(n4789), .n4788(n4788), .\REG.mem_6_6 (\REG.mem_6_6 ), 
            .n4787(n4787), .\REG.mem_6_5 (\REG.mem_6_5 ), .n4786(n4786), 
            .\REG.mem_6_4 (\REG.mem_6_4 ), .n4785(n4785), .n4784(n4784), 
            .n4783(n4783), .n4779(n4779), .\REG.mem_6_0 (\REG.mem_6_0 ), 
            .n4778(n4778), .n4777(n4777), .n4776(n4776), .\REG.mem_5_13 (\REG.mem_5_13 ), 
            .n4775(n4775), .n4774(n4774), .n4773(n4773), .n4772(n4772), 
            .\REG.mem_5_9 (\REG.mem_5_9 ), .n4771(n4771), .n4770(n4770), 
            .n4769(n4769), .\REG.mem_5_6 (\REG.mem_5_6 ), .n4768(n4768), 
            .\REG.mem_5_5 (\REG.mem_5_5 ), .n4767(n4767), .\REG.mem_5_4 (\REG.mem_5_4 ), 
            .n4766(n4766), .n4765(n4765), .n4764(n4764), .n4763(n4763), 
            .\REG.mem_5_0 (\REG.mem_5_0 ), .n4762(n4762), .n4761(n4761), 
            .n4760(n4760), .\REG.mem_4_13 (\REG.mem_4_13 ), .n4759(n4759), 
            .n4758(n4758), .n4757(n4757), .n4756(n4756), .\REG.mem_4_9 (\REG.mem_4_9 ), 
            .n4755(n4755), .n4754(n4754), .n4753(n4753), .\REG.mem_4_6 (\REG.mem_4_6 ), 
            .n4752(n4752), .\REG.mem_4_5 (\REG.mem_4_5 ), .n4751(n4751), 
            .\REG.mem_4_4 (\REG.mem_4_4 ), .n4750(n4750), .n4749(n4749), 
            .n4748(n4748), .n4747(n4747), .\REG.mem_4_0 (\REG.mem_4_0 ), 
            .n4612(n4612), .n57(n57), .n25(n25), .n42(n42), .n10(n10), 
            .n49(n49), .n17(n17), .n48(n48), .n16(n16), .n55(n55), 
            .n23(n23), .n59(n59), .n27(n27)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(537[21] 552[2])
    SB_LUT4 i3693_3_lut (.I0(\REG.mem_13_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n52), .I3(GND_net), .O(n4895));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3692_3_lut (.I0(\REG.mem_13_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n52), .I3(GND_net), .O(n4894));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3691_3_lut (.I0(\REG.mem_12_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n53), .I3(GND_net), .O(n4893));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3477_2_lut_3_lut (.I0(reset_all_w), .I1(fifo_read_cmd), .I2(is_fifo_empty_flag), 
            .I3(GND_net), .O(n4679));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    defparam i3477_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i3690_3_lut (.I0(\REG.mem_12_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n53), .I3(GND_net), .O(n4892));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1138_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(reset_all_w), .I3(GND_net), .O(n2207));
    defparam i1138_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i3689_3_lut (.I0(\REG.mem_12_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n53), .I3(GND_net), .O(n4891));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3688_3_lut (.I0(\REG.mem_12_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n53), .I3(GND_net), .O(n4890));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3687_3_lut (.I0(\REG.mem_12_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n53), .I3(GND_net), .O(n4889));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3686_3_lut (.I0(\REG.mem_12_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n53), .I3(GND_net), .O(n4888));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3685_3_lut (.I0(\REG.mem_12_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n53), .I3(GND_net), .O(n4887));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3684_3_lut (.I0(\REG.mem_12_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n53), .I3(GND_net), .O(n4886));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3683_3_lut (.I0(\REG.mem_12_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n53), .I3(GND_net), .O(n4885));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3682_3_lut (.I0(\REG.mem_12_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n53), .I3(GND_net), .O(n4884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3681_3_lut (.I0(\REG.mem_12_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n53), .I3(GND_net), .O(n4883));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3680_3_lut (.I0(\REG.mem_12_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n53), .I3(GND_net), .O(n4882));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3679_3_lut (.I0(\REG.mem_12_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n53), .I3(GND_net), .O(n4881));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3678_3_lut (.I0(\REG.mem_12_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n53), .I3(GND_net), .O(n4880));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3677_3_lut (.I0(\REG.mem_12_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n53), .I3(GND_net), .O(n4879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3676_3_lut (.I0(\REG.mem_12_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n53), .I3(GND_net), .O(n4878));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3676_3_lut.LUT_INIT = 16'hcaca;
    \uart_rx(CLKS_PER_BIT=20)  pc_rx (.SLM_CLK_c(SLM_CLK_c), .r_Rx_Data(r_Rx_Data), 
            .UART_RX_c(UART_RX_c), .GND_net(GND_net), .n4(n4), .n4_adj_1(n4_adj_1205), 
            .n7455(n7455), .n4_adj_2(n4_adj_1206), .n10847(n10847), .debug_led3(debug_led3), 
            .n5869(n5869), .pc_data_rx({pc_data_rx}), .VCC_net(VCC_net), 
            .n5844(n5844), .n5843(n5843), .n5842(n5842), .n5841(n5841), 
            .n5840(n5840), .n5839(n5839), .n5838(n5838), .n3997(n3997), 
            .n4002(n4002)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(689[42] 694[3])
    SB_LUT4 i3444_2_lut (.I0(reset_all), .I1(wp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4646));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i3444_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4691_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [5]), 
            .I3(fifo_data_out[5]), .O(n5893));
    defparam i4691_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3442_2_lut (.I0(reset_all), .I1(wr_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4644));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    defparam i3442_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i12_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [7]), 
            .I3(fifo_data_out[7]), .O(n11119));
    defparam i12_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i914_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(n63), 
            .I3(state[2]), .O(n1876));   // src/timing_controller.v(48[11:16])
    defparam i914_4_lut_4_lut.LUT_INIT = 16'h0806;
    SB_LUT4 i12_4_lut_4_lut_adj_94 (.I0(t_rd_fifo_en_w), .I1(reset_all), 
            .I2(\REG.out_raw [3]), .I3(fifo_data_out[3]), .O(n11139));
    defparam i12_4_lut_4_lut_adj_94.LUT_INIT = 16'h3120;
    SB_LUT4 i3437_2_lut (.I0(reset_all), .I1(rp_sync1_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4639));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i3437_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3675_3_lut (.I0(\REG.mem_11_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n54), .I3(GND_net), .O(n4877));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_95 (.I0(t_rd_fifo_en_w), .I1(reset_all), 
            .I2(\REG.out_raw [8]), .I3(fifo_data_out[8]), .O(n11097));
    defparam i12_4_lut_4_lut_adj_95.LUT_INIT = 16'h3120;
    SB_LUT4 i4206_2_lut_4_lut (.I0(reset_all), .I1(wr_grey_sync_r[6]), .I2(wr_addr_p1_w[6]), 
            .I3(n7596), .O(n5408));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    defparam i4206_2_lut_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i3674_3_lut (.I0(\REG.mem_11_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n54), .I3(GND_net), .O(n4876));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3673_3_lut (.I0(\REG.mem_11_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n54), .I3(GND_net), .O(n4875));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3672_3_lut (.I0(\REG.mem_11_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n54), .I3(GND_net), .O(n4874));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3671_3_lut (.I0(\REG.mem_11_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n54), .I3(GND_net), .O(n4873));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3670_3_lut (.I0(\REG.mem_11_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n54), .I3(GND_net), .O(n4872));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3669_3_lut (.I0(\REG.mem_11_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n54), .I3(GND_net), .O(n4871));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3668_3_lut (.I0(\REG.mem_11_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n54), .I3(GND_net), .O(n4870));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3667_3_lut (.I0(\REG.mem_11_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n54), .I3(GND_net), .O(n4869));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4652_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [0]), 
            .I3(fifo_data_out[0]), .O(n5854));
    defparam i4652_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i3436_2_lut (.I0(reset_all), .I1(rd_grey_sync_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4638));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    defparam i3436_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3435_3_lut (.I0(rx_buf_byte[0]), .I1(rx_shift_reg[0]), .I2(n3204), 
            .I3(GND_net), .O(n4637));   // src/spi.v(76[8] 221[4])
    defparam i3435_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3430_3_lut (.I0(r_Tx_Data[0]), .I1(fifo_temp_output[0]), .I2(n3710), 
            .I3(GND_net), .O(n4632));   // src/uart_tx.v(38[10] 141[8])
    defparam i3430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3666_3_lut (.I0(\REG.mem_11_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n54), .I3(GND_net), .O(n4868));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3665_3_lut (.I0(\REG.mem_11_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n54), .I3(GND_net), .O(n4867));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3664_3_lut (.I0(\REG.mem_11_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n54), .I3(GND_net), .O(n4866));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3663_3_lut (.I0(\REG.mem_11_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n54), .I3(GND_net), .O(n4865));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3662_3_lut (.I0(\REG.mem_11_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n54), .I3(GND_net), .O(n4864));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3661_3_lut (.I0(\REG.mem_11_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n54), .I3(GND_net), .O(n4863));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3660_3_lut (.I0(\REG.mem_11_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n54), .I3(GND_net), .O(n4862));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3659_3_lut (.I0(\REG.mem_10_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n55), .I3(GND_net), .O(n4861));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_96 (.I0(t_rd_fifo_en_w), .I1(reset_all), 
            .I2(\REG.out_raw [15]), .I3(fifo_data_out[15]), .O(n11069));
    defparam i12_4_lut_4_lut_adj_96.LUT_INIT = 16'h3120;
    SB_LUT4 i1_2_lut_4_lut (.I0(reset_clk_counter[2]), .I1(reset_all_w_N_61), 
            .I2(reset_clk_counter[0]), .I3(reset_clk_counter[1]), .O(n10800));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'haaa6;
    SB_LUT4 i3658_3_lut (.I0(\REG.mem_10_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n55), .I3(GND_net), .O(n4860));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3657_3_lut (.I0(\REG.mem_10_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n55), .I3(GND_net), .O(n4859));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3656_3_lut (.I0(\REG.mem_10_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n55), .I3(GND_net), .O(n4858));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3655_3_lut (.I0(\REG.mem_10_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n55), .I3(GND_net), .O(n4857));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3654_3_lut (.I0(\REG.mem_10_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n55), .I3(GND_net), .O(n4856));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3653_3_lut (.I0(\REG.mem_10_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n55), .I3(GND_net), .O(n4855));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3652_3_lut (.I0(\REG.mem_10_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n55), .I3(GND_net), .O(n4854));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3651_3_lut (.I0(\REG.mem_10_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n55), .I3(GND_net), .O(n4853));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3650_3_lut (.I0(\REG.mem_10_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n55), .I3(GND_net), .O(n4852));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3649_3_lut (.I0(\REG.mem_10_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n55), .I3(GND_net), .O(n4851));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3648_3_lut (.I0(\REG.mem_10_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n55), .I3(GND_net), .O(n4850));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3647_3_lut (.I0(\REG.mem_10_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n55), .I3(GND_net), .O(n4849));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3646_3_lut (.I0(\REG.mem_10_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n55), .I3(GND_net), .O(n4848));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3645_3_lut (.I0(\REG.mem_10_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n55), .I3(GND_net), .O(n4847));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3644_3_lut (.I0(\REG.mem_10_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n55), .I3(GND_net), .O(n4846));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3643_3_lut (.I0(\REG.mem_9_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n56), .I3(GND_net), .O(n4845));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_97 (.I0(t_rd_fifo_en_w), .I1(reset_all), 
            .I2(\REG.out_raw [11]), .I3(fifo_data_out[11]), .O(n11135));
    defparam i12_4_lut_4_lut_adj_97.LUT_INIT = 16'h3120;
    SB_LUT4 i3642_3_lut (.I0(\REG.mem_9_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n56), .I3(GND_net), .O(n4844));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3641_3_lut (.I0(\REG.mem_9_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n56), .I3(GND_net), .O(n4843));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3640_3_lut (.I0(\REG.mem_9_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n56), .I3(GND_net), .O(n4842));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3639_3_lut (.I0(\REG.mem_9_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n56), .I3(GND_net), .O(n4841));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3638_3_lut (.I0(\REG.mem_9_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n56), .I3(GND_net), .O(n4840));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3637_3_lut (.I0(\REG.mem_9_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n56), .I3(GND_net), .O(n4839));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_4_lut (.I0(is_tx_fifo_full_flag), .I1(n11424), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3636_3_lut (.I0(\REG.mem_9_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n56), .I3(GND_net), .O(n4838));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3635_3_lut (.I0(\REG.mem_9_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n56), .I3(GND_net), .O(n4837));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3634_3_lut (.I0(\REG.mem_9_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n56), .I3(GND_net), .O(n4836));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3633_3_lut (.I0(\REG.mem_9_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n56), .I3(GND_net), .O(n4835));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3632_3_lut (.I0(\REG.mem_9_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n56), .I3(GND_net), .O(n4834));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3631_3_lut (.I0(\REG.mem_9_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n56), .I3(GND_net), .O(n4833));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3630_3_lut (.I0(\REG.mem_9_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n56), .I3(GND_net), .O(n4832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3629_3_lut (.I0(\REG.mem_9_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n56), .I3(GND_net), .O(n4831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3628_3_lut (.I0(\REG.mem_9_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n56), .I3(GND_net), .O(n4830));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3627_3_lut (.I0(\REG.mem_8_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n57), .I3(GND_net), .O(n4829));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_98 (.I0(t_rd_fifo_en_w), .I1(reset_all), 
            .I2(\REG.out_raw [10]), .I3(fifo_data_out[10]), .O(n11089));
    defparam i12_4_lut_4_lut_adj_98.LUT_INIT = 16'h3120;
    SB_LUT4 i3468_4_lut_4_lut (.I0(reset_all_w), .I1(rd_addr_r_adj_1252[1]), 
            .I2(rd_addr_r_adj_1252[0]), .I3(rd_fifo_en_w), .O(n4670));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i3468_4_lut_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i3626_3_lut (.I0(\REG.mem_8_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n57), .I3(GND_net), .O(n4828));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3625_3_lut (.I0(\REG.mem_8_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n57), .I3(GND_net), .O(n4827));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3624_3_lut (.I0(\REG.mem_8_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n57), .I3(GND_net), .O(n4826));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3623_3_lut (.I0(\REG.mem_8_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n57), .I3(GND_net), .O(n4825));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3622_3_lut (.I0(\REG.mem_8_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n57), .I3(GND_net), .O(n4824));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3621_3_lut (.I0(\REG.mem_8_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n57), .I3(GND_net), .O(n4823));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3620_3_lut (.I0(\REG.mem_8_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n57), .I3(GND_net), .O(n4822));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3619_3_lut (.I0(\REG.mem_8_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n57), .I3(GND_net), .O(n4821));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3618_3_lut (.I0(\REG.mem_8_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n57), .I3(GND_net), .O(n4820));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3617_3_lut (.I0(\REG.mem_8_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n57), .I3(GND_net), .O(n4819));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3616_3_lut (.I0(\REG.mem_8_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n57), .I3(GND_net), .O(n4818));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3615_3_lut (.I0(\REG.mem_8_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n57), .I3(GND_net), .O(n4817));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3614_3_lut (.I0(\REG.mem_8_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n57), .I3(GND_net), .O(n4816));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3613_3_lut (.I0(\REG.mem_8_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n57), .I3(GND_net), .O(n4815));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3612_3_lut (.I0(\REG.mem_8_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n57), .I3(GND_net), .O(n4814));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3611_3_lut (.I0(\REG.mem_7_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n58), .I3(GND_net), .O(n4813));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_99 (.I0(t_rd_fifo_en_w), .I1(reset_all), 
            .I2(\REG.out_raw [2]), .I3(fifo_data_out[2]), .O(n11141));
    defparam i12_4_lut_4_lut_adj_99.LUT_INIT = 16'h3120;
    SB_LUT4 i3610_3_lut (.I0(\REG.mem_7_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n58), .I3(GND_net), .O(n4812));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3609_3_lut (.I0(\REG.mem_7_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n58), .I3(GND_net), .O(n4811));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3608_3_lut (.I0(\REG.mem_7_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n58), .I3(GND_net), .O(n4810));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3607_3_lut (.I0(\REG.mem_7_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n58), .I3(GND_net), .O(n4809));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3606_3_lut (.I0(\REG.mem_7_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n58), .I3(GND_net), .O(n4808));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3605_3_lut (.I0(\REG.mem_7_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n58), .I3(GND_net), .O(n4807));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3604_3_lut (.I0(\REG.mem_7_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n58), .I3(GND_net), .O(n4806));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3603_3_lut (.I0(\REG.mem_7_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n58), .I3(GND_net), .O(n4805));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3602_3_lut (.I0(\REG.mem_7_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n58), .I3(GND_net), .O(n4804));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3601_3_lut (.I0(\REG.mem_7_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n58), .I3(GND_net), .O(n4803));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3600_3_lut (.I0(\REG.mem_7_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n58), .I3(GND_net), .O(n4802));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3599_3_lut (.I0(\REG.mem_7_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n58), .I3(GND_net), .O(n4801));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3598_3_lut (.I0(\REG.mem_7_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n58), .I3(GND_net), .O(n4800));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3597_3_lut (.I0(\REG.mem_7_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n58), .I3(GND_net), .O(n4799));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3596_3_lut (.I0(\REG.mem_7_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n58), .I3(GND_net), .O(n4798));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3595_3_lut (.I0(\REG.mem_6_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n59), .I3(GND_net), .O(n4797));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_100 (.I0(t_rd_fifo_en_w), .I1(reset_all), 
            .I2(\REG.out_raw [14]), .I3(fifo_data_out[14]), .O(n11071));
    defparam i12_4_lut_4_lut_adj_100.LUT_INIT = 16'h3120;
    SB_LUT4 i4668_2_lut_3_lut (.I0(fifo_data_out[0]), .I1(bluejay_data_out_31__N_703), 
            .I2(bluejay_data_out_31__N_704), .I3(GND_net), .O(n5870));   // src/bluejay_data.v(126[8] 148[4])
    defparam i4668_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i3594_3_lut (.I0(\REG.mem_6_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n59), .I3(GND_net), .O(n4796));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3593_3_lut (.I0(\REG.mem_6_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n59), .I3(GND_net), .O(n4795));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3592_3_lut (.I0(\REG.mem_6_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n59), .I3(GND_net), .O(n4794));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3591_3_lut (.I0(\REG.mem_6_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n59), .I3(GND_net), .O(n4793));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3590_3_lut (.I0(\REG.mem_6_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n59), .I3(GND_net), .O(n4792));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3589_3_lut (.I0(\REG.mem_6_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n59), .I3(GND_net), .O(n4791));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3588_3_lut (.I0(\REG.mem_6_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n59), .I3(GND_net), .O(n4790));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3587_3_lut (.I0(\REG.mem_6_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n59), .I3(GND_net), .O(n4789));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3586_3_lut (.I0(\REG.mem_6_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n59), .I3(GND_net), .O(n4788));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3585_3_lut (.I0(\REG.mem_6_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n59), .I3(GND_net), .O(n4787));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3584_3_lut (.I0(\REG.mem_6_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n59), .I3(GND_net), .O(n4786));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3583_3_lut (.I0(\REG.mem_6_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n59), .I3(GND_net), .O(n4785));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3582_3_lut (.I0(\REG.mem_6_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n59), .I3(GND_net), .O(n4784));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3581_3_lut (.I0(\REG.mem_6_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n59), .I3(GND_net), .O(n4783));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3577_3_lut (.I0(\REG.mem_6_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n59), .I3(GND_net), .O(n4779));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3576_3_lut (.I0(\REG.mem_5_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n60), .I3(GND_net), .O(n4778));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_4_lut_adj_101 (.I0(t_rd_fifo_en_w), .I1(reset_all), 
            .I2(\REG.out_raw [13]), .I3(fifo_data_out[13]), .O(n11073));
    defparam i12_4_lut_4_lut_adj_101.LUT_INIT = 16'h3120;
    SB_LUT4 i1_2_lut_4_lut_adj_102 (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(wr_addr_r_adj_1249[0]), .I3(rd_addr_r_adj_1252[0]), .O(n4_adj_1186));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1_2_lut_4_lut_adj_102.LUT_INIT = 16'h0220;
    SB_LUT4 i3575_3_lut (.I0(\REG.mem_5_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n60), .I3(GND_net), .O(n4777));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3574_3_lut (.I0(\REG.mem_5_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n60), .I3(GND_net), .O(n4776));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3573_3_lut (.I0(\REG.mem_5_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n60), .I3(GND_net), .O(n4775));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3572_3_lut (.I0(\REG.mem_5_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n60), .I3(GND_net), .O(n4774));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3571_3_lut (.I0(\REG.mem_5_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n60), .I3(GND_net), .O(n4773));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3570_3_lut (.I0(\REG.mem_5_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n60), .I3(GND_net), .O(n4772));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3569_3_lut (.I0(\REG.mem_5_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n60), .I3(GND_net), .O(n4771));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3568_3_lut (.I0(\REG.mem_5_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n60), .I3(GND_net), .O(n4770));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3567_3_lut (.I0(\REG.mem_5_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n60), .I3(GND_net), .O(n4769));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3566_3_lut (.I0(\REG.mem_5_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n60), .I3(GND_net), .O(n4768));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3566_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3565_3_lut (.I0(\REG.mem_5_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n60), .I3(GND_net), .O(n4767));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3564_3_lut (.I0(\REG.mem_5_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n60), .I3(GND_net), .O(n4766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3564_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3563_3_lut (.I0(\REG.mem_5_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n60), .I3(GND_net), .O(n4765));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3562_3_lut (.I0(\REG.mem_5_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n60), .I3(GND_net), .O(n4764));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3561_3_lut (.I0(\REG.mem_5_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n60), .I3(GND_net), .O(n4763));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3560_3_lut (.I0(\REG.mem_4_15 ), .I1(dc32_fifo_data_in[15]), 
            .I2(n61), .I3(GND_net), .O(n4762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4656_3_lut_4_lut (.I0(r_SM_Main_2__N_811[0]), .I1(fifo_read_cmd), 
            .I2(is_fifo_empty_flag), .I3(tx_uart_active_flag), .O(n5858));   // src/top.v(900[8] 918[4])
    defparam i4656_3_lut_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i3559_3_lut (.I0(\REG.mem_4_14 ), .I1(dc32_fifo_data_in[14]), 
            .I2(n61), .I3(GND_net), .O(n4761));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3558_3_lut (.I0(\REG.mem_4_13 ), .I1(dc32_fifo_data_in[13]), 
            .I2(n61), .I3(GND_net), .O(n4760));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3557_3_lut (.I0(\REG.mem_4_12 ), .I1(dc32_fifo_data_in[12]), 
            .I2(n61), .I3(GND_net), .O(n4759));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3556_3_lut (.I0(\REG.mem_4_11 ), .I1(dc32_fifo_data_in[11]), 
            .I2(n61), .I3(GND_net), .O(n4758));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3555_3_lut (.I0(\REG.mem_4_10 ), .I1(dc32_fifo_data_in[10]), 
            .I2(n61), .I3(GND_net), .O(n4757));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3554_3_lut (.I0(\REG.mem_4_9 ), .I1(dc32_fifo_data_in[9]), 
            .I2(n61), .I3(GND_net), .O(n4756));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3553_3_lut (.I0(\REG.mem_4_8 ), .I1(dc32_fifo_data_in[8]), 
            .I2(n61), .I3(GND_net), .O(n4755));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3552_3_lut (.I0(\REG.mem_4_7 ), .I1(dc32_fifo_data_in[7]), 
            .I2(n61), .I3(GND_net), .O(n4754));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3551_3_lut (.I0(\REG.mem_4_6 ), .I1(dc32_fifo_data_in[6]), 
            .I2(n61), .I3(GND_net), .O(n4753));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3550_3_lut (.I0(\REG.mem_4_5 ), .I1(dc32_fifo_data_in[5]), 
            .I2(n61), .I3(GND_net), .O(n4752));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3549_3_lut (.I0(\REG.mem_4_4 ), .I1(dc32_fifo_data_in[4]), 
            .I2(n61), .I3(GND_net), .O(n4751));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3548_3_lut (.I0(\REG.mem_4_3 ), .I1(dc32_fifo_data_in[3]), 
            .I2(n61), .I3(GND_net), .O(n4750));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3547_3_lut (.I0(\REG.mem_4_2 ), .I1(dc32_fifo_data_in[2]), 
            .I2(n61), .I3(GND_net), .O(n4749));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3546_3_lut (.I0(\REG.mem_4_1 ), .I1(dc32_fifo_data_in[1]), 
            .I2(n61), .I3(GND_net), .O(n4748));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3545_3_lut (.I0(\REG.mem_4_0 ), .I1(dc32_fifo_data_in[0]), 
            .I2(n61), .I3(GND_net), .O(n4747));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    defparam i3545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_1225[1]), .I1(r_SM_Main_2__N_808[1]), 
            .I2(r_SM_Main_adj_1225[0]), .I3(r_SM_Main_adj_1225[2]), .O(n14415));   // src/uart_tx.v(38[10] 141[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i4694_4_lut_4_lut (.I0(t_rd_fifo_en_w), .I1(reset_all), .I2(\REG.out_raw [6]), 
            .I3(fifo_data_out[6]), .O(n5896));
    defparam i4694_4_lut_4_lut.LUT_INIT = 16'h3120;
    SB_LUT4 i12_4_lut_4_lut_adj_103 (.I0(t_rd_fifo_en_w), .I1(reset_all), 
            .I2(\REG.out_raw [4]), .I3(fifo_data_out[4]), .O(n11137));
    defparam i12_4_lut_4_lut_adj_103.LUT_INIT = 16'h3120;
    SB_LUT4 i12_4_lut_4_lut_adj_104 (.I0(t_rd_fifo_en_w), .I1(reset_all), 
            .I2(\REG.out_raw [12]), .I3(fifo_data_out[12]), .O(n11133));
    defparam i12_4_lut_4_lut_adj_104.LUT_INIT = 16'h3120;
    SB_LUT4 i12_4_lut_4_lut_adj_105 (.I0(t_rd_fifo_en_w), .I1(reset_all), 
            .I2(\REG.out_raw [1]), .I3(fifo_data_out[1]), .O(n11143));
    defparam i12_4_lut_4_lut_adj_105.LUT_INIT = 16'h3120;
    SB_LUT4 i12_4_lut_4_lut_adj_106 (.I0(t_rd_fifo_en_w), .I1(reset_all), 
            .I2(\REG.out_raw [9]), .I3(fifo_data_out[9]), .O(n11095));
    defparam i12_4_lut_4_lut_adj_106.LUT_INIT = 16'h3120;
    SB_LUT4 i4625_2_lut_3_lut (.I0(fifo_data_out[6]), .I1(bluejay_data_out_31__N_703), 
            .I2(bluejay_data_out_31__N_704), .I3(GND_net), .O(n5827));   // src/bluejay_data.v(126[8] 148[4])
    defparam i4625_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i4624_2_lut_3_lut (.I0(fifo_data_out[5]), .I1(bluejay_data_out_31__N_703), 
            .I2(bluejay_data_out_31__N_704), .I3(GND_net), .O(n5826));   // src/bluejay_data.v(126[8] 148[4])
    defparam i4624_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i3407_3_lut (.I0(tx_data_byte[0]), .I1(pc_data_rx[0]), .I2(uart_rx_complete_rising_edge), 
            .I3(GND_net), .O(n4609));   // src/top.v(1064[8] 1131[4])
    defparam i3407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3544_3_lut (.I0(r_Tx_Data[1]), .I1(fifo_temp_output[1]), .I2(n3710), 
            .I3(GND_net), .O(n4746));   // src/uart_tx.v(38[10] 141[8])
    defparam i3544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3543_3_lut (.I0(r_Tx_Data[2]), .I1(fifo_temp_output[2]), .I2(n3710), 
            .I3(GND_net), .O(n4745));   // src/uart_tx.v(38[10] 141[8])
    defparam i3543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11065_4_lut (.I0(tx_data_byte[0]), .I1(tx_data_byte[1]), .I2(tx_data_byte[6]), 
            .I3(n11471), .O(multi_byte_spi_trans_flag_r_N_72));   // src/top.v(1113[10:31])
    defparam i11065_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i9823_4_lut (.I0(tx_data_byte[3]), .I1(tx_data_byte[2]), .I2(tx_data_byte[4]), 
            .I3(n11412), .O(n11471));
    defparam i9823_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i9764_2_lut (.I0(tx_data_byte[5]), .I1(tx_data_byte[7]), .I2(GND_net), 
            .I3(GND_net), .O(n11412));
    defparam i9764_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3542_3_lut (.I0(r_Tx_Data[3]), .I1(fifo_temp_output[3]), .I2(n3710), 
            .I3(GND_net), .O(n4744));   // src/uart_tx.v(38[10] 141[8])
    defparam i3542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3541_3_lut (.I0(r_Tx_Data[4]), .I1(fifo_temp_output[4]), .I2(n3710), 
            .I3(GND_net), .O(n4743));   // src/uart_tx.v(38[10] 141[8])
    defparam i3541_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3540_3_lut (.I0(r_Tx_Data[5]), .I1(fifo_temp_output[5]), .I2(n3710), 
            .I3(GND_net), .O(n4742));   // src/uart_tx.v(38[10] 141[8])
    defparam i3540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3538_3_lut (.I0(r_Tx_Data[6]), .I1(fifo_temp_output[6]), .I2(n3710), 
            .I3(GND_net), .O(n4740));   // src/uart_tx.v(38[10] 141[8])
    defparam i3538_3_lut.LUT_INIT = 16'hcaca;
    clock clock_inst (.GND_net(GND_net), .VCC_net(VCC_net), .ICE_SYSCLK_c(ICE_SYSCLK_c), 
          .pll_clk_unbuf(pll_clk_unbuf)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(222[7] 228[3])
    spi spi0 (.\tx_data_byte[1] (tx_data_byte[1]), .\tx_shift_reg[0] (tx_shift_reg[0]), 
        .n1928(n1928), .GND_net(GND_net), .\tx_data_byte[2] (tx_data_byte[2]), 
        .\tx_data_byte[3] (tx_data_byte[3]), .VCC_net(VCC_net), .SEN_c_1(SEN_c_1), 
        .SLM_CLK_c(SLM_CLK_c), .SOUT_c(SOUT_c), .n4093(n4093), .\rx_shift_reg[0] (rx_shift_reg[0]), 
        .\tx_data_byte[4] (tx_data_byte[4]), .\tx_data_byte[5] (tx_data_byte[5]), 
        .\tx_data_byte[6] (tx_data_byte[6]), .\tx_data_byte[7] (tx_data_byte[7]), 
        .tx_addr_byte({tx_addr_byte}), .n4070(n4070), .SDAT_c_15(SDAT_c_15), 
        .multi_byte_spi_trans_flag_r(multi_byte_spi_trans_flag_r), .n11007(n11007), 
        .n5756(n5756), .\rx_shift_reg[1] (rx_shift_reg[1]), .n5755(n5755), 
        .\rx_shift_reg[2] (rx_shift_reg[2]), .n5754(n5754), .\rx_shift_reg[3] (rx_shift_reg[3]), 
        .n5753(n5753), .\rx_shift_reg[4] (rx_shift_reg[4]), .n5752(n5752), 
        .\rx_shift_reg[5] (rx_shift_reg[5]), .n5751(n5751), .\rx_shift_reg[6] (rx_shift_reg[6]), 
        .n5750(n5750), .\rx_shift_reg[7] (rx_shift_reg[7]), .n5733(n5733), 
        .rx_buf_byte({rx_buf_byte}), .n5732(n5732), .n5731(n5731), .n5730(n5730), 
        .n5729(n5729), .n5728(n5728), .n5727(n5727), .spi_rx_byte_ready(spi_rx_byte_ready), 
        .SCK_c_0(SCK_c_0), .spi_start_transfer_r(spi_start_transfer_r), 
        .n4637(n4637), .n3204(n3204)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(823[5] 847[2])
    \uart_tx(CLKS_PER_BIT=20)  pc_tx (.UART_TX_c(UART_TX_c), .SLM_CLK_c(SLM_CLK_c), 
            .r_SM_Main({r_SM_Main_adj_1225}), .n4724(n4724), .r_Tx_Data({r_Tx_Data}), 
            .n5861(n5861), .VCC_net(VCC_net), .r_Bit_Index({Open_0, Open_1, 
            r_Bit_Index_adj_1227[0]}), .n14415(n14415), .\r_SM_Main_2__N_808[1] (r_SM_Main_2__N_808[1]), 
            .GND_net(GND_net), .n4133(n4133), .\r_SM_Main_2__N_811[0] (r_SM_Main_2__N_811[0]), 
            .n4632(n4632), .n4631(n4631), .tx_uart_active_flag(tx_uart_active_flag), 
            .n11319(n11319), .n3710(n3710), .n4746(n4746), .n4745(n4745), 
            .n4744(n4744), .n4743(n4743), .n4742(n4742), .n4740(n4740), 
            .n11339(n11339)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(758[42] 767[3])
    FIFO_Quad_Word tx_fifo (.rd_fifo_en_w(rd_fifo_en_w), .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r [0]), 
            .SLM_CLK_c(SLM_CLK_c), .rd_addr_r({rd_addr_r_adj_1252}), .reset_all_w(reset_all_w), 
            .wr_addr_r({wr_addr_r_adj_1249}), .n5905(n5905), .VCC_net(VCC_net), 
            .\fifo_temp_output[7] (fifo_temp_output[7]), .\rd_addr_p1_w[2] (rd_addr_p1_w_adj_1254[2]), 
            .GND_net(GND_net), .n5902(n5902), .\fifo_temp_output[6] (fifo_temp_output[6]), 
            .n5899(n5899), .\fifo_temp_output[5] (fifo_temp_output[5]), 
            .n5890(n5890), .\fifo_temp_output[4] (fifo_temp_output[4]), 
            .n5887(n5887), .\fifo_temp_output[3] (fifo_temp_output[3]), 
            .n5884(n5884), .\fifo_temp_output[2] (fifo_temp_output[2]), 
            .n1(n1), .n5881(n5881), .\fifo_temp_output[1] (fifo_temp_output[1]), 
            .n10921(n10921), .is_tx_fifo_full_flag(is_tx_fifo_full_flag), 
            .\wr_addr_p1_w[2] (wr_addr_p1_w_adj_1251[2]), .n5857(n5857), 
            .\fifo_temp_output[0] (fifo_temp_output[0]), .n10727(n10727), 
            .\rd_addr_p1_w[1] (rd_addr_p1_w_adj_1254[1]), .n4679(n4679), 
            .rx_buf_byte({rx_buf_byte}), .n4670(n4670), .n11324(n11324), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .n4674(n4674), .n4697(n4697), 
            .fifo_write_cmd(fifo_write_cmd), .full_nxt_r(full_nxt_r), .n2207(n2207), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r [7]), .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r [6]), 
            .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r [5]), .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r [4]), 
            .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r [3]), .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r [2]), 
            .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r [1]), .n4700(n4700), 
            .fifo_read_cmd(fifo_read_cmd), .n4249(n4249), .empty_o_N_1116(empty_o_N_1116)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(923[16] 939[2])
    usb3_if usb3_if_inst (.VCC_net(VCC_net), .GND_net(GND_net), .\dc32_fifo_data_in[13] (dc32_fifo_data_in[13]), 
            .DEBUG_6_c_c(DEBUG_6_c_c), .\dc32_fifo_data_in[12] (dc32_fifo_data_in[12]), 
            .\dc32_fifo_data_in[11] (dc32_fifo_data_in[11]), .\dc32_fifo_data_in[10] (dc32_fifo_data_in[10]), 
            .\dc32_fifo_data_in[9] (dc32_fifo_data_in[9]), .\dc32_fifo_data_in[8] (dc32_fifo_data_in[8]), 
            .\dc32_fifo_data_in[7] (dc32_fifo_data_in[7]), .\dc32_fifo_data_in[6] (dc32_fifo_data_in[6]), 
            .\dc32_fifo_data_in[5] (dc32_fifo_data_in[5]), .\dc32_fifo_data_in[4] (dc32_fifo_data_in[4]), 
            .DEBUG_3_c(DEBUG_3_c), .\dc32_fifo_data_in[0] (dc32_fifo_data_in[0]), 
            .buffer_switch_done(buffer_switch_done), .buffer_switch_done_latched(buffer_switch_done_latched), 
            .SLM_CLK_c(SLM_CLK_c), .reset_per_frame(reset_per_frame), .FT_OE_c(FT_OE_c), 
            .\dc32_fifo_data_in[3] (dc32_fifo_data_in[3]), .DEBUG_9_c(DEBUG_9_c), 
            .\dc32_fifo_data_in[2] (dc32_fifo_data_in[2]), .\dc32_fifo_data_in[1] (dc32_fifo_data_in[1]), 
            .DEBUG_2_c_c(DEBUG_2_c_c), .\dc32_fifo_data_in[15] (dc32_fifo_data_in[15]), 
            .DEBUG_5_c(DEBUG_5_c), .FIFO_D15_c_15(FIFO_D15_c_15), .FIFO_D14_c_14(FIFO_D14_c_14), 
            .FIFO_D13_c_13(FIFO_D13_c_13), .FIFO_D12_c_12(FIFO_D12_c_12), 
            .FIFO_D11_c_11(FIFO_D11_c_11), .FIFO_D10_c_10(FIFO_D10_c_10), 
            .FIFO_D9_c_9(FIFO_D9_c_9), .FIFO_D8_c_8(FIFO_D8_c_8), .FIFO_D7_c_7(FIFO_D7_c_7), 
            .FIFO_D6_c_6(FIFO_D6_c_6), .FIFO_D5_c_5(FIFO_D5_c_5), .FIFO_D4_c_4(FIFO_D4_c_4), 
            .FIFO_D3_c_3(FIFO_D3_c_3), .FIFO_D2_c_2(FIFO_D2_c_2), .FIFO_D1_c_1(FIFO_D1_c_1), 
            .\afull_flag_impl.af_flag_p_w_N_603[3] (\afull_flag_impl.af_flag_p_w_N_603 [3]), 
            .\dc32_fifo_data_in[14] (dc32_fifo_data_in[14]), .DEBUG_1_c_0_c(DEBUG_1_c_0_c)) /* synthesis syn_module_defined=1 */ ;   // src/top.v(503[9] 520[3])
    
endmodule
//
// Verilog Description of module timing_controller
//

module timing_controller (state, SLM_CLK_c, n1721, GND_net, VCC_net, 
            n63, n4, n11342, reset_per_frame, n1616, n7383, INVERT_c_4, 
            reset_all, n7495, buffer_switch_done, n11015, n3514, n7566, 
            n11376, UPDATE_c_3, n3929) /* synthesis syn_module_defined=1 */ ;
    output [3:0]state;
    input SLM_CLK_c;
    input n1721;
    input GND_net;
    input VCC_net;
    output n63;
    output n4;
    input n11342;
    output reset_per_frame;
    input n1616;
    input n7383;
    output INVERT_c_4;
    output reset_all;
    input n7495;
    output buffer_switch_done;
    input n11015;
    output n3514;
    output n7566;
    output n11376;
    output UPDATE_c_3;
    output n3929;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [3:0]state_3__N_80;
    
    wire n11377, n12554;
    wire [31:0]n1722;
    
    wire n12553, n11368, n1793;
    wire [31:0]n1794;
    
    wire n10591;
    wire [31:0]state_timeout_counter;   // src/timing_controller.v(49[12:33])
    
    wire n10592, n10609, n10610;
    wire [31:0]n506;
    
    wire n10608, n12552, n10590, n12542, n10607, n12544, n10606, 
        n10589, n12545, n10605, n10604, n10588, n10603, n12547, 
        n10602, n12532, n12548, n10601, n10600, n12549, n10599, 
        n10618, n10617, n10598, n10616, n4301, n4589, n4586;
    wire [4:0]n858;
    
    wire n11353, n10615, n12550, n10597, n10614, n12551, n10596, 
        n10613, n10595, n4200, n11347, n1875, n11354, n10612, 
        n10594, n12539, n10611, n10593, n11375, n38, n52, n56, 
        n54, n12555, n55, n53, n50, n58, n62, n49, n7592, 
        n12604, n7, n12540, n12698, n5, n12541;
    
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n11377), .D(state_3__N_80[0]));   // src/timing_controller.v(53[8] 129[4])
    SB_LUT4 state_3__I_0_59_Mux_2_i15_4_lut (.I0(state[1]), .I1(state[2]), 
            .I2(state[3]), .I3(state[0]), .O(state_3__N_80[2]));   // src/timing_controller.v(59[5] 128[12])
    defparam state_3__I_0_59_Mux_2_i15_4_lut.LUT_INIT = 16'hc2ce;
    SB_LUT4 mux_855_i2_3_lut (.I0(n12554), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[1]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_855_i3_3_lut (.I0(n12553), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[2]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_863_i25_3_lut_4_lut (.I0(state[1]), .I1(n11368), .I2(n1793), 
            .I3(n1722[24]), .O(n1794[24]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_863_i25_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_863_i24_3_lut_4_lut (.I0(state[1]), .I1(n11368), .I2(n1793), 
            .I3(n1722[23]), .O(n1794[23]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_863_i24_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_863_i23_3_lut_4_lut (.I0(state[1]), .I1(n11368), .I2(n1793), 
            .I3(n1722[22]), .O(n1794[22]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_863_i23_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_863_i21_3_lut_4_lut (.I0(state[1]), .I1(n11368), .I2(n1793), 
            .I3(n1722[20]), .O(n1794[20]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_863_i21_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_863_i20_3_lut_4_lut (.I0(state[1]), .I1(n11368), .I2(n1793), 
            .I3(n1722[19]), .O(n1794[19]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_863_i20_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_863_i19_3_lut_4_lut (.I0(state[1]), .I1(n11368), .I2(n1793), 
            .I3(n1722[18]), .O(n1794[18]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_863_i19_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_863_i16_3_lut_4_lut (.I0(state[1]), .I1(n11368), .I2(n1793), 
            .I3(n1722[15]), .O(n1794[15]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_863_i16_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_CARRY sub_31_add_2_6 (.CI(n10591), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n10592));
    SB_LUT4 mux_863_i15_3_lut_4_lut (.I0(state[1]), .I1(n11368), .I2(n1793), 
            .I3(n1722[14]), .O(n1794[14]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_863_i15_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_863_i13_3_lut_4_lut (.I0(state[1]), .I1(n11368), .I2(n1793), 
            .I3(n1722[12]), .O(n1794[12]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_863_i13_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_863_i10_3_lut_4_lut (.I0(state[1]), .I1(n11368), .I2(n1793), 
            .I3(n1722[9]), .O(n1794[9]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_863_i10_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_863_i11_3_lut_4_lut (.I0(state[1]), .I1(n11368), .I2(n1793), 
            .I3(n1722[10]), .O(n1794[10]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_863_i11_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 mux_863_i4_3_lut_4_lut (.I0(state[1]), .I1(n11368), .I2(n1793), 
            .I3(n1722[3]), .O(n1794[3]));   // src/timing_controller.v(53[8] 129[4])
    defparam mux_863_i4_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i1_2_lut (.I0(state[2]), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n4));   // src/timing_controller.v(59[5] 128[12])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_DFF invert_55_i1 (.Q(reset_per_frame), .C(SLM_CLK_c), .D(n11342));   // src/timing_controller.v(59[5] 128[12])
    SB_CARRY sub_31_add_2_24 (.CI(n10609), .I0(state_timeout_counter[22]), 
            .I1(VCC_net), .CO(n10610));
    SB_LUT4 sub_31_add_2_23_lut (.I0(GND_net), .I1(state_timeout_counter[21]), 
            .I2(VCC_net), .I3(n10608), .O(n506[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_23 (.CI(n10608), .I0(state_timeout_counter[21]), 
            .I1(VCC_net), .CO(n10609));
    SB_LUT4 sub_31_add_2_5_lut (.I0(n1616), .I1(state_timeout_counter[3]), 
            .I2(VCC_net), .I3(n10590), .O(n12552)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_5 (.CI(n10590), .I0(state_timeout_counter[3]), 
            .I1(VCC_net), .CO(n10591));
    SB_LUT4 sub_31_add_2_22_lut (.I0(n1616), .I1(state_timeout_counter[20]), 
            .I2(VCC_net), .I3(n10607), .O(n12542)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_22 (.CI(n10607), .I0(state_timeout_counter[20]), 
            .I1(VCC_net), .CO(n10608));
    SB_LUT4 sub_31_add_2_21_lut (.I0(n1616), .I1(state_timeout_counter[19]), 
            .I2(VCC_net), .I3(n10606), .O(n12544)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_21 (.CI(n10606), .I0(state_timeout_counter[19]), 
            .I1(VCC_net), .CO(n10607));
    SB_LUT4 sub_31_add_2_4_lut (.I0(n7383), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n10589), .O(n12553)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_4_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_31_add_2_4 (.CI(n10589), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n10590));
    SB_LUT4 sub_31_add_2_20_lut (.I0(n1616), .I1(state_timeout_counter[18]), 
            .I2(VCC_net), .I3(n10605), .O(n12545)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_20 (.CI(n10605), .I0(state_timeout_counter[18]), 
            .I1(VCC_net), .CO(n10606));
    SB_LUT4 sub_31_add_2_19_lut (.I0(GND_net), .I1(state_timeout_counter[17]), 
            .I2(VCC_net), .I3(n10604), .O(n506[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_19 (.CI(n10604), .I0(state_timeout_counter[17]), 
            .I1(VCC_net), .CO(n10605));
    SB_LUT4 sub_31_add_2_3_lut (.I0(n1616), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n10588), .O(n12554)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_3 (.CI(n10588), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n10589));
    SB_LUT4 sub_31_add_2_18_lut (.I0(GND_net), .I1(state_timeout_counter[16]), 
            .I2(VCC_net), .I3(n10603), .O(n506[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_18 (.CI(n10603), .I0(state_timeout_counter[16]), 
            .I1(VCC_net), .CO(n10604));
    SB_LUT4 sub_31_add_2_17_lut (.I0(n1616), .I1(state_timeout_counter[15]), 
            .I2(VCC_net), .I3(n10602), .O(n12547)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_17 (.CI(n10602), .I0(state_timeout_counter[15]), 
            .I1(VCC_net), .CO(n10603));
    SB_LUT4 sub_31_add_2_2_lut (.I0(n7383), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n12532)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_31_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n10588));
    SB_LUT4 sub_31_add_2_16_lut (.I0(n1616), .I1(state_timeout_counter[14]), 
            .I2(VCC_net), .I3(n10601), .O(n12548)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_16 (.CI(n10601), .I0(state_timeout_counter[14]), 
            .I1(VCC_net), .CO(n10602));
    SB_LUT4 sub_31_add_2_15_lut (.I0(GND_net), .I1(state_timeout_counter[13]), 
            .I2(VCC_net), .I3(n10600), .O(n506[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_15 (.CI(n10600), .I0(state_timeout_counter[13]), 
            .I1(VCC_net), .CO(n10601));
    SB_LUT4 sub_31_add_2_14_lut (.I0(n1616), .I1(state_timeout_counter[12]), 
            .I2(VCC_net), .I3(n10599), .O(n12549)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_33_lut (.I0(GND_net), .I1(state_timeout_counter[31]), 
            .I2(VCC_net), .I3(n10618), .O(n506[31])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_32_lut (.I0(GND_net), .I1(state_timeout_counter[30]), 
            .I2(VCC_net), .I3(n10617), .O(n506[30])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_14 (.CI(n10599), .I0(state_timeout_counter[12]), 
            .I1(VCC_net), .CO(n10600));
    SB_LUT4 sub_31_add_2_13_lut (.I0(GND_net), .I1(state_timeout_counter[11]), 
            .I2(VCC_net), .I3(n10598), .O(n506[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_32 (.CI(n10617), .I0(state_timeout_counter[30]), 
            .I1(VCC_net), .CO(n10618));
    SB_LUT4 sub_31_add_2_31_lut (.I0(GND_net), .I1(state_timeout_counter[29]), 
            .I2(VCC_net), .I3(n10616), .O(n506[29])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_13 (.CI(n10598), .I0(state_timeout_counter[11]), 
            .I1(VCC_net), .CO(n10599));
    SB_DFFESR state_timeout_counter_i0_i31 (.Q(state_timeout_counter[31]), 
            .C(SLM_CLK_c), .E(n4301), .D(n506[31]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i30 (.Q(state_timeout_counter[30]), 
            .C(SLM_CLK_c), .E(n4301), .D(n506[30]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i29 (.Q(state_timeout_counter[29]), 
            .C(SLM_CLK_c), .E(n4301), .D(n506[29]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_CARRY sub_31_add_2_31 (.CI(n10616), .I0(state_timeout_counter[29]), 
            .I1(VCC_net), .CO(n10617));
    SB_DFFESR state_timeout_counter_i0_i28 (.Q(state_timeout_counter[28]), 
            .C(SLM_CLK_c), .E(n4301), .D(n506[28]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i27 (.Q(state_timeout_counter[27]), 
            .C(SLM_CLK_c), .E(n4301), .D(n506[27]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i26 (.Q(state_timeout_counter[26]), 
            .C(SLM_CLK_c), .E(n4301), .D(n506[26]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i25 (.Q(state_timeout_counter[25]), 
            .C(SLM_CLK_c), .E(n4301), .D(n506[25]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i21 (.Q(state_timeout_counter[21]), 
            .C(SLM_CLK_c), .E(n4301), .D(n506[21]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i17 (.Q(state_timeout_counter[17]), 
            .C(SLM_CLK_c), .E(n4301), .D(n506[17]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i16 (.Q(state_timeout_counter[16]), 
            .C(SLM_CLK_c), .E(n4301), .D(n506[16]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i13 (.Q(state_timeout_counter[13]), 
            .C(SLM_CLK_c), .E(n4301), .D(n506[13]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i11 (.Q(state_timeout_counter[11]), 
            .C(SLM_CLK_c), .E(n4301), .D(n506[11]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i8 (.Q(state_timeout_counter[8]), .C(SLM_CLK_c), 
            .E(n4301), .D(n506[8]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(SLM_CLK_c), 
            .E(n4301), .D(n506[7]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n4301), .D(n506[6]), .R(n4589));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1722[2]), .R(n4586));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFESR state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1722[1]), .R(n4586));   // src/timing_controller.v(53[8] 129[4])
    SB_DFF invert_55_i4 (.Q(INVERT_c_4), .C(SLM_CLK_c), .D(n858[4]));   // src/timing_controller.v(59[5] 128[12])
    SB_DFF invert_55_i0 (.Q(reset_all), .C(SLM_CLK_c), .D(n11353));   // src/timing_controller.v(59[5] 128[12])
    SB_LUT4 sub_31_add_2_30_lut (.I0(GND_net), .I1(state_timeout_counter[28]), 
            .I2(VCC_net), .I3(n10615), .O(n506[28])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_12_lut (.I0(n1616), .I1(state_timeout_counter[10]), 
            .I2(VCC_net), .I3(n10597), .O(n12550)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_12 (.CI(n10597), .I0(state_timeout_counter[10]), 
            .I1(VCC_net), .CO(n10598));
    SB_CARRY sub_31_add_2_30 (.CI(n10615), .I0(state_timeout_counter[28]), 
            .I1(VCC_net), .CO(n10616));
    SB_LUT4 sub_31_add_2_29_lut (.I0(GND_net), .I1(state_timeout_counter[27]), 
            .I2(VCC_net), .I3(n10614), .O(n506[27])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_11_lut (.I0(n1616), .I1(state_timeout_counter[9]), 
            .I2(VCC_net), .I3(n10596), .O(n12551)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_31_add_2_11 (.CI(n10596), .I0(state_timeout_counter[9]), 
            .I1(VCC_net), .CO(n10597));
    SB_CARRY sub_31_add_2_29 (.CI(n10614), .I0(state_timeout_counter[27]), 
            .I1(VCC_net), .CO(n10615));
    SB_LUT4 sub_31_add_2_28_lut (.I0(GND_net), .I1(state_timeout_counter[26]), 
            .I2(VCC_net), .I3(n10613), .O(n506[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_10_lut (.I0(GND_net), .I1(state_timeout_counter[8]), 
            .I2(VCC_net), .I3(n10595), .O(n506[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n4200), .D(state_3__N_80[2]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n4200), .D(state_3__N_80[1]));   // src/timing_controller.v(53[8] 129[4])
    SB_LUT4 i1_2_lut_adj_86 (.I0(n1616), .I1(n1721), .I2(GND_net), .I3(GND_net), 
            .O(n11347));   // src/timing_controller.v(59[5] 128[12])
    defparam i1_2_lut_adj_86.LUT_INIT = 16'h2222;
    SB_LUT4 i924_4_lut (.I0(state[3]), .I1(n1875), .I2(n7495), .I3(state[2]), 
            .O(n1793));   // src/timing_controller.v(53[8] 129[4])
    defparam i924_4_lut.LUT_INIT = 16'h0544;
    SB_DFF invert_55_i2 (.Q(buffer_switch_done), .C(SLM_CLK_c), .D(n11354));   // src/timing_controller.v(59[5] 128[12])
    SB_CARRY sub_31_add_2_10 (.CI(n10595), .I0(state_timeout_counter[8]), 
            .I1(VCC_net), .CO(n10596));
    SB_CARRY sub_31_add_2_28 (.CI(n10613), .I0(state_timeout_counter[26]), 
            .I1(VCC_net), .CO(n10614));
    SB_LUT4 sub_31_add_2_27_lut (.I0(GND_net), .I1(state_timeout_counter[25]), 
            .I2(VCC_net), .I3(n10612), .O(n506[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_31_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n10594), .O(n506[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_9 (.CI(n10594), .I0(state_timeout_counter[7]), 
            .I1(VCC_net), .CO(n10595));
    SB_DFF state_i3 (.Q(state[3]), .C(SLM_CLK_c), .D(n11015));   // src/timing_controller.v(53[8] 129[4])
    SB_CARRY sub_31_add_2_27 (.CI(n10612), .I0(state_timeout_counter[25]), 
            .I1(VCC_net), .CO(n10613));
    SB_LUT4 sub_31_add_2_26_lut (.I0(n1616), .I1(state_timeout_counter[24]), 
            .I2(VCC_net), .I3(n10611), .O(n12539)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_31_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n10593), .O(n506[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_31_add_2_26 (.CI(n10611), .I0(state_timeout_counter[24]), 
            .I1(VCC_net), .CO(n10612));
    SB_DFFE state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[0]));   // src/timing_controller.v(53[8] 129[4])
    SB_LUT4 i1_2_lut_3_lut (.I0(state[2]), .I1(state[0]), .I2(n63), .I3(GND_net), 
            .O(n11375));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2319_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n3514));   // src/timing_controller.v(59[5] 128[12])
    defparam i2319_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6388_3_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n7566));
    defparam i6388_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY sub_31_add_2_8 (.CI(n10593), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n10594));
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(state[3]), 
            .I3(state[2]), .O(n11354));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_4_lut_adj_87 (.I0(state[0]), .I1(state[1]), .I2(state[3]), 
            .I3(state[2]), .O(n11353));
    defparam i1_2_lut_4_lut_adj_87.LUT_INIT = 16'h0002;
    SB_DFFE state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[3]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[4]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[5]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i9 (.Q(state_timeout_counter[9]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[9]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i10 (.Q(state_timeout_counter[10]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[10]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i12 (.Q(state_timeout_counter[12]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[12]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i14 (.Q(state_timeout_counter[14]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[14]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i15 (.Q(state_timeout_counter[15]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[15]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i18 (.Q(state_timeout_counter[18]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[18]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i19 (.Q(state_timeout_counter[19]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[19]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i20 (.Q(state_timeout_counter[20]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[20]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i22 (.Q(state_timeout_counter[22]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[22]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i23 (.Q(state_timeout_counter[23]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[23]));   // src/timing_controller.v(53[8] 129[4])
    SB_DFFE state_timeout_counter_i0_i24 (.Q(state_timeout_counter[24]), .C(SLM_CLK_c), 
            .E(n4301), .D(n1794[24]));   // src/timing_controller.v(53[8] 129[4])
    SB_LUT4 i6_2_lut (.I0(state_timeout_counter[9]), .I1(state_timeout_counter[12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // src/timing_controller.v(81[17:45])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut (.I0(state_timeout_counter[17]), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[24]), .I3(state_timeout_counter[4]), 
            .O(n52));   // src/timing_controller.v(81[17:45])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(state_timeout_counter[29]), .I1(state_timeout_counter[3]), 
            .I2(state_timeout_counter[13]), .I3(state_timeout_counter[31]), 
            .O(n56));   // src/timing_controller.v(81[17:45])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(state_timeout_counter[19]), .I1(state_timeout_counter[5]), 
            .I2(state_timeout_counter[22]), .I3(state_timeout_counter[6]), 
            .O(n54));   // src/timing_controller.v(81[17:45])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_31_add_2_7_lut (.I0(n11347), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n10592), .O(n12555)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i23_4_lut (.I0(state_timeout_counter[10]), .I1(state_timeout_counter[15]), 
            .I2(state_timeout_counter[20]), .I3(state_timeout_counter[23]), 
            .O(n55));   // src/timing_controller.v(81[17:45])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(state_timeout_counter[27]), .I1(state_timeout_counter[7]), 
            .I2(state_timeout_counter[30]), .I3(state_timeout_counter[14]), 
            .O(n53));   // src/timing_controller.v(81[17:45])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(state_timeout_counter[8]), .I1(state_timeout_counter[11]), 
            .I2(state_timeout_counter[16]), .I3(state_timeout_counter[21]), 
            .O(n50));   // src/timing_controller.v(81[17:45])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i913_2_lut_3_lut (.I0(state[0]), .I1(n63), .I2(state[1]), 
            .I3(GND_net), .O(n1875));   // src/timing_controller.v(53[8] 129[4])
    defparam i913_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i26_4_lut (.I0(state_timeout_counter[25]), .I1(n52), .I2(n38), 
            .I3(state_timeout_counter[26]), .O(n58));   // src/timing_controller.v(81[17:45])
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 state_3__I_0_59_Mux_1_i15_4_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[3]), .I3(n11375), .O(state_3__N_80[1]));   // src/timing_controller.v(59[5] 128[12])
    defparam state_3__I_0_59_Mux_1_i15_4_lut_4_lut.LUT_INIT = 16'hc6f6;
    SB_LUT4 i30_4_lut (.I0(n53), .I1(n55), .I2(n54), .I3(n56), .O(n62));   // src/timing_controller.v(81[17:45])
    defparam i30_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(state_timeout_counter[0]), .I1(state_timeout_counter[18]), 
            .I2(state_timeout_counter[28]), .I3(state_timeout_counter[2]), 
            .O(n49));   // src/timing_controller.v(81[17:45])
    defparam i17_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i31_4_lut (.I0(n49), .I1(n62), .I2(n58), .I3(n50), .O(n63));   // src/timing_controller.v(81[17:45])
    defparam i31_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_88 (.I0(state[3]), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n11376));
    defparam i1_2_lut_adj_88.LUT_INIT = 16'hbbbb;
    SB_CARRY sub_31_add_2_7 (.CI(n10592), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n10593));
    SB_LUT4 i6413_3_lut (.I0(n63), .I1(state[1]), .I2(state[2]), .I3(GND_net), 
            .O(n7592));
    defparam i6413_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 sub_31_add_2_6_lut (.I0(n1616), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n10591), .O(n12604)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 state_3__I_0_59_Mux_0_i7_4_lut (.I0(state[1]), .I1(n63), .I2(state[2]), 
            .I3(state[0]), .O(n7));   // src/timing_controller.v(59[5] 128[12])
    defparam state_3__I_0_59_Mux_0_i7_4_lut.LUT_INIT = 16'hc535;
    SB_LUT4 state_3__I_0_59_Mux_0_i15_4_lut (.I0(n7), .I1(n7592), .I2(state[3]), 
            .I3(state[0]), .O(state_3__N_80[0]));   // src/timing_controller.v(59[5] 128[12])
    defparam state_3__I_0_59_Mux_0_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 sub_31_add_2_25_lut (.I0(n1616), .I1(state_timeout_counter[23]), 
            .I2(VCC_net), .I3(n10610), .O(n12540)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_25_lut.LUT_INIT = 16'h8228;
    SB_DFFESR invert_55_i3 (.Q(UPDATE_c_3), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n12698), .R(n5));   // src/timing_controller.v(59[5] 128[12])
    SB_CARRY sub_31_add_2_25 (.CI(n10610), .I0(state_timeout_counter[23]), 
            .I1(VCC_net), .CO(n10611));
    SB_LUT4 sub_31_add_2_24_lut (.I0(n1616), .I1(state_timeout_counter[22]), 
            .I2(VCC_net), .I3(n10609), .O(n12541)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_31_add_2_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11069_2_lut_3_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(state[1]), 
            .I3(state[0]), .O(n4301));   // src/timing_controller.v(59[5] 128[12])
    defparam i11069_2_lut_3_lut_4_lut.LUT_INIT = 16'h5557;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[3]), .I1(n63), .I2(state[1]), .I3(state[2]), 
            .O(n11377));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[0]), .I1(n63), .I2(state[3]), 
            .I3(state[2]), .O(n11368));   // src/timing_controller.v(53[8] 129[4])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_adj_89 (.I0(state[2]), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n3929));   // src/timing_controller.v(59[5] 128[12])
    defparam i1_2_lut_3_lut_adj_89.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_863_i1_4_lut (.I0(n1722[0]), .I1(state[1]), .I2(n1793), 
            .I3(n11368), .O(n1794[0]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_863_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 mux_855_i1_3_lut (.I0(n12532), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[0]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i1_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i11088_2_lut (.I0(state[3]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // src/timing_controller.v(53[8] 129[4])
    defparam i11088_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i11121_3_lut_4_lut (.I0(state[3]), .I1(n3929), .I2(n1793), 
            .I3(n11347), .O(n4589));
    defparam i11121_3_lut_4_lut.LUT_INIT = 16'h7077;
    SB_LUT4 mux_855_i4_3_lut (.I0(n12552), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[3]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9812_4_lut (.I0(n12604), .I1(state[1]), .I2(n1721), .I3(n1793), 
            .O(n1794[4]));   // src/timing_controller.v(59[5] 128[12])
    defparam i9812_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_863_i6_3_lut (.I0(n12555), .I1(state[1]), .I2(n1793), 
            .I3(GND_net), .O(n1794[5]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_863_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_855_i10_3_lut (.I0(n12551), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[9]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_855_i11_3_lut (.I0(n12550), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[10]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i11_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_855_i13_3_lut (.I0(n12549), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[12]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i13_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_855_i15_3_lut (.I0(n12548), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[14]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i15_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_855_i16_3_lut (.I0(n12547), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[15]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_855_i19_3_lut (.I0(n12545), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[18]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i19_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_855_i20_3_lut (.I0(n12544), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[19]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_855_i21_3_lut (.I0(n12542), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[20]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i21_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_855_i23_3_lut (.I0(n12541), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[22]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i23_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_855_i24_3_lut (.I0(n12540), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[23]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_855_i25_3_lut (.I0(n12539), .I1(state[1]), .I2(n1721), 
            .I3(GND_net), .O(n1722[24]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_855_i25_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i11049_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n12698));   // src/timing_controller.v(59[5] 128[12])
    defparam i11049_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i3384_2_lut_3_lut (.I0(state[3]), .I1(n3929), .I2(n1793), 
            .I3(GND_net), .O(n4586));   // src/timing_controller.v(53[8] 129[4])
    defparam i3384_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 mux_321_Mux_4_i15_4_lut_4_lut (.I0(state[2]), .I1(state[0]), 
            .I2(state[1]), .I3(state[3]), .O(n858[4]));   // src/timing_controller.v(59[5] 128[12])
    defparam mux_321_Mux_4_i15_4_lut_4_lut.LUT_INIT = 16'h01a0;
    SB_LUT4 i1_2_lut_4_lut_adj_90 (.I0(state[2]), .I1(state[0]), .I2(state[1]), 
            .I3(n11376), .O(n4200));
    defparam i1_2_lut_4_lut_adj_90.LUT_INIT = 16'hff01;
    
endmodule
//
// Verilog Description of module bluejay_data
//

module bluejay_data (VCC_net, VALID_c, SLM_CLK_c, \state_timeout_counter[3] , 
            buffer_switch_done_latched, bluejay_data_out_31__N_704, n5870, 
            DATA16_c, DATA15_c, DATA14_c, DATA13_c, DATA12_c, DATA11_c, 
            DATA10_c, DATA9_c, DATA8_c, DATA7_c, n5827, DATA6_c, 
            n5826, DATA5_c, DATA20_c, DATA19_c, DATA18_c, DATA17_c, 
            GND_net, SYNC_c, buffer_switch_done, bluejay_data_out_31__N_703, 
            n14424, n718, n7, n5, \rd_sig_diff0_w[0] , \rd_sig_diff0_w[1] , 
            get_next_word, \aempty_flag_impl.ae_flag_nxt_w , DEBUG_9_c, 
            dc32_fifo_almost_empty, DEBUG_5_c, reset_all, n4667, \fifo_data_out[15] , 
            \fifo_data_out[14] , \fifo_data_out[13] , \fifo_data_out[12] , 
            \fifo_data_out[11] , \fifo_data_out[10] , \fifo_data_out[9] , 
            \fifo_data_out[8] , \fifo_data_out[7] , \fifo_data_out[4] , 
            \fifo_data_out[3] , \fifo_data_out[2] , \fifo_data_out[1] ) /* synthesis syn_module_defined=1 */ ;
    input VCC_net;
    output VALID_c;
    input SLM_CLK_c;
    output \state_timeout_counter[3] ;
    input buffer_switch_done_latched;
    output bluejay_data_out_31__N_704;
    input n5870;
    output DATA16_c;
    output DATA15_c;
    output DATA14_c;
    output DATA13_c;
    output DATA12_c;
    output DATA11_c;
    output DATA10_c;
    output DATA9_c;
    output DATA8_c;
    output DATA7_c;
    input n5827;
    output DATA6_c;
    input n5826;
    output DATA5_c;
    output DATA20_c;
    output DATA19_c;
    output DATA18_c;
    output DATA17_c;
    input GND_net;
    output SYNC_c;
    input buffer_switch_done;
    output bluejay_data_out_31__N_703;
    input n14424;
    output n718;
    output n7;
    input n5;
    input \rd_sig_diff0_w[0] ;
    input \rd_sig_diff0_w[1] ;
    output get_next_word;
    output \aempty_flag_impl.ae_flag_nxt_w ;
    input DEBUG_9_c;
    input dc32_fifo_almost_empty;
    input DEBUG_5_c;
    input reset_all;
    output n4667;
    input \fifo_data_out[15] ;
    input \fifo_data_out[14] ;
    input \fifo_data_out[13] ;
    input \fifo_data_out[12] ;
    input \fifo_data_out[11] ;
    input \fifo_data_out[10] ;
    input \fifo_data_out[9] ;
    input \fifo_data_out[8] ;
    input \fifo_data_out[7] ;
    input \fifo_data_out[4] ;
    input \fifo_data_out[3] ;
    input \fifo_data_out[2] ;
    input \fifo_data_out[1] ;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n1;
    wire [7:0]state_timeout_counter;   // src/bluejay_data.v(52[11:32])
    
    wire n10581, n1137, valid_N_707, n4062, n4442, n4, n4522, 
        n1_adj_1175, n4519, n1_adj_1176, n11177, n1_adj_1177;
    wire [8:0]n62;
    
    wire n7424, n10583, n21;
    wire [15:0]n703;
    
    wire n2779, n5836, n5835, n5834, n5833, n5832, n5831, n5830, 
        n5829, n5828, n5825, n5824, n5823, n5822, n10584, n10585, 
        n10587, n10586, bluejay_data_out_31__N_701, n770, n2777, n766, 
        bluejay_data_out_31__N_702, n2775, n2773, n3955, n3961;
    wire [10:0]v_counter_10__N_682;
    
    wire n4162;
    wire [10:0]v_counter;   // src/bluejay_data.v(51[12:21])
    
    wire n108, n10582, n86, n1_adj_1178, n10652, n10651, n10650, 
        n12, n10649, n10648, n10, n11418, n11330, n12_adj_1179, 
        n8, n10_adj_1180, n14, n10781, n10745, n6, n10647, n4618, 
        n10646, n10645, n10644, n10643;
    
    SB_LUT4 sub_116_add_2_3_lut (.I0(n1137), .I1(state_timeout_counter[1]), 
            .I2(VCC_net), .I3(n10581), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_DFFN valid_56 (.Q(VALID_c), .C(SLM_CLK_c), .D(valid_N_707));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFESS state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(SLM_CLK_c), 
            .E(n4062), .D(n1), .S(n4442));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(SLM_CLK_c), 
            .E(n4062), .D(n4), .S(n4522));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS state_timeout_counter_i0_i3 (.Q(\state_timeout_counter[3] ), 
            .C(SLM_CLK_c), .E(n4062), .D(n1_adj_1175), .S(n4519));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS state_timeout_counter_i0_i4 (.Q(state_timeout_counter[4]), .C(SLM_CLK_c), 
            .E(n4062), .D(n1_adj_1176), .S(n11177));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS state_timeout_counter_i0_i5 (.Q(state_timeout_counter[5]), .C(SLM_CLK_c), 
            .E(n4062), .D(n1_adj_1177), .S(n4519));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR state_timeout_counter_i0_i6 (.Q(state_timeout_counter[6]), .C(SLM_CLK_c), 
            .E(n4062), .D(n62[6]), .R(n7424));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR state_timeout_counter_i0_i7 (.Q(state_timeout_counter[7]), .C(SLM_CLK_c), 
            .E(n4062), .D(n62[7]), .R(n7424));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 sub_116_add_2_5_lut (.I0(n1137), .I1(\state_timeout_counter[3] ), 
            .I2(VCC_net), .I3(n10583), .O(n1_adj_1175)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i133_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n21), 
            .I2(bluejay_data_out_31__N_704), .I3(n703[9]), .O(n2779));   // src/bluejay_data.v(66[9] 121[16])
    defparam i133_3_lut_4_lut.LUT_INIT = 16'hf4f0;
    SB_DFFN bluejay_data_out_i1 (.Q(DATA16_c), .C(SLM_CLK_c), .D(n5870));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i16 (.Q(DATA15_c), .C(SLM_CLK_c), .D(n5836));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i15 (.Q(DATA14_c), .C(SLM_CLK_c), .D(n5835));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i14 (.Q(DATA13_c), .C(SLM_CLK_c), .D(n5834));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i13 (.Q(DATA12_c), .C(SLM_CLK_c), .D(n5833));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i12 (.Q(DATA11_c), .C(SLM_CLK_c), .D(n5832));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i11 (.Q(DATA10_c), .C(SLM_CLK_c), .D(n5831));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i10 (.Q(DATA9_c), .C(SLM_CLK_c), .D(n5830));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i9 (.Q(DATA8_c), .C(SLM_CLK_c), .D(n5829));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i8 (.Q(DATA7_c), .C(SLM_CLK_c), .D(n5828));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i7 (.Q(DATA6_c), .C(SLM_CLK_c), .D(n5827));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i6 (.Q(DATA5_c), .C(SLM_CLK_c), .D(n5826));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i5 (.Q(DATA20_c), .C(SLM_CLK_c), .D(n5825));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i4 (.Q(DATA19_c), .C(SLM_CLK_c), .D(n5824));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i3 (.Q(DATA18_c), .C(SLM_CLK_c), .D(n5823));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFN bluejay_data_out_i2 (.Q(DATA17_c), .C(SLM_CLK_c), .D(n5822));   // src/bluejay_data.v(126[8] 148[4])
    SB_CARRY sub_116_add_2_6 (.CI(n10584), .I0(state_timeout_counter[4]), 
            .I1(VCC_net), .CO(n10585));
    SB_LUT4 sub_116_add_2_9_lut (.I0(GND_net), .I1(state_timeout_counter[7]), 
            .I2(VCC_net), .I3(n10587), .O(n62[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_116_add_2_8_lut (.I0(GND_net), .I1(state_timeout_counter[6]), 
            .I2(VCC_net), .I3(n10586), .O(n62[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_116_add_2_8 (.CI(n10586), .I0(state_timeout_counter[6]), 
            .I1(VCC_net), .CO(n10587));
    SB_CARRY sub_116_add_2_7 (.CI(n10585), .I0(state_timeout_counter[5]), 
            .I1(VCC_net), .CO(n10586));
    SB_LUT4 sub_116_add_2_7_lut (.I0(n1137), .I1(state_timeout_counter[5]), 
            .I2(VCC_net), .I3(n10585), .O(n1_adj_1177)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_DFFN sync_58 (.Q(SYNC_c), .C(SLM_CLK_c), .D(bluejay_data_out_31__N_701));   // src/bluejay_data.v(126[8] 148[4])
    SB_DFFSR state_FSM_i10 (.Q(n703[9]), .C(SLM_CLK_c), .D(n2779), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i9 (.Q(bluejay_data_out_31__N_704), .C(SLM_CLK_c), 
            .D(n770), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i8 (.Q(bluejay_data_out_31__N_703), .C(SLM_CLK_c), 
            .D(n2777), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i7 (.Q(bluejay_data_out_31__N_702), .C(SLM_CLK_c), 
            .D(n766), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i6 (.Q(n703[5]), .C(SLM_CLK_c), .D(n2775), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i5 (.Q(n703[4]), .C(SLM_CLK_c), .D(n2773), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i4 (.Q(bluejay_data_out_31__N_701), .C(SLM_CLK_c), 
            .D(n14424), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i3 (.Q(n703[2]), .C(SLM_CLK_c), .D(n3955), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_DFFSR state_FSM_i2 (.Q(n718), .C(SLM_CLK_c), .D(n3961), .R(buffer_switch_done));   // src/bluejay_data.v(66[9] 121[16])
    SB_LUT4 i11075_2_lut (.I0(n4062), .I1(n1137), .I2(GND_net), .I3(GND_net), 
            .O(n7424));
    defparam i11075_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut (.I0(buffer_switch_done_latched), .I1(buffer_switch_done), 
            .I2(GND_net), .I3(GND_net), .O(n11177));   // src/bluejay_data.v(61[10] 122[8])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESR v_counter_i1 (.Q(v_counter[1]), .C(SLM_CLK_c), .E(n4162), 
            .D(v_counter_10__N_682[1]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 i1_2_lut_adj_58 (.I0(n4062), .I1(bluejay_data_out_31__N_704), 
            .I2(GND_net), .I3(GND_net), .O(n4522));   // src/bluejay_data.v(61[10] 122[8])
    defparam i1_2_lut_adj_58.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(n703[5]), .I1(n703[2]), .I2(bluejay_data_out_31__N_703), 
            .I3(GND_net), .O(n108));   // src/bluejay_data.v(66[9] 121[16])
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3240_2_lut (.I0(n4062), .I1(bluejay_data_out_31__N_701), .I2(GND_net), 
            .I3(GND_net), .O(n4442));   // src/bluejay_data.v(56[8] 123[4])
    defparam i3240_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11119_3_lut (.I0(buffer_switch_done_latched), .I1(buffer_switch_done), 
            .I2(n108), .I3(GND_net), .O(n4062));   // src/bluejay_data.v(61[10] 122[8])
    defparam i11119_3_lut.LUT_INIT = 16'h2323;
    SB_CARRY sub_116_add_2_5 (.CI(n10583), .I0(\state_timeout_counter[3] ), 
            .I1(VCC_net), .CO(n10584));
    SB_LUT4 sub_116_add_2_6_lut (.I0(n1137), .I1(state_timeout_counter[4]), 
            .I2(VCC_net), .I3(n10584), .O(n1_adj_1176)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_116_add_2_3 (.CI(n10581), .I0(state_timeout_counter[1]), 
            .I1(VCC_net), .CO(n10582));
    SB_LUT4 sub_116_add_2_4_lut (.I0(n1137), .I1(state_timeout_counter[2]), 
            .I2(VCC_net), .I3(n10582), .O(n86)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_116_add_2_2_lut (.I0(n1137), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(VCC_net), .O(n1_adj_1178)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_116_add_2_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_116_add_2_2 (.CI(VCC_net), .I0(state_timeout_counter[0]), 
            .I1(GND_net), .CO(n10581));
    SB_LUT4 sub_118_add_2_12_lut (.I0(GND_net), .I1(v_counter[10]), .I2(VCC_net), 
            .I3(n10652), .O(v_counter_10__N_682[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_118_add_2_11_lut (.I0(GND_net), .I1(v_counter[9]), .I2(VCC_net), 
            .I3(n10651), .O(v_counter_10__N_682[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_11 (.CI(n10651), .I0(v_counter[9]), .I1(VCC_net), 
            .CO(n10652));
    SB_LUT4 sub_118_add_2_10_lut (.I0(GND_net), .I1(v_counter[8]), .I2(VCC_net), 
            .I3(n10650), .O(v_counter_10__N_682[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_10 (.CI(n10650), .I0(v_counter[8]), .I1(VCC_net), 
            .CO(n10651));
    SB_LUT4 i1_2_lut_3_lut (.I0(n12), .I1(state_timeout_counter[0]), .I2(state_timeout_counter[4]), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_DFFESR v_counter_i2 (.Q(v_counter[2]), .C(SLM_CLK_c), .E(n4162), 
            .D(v_counter_10__N_682[2]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 sub_118_add_2_9_lut (.I0(GND_net), .I1(v_counter[7]), .I2(VCC_net), 
            .I3(n10649), .O(v_counter_10__N_682[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_9 (.CI(n10649), .I0(v_counter[7]), .I1(VCC_net), 
            .CO(n10650));
    SB_LUT4 sub_118_add_2_8_lut (.I0(GND_net), .I1(v_counter[6]), .I2(VCC_net), 
            .I3(n10648), .O(v_counter_10__N_682[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_59 (.I0(n703[9]), .I1(buffer_switch_done), .I2(GND_net), 
            .I3(GND_net), .O(n4162));
    defparam i1_2_lut_adj_59.LUT_INIT = 16'heeee;
    SB_CARRY sub_118_add_2_8 (.CI(n10648), .I0(v_counter[6]), .I1(VCC_net), 
            .CO(n10649));
    SB_DFFESS v_counter_i3 (.Q(v_counter[3]), .C(SLM_CLK_c), .E(n4162), 
            .D(v_counter_10__N_682[3]), .S(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 i1_4_lut (.I0(n5), .I1(\rd_sig_diff0_w[0] ), .I2(\rd_sig_diff0_w[1] ), 
            .I3(get_next_word), .O(\aempty_flag_impl.ae_flag_nxt_w ));   // src/fifo_dc_32_lut_gen.v(233[30:44])
    defparam i1_4_lut.LUT_INIT = 16'h1505;
    SB_DFFESR v_counter_i4 (.Q(v_counter[4]), .C(SLM_CLK_c), .E(n4162), 
            .D(v_counter_10__N_682[4]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESS v_counter_i5 (.Q(v_counter[5]), .C(SLM_CLK_c), .E(n4162), 
            .D(v_counter_10__N_682[5]), .S(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i6 (.Q(v_counter[6]), .C(SLM_CLK_c), .E(n4162), 
            .D(v_counter_10__N_682[6]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i7 (.Q(v_counter[7]), .C(SLM_CLK_c), .E(n4162), 
            .D(v_counter_10__N_682[7]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i8 (.Q(v_counter[8]), .C(SLM_CLK_c), .E(n4162), 
            .D(v_counter_10__N_682[8]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i9 (.Q(v_counter[9]), .C(SLM_CLK_c), .E(n4162), 
            .D(v_counter_10__N_682[9]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_DFFESR v_counter_i10 (.Q(v_counter[10]), .C(SLM_CLK_c), .E(n4162), 
            .D(v_counter_10__N_682[10]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 i9770_2_lut (.I0(n10), .I1(v_counter[6]), .I2(GND_net), .I3(GND_net), 
            .O(n11418));
    defparam i9770_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_60 (.I0(n703[9]), .I1(v_counter[5]), .I2(n11418), 
            .I3(v_counter[3]), .O(n11330));   // src/top.v(122[12:19])
    defparam i1_4_lut_adj_60.LUT_INIT = 16'h0002;
    SB_LUT4 i1_4_lut_adj_61 (.I0(\state_timeout_counter[3] ), .I1(n718), 
            .I2(n11330), .I3(DEBUG_9_c), .O(n12_adj_1179));   // src/top.v(122[12:19])
    defparam i1_4_lut_adj_61.LUT_INIT = 16'h5054;
    SB_LUT4 i1_4_lut_adj_62 (.I0(n703[2]), .I1(n8), .I2(n12_adj_1179), 
            .I3(n12), .O(n3955));   // src/top.v(122[12:19])
    defparam i1_4_lut_adj_62.LUT_INIT = 16'haaba;
    SB_LUT4 i2_2_lut (.I0(v_counter[4]), .I1(v_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_1180));   // src/bluejay_data.v(56[8] 123[4])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(v_counter[1]), .I1(v_counter[7]), .I2(v_counter[10]), 
            .I3(v_counter[9]), .O(n14));   // src/bluejay_data.v(56[8] 123[4])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(v_counter[8]), .I1(n14), .I2(n10_adj_1180), 
            .I3(v_counter[0]), .O(n10));   // src/bluejay_data.v(56[8] 123[4])
    defparam i7_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i3_4_lut (.I0(n10), .I1(v_counter[6]), .I2(v_counter[5]), 
            .I3(v_counter[3]), .O(n10781));   // src/bluejay_data.v(56[8] 123[4])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1591_4_lut (.I0(buffer_switch_done_latched), .I1(n10745), .I2(n703[5]), 
            .I3(DEBUG_9_c), .O(n2775));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1591_4_lut.LUT_INIT = 16'hccdc;
    SB_LUT4 i135_4_lut (.I0(DEBUG_9_c), .I1(n703[4]), .I2(n703[5]), .I3(n21), 
            .O(n766));   // src/top.v(122[12:19])
    defparam i135_4_lut.LUT_INIT = 16'ha0ec;
    SB_LUT4 i1_4_lut_adj_63 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_702), 
            .I2(dc32_fifo_almost_empty), .I3(buffer_switch_done_latched), 
            .O(n2777));   // src/bluejay_data.v(62[9] 65[12])
    defparam i1_4_lut_adj_63.LUT_INIT = 16'hccce;
    SB_LUT4 i1_2_lut_adj_64 (.I0(bluejay_data_out_31__N_703), .I1(dc32_fifo_almost_empty), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_2_lut_adj_64.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_65 (.I0(state_timeout_counter[0]), .I1(state_timeout_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // src/bluejay_data.v(56[8] 123[4])
    defparam i1_2_lut_adj_65.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_66 (.I0(state_timeout_counter[5]), .I1(state_timeout_counter[6]), 
            .I2(GND_net), .I3(GND_net), .O(n6));
    defparam i1_2_lut_adj_66.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(state_timeout_counter[2]), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[7]), .I3(n6), .O(n12));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_118_add_2_7_lut (.I0(GND_net), .I1(v_counter[5]), .I2(VCC_net), 
            .I3(n10647), .O(v_counter_10__N_682[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_7 (.CI(n10647), .I0(v_counter[5]), .I1(VCC_net), 
            .CO(n10648));
    SB_LUT4 i1_2_lut_adj_67 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(GND_net), .I3(GND_net), .O(valid_N_707));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_2_lut_adj_67.LUT_INIT = 16'heeee;
    SB_DFFN get_next_word_57 (.Q(get_next_word), .C(SLM_CLK_c), .D(n4618));   // src/bluejay_data.v(126[8] 148[4])
    SB_LUT4 i2_3_lut_adj_68 (.I0(n703[4]), .I1(n718), .I2(n703[9]), .I3(GND_net), 
            .O(n1137));   // src/bluejay_data.v(66[9] 121[16])
    defparam i2_3_lut_adj_68.LUT_INIT = 16'hfefe;
    SB_DFFESR v_counter_i0 (.Q(v_counter[0]), .C(SLM_CLK_c), .E(n4162), 
            .D(v_counter_10__N_682[0]), .R(buffer_switch_done));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 sub_118_add_2_6_lut (.I0(GND_net), .I1(v_counter[4]), .I2(VCC_net), 
            .I3(n10646), .O(v_counter_10__N_682[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1589_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n21), 
            .I2(bluejay_data_out_31__N_701), .I3(n703[4]), .O(n2773));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1589_3_lut_4_lut.LUT_INIT = 16'hf4f0;
    SB_CARRY sub_118_add_2_6 (.CI(n10646), .I0(v_counter[4]), .I1(VCC_net), 
            .CO(n10647));
    SB_LUT4 sub_118_add_2_5_lut (.I0(GND_net), .I1(v_counter[3]), .I2(VCC_net), 
            .I3(n10645), .O(v_counter_10__N_682[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut (.I0(buffer_switch_done_latched), .I1(n108), 
            .I2(bluejay_data_out_31__N_702), .I3(n4062), .O(n4519));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_69 (.I0(buffer_switch_done_latched), .I1(n108), 
            .I2(n86), .I3(GND_net), .O(n4));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_2_lut_3_lut_adj_69.LUT_INIT = 16'hfefe;
    SB_CARRY sub_118_add_2_5 (.CI(n10645), .I0(v_counter[3]), .I1(VCC_net), 
            .CO(n10646));
    SB_LUT4 sub_118_add_2_4_lut (.I0(GND_net), .I1(v_counter[2]), .I2(VCC_net), 
            .I3(n10644), .O(v_counter_10__N_682[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_4 (.CI(n10644), .I0(v_counter[2]), .I1(VCC_net), 
            .CO(n10645));
    SB_DFFESS state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(SLM_CLK_c), 
            .E(n4062), .D(n1_adj_1178), .S(n4442));   // src/bluejay_data.v(56[8] 123[4])
    SB_LUT4 sub_118_add_2_3_lut (.I0(GND_net), .I1(v_counter[1]), .I2(VCC_net), 
            .I3(n10643), .O(v_counter_10__N_682[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_3 (.CI(n10643), .I0(v_counter[1]), .I1(VCC_net), 
            .CO(n10644));
    SB_CARRY sub_116_add_2_4 (.CI(n10582), .I0(state_timeout_counter[2]), 
            .I1(VCC_net), .CO(n10583));
    SB_LUT4 sub_118_add_2_2_lut (.I0(GND_net), .I1(v_counter[0]), .I2(n21), 
            .I3(VCC_net), .O(v_counter_10__N_682[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_118_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_118_add_2_2 (.CI(VCC_net), .I0(v_counter[0]), .I1(n21), 
            .CO(n10643));
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\state_timeout_counter[3] ), .I1(n12), 
            .I2(state_timeout_counter[0]), .I3(state_timeout_counter[4]), 
            .O(n21));   // src/bluejay_data.v(56[8] 123[4])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state_timeout_counter[3] ), .I1(n7), .I2(n10781), 
            .I3(n703[9]), .O(n10745));   // src/bluejay_data.v(66[9] 121[16])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_3_lut_4_lut_adj_70 (.I0(buffer_switch_done_latched), .I1(\state_timeout_counter[3] ), 
            .I2(n7), .I3(n718), .O(n3961));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_3_lut_4_lut_adj_70.LUT_INIT = 16'hfeaa;
    SB_LUT4 i1_2_lut_adj_71 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_702), 
            .I2(GND_net), .I3(GND_net), .O(n4618));   // src/bluejay_data.v(66[9] 121[16])
    defparam i1_2_lut_adj_71.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_72 (.I0(DEBUG_5_c), .I1(get_next_word), .I2(reset_all), 
            .I3(GND_net), .O(n4667));
    defparam i1_2_lut_3_lut_adj_72.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_3_lut_adj_73 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[15] ), .I3(GND_net), .O(n5836));
    defparam i1_2_lut_3_lut_adj_73.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_74 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[14] ), .I3(GND_net), .O(n5835));
    defparam i1_2_lut_3_lut_adj_74.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_75 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[13] ), .I3(GND_net), .O(n5834));
    defparam i1_2_lut_3_lut_adj_75.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_76 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[12] ), .I3(GND_net), .O(n5833));
    defparam i1_2_lut_3_lut_adj_76.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_77 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[11] ), .I3(GND_net), .O(n5832));
    defparam i1_2_lut_3_lut_adj_77.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_78 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[10] ), .I3(GND_net), .O(n5831));
    defparam i1_2_lut_3_lut_adj_78.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_79 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[9] ), .I3(GND_net), .O(n5830));
    defparam i1_2_lut_3_lut_adj_79.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_80 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[8] ), .I3(GND_net), .O(n5829));
    defparam i1_2_lut_3_lut_adj_80.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_81 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[7] ), .I3(GND_net), .O(n5828));
    defparam i1_2_lut_3_lut_adj_81.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_82 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[4] ), .I3(GND_net), .O(n5825));
    defparam i1_2_lut_3_lut_adj_82.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_83 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[3] ), .I3(GND_net), .O(n5824));
    defparam i1_2_lut_3_lut_adj_83.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_84 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[2] ), .I3(GND_net), .O(n5823));
    defparam i1_2_lut_3_lut_adj_84.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_85 (.I0(bluejay_data_out_31__N_703), .I1(bluejay_data_out_31__N_704), 
            .I2(\fifo_data_out[1] ), .I3(GND_net), .O(n5822));
    defparam i1_2_lut_3_lut_adj_85.LUT_INIT = 16'he0e0;
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen2
//

module fifo_dc_32_lut_gen2 (\REG.mem_58_4 , GND_net, \REG.mem_14_8 , \REG.mem_15_8 , 
            \dc32_fifo_data_in[10] , \dc32_fifo_data_in[9] , DEBUG_6_c_c, 
            \REG.mem_13_8 , \REG.mem_12_8 , \dc32_fifo_data_in[8] , \REG.mem_10_10 , 
            \REG.mem_11_10 , \REG.mem_9_10 , \REG.mem_8_10 , t_rd_fifo_en_w, 
            \REG.out_raw[0] , SLM_CLK_c, \dc32_fifo_data_in[7] , \REG.mem_10_13 , 
            \REG.mem_11_13 , \REG.mem_9_13 , \REG.mem_8_13 , \dc32_fifo_data_in[6] , 
            DEBUG_9_c, n7596, \wr_addr_nxt_c[4] , \REG.mem_26_14 , \dc32_fifo_data_in[5] , 
            \REG.mem_42_2 , \REG.mem_43_2 , \REG.mem_41_2 , \REG.mem_40_2 , 
            \REG.mem_14_10 , \REG.mem_15_10 , reset_all, \REG.mem_55_8 , 
            \REG.mem_13_10 , \REG.mem_12_10 , \dc32_fifo_data_in[4] , 
            \REG.mem_42_3 , \REG.mem_43_3 , \REG.mem_41_3 , \REG.mem_40_3 , 
            \rd_grey_sync_r[0] , \dc32_fifo_data_in[3] , \REG.mem_58_8 , 
            DEBUG_5_c, wr_grey_sync_r, \REG.mem_48_5 , \REG.mem_49_5 , 
            \aempty_flag_impl.ae_flag_nxt_w , dc32_fifo_almost_empty, \dc32_fifo_data_in[2] , 
            \REG.mem_55_11 , \REG.mem_50_5 , \REG.mem_51_5 , \dc32_fifo_data_in[1] , 
            \REG.mem_55_5 , \REG.mem_63_4 , \REG.mem_23_11 , \dc32_fifo_data_in[0] , 
            \REG.mem_10_12 , \REG.mem_11_12 , \REG.mem_9_12 , \REG.mem_8_12 , 
            \REG.mem_38_11 , \REG.mem_39_11 , \REG.mem_37_11 , \REG.mem_36_11 , 
            \REG.mem_14_12 , \REG.mem_15_12 , \REG.mem_14_13 , \REG.mem_15_13 , 
            \REG.mem_6_12 , \REG.mem_7_12 , \REG.mem_4_12 , \REG.mem_5_12 , 
            \REG.mem_13_13 , \REG.mem_12_13 , \REG.mem_13_12 , \REG.mem_12_12 , 
            \REG.mem_23_15 , \REG.mem_18_12 , \REG.mem_19_12 , \REG.mem_6_8 , 
            \REG.mem_7_8 , \REG.mem_17_12 , \REG.mem_16_12 , \wr_addr_nxt_c[2] , 
            \REG.mem_26_0 , \REG.mem_42_10 , \REG.mem_43_10 , \REG.mem_18_8 , 
            \REG.mem_19_8 , \REG.mem_14_15 , \REG.mem_15_15 , \REG.mem_17_8 , 
            \REG.mem_16_8 , \REG.mem_41_10 , \REG.mem_40_10 , n60, \REG.mem_18_13 , 
            \REG.mem_19_13 , \REG.mem_17_13 , \REG.mem_16_13 , n28, 
            \REG.mem_13_15 , \REG.mem_12_15 , \REG.mem_26_3 , \REG.mem_46_6 , 
            \REG.mem_47_6 , \REG.mem_45_6 , \REG.mem_44_6 , \REG.mem_63_8 , 
            \REG.mem_46_2 , \REG.mem_47_2 , \REG.mem_45_2 , \REG.mem_44_2 , 
            \dc32_fifo_data_in[15] , \dc32_fifo_data_in[14] , \REG.mem_6_7 , 
            \REG.mem_7_7 , \dc32_fifo_data_in[13] , \REG.mem_46_11 , \REG.mem_47_11 , 
            \dc32_fifo_data_in[12] , \REG.mem_5_7 , \REG.mem_4_7 , \dc32_fifo_data_in[11] , 
            \REG.mem_45_11 , \REG.mem_44_11 , \REG.mem_23_13 , \REG.mem_58_5 , 
            \REG.mem_23_8 , \REG.mem_46_3 , \REG.mem_47_3 , \REG.mem_10_7 , 
            \REG.mem_11_7 , \REG.mem_45_3 , \REG.mem_44_3 , \REG.mem_8_2 , 
            \REG.mem_9_2 , \REG.mem_9_7 , \REG.mem_8_7 , \REG.mem_31_14 , 
            \REG.mem_10_2 , \REG.mem_11_2 , \REG.mem_58_13 , \REG.mem_26_8 , 
            \REG.mem_14_2 , \REG.mem_15_2 , \REG.mem_12_2 , \REG.mem_13_2 , 
            \REG.mem_14_7 , \REG.mem_15_7 , \REG.mem_13_7 , \REG.mem_12_7 , 
            \REG.mem_26_13 , \REG.mem_6_3 , \REG.mem_7_3 , \REG.mem_5_3 , 
            \REG.mem_4_3 , \REG.mem_40_1 , \REG.mem_41_1 , \REG.mem_14_5 , 
            \REG.mem_15_5 , \REG.mem_13_5 , \REG.mem_12_5 , \REG.mem_42_1 , 
            \REG.mem_43_1 , \REG.mem_46_1 , \REG.mem_47_1 , \REG.mem_44_1 , 
            \REG.mem_45_1 , \REG.mem_31_8 , \REG.mem_26_10 , \REG.mem_18_2 , 
            \REG.mem_19_2 , \REG.mem_31_3 , \REG.mem_17_2 , \REG.mem_16_2 , 
            n61, \REG.mem_63_13 , n34, n29, \REG.mem_50_6 , \REG.mem_51_6 , 
            n58, \REG.mem_6_14 , \REG.mem_7_14 , n26, \REG.mem_6_10 , 
            \REG.mem_7_10 , \REG.mem_4_10 , \REG.mem_5_10 , \REG.mem_4_14 , 
            \REG.mem_5_14 , n5896, VCC_net, \fifo_data_out[6] , n5893, 
            \fifo_data_out[5] , \REG.mem_16_10 , \REG.mem_17_10 , \REG.mem_18_10 , 
            \REG.mem_19_10 , n11119, \fifo_data_out[7] , \REG.mem_18_7 , 
            \REG.mem_19_7 , n11139, \fifo_data_out[3] , \REG.mem_17_7 , 
            \REG.mem_16_7 , \REG.mem_50_2 , \REG.mem_51_2 , \REG.mem_46_0 , 
            \REG.mem_47_0 , \REG.mem_46_9 , \REG.mem_47_9 , \REG.mem_45_9 , 
            \REG.mem_44_9 , \REG.mem_49_6 , \REG.mem_48_6 , \REG.mem_49_2 , 
            \REG.mem_48_2 , n11097, \fifo_data_out[8] , n5854, \fifo_data_out[0] , 
            \REG.mem_5_8 , \REG.mem_4_8 , \REG.mem_6_11 , \REG.mem_7_11 , 
            \REG.mem_58_1 , \REG.mem_26_15 , n11095, \fifo_data_out[9] , 
            \REG.mem_23_7 , n11143, \fifo_data_out[1] , n11141, \fifo_data_out[2] , 
            n11089, \fifo_data_out[10] , n11135, \fifo_data_out[11] , 
            \REG.mem_50_3 , \REG.mem_51_3 , \REG.mem_31_13 , \REG.mem_49_3 , 
            \REG.mem_48_3 , \REG.mem_10_9 , \REG.mem_11_9 , \REG.mem_9_9 , 
            \REG.mem_8_9 , \REG.mem_23_10 , \REG.mem_26_1 , n47, n5789, 
            \REG.mem_63_15 , n5788, \REG.mem_63_14 , n5787, \REG.mem_31_11 , 
            \REG.mem_5_11 , \REG.mem_4_11 , \REG.mem_31_1 , \REG.mem_23_12 , 
            n5786, \REG.mem_63_12 , n5785, \REG.mem_63_11 , n5784, 
            \REG.mem_63_10 , n5783, \REG.mem_63_9 , \REG.mem_14_9 , 
            \REG.mem_15_9 , n5782, n5781, \REG.mem_63_7 , n5780, \REG.mem_63_6 , 
            n5779, \REG.mem_63_5 , n5778, n5777, \REG.mem_63_3 , n5776, 
            \REG.mem_63_2 , n5775, \REG.mem_63_1 , n11133, \fifo_data_out[12] , 
            n5773, \REG.mem_63_0 , \REG.mem_13_9 , \REG.mem_12_9 , \REG.mem_38_10 , 
            \REG.mem_39_10 , n15, \REG.mem_36_10 , \REG.mem_37_10 , 
            \REG.mem_8_1 , \REG.mem_9_1 , \REG.mem_10_1 , \REG.mem_11_1 , 
            n11137, \fifo_data_out[4] , \REG.mem_14_1 , \REG.mem_15_1 , 
            \REG.mem_12_1 , \REG.mem_13_1 , \REG.mem_38_12 , \REG.mem_39_12 , 
            \REG.mem_36_12 , \REG.mem_37_12 , \REG.mem_38_5 , \REG.mem_39_5 , 
            n5709, rp_sync1_r, n5708, n5707, n5706, n5705, \REG.mem_36_5 , 
            \REG.mem_37_5 , \REG.mem_48_12 , \REG.mem_49_12 , \wr_addr_r[0] , 
            \REG.mem_50_12 , \REG.mem_51_12 , \REG.mem_55_12 , \wr_addr_p1_w[6] , 
            n5704, \rd_sig_diff0_w[1] , n5686, n5685, n5684, n5683, 
            n5682, \REG.mem_58_15 , n5681, \REG.mem_58_14 , n5680, 
            n5679, \REG.mem_58_12 , n5678, \REG.mem_58_11 , n5677, 
            \REG.mem_58_10 , n5676, \REG.mem_58_9 , n5675, n5674, 
            \REG.mem_58_7 , n5673, \REG.mem_58_6 , \REG.mem_26_7 , \rd_sig_diff0_w[0] , 
            n5672, n5671, n5670, \REG.mem_58_3 , n5669, \REG.mem_58_2 , 
            n5668, n5667, \REG.mem_58_0 , n5666, n5665, n5664, n5662, 
            n5660, \rd_addr_r[6] , \REG.out_raw[15] , \REG.out_raw[14] , 
            \REG.out_raw[13] , \REG.out_raw[12] , \REG.out_raw[11] , \REG.out_raw[10] , 
            \REG.out_raw[9] , \REG.out_raw[8] , \REG.out_raw[7] , \REG.out_raw[6] , 
            \REG.out_raw[5] , \REG.out_raw[4] , \REG.out_raw[3] , \REG.out_raw[2] , 
            \REG.out_raw[1] , \REG.mem_31_7 , \REG.mem_42_11 , \REG.mem_43_11 , 
            \REG.mem_41_11 , \REG.mem_40_11 , n2, \REG.mem_6_1 , \REG.mem_7_1 , 
            \REG.mem_4_1 , \REG.mem_5_1 , \REG.mem_38_4 , \REG.mem_39_4 , 
            \REG.mem_16_1 , \REG.mem_17_1 , \REG.mem_37_4 , \REG.mem_36_4 , 
            \REG.mem_55_2 , \REG.mem_18_1 , \REG.mem_19_1 , n5626, \REG.mem_55_15 , 
            \REG.mem_23_1 , \REG.mem_31_10 , n5625, \REG.mem_55_14 , 
            n5624, \REG.mem_55_13 , n5623, n5622, n5621, \REG.mem_55_10 , 
            n5620, \REG.mem_55_9 , n5619, n5618, \REG.mem_55_7 , n5617, 
            \REG.mem_55_6 , n5616, n5615, \REG.mem_55_4 , n5614, \REG.mem_55_3 , 
            n5613, n5612, \REG.mem_55_1 , n11073, \fifo_data_out[13] , 
            n5610, \REG.mem_55_0 , n5609, wp_sync1_r, n5608, n5607, 
            n5606, n5605, n5604, n5603, n5586, n5585, n5584, n5583, 
            n5582, n11071, \fifo_data_out[14] , \REG.mem_38_1 , \REG.mem_39_1 , 
            \REG.mem_36_1 , \REG.mem_37_1 , \REG.mem_6_2 , \REG.mem_7_2 , 
            \REG.mem_5_2 , \REG.mem_4_2 , n5548, \REG.mem_51_15 , n5547, 
            \REG.mem_51_14 , n5546, \REG.mem_51_13 , n5545, n5544, 
            \REG.mem_51_11 , n5543, \REG.mem_51_10 , n5542, \REG.mem_51_9 , 
            n5541, \REG.mem_51_8 , n5540, \REG.mem_51_7 , n5539, n5538, 
            n5537, \REG.mem_51_4 , n5536, n5535, n5534, \REG.mem_51_1 , 
            n5533, \REG.mem_51_0 , n5532, \REG.mem_50_15 , \REG.mem_48_1 , 
            \REG.mem_49_1 , n5531, \REG.mem_50_14 , n5530, \REG.mem_50_13 , 
            n5529, n5528, \REG.mem_50_11 , n5527, \REG.mem_50_10 , 
            n5526, \REG.mem_50_9 , n5525, \REG.mem_50_8 , n5524, \REG.mem_50_7 , 
            n5523, n5522, n5521, \REG.mem_50_4 , n5520, n5519, n5518, 
            \REG.mem_50_1 , n5517, \REG.mem_50_0 , n5516, \REG.mem_49_15 , 
            n5515, \REG.mem_49_14 , \REG.mem_31_12 , \REG.mem_26_11 , 
            n5514, \REG.mem_49_13 , n5513, n5512, \REG.mem_49_11 , 
            n5511, \REG.mem_49_10 , n5510, \REG.mem_49_9 , n5509, 
            \REG.mem_49_8 , n5508, \REG.mem_49_7 , n5507, n5506, n5505, 
            \REG.mem_49_4 , n5504, n5503, n5502, n5501, \REG.mem_49_0 , 
            \REG.mem_31_0 , \REG.mem_26_4 , n5492, \REG.mem_48_15 , 
            n5491, n5490, \REG.mem_48_14 , n5489, \REG.mem_48_13 , 
            n5488, n5487, \REG.mem_48_11 , n5486, \REG.mem_48_10 , 
            n5485, \REG.mem_48_9 , n5484, \REG.mem_48_8 , n5483, \REG.mem_48_7 , 
            \REG.mem_46_10 , \REG.mem_47_10 , n5482, n5481, n5480, 
            \REG.mem_48_4 , n5479, n5478, n5477, n5476, \REG.mem_48_0 , 
            n5474, n5472, \REG.mem_47_15 , n5471, \REG.mem_47_14 , 
            n5470, \REG.mem_47_13 , n5469, \REG.mem_47_12 , n5468, 
            n5467, \REG.mem_45_0 , \REG.mem_44_0 , \REG.mem_45_10 , 
            \REG.mem_44_10 , n5466, n5465, \REG.mem_47_8 , n5464, 
            \REG.mem_47_7 , n5463, n5462, \REG.mem_47_5 , n5461, \REG.mem_47_4 , 
            n5460, n5459, n5458, n5457, n5456, \REG.mem_46_15 , 
            n5455, \REG.mem_46_14 , n5454, \REG.mem_46_13 , n5453, 
            \REG.mem_46_12 , n5452, n5451, n5450, n5449, \REG.mem_46_8 , 
            n5448, \REG.mem_46_7 , n5447, n5446, \REG.mem_46_5 , n5445, 
            \REG.mem_46_4 , n5444, n5443, n5442, n5441, n5440, \REG.mem_45_15 , 
            n5439, \REG.mem_45_14 , n5438, \REG.mem_45_13 , n5437, 
            \REG.mem_45_12 , n5436, n5435, n5434, \REG.mem_38_7 , 
            \REG.mem_39_7 , \REG.mem_37_7 , \REG.mem_36_7 , n5433, \REG.mem_45_8 , 
            n5432, \REG.mem_45_7 , n5431, n5430, \REG.mem_45_5 , n5429, 
            \REG.mem_45_4 , n5428, n5427, n5426, n5425, n5424, \REG.mem_44_15 , 
            n5423, \REG.mem_44_14 , n5422, \REG.mem_44_13 , n5421, 
            \REG.mem_44_12 , n5420, n5419, \REG.mem_10_0 , \REG.mem_11_0 , 
            n5418, \REG.mem_9_0 , \REG.mem_8_0 , n5417, \REG.mem_44_8 , 
            n5416, \REG.mem_44_7 , n5415, n5414, \REG.mem_44_5 , n5413, 
            \REG.mem_44_4 , n5412, n5411, n5410, n5409, n5408, n5407, 
            \REG.mem_43_15 , n5406, \REG.mem_43_14 , n5405, \REG.mem_43_13 , 
            n5404, \REG.mem_43_12 , n5403, n5402, \REG.mem_10_5 , 
            \REG.mem_11_5 , \REG.mem_9_5 , \REG.mem_8_5 , \wr_addr_p1_w[0] , 
            n5401, \REG.mem_43_9 , n5400, \REG.mem_43_8 , n5399, \REG.mem_43_7 , 
            n5398, \REG.mem_43_6 , n5397, \REG.mem_43_5 , n5396, \REG.mem_43_4 , 
            n5395, n5394, n5393, n5392, \REG.mem_43_0 , n11069, 
            \fifo_data_out[15] , n5390, \REG.mem_42_15 , n5389, \REG.mem_42_14 , 
            n5388, \REG.mem_42_13 , n5387, \REG.mem_42_12 , n5386, 
            \REG.mem_42_4 , \REG.mem_41_4 , \REG.mem_40_4 , n5385, n5384, 
            \REG.mem_42_9 , n5383, \REG.mem_42_8 , n5382, \REG.mem_42_7 , 
            n5381, \REG.mem_42_6 , n5380, \REG.mem_42_5 , n5379, n5378, 
            n5377, n5376, n5375, \REG.mem_42_0 , n5374, \REG.mem_41_15 , 
            n5373, \REG.mem_41_14 , n5372, \REG.mem_41_13 , n5371, 
            \REG.mem_41_12 , n4667, n5370, n5369, n5368, \REG.mem_41_9 , 
            n5367, \REG.mem_41_8 , n5366, \REG.mem_41_7 , n5365, \REG.mem_41_6 , 
            n5364, \REG.mem_41_5 , n5363, n5362, n5361, n5360, n5358, 
            \REG.mem_41_0 , n5357, \REG.mem_40_15 , n5356, \REG.mem_40_14 , 
            n5355, \REG.mem_40_13 , n5354, \REG.mem_40_12 , \REG.mem_38_13 , 
            \REG.mem_39_13 , \REG.mem_37_13 , \REG.mem_36_13 , n5353, 
            n5352, n5351, \REG.mem_40_9 , n5350, \REG.mem_40_8 , n5349, 
            \REG.mem_40_7 , n5348, \REG.mem_40_6 , n5347, \REG.mem_40_5 , 
            n5346, n5345, n5344, n5343, n5342, \REG.mem_40_0 , n5341, 
            \REG.mem_39_15 , n5340, \REG.mem_39_14 , n5339, \REG.mem_23_5 , 
            \REG.mem_14_0 , \REG.mem_15_0 , \REG.mem_13_0 , \REG.mem_12_0 , 
            n5338, n5337, n5336, n5335, \REG.mem_39_9 , n5334, \REG.mem_39_8 , 
            n5333, n5332, \REG.mem_39_6 , n5331, n5330, n5329, \REG.mem_39_3 , 
            n5328, \REG.mem_39_2 , n5327, n5326, \REG.mem_39_0 , n5323, 
            \REG.mem_38_15 , n5322, \REG.mem_38_14 , n5321, n5320, 
            n5319, n5318, n5317, \REG.mem_38_9 , n5316, \REG.mem_38_8 , 
            n5315, n5314, \REG.mem_38_6 , n5313, n5312, n5311, \REG.mem_38_3 , 
            n5310, \REG.mem_38_2 , n5309, n5308, \REG.mem_38_0 , n5302, 
            \REG.mem_37_15 , n5301, \REG.mem_37_14 , n5300, n5299, 
            n5298, n5297, n5296, \REG.mem_37_9 , n5295, \REG.mem_37_8 , 
            n5294, n5293, \REG.mem_37_6 , n5292, n5291, n5290, \REG.mem_37_3 , 
            n5289, \REG.mem_37_2 , n5288, n5286, \REG.mem_37_0 , n5285, 
            \REG.mem_36_15 , n5284, \REG.mem_36_14 , n5283, n5282, 
            n5281, n5280, n5279, \REG.mem_36_9 , n5278, \REG.mem_36_8 , 
            n5277, n5276, \REG.mem_36_6 , n5275, n5274, n5273, \REG.mem_36_3 , 
            n5272, \REG.mem_36_2 , n5271, n5270, \REG.mem_36_0 , \REG.mem_26_12 , 
            \REG.mem_10_3 , \REG.mem_11_3 , n5202, \REG.mem_31_15 , 
            n5201, n5200, n5199, n5198, n5197, n5196, \REG.mem_31_9 , 
            n5195, n5194, n5193, \REG.mem_31_6 , n5192, \REG.mem_31_5 , 
            n5191, \REG.mem_31_4 , n5190, n5189, \REG.mem_31_2 , \REG.mem_9_3 , 
            \REG.mem_8_3 , n5188, n5187, \REG.mem_10_14 , \REG.mem_11_14 , 
            \REG.mem_9_14 , \REG.mem_8_14 , \REG.mem_23_2 , n5121, n5120, 
            n5119, n5118, n5117, n5116, n5115, \REG.mem_26_9 , n5114, 
            n5113, n5112, \REG.mem_26_6 , n5111, \REG.mem_26_5 , n5110, 
            n5109, n5108, \REG.mem_26_2 , n5107, n5106, n5073, n5072, 
            \REG.mem_23_14 , n5071, n5070, n5069, n5068, n5067, 
            \REG.mem_23_9 , n5066, \rd_grey_sync_r[5] , \rd_grey_sync_r[4] , 
            \REG.mem_10_6 , \REG.mem_11_6 , \rd_grey_sync_r[3] , \rd_grey_sync_r[2] , 
            \rd_grey_sync_r[1] , n5065, n5064, \REG.mem_23_6 , n5063, 
            n5062, \REG.mem_23_4 , n5061, \REG.mem_23_3 , n5060, n5059, 
            n5058, \REG.mem_23_0 , \REG.mem_9_6 , \REG.mem_8_6 , n5, 
            \REG.mem_14_6 , \REG.mem_15_6 , \REG.mem_13_6 , \REG.mem_12_6 , 
            n5006, \REG.mem_19_15 , n5005, \REG.mem_19_14 , n5004, 
            n5003, n5002, \REG.mem_19_11 , n5001, n5000, \REG.mem_19_9 , 
            n4999, n4998, n4997, \REG.mem_19_6 , n4996, \REG.mem_19_5 , 
            n4995, \REG.mem_19_4 , n4994, \REG.mem_19_3 , n4993, n4992, 
            n4991, \REG.mem_19_0 , n4990, \REG.mem_18_15 , n4989, 
            \REG.mem_18_14 , n4988, n4987, n4986, \REG.mem_18_11 , 
            n4985, n4984, \REG.mem_18_9 , n4983, n4982, n4981, \REG.mem_18_6 , 
            n4980, \REG.mem_18_5 , n4979, \REG.mem_18_4 , n4978, \REG.mem_18_3 , 
            n4977, n4976, n4975, \REG.mem_18_0 , n4974, \REG.mem_17_15 , 
            n4973, \REG.mem_17_14 , n4972, n4971, n4970, \REG.mem_17_11 , 
            n4969, n4968, \REG.mem_17_9 , n4967, n4966, n4965, \REG.mem_17_6 , 
            n4964, \REG.mem_17_5 , n4963, \REG.mem_17_4 , n4962, \REG.mem_17_3 , 
            n4961, n4960, n4958, \REG.mem_17_0 , n4957, \REG.mem_16_15 , 
            n4956, \REG.mem_16_14 , n4955, n4954, n4953, \REG.mem_16_11 , 
            n4952, n51, n4951, \REG.mem_16_9 , n4950, n4949, n4948, 
            \REG.mem_16_6 , n4947, \REG.mem_16_5 , n4946, \REG.mem_16_4 , 
            n4945, \REG.mem_16_3 , n4944, n4943, n4942, \REG.mem_16_0 , 
            n4941, n4940, \REG.mem_15_14 , n4939, n4938, n4937, 
            \REG.mem_15_11 , \rd_addr_nxt_c_6__N_465[5] , n19, n4936, 
            n4935, get_next_word, \rd_addr_nxt_c_6__N_465[3] , n4934, 
            n4933, n4932, n4931, n4930, \REG.mem_15_4 , n4929, \REG.mem_15_3 , 
            n4928, n4927, n4926, n4925, n4924, \REG.mem_14_14 , 
            n4923, n4922, n4921, \REG.mem_14_11 , n4920, n4919, 
            n4918, \rd_addr_nxt_c_6__N_465[1] , \state_timeout_counter[3] , 
            n718, n7, n14424, n4917, n4916, n4915, n4914, \REG.mem_14_4 , 
            n4913, \REG.mem_14_3 , n4912, n4911, n4910, \REG.mem_6_15 , 
            \REG.mem_7_15 , \REG.mem_5_15 , \REG.mem_4_15 , \REG.mem_10_15 , 
            \REG.mem_11_15 , \REG.mem_9_15 , \REG.mem_8_15 , n50, n52, 
            n20, n18, n4909, n4908, \REG.mem_13_14 , n4907, n4906, 
            n4905, \REG.mem_13_11 , n4904, n4903, n4902, n4901, 
            n46, n4900, n4899, n14, \REG.mem_10_11 , \REG.mem_11_11 , 
            n4898, \REG.mem_13_4 , n4897, \REG.mem_13_3 , \REG.mem_9_11 , 
            \REG.mem_8_11 , \REG.mem_12_14 , \REG.mem_12_11 , n4896, 
            n4895, n4894, n4893, n4892, n53, n4891, n4890, n21, 
            n4889, n4888, n4887, n4886, n4885, n4884, n4883, n4882, 
            \REG.mem_12_4 , n4881, \REG.mem_12_3 , n4880, n4879, n4878, 
            n4646, n4644, n4639, n4877, n4876, n4875, n4874, n4873, 
            n4872, n4871, n4870, \REG.mem_11_8 , n4869, n4638, n4868, 
            n4867, n4866, \REG.mem_11_4 , n4865, n4864, n4863, n4862, 
            n4861, n4860, n4859, n54, n22, n39, n7_adj_4, n4858, 
            n4857, n4856, n4855, n4854, \REG.mem_10_8 , n4853, n4852, 
            n4851, n56, n24, n4850, \REG.mem_10_4 , n4849, n4848, 
            n4847, n4846, n4845, n4844, n4843, n4842, n4841, n4840, 
            n4839, \afull_flag_impl.af_flag_p_w_N_603[3] , n4838, \REG.mem_9_8 , 
            n4837, n4836, n4835, n4834, \REG.mem_9_4 , n4833, n4832, 
            n4831, n4830, n4829, n4828, n4827, n4826, n4825, n4824, 
            n4823, n4822, \REG.mem_8_8 , n4821, n4820, n4819, n4818, 
            \REG.mem_8_4 , n4817, n4816, n4815, n4814, n4813, n4812, 
            n4811, \REG.mem_7_13 , n4810, n4809, n4808, n4807, \REG.mem_7_9 , 
            n4806, n4805, n4804, \REG.mem_7_6 , n4803, \REG.mem_7_5 , 
            n4802, \REG.mem_7_4 , n4801, n4800, n4799, n4798, \REG.mem_7_0 , 
            n4797, n4796, n4795, \REG.mem_6_13 , n4794, n4793, n4792, 
            n4791, \REG.mem_6_9 , n4790, n4789, n4788, \REG.mem_6_6 , 
            n4787, \REG.mem_6_5 , n4786, \REG.mem_6_4 , n4785, n4784, 
            n4783, n4779, \REG.mem_6_0 , n4778, n4777, n4776, \REG.mem_5_13 , 
            n4775, n4774, n4773, n4772, \REG.mem_5_9 , n4771, n4770, 
            n4769, \REG.mem_5_6 , n4768, \REG.mem_5_5 , n4767, \REG.mem_5_4 , 
            n4766, n4765, n4764, n4763, \REG.mem_5_0 , n4762, n4761, 
            n4760, \REG.mem_4_13 , n4759, n4758, n4757, n4756, \REG.mem_4_9 , 
            n4755, n4754, n4753, \REG.mem_4_6 , n4752, \REG.mem_4_5 , 
            n4751, \REG.mem_4_4 , n4750, n4749, n4748, n4747, \REG.mem_4_0 , 
            n4612, n57, n25, n42, n10, n49, n17, n48, n16, 
            n55, n23, n59, n27) /* synthesis syn_module_defined=1 */ ;
    output \REG.mem_58_4 ;
    input GND_net;
    output \REG.mem_14_8 ;
    output \REG.mem_15_8 ;
    input \dc32_fifo_data_in[10] ;
    input \dc32_fifo_data_in[9] ;
    input DEBUG_6_c_c;
    output \REG.mem_13_8 ;
    output \REG.mem_12_8 ;
    input \dc32_fifo_data_in[8] ;
    output \REG.mem_10_10 ;
    output \REG.mem_11_10 ;
    output \REG.mem_9_10 ;
    output \REG.mem_8_10 ;
    output t_rd_fifo_en_w;
    output \REG.out_raw[0] ;
    input SLM_CLK_c;
    input \dc32_fifo_data_in[7] ;
    output \REG.mem_10_13 ;
    output \REG.mem_11_13 ;
    output \REG.mem_9_13 ;
    output \REG.mem_8_13 ;
    input \dc32_fifo_data_in[6] ;
    output DEBUG_9_c;
    output n7596;
    output \wr_addr_nxt_c[4] ;
    output \REG.mem_26_14 ;
    input \dc32_fifo_data_in[5] ;
    output \REG.mem_42_2 ;
    output \REG.mem_43_2 ;
    output \REG.mem_41_2 ;
    output \REG.mem_40_2 ;
    output \REG.mem_14_10 ;
    output \REG.mem_15_10 ;
    input reset_all;
    output \REG.mem_55_8 ;
    output \REG.mem_13_10 ;
    output \REG.mem_12_10 ;
    input \dc32_fifo_data_in[4] ;
    output \REG.mem_42_3 ;
    output \REG.mem_43_3 ;
    output \REG.mem_41_3 ;
    output \REG.mem_40_3 ;
    output \rd_grey_sync_r[0] ;
    input \dc32_fifo_data_in[3] ;
    output \REG.mem_58_8 ;
    output DEBUG_5_c;
    output [6:0]wr_grey_sync_r;
    output \REG.mem_48_5 ;
    output \REG.mem_49_5 ;
    input \aempty_flag_impl.ae_flag_nxt_w ;
    output dc32_fifo_almost_empty;
    input \dc32_fifo_data_in[2] ;
    output \REG.mem_55_11 ;
    output \REG.mem_50_5 ;
    output \REG.mem_51_5 ;
    input \dc32_fifo_data_in[1] ;
    output \REG.mem_55_5 ;
    output \REG.mem_63_4 ;
    output \REG.mem_23_11 ;
    input \dc32_fifo_data_in[0] ;
    output \REG.mem_10_12 ;
    output \REG.mem_11_12 ;
    output \REG.mem_9_12 ;
    output \REG.mem_8_12 ;
    output \REG.mem_38_11 ;
    output \REG.mem_39_11 ;
    output \REG.mem_37_11 ;
    output \REG.mem_36_11 ;
    output \REG.mem_14_12 ;
    output \REG.mem_15_12 ;
    output \REG.mem_14_13 ;
    output \REG.mem_15_13 ;
    output \REG.mem_6_12 ;
    output \REG.mem_7_12 ;
    output \REG.mem_4_12 ;
    output \REG.mem_5_12 ;
    output \REG.mem_13_13 ;
    output \REG.mem_12_13 ;
    output \REG.mem_13_12 ;
    output \REG.mem_12_12 ;
    output \REG.mem_23_15 ;
    output \REG.mem_18_12 ;
    output \REG.mem_19_12 ;
    output \REG.mem_6_8 ;
    output \REG.mem_7_8 ;
    output \REG.mem_17_12 ;
    output \REG.mem_16_12 ;
    output \wr_addr_nxt_c[2] ;
    output \REG.mem_26_0 ;
    output \REG.mem_42_10 ;
    output \REG.mem_43_10 ;
    output \REG.mem_18_8 ;
    output \REG.mem_19_8 ;
    output \REG.mem_14_15 ;
    output \REG.mem_15_15 ;
    output \REG.mem_17_8 ;
    output \REG.mem_16_8 ;
    output \REG.mem_41_10 ;
    output \REG.mem_40_10 ;
    output n60;
    output \REG.mem_18_13 ;
    output \REG.mem_19_13 ;
    output \REG.mem_17_13 ;
    output \REG.mem_16_13 ;
    output n28;
    output \REG.mem_13_15 ;
    output \REG.mem_12_15 ;
    output \REG.mem_26_3 ;
    output \REG.mem_46_6 ;
    output \REG.mem_47_6 ;
    output \REG.mem_45_6 ;
    output \REG.mem_44_6 ;
    output \REG.mem_63_8 ;
    output \REG.mem_46_2 ;
    output \REG.mem_47_2 ;
    output \REG.mem_45_2 ;
    output \REG.mem_44_2 ;
    input \dc32_fifo_data_in[15] ;
    input \dc32_fifo_data_in[14] ;
    output \REG.mem_6_7 ;
    output \REG.mem_7_7 ;
    input \dc32_fifo_data_in[13] ;
    output \REG.mem_46_11 ;
    output \REG.mem_47_11 ;
    input \dc32_fifo_data_in[12] ;
    output \REG.mem_5_7 ;
    output \REG.mem_4_7 ;
    input \dc32_fifo_data_in[11] ;
    output \REG.mem_45_11 ;
    output \REG.mem_44_11 ;
    output \REG.mem_23_13 ;
    output \REG.mem_58_5 ;
    output \REG.mem_23_8 ;
    output \REG.mem_46_3 ;
    output \REG.mem_47_3 ;
    output \REG.mem_10_7 ;
    output \REG.mem_11_7 ;
    output \REG.mem_45_3 ;
    output \REG.mem_44_3 ;
    output \REG.mem_8_2 ;
    output \REG.mem_9_2 ;
    output \REG.mem_9_7 ;
    output \REG.mem_8_7 ;
    output \REG.mem_31_14 ;
    output \REG.mem_10_2 ;
    output \REG.mem_11_2 ;
    output \REG.mem_58_13 ;
    output \REG.mem_26_8 ;
    output \REG.mem_14_2 ;
    output \REG.mem_15_2 ;
    output \REG.mem_12_2 ;
    output \REG.mem_13_2 ;
    output \REG.mem_14_7 ;
    output \REG.mem_15_7 ;
    output \REG.mem_13_7 ;
    output \REG.mem_12_7 ;
    output \REG.mem_26_13 ;
    output \REG.mem_6_3 ;
    output \REG.mem_7_3 ;
    output \REG.mem_5_3 ;
    output \REG.mem_4_3 ;
    output \REG.mem_40_1 ;
    output \REG.mem_41_1 ;
    output \REG.mem_14_5 ;
    output \REG.mem_15_5 ;
    output \REG.mem_13_5 ;
    output \REG.mem_12_5 ;
    output \REG.mem_42_1 ;
    output \REG.mem_43_1 ;
    output \REG.mem_46_1 ;
    output \REG.mem_47_1 ;
    output \REG.mem_44_1 ;
    output \REG.mem_45_1 ;
    output \REG.mem_31_8 ;
    output \REG.mem_26_10 ;
    output \REG.mem_18_2 ;
    output \REG.mem_19_2 ;
    output \REG.mem_31_3 ;
    output \REG.mem_17_2 ;
    output \REG.mem_16_2 ;
    output n61;
    output \REG.mem_63_13 ;
    output n34;
    output n29;
    output \REG.mem_50_6 ;
    output \REG.mem_51_6 ;
    output n58;
    output \REG.mem_6_14 ;
    output \REG.mem_7_14 ;
    output n26;
    output \REG.mem_6_10 ;
    output \REG.mem_7_10 ;
    output \REG.mem_4_10 ;
    output \REG.mem_5_10 ;
    output \REG.mem_4_14 ;
    output \REG.mem_5_14 ;
    input n5896;
    input VCC_net;
    output \fifo_data_out[6] ;
    input n5893;
    output \fifo_data_out[5] ;
    output \REG.mem_16_10 ;
    output \REG.mem_17_10 ;
    output \REG.mem_18_10 ;
    output \REG.mem_19_10 ;
    input n11119;
    output \fifo_data_out[7] ;
    output \REG.mem_18_7 ;
    output \REG.mem_19_7 ;
    input n11139;
    output \fifo_data_out[3] ;
    output \REG.mem_17_7 ;
    output \REG.mem_16_7 ;
    output \REG.mem_50_2 ;
    output \REG.mem_51_2 ;
    output \REG.mem_46_0 ;
    output \REG.mem_47_0 ;
    output \REG.mem_46_9 ;
    output \REG.mem_47_9 ;
    output \REG.mem_45_9 ;
    output \REG.mem_44_9 ;
    output \REG.mem_49_6 ;
    output \REG.mem_48_6 ;
    output \REG.mem_49_2 ;
    output \REG.mem_48_2 ;
    input n11097;
    output \fifo_data_out[8] ;
    input n5854;
    output \fifo_data_out[0] ;
    output \REG.mem_5_8 ;
    output \REG.mem_4_8 ;
    output \REG.mem_6_11 ;
    output \REG.mem_7_11 ;
    output \REG.mem_58_1 ;
    output \REG.mem_26_15 ;
    input n11095;
    output \fifo_data_out[9] ;
    output \REG.mem_23_7 ;
    input n11143;
    output \fifo_data_out[1] ;
    input n11141;
    output \fifo_data_out[2] ;
    input n11089;
    output \fifo_data_out[10] ;
    input n11135;
    output \fifo_data_out[11] ;
    output \REG.mem_50_3 ;
    output \REG.mem_51_3 ;
    output \REG.mem_31_13 ;
    output \REG.mem_49_3 ;
    output \REG.mem_48_3 ;
    output \REG.mem_10_9 ;
    output \REG.mem_11_9 ;
    output \REG.mem_9_9 ;
    output \REG.mem_8_9 ;
    output \REG.mem_23_10 ;
    output \REG.mem_26_1 ;
    output n47;
    input n5789;
    output \REG.mem_63_15 ;
    input n5788;
    output \REG.mem_63_14 ;
    input n5787;
    output \REG.mem_31_11 ;
    output \REG.mem_5_11 ;
    output \REG.mem_4_11 ;
    output \REG.mem_31_1 ;
    output \REG.mem_23_12 ;
    input n5786;
    output \REG.mem_63_12 ;
    input n5785;
    output \REG.mem_63_11 ;
    input n5784;
    output \REG.mem_63_10 ;
    input n5783;
    output \REG.mem_63_9 ;
    output \REG.mem_14_9 ;
    output \REG.mem_15_9 ;
    input n5782;
    input n5781;
    output \REG.mem_63_7 ;
    input n5780;
    output \REG.mem_63_6 ;
    input n5779;
    output \REG.mem_63_5 ;
    input n5778;
    input n5777;
    output \REG.mem_63_3 ;
    input n5776;
    output \REG.mem_63_2 ;
    input n5775;
    output \REG.mem_63_1 ;
    input n11133;
    output \fifo_data_out[12] ;
    input n5773;
    output \REG.mem_63_0 ;
    output \REG.mem_13_9 ;
    output \REG.mem_12_9 ;
    output \REG.mem_38_10 ;
    output \REG.mem_39_10 ;
    output n15;
    output \REG.mem_36_10 ;
    output \REG.mem_37_10 ;
    output \REG.mem_8_1 ;
    output \REG.mem_9_1 ;
    output \REG.mem_10_1 ;
    output \REG.mem_11_1 ;
    input n11137;
    output \fifo_data_out[4] ;
    output \REG.mem_14_1 ;
    output \REG.mem_15_1 ;
    output \REG.mem_12_1 ;
    output \REG.mem_13_1 ;
    output \REG.mem_38_12 ;
    output \REG.mem_39_12 ;
    output \REG.mem_36_12 ;
    output \REG.mem_37_12 ;
    output \REG.mem_38_5 ;
    output \REG.mem_39_5 ;
    input n5709;
    output [6:0]rp_sync1_r;
    input n5708;
    input n5707;
    input n5706;
    input n5705;
    output \REG.mem_36_5 ;
    output \REG.mem_37_5 ;
    output \REG.mem_48_12 ;
    output \REG.mem_49_12 ;
    output \wr_addr_r[0] ;
    output \REG.mem_50_12 ;
    output \REG.mem_51_12 ;
    output \REG.mem_55_12 ;
    output \wr_addr_p1_w[6] ;
    input n5704;
    output \rd_sig_diff0_w[1] ;
    input n5686;
    input n5685;
    input n5684;
    input n5683;
    input n5682;
    output \REG.mem_58_15 ;
    input n5681;
    output \REG.mem_58_14 ;
    input n5680;
    input n5679;
    output \REG.mem_58_12 ;
    input n5678;
    output \REG.mem_58_11 ;
    input n5677;
    output \REG.mem_58_10 ;
    input n5676;
    output \REG.mem_58_9 ;
    input n5675;
    input n5674;
    output \REG.mem_58_7 ;
    input n5673;
    output \REG.mem_58_6 ;
    output \REG.mem_26_7 ;
    output \rd_sig_diff0_w[0] ;
    input n5672;
    input n5671;
    input n5670;
    output \REG.mem_58_3 ;
    input n5669;
    output \REG.mem_58_2 ;
    input n5668;
    input n5667;
    output \REG.mem_58_0 ;
    input n5666;
    input n5665;
    input n5664;
    input n5662;
    input n5660;
    output \rd_addr_r[6] ;
    output \REG.out_raw[15] ;
    output \REG.out_raw[14] ;
    output \REG.out_raw[13] ;
    output \REG.out_raw[12] ;
    output \REG.out_raw[11] ;
    output \REG.out_raw[10] ;
    output \REG.out_raw[9] ;
    output \REG.out_raw[8] ;
    output \REG.out_raw[7] ;
    output \REG.out_raw[6] ;
    output \REG.out_raw[5] ;
    output \REG.out_raw[4] ;
    output \REG.out_raw[3] ;
    output \REG.out_raw[2] ;
    output \REG.out_raw[1] ;
    output \REG.mem_31_7 ;
    output \REG.mem_42_11 ;
    output \REG.mem_43_11 ;
    output \REG.mem_41_11 ;
    output \REG.mem_40_11 ;
    output n2;
    output \REG.mem_6_1 ;
    output \REG.mem_7_1 ;
    output \REG.mem_4_1 ;
    output \REG.mem_5_1 ;
    output \REG.mem_38_4 ;
    output \REG.mem_39_4 ;
    output \REG.mem_16_1 ;
    output \REG.mem_17_1 ;
    output \REG.mem_37_4 ;
    output \REG.mem_36_4 ;
    output \REG.mem_55_2 ;
    output \REG.mem_18_1 ;
    output \REG.mem_19_1 ;
    input n5626;
    output \REG.mem_55_15 ;
    output \REG.mem_23_1 ;
    output \REG.mem_31_10 ;
    input n5625;
    output \REG.mem_55_14 ;
    input n5624;
    output \REG.mem_55_13 ;
    input n5623;
    input n5622;
    input n5621;
    output \REG.mem_55_10 ;
    input n5620;
    output \REG.mem_55_9 ;
    input n5619;
    input n5618;
    output \REG.mem_55_7 ;
    input n5617;
    output \REG.mem_55_6 ;
    input n5616;
    input n5615;
    output \REG.mem_55_4 ;
    input n5614;
    output \REG.mem_55_3 ;
    input n5613;
    input n5612;
    output \REG.mem_55_1 ;
    input n11073;
    output \fifo_data_out[13] ;
    input n5610;
    output \REG.mem_55_0 ;
    input n5609;
    output [6:0]wp_sync1_r;
    input n5608;
    input n5607;
    input n5606;
    input n5605;
    input n5604;
    input n5603;
    input n5586;
    input n5585;
    input n5584;
    input n5583;
    input n5582;
    input n11071;
    output \fifo_data_out[14] ;
    output \REG.mem_38_1 ;
    output \REG.mem_39_1 ;
    output \REG.mem_36_1 ;
    output \REG.mem_37_1 ;
    output \REG.mem_6_2 ;
    output \REG.mem_7_2 ;
    output \REG.mem_5_2 ;
    output \REG.mem_4_2 ;
    input n5548;
    output \REG.mem_51_15 ;
    input n5547;
    output \REG.mem_51_14 ;
    input n5546;
    output \REG.mem_51_13 ;
    input n5545;
    input n5544;
    output \REG.mem_51_11 ;
    input n5543;
    output \REG.mem_51_10 ;
    input n5542;
    output \REG.mem_51_9 ;
    input n5541;
    output \REG.mem_51_8 ;
    input n5540;
    output \REG.mem_51_7 ;
    input n5539;
    input n5538;
    input n5537;
    output \REG.mem_51_4 ;
    input n5536;
    input n5535;
    input n5534;
    output \REG.mem_51_1 ;
    input n5533;
    output \REG.mem_51_0 ;
    input n5532;
    output \REG.mem_50_15 ;
    output \REG.mem_48_1 ;
    output \REG.mem_49_1 ;
    input n5531;
    output \REG.mem_50_14 ;
    input n5530;
    output \REG.mem_50_13 ;
    input n5529;
    input n5528;
    output \REG.mem_50_11 ;
    input n5527;
    output \REG.mem_50_10 ;
    input n5526;
    output \REG.mem_50_9 ;
    input n5525;
    output \REG.mem_50_8 ;
    input n5524;
    output \REG.mem_50_7 ;
    input n5523;
    input n5522;
    input n5521;
    output \REG.mem_50_4 ;
    input n5520;
    input n5519;
    input n5518;
    output \REG.mem_50_1 ;
    input n5517;
    output \REG.mem_50_0 ;
    input n5516;
    output \REG.mem_49_15 ;
    input n5515;
    output \REG.mem_49_14 ;
    output \REG.mem_31_12 ;
    output \REG.mem_26_11 ;
    input n5514;
    output \REG.mem_49_13 ;
    input n5513;
    input n5512;
    output \REG.mem_49_11 ;
    input n5511;
    output \REG.mem_49_10 ;
    input n5510;
    output \REG.mem_49_9 ;
    input n5509;
    output \REG.mem_49_8 ;
    input n5508;
    output \REG.mem_49_7 ;
    input n5507;
    input n5506;
    input n5505;
    output \REG.mem_49_4 ;
    input n5504;
    input n5503;
    input n5502;
    input n5501;
    output \REG.mem_49_0 ;
    output \REG.mem_31_0 ;
    output \REG.mem_26_4 ;
    input n5492;
    output \REG.mem_48_15 ;
    input n5491;
    input n5490;
    output \REG.mem_48_14 ;
    input n5489;
    output \REG.mem_48_13 ;
    input n5488;
    input n5487;
    output \REG.mem_48_11 ;
    input n5486;
    output \REG.mem_48_10 ;
    input n5485;
    output \REG.mem_48_9 ;
    input n5484;
    output \REG.mem_48_8 ;
    input n5483;
    output \REG.mem_48_7 ;
    output \REG.mem_46_10 ;
    output \REG.mem_47_10 ;
    input n5482;
    input n5481;
    input n5480;
    output \REG.mem_48_4 ;
    input n5479;
    input n5478;
    input n5477;
    input n5476;
    output \REG.mem_48_0 ;
    input n5474;
    input n5472;
    output \REG.mem_47_15 ;
    input n5471;
    output \REG.mem_47_14 ;
    input n5470;
    output \REG.mem_47_13 ;
    input n5469;
    output \REG.mem_47_12 ;
    input n5468;
    input n5467;
    output \REG.mem_45_0 ;
    output \REG.mem_44_0 ;
    output \REG.mem_45_10 ;
    output \REG.mem_44_10 ;
    input n5466;
    input n5465;
    output \REG.mem_47_8 ;
    input n5464;
    output \REG.mem_47_7 ;
    input n5463;
    input n5462;
    output \REG.mem_47_5 ;
    input n5461;
    output \REG.mem_47_4 ;
    input n5460;
    input n5459;
    input n5458;
    input n5457;
    input n5456;
    output \REG.mem_46_15 ;
    input n5455;
    output \REG.mem_46_14 ;
    input n5454;
    output \REG.mem_46_13 ;
    input n5453;
    output \REG.mem_46_12 ;
    input n5452;
    input n5451;
    input n5450;
    input n5449;
    output \REG.mem_46_8 ;
    input n5448;
    output \REG.mem_46_7 ;
    input n5447;
    input n5446;
    output \REG.mem_46_5 ;
    input n5445;
    output \REG.mem_46_4 ;
    input n5444;
    input n5443;
    input n5442;
    input n5441;
    input n5440;
    output \REG.mem_45_15 ;
    input n5439;
    output \REG.mem_45_14 ;
    input n5438;
    output \REG.mem_45_13 ;
    input n5437;
    output \REG.mem_45_12 ;
    input n5436;
    input n5435;
    input n5434;
    output \REG.mem_38_7 ;
    output \REG.mem_39_7 ;
    output \REG.mem_37_7 ;
    output \REG.mem_36_7 ;
    input n5433;
    output \REG.mem_45_8 ;
    input n5432;
    output \REG.mem_45_7 ;
    input n5431;
    input n5430;
    output \REG.mem_45_5 ;
    input n5429;
    output \REG.mem_45_4 ;
    input n5428;
    input n5427;
    input n5426;
    input n5425;
    input n5424;
    output \REG.mem_44_15 ;
    input n5423;
    output \REG.mem_44_14 ;
    input n5422;
    output \REG.mem_44_13 ;
    input n5421;
    output \REG.mem_44_12 ;
    input n5420;
    input n5419;
    output \REG.mem_10_0 ;
    output \REG.mem_11_0 ;
    input n5418;
    output \REG.mem_9_0 ;
    output \REG.mem_8_0 ;
    input n5417;
    output \REG.mem_44_8 ;
    input n5416;
    output \REG.mem_44_7 ;
    input n5415;
    input n5414;
    output \REG.mem_44_5 ;
    input n5413;
    output \REG.mem_44_4 ;
    input n5412;
    input n5411;
    input n5410;
    input n5409;
    input n5408;
    input n5407;
    output \REG.mem_43_15 ;
    input n5406;
    output \REG.mem_43_14 ;
    input n5405;
    output \REG.mem_43_13 ;
    input n5404;
    output \REG.mem_43_12 ;
    input n5403;
    input n5402;
    output \REG.mem_10_5 ;
    output \REG.mem_11_5 ;
    output \REG.mem_9_5 ;
    output \REG.mem_8_5 ;
    output \wr_addr_p1_w[0] ;
    input n5401;
    output \REG.mem_43_9 ;
    input n5400;
    output \REG.mem_43_8 ;
    input n5399;
    output \REG.mem_43_7 ;
    input n5398;
    output \REG.mem_43_6 ;
    input n5397;
    output \REG.mem_43_5 ;
    input n5396;
    output \REG.mem_43_4 ;
    input n5395;
    input n5394;
    input n5393;
    input n5392;
    output \REG.mem_43_0 ;
    input n11069;
    output \fifo_data_out[15] ;
    input n5390;
    output \REG.mem_42_15 ;
    input n5389;
    output \REG.mem_42_14 ;
    input n5388;
    output \REG.mem_42_13 ;
    input n5387;
    output \REG.mem_42_12 ;
    input n5386;
    output \REG.mem_42_4 ;
    output \REG.mem_41_4 ;
    output \REG.mem_40_4 ;
    input n5385;
    input n5384;
    output \REG.mem_42_9 ;
    input n5383;
    output \REG.mem_42_8 ;
    input n5382;
    output \REG.mem_42_7 ;
    input n5381;
    output \REG.mem_42_6 ;
    input n5380;
    output \REG.mem_42_5 ;
    input n5379;
    input n5378;
    input n5377;
    input n5376;
    input n5375;
    output \REG.mem_42_0 ;
    input n5374;
    output \REG.mem_41_15 ;
    input n5373;
    output \REG.mem_41_14 ;
    input n5372;
    output \REG.mem_41_13 ;
    input n5371;
    output \REG.mem_41_12 ;
    input n4667;
    input n5370;
    input n5369;
    input n5368;
    output \REG.mem_41_9 ;
    input n5367;
    output \REG.mem_41_8 ;
    input n5366;
    output \REG.mem_41_7 ;
    input n5365;
    output \REG.mem_41_6 ;
    input n5364;
    output \REG.mem_41_5 ;
    input n5363;
    input n5362;
    input n5361;
    input n5360;
    input n5358;
    output \REG.mem_41_0 ;
    input n5357;
    output \REG.mem_40_15 ;
    input n5356;
    output \REG.mem_40_14 ;
    input n5355;
    output \REG.mem_40_13 ;
    input n5354;
    output \REG.mem_40_12 ;
    output \REG.mem_38_13 ;
    output \REG.mem_39_13 ;
    output \REG.mem_37_13 ;
    output \REG.mem_36_13 ;
    input n5353;
    input n5352;
    input n5351;
    output \REG.mem_40_9 ;
    input n5350;
    output \REG.mem_40_8 ;
    input n5349;
    output \REG.mem_40_7 ;
    input n5348;
    output \REG.mem_40_6 ;
    input n5347;
    output \REG.mem_40_5 ;
    input n5346;
    input n5345;
    input n5344;
    input n5343;
    input n5342;
    output \REG.mem_40_0 ;
    input n5341;
    output \REG.mem_39_15 ;
    input n5340;
    output \REG.mem_39_14 ;
    input n5339;
    output \REG.mem_23_5 ;
    output \REG.mem_14_0 ;
    output \REG.mem_15_0 ;
    output \REG.mem_13_0 ;
    output \REG.mem_12_0 ;
    input n5338;
    input n5337;
    input n5336;
    input n5335;
    output \REG.mem_39_9 ;
    input n5334;
    output \REG.mem_39_8 ;
    input n5333;
    input n5332;
    output \REG.mem_39_6 ;
    input n5331;
    input n5330;
    input n5329;
    output \REG.mem_39_3 ;
    input n5328;
    output \REG.mem_39_2 ;
    input n5327;
    input n5326;
    output \REG.mem_39_0 ;
    input n5323;
    output \REG.mem_38_15 ;
    input n5322;
    output \REG.mem_38_14 ;
    input n5321;
    input n5320;
    input n5319;
    input n5318;
    input n5317;
    output \REG.mem_38_9 ;
    input n5316;
    output \REG.mem_38_8 ;
    input n5315;
    input n5314;
    output \REG.mem_38_6 ;
    input n5313;
    input n5312;
    input n5311;
    output \REG.mem_38_3 ;
    input n5310;
    output \REG.mem_38_2 ;
    input n5309;
    input n5308;
    output \REG.mem_38_0 ;
    input n5302;
    output \REG.mem_37_15 ;
    input n5301;
    output \REG.mem_37_14 ;
    input n5300;
    input n5299;
    input n5298;
    input n5297;
    input n5296;
    output \REG.mem_37_9 ;
    input n5295;
    output \REG.mem_37_8 ;
    input n5294;
    input n5293;
    output \REG.mem_37_6 ;
    input n5292;
    input n5291;
    input n5290;
    output \REG.mem_37_3 ;
    input n5289;
    output \REG.mem_37_2 ;
    input n5288;
    input n5286;
    output \REG.mem_37_0 ;
    input n5285;
    output \REG.mem_36_15 ;
    input n5284;
    output \REG.mem_36_14 ;
    input n5283;
    input n5282;
    input n5281;
    input n5280;
    input n5279;
    output \REG.mem_36_9 ;
    input n5278;
    output \REG.mem_36_8 ;
    input n5277;
    input n5276;
    output \REG.mem_36_6 ;
    input n5275;
    input n5274;
    input n5273;
    output \REG.mem_36_3 ;
    input n5272;
    output \REG.mem_36_2 ;
    input n5271;
    input n5270;
    output \REG.mem_36_0 ;
    output \REG.mem_26_12 ;
    output \REG.mem_10_3 ;
    output \REG.mem_11_3 ;
    input n5202;
    output \REG.mem_31_15 ;
    input n5201;
    input n5200;
    input n5199;
    input n5198;
    input n5197;
    input n5196;
    output \REG.mem_31_9 ;
    input n5195;
    input n5194;
    input n5193;
    output \REG.mem_31_6 ;
    input n5192;
    output \REG.mem_31_5 ;
    input n5191;
    output \REG.mem_31_4 ;
    input n5190;
    input n5189;
    output \REG.mem_31_2 ;
    output \REG.mem_9_3 ;
    output \REG.mem_8_3 ;
    input n5188;
    input n5187;
    output \REG.mem_10_14 ;
    output \REG.mem_11_14 ;
    output \REG.mem_9_14 ;
    output \REG.mem_8_14 ;
    output \REG.mem_23_2 ;
    input n5121;
    input n5120;
    input n5119;
    input n5118;
    input n5117;
    input n5116;
    input n5115;
    output \REG.mem_26_9 ;
    input n5114;
    input n5113;
    input n5112;
    output \REG.mem_26_6 ;
    input n5111;
    output \REG.mem_26_5 ;
    input n5110;
    input n5109;
    input n5108;
    output \REG.mem_26_2 ;
    input n5107;
    input n5106;
    input n5073;
    input n5072;
    output \REG.mem_23_14 ;
    input n5071;
    input n5070;
    input n5069;
    input n5068;
    input n5067;
    output \REG.mem_23_9 ;
    input n5066;
    output \rd_grey_sync_r[5] ;
    output \rd_grey_sync_r[4] ;
    output \REG.mem_10_6 ;
    output \REG.mem_11_6 ;
    output \rd_grey_sync_r[3] ;
    output \rd_grey_sync_r[2] ;
    output \rd_grey_sync_r[1] ;
    input n5065;
    input n5064;
    output \REG.mem_23_6 ;
    input n5063;
    input n5062;
    output \REG.mem_23_4 ;
    input n5061;
    output \REG.mem_23_3 ;
    input n5060;
    input n5059;
    input n5058;
    output \REG.mem_23_0 ;
    output \REG.mem_9_6 ;
    output \REG.mem_8_6 ;
    output n5;
    output \REG.mem_14_6 ;
    output \REG.mem_15_6 ;
    output \REG.mem_13_6 ;
    output \REG.mem_12_6 ;
    input n5006;
    output \REG.mem_19_15 ;
    input n5005;
    output \REG.mem_19_14 ;
    input n5004;
    input n5003;
    input n5002;
    output \REG.mem_19_11 ;
    input n5001;
    input n5000;
    output \REG.mem_19_9 ;
    input n4999;
    input n4998;
    input n4997;
    output \REG.mem_19_6 ;
    input n4996;
    output \REG.mem_19_5 ;
    input n4995;
    output \REG.mem_19_4 ;
    input n4994;
    output \REG.mem_19_3 ;
    input n4993;
    input n4992;
    input n4991;
    output \REG.mem_19_0 ;
    input n4990;
    output \REG.mem_18_15 ;
    input n4989;
    output \REG.mem_18_14 ;
    input n4988;
    input n4987;
    input n4986;
    output \REG.mem_18_11 ;
    input n4985;
    input n4984;
    output \REG.mem_18_9 ;
    input n4983;
    input n4982;
    input n4981;
    output \REG.mem_18_6 ;
    input n4980;
    output \REG.mem_18_5 ;
    input n4979;
    output \REG.mem_18_4 ;
    input n4978;
    output \REG.mem_18_3 ;
    input n4977;
    input n4976;
    input n4975;
    output \REG.mem_18_0 ;
    input n4974;
    output \REG.mem_17_15 ;
    input n4973;
    output \REG.mem_17_14 ;
    input n4972;
    input n4971;
    input n4970;
    output \REG.mem_17_11 ;
    input n4969;
    input n4968;
    output \REG.mem_17_9 ;
    input n4967;
    input n4966;
    input n4965;
    output \REG.mem_17_6 ;
    input n4964;
    output \REG.mem_17_5 ;
    input n4963;
    output \REG.mem_17_4 ;
    input n4962;
    output \REG.mem_17_3 ;
    input n4961;
    input n4960;
    input n4958;
    output \REG.mem_17_0 ;
    input n4957;
    output \REG.mem_16_15 ;
    input n4956;
    output \REG.mem_16_14 ;
    input n4955;
    input n4954;
    input n4953;
    output \REG.mem_16_11 ;
    input n4952;
    output n51;
    input n4951;
    output \REG.mem_16_9 ;
    input n4950;
    input n4949;
    input n4948;
    output \REG.mem_16_6 ;
    input n4947;
    output \REG.mem_16_5 ;
    input n4946;
    output \REG.mem_16_4 ;
    input n4945;
    output \REG.mem_16_3 ;
    input n4944;
    input n4943;
    input n4942;
    output \REG.mem_16_0 ;
    input n4941;
    input n4940;
    output \REG.mem_15_14 ;
    input n4939;
    input n4938;
    input n4937;
    output \REG.mem_15_11 ;
    output \rd_addr_nxt_c_6__N_465[5] ;
    output n19;
    input n4936;
    input n4935;
    input get_next_word;
    output \rd_addr_nxt_c_6__N_465[3] ;
    input n4934;
    input n4933;
    input n4932;
    input n4931;
    input n4930;
    output \REG.mem_15_4 ;
    input n4929;
    output \REG.mem_15_3 ;
    input n4928;
    input n4927;
    input n4926;
    input n4925;
    input n4924;
    output \REG.mem_14_14 ;
    input n4923;
    input n4922;
    input n4921;
    output \REG.mem_14_11 ;
    input n4920;
    input n4919;
    input n4918;
    output \rd_addr_nxt_c_6__N_465[1] ;
    input \state_timeout_counter[3] ;
    input n718;
    input n7;
    output n14424;
    input n4917;
    input n4916;
    input n4915;
    input n4914;
    output \REG.mem_14_4 ;
    input n4913;
    output \REG.mem_14_3 ;
    input n4912;
    input n4911;
    input n4910;
    output \REG.mem_6_15 ;
    output \REG.mem_7_15 ;
    output \REG.mem_5_15 ;
    output \REG.mem_4_15 ;
    output \REG.mem_10_15 ;
    output \REG.mem_11_15 ;
    output \REG.mem_9_15 ;
    output \REG.mem_8_15 ;
    output n50;
    output n52;
    output n20;
    output n18;
    input n4909;
    input n4908;
    output \REG.mem_13_14 ;
    input n4907;
    input n4906;
    input n4905;
    output \REG.mem_13_11 ;
    input n4904;
    input n4903;
    input n4902;
    input n4901;
    output n46;
    input n4900;
    input n4899;
    output n14;
    output \REG.mem_10_11 ;
    output \REG.mem_11_11 ;
    input n4898;
    output \REG.mem_13_4 ;
    input n4897;
    output \REG.mem_13_3 ;
    output \REG.mem_9_11 ;
    output \REG.mem_8_11 ;
    output \REG.mem_12_14 ;
    output \REG.mem_12_11 ;
    input n4896;
    input n4895;
    input n4894;
    input n4893;
    input n4892;
    output n53;
    input n4891;
    input n4890;
    output n21;
    input n4889;
    input n4888;
    input n4887;
    input n4886;
    input n4885;
    input n4884;
    input n4883;
    input n4882;
    output \REG.mem_12_4 ;
    input n4881;
    output \REG.mem_12_3 ;
    input n4880;
    input n4879;
    input n4878;
    input n4646;
    input n4644;
    input n4639;
    input n4877;
    input n4876;
    input n4875;
    input n4874;
    input n4873;
    input n4872;
    input n4871;
    input n4870;
    output \REG.mem_11_8 ;
    input n4869;
    input n4638;
    input n4868;
    input n4867;
    input n4866;
    output \REG.mem_11_4 ;
    input n4865;
    input n4864;
    input n4863;
    input n4862;
    input n4861;
    input n4860;
    input n4859;
    output n54;
    output n22;
    output n39;
    output n7_adj_4;
    input n4858;
    input n4857;
    input n4856;
    input n4855;
    input n4854;
    output \REG.mem_10_8 ;
    input n4853;
    input n4852;
    input n4851;
    output n56;
    output n24;
    input n4850;
    output \REG.mem_10_4 ;
    input n4849;
    input n4848;
    input n4847;
    input n4846;
    input n4845;
    input n4844;
    input n4843;
    input n4842;
    input n4841;
    input n4840;
    input n4839;
    input \afull_flag_impl.af_flag_p_w_N_603[3] ;
    input n4838;
    output \REG.mem_9_8 ;
    input n4837;
    input n4836;
    input n4835;
    input n4834;
    output \REG.mem_9_4 ;
    input n4833;
    input n4832;
    input n4831;
    input n4830;
    input n4829;
    input n4828;
    input n4827;
    input n4826;
    input n4825;
    input n4824;
    input n4823;
    input n4822;
    output \REG.mem_8_8 ;
    input n4821;
    input n4820;
    input n4819;
    input n4818;
    output \REG.mem_8_4 ;
    input n4817;
    input n4816;
    input n4815;
    input n4814;
    input n4813;
    input n4812;
    input n4811;
    output \REG.mem_7_13 ;
    input n4810;
    input n4809;
    input n4808;
    input n4807;
    output \REG.mem_7_9 ;
    input n4806;
    input n4805;
    input n4804;
    output \REG.mem_7_6 ;
    input n4803;
    output \REG.mem_7_5 ;
    input n4802;
    output \REG.mem_7_4 ;
    input n4801;
    input n4800;
    input n4799;
    input n4798;
    output \REG.mem_7_0 ;
    input n4797;
    input n4796;
    input n4795;
    output \REG.mem_6_13 ;
    input n4794;
    input n4793;
    input n4792;
    input n4791;
    output \REG.mem_6_9 ;
    input n4790;
    input n4789;
    input n4788;
    output \REG.mem_6_6 ;
    input n4787;
    output \REG.mem_6_5 ;
    input n4786;
    output \REG.mem_6_4 ;
    input n4785;
    input n4784;
    input n4783;
    input n4779;
    output \REG.mem_6_0 ;
    input n4778;
    input n4777;
    input n4776;
    output \REG.mem_5_13 ;
    input n4775;
    input n4774;
    input n4773;
    input n4772;
    output \REG.mem_5_9 ;
    input n4771;
    input n4770;
    input n4769;
    output \REG.mem_5_6 ;
    input n4768;
    output \REG.mem_5_5 ;
    input n4767;
    output \REG.mem_5_4 ;
    input n4766;
    input n4765;
    input n4764;
    input n4763;
    output \REG.mem_5_0 ;
    input n4762;
    input n4761;
    input n4760;
    output \REG.mem_4_13 ;
    input n4759;
    input n4758;
    input n4757;
    input n4756;
    output \REG.mem_4_9 ;
    input n4755;
    input n4754;
    input n4753;
    output \REG.mem_4_6 ;
    input n4752;
    output \REG.mem_4_5 ;
    input n4751;
    output \REG.mem_4_4 ;
    input n4750;
    input n4749;
    input n4748;
    input n4747;
    output \REG.mem_4_0 ;
    input n4612;
    output n57;
    output n25;
    output n42;
    output n10;
    output n49;
    output n17;
    output n48;
    output n16;
    output n55;
    output n23;
    output n59;
    output n27;
    
    wire DEBUG_6_c_c /* synthesis is_clock=1, SET_AS_NETWORK=DEBUG_6_c_c */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 lscc_fifo_dc_inst (.\REG.mem_58_4 (\REG.mem_58_4 ), 
            .GND_net(GND_net), .\REG.mem_14_8 (\REG.mem_14_8 ), .\REG.mem_15_8 (\REG.mem_15_8 ), 
            .\dc32_fifo_data_in[10] (\dc32_fifo_data_in[10] ), .\dc32_fifo_data_in[9] (\dc32_fifo_data_in[9] ), 
            .DEBUG_6_c_c(DEBUG_6_c_c), .\REG.mem_13_8 (\REG.mem_13_8 ), 
            .\REG.mem_12_8 (\REG.mem_12_8 ), .\dc32_fifo_data_in[8] (\dc32_fifo_data_in[8] ), 
            .\REG.mem_10_10 (\REG.mem_10_10 ), .\REG.mem_11_10 (\REG.mem_11_10 ), 
            .\REG.mem_9_10 (\REG.mem_9_10 ), .\REG.mem_8_10 (\REG.mem_8_10 ), 
            .t_rd_fifo_en_w(t_rd_fifo_en_w), .\REG.out_raw[0] (\REG.out_raw[0] ), 
            .SLM_CLK_c(SLM_CLK_c), .\dc32_fifo_data_in[7] (\dc32_fifo_data_in[7] ), 
            .\REG.mem_10_13 (\REG.mem_10_13 ), .\REG.mem_11_13 (\REG.mem_11_13 ), 
            .\REG.mem_9_13 (\REG.mem_9_13 ), .\REG.mem_8_13 (\REG.mem_8_13 ), 
            .\dc32_fifo_data_in[6] (\dc32_fifo_data_in[6] ), .DEBUG_9_c(DEBUG_9_c), 
            .n7596(n7596), .\wr_addr_nxt_c[4] (\wr_addr_nxt_c[4] ), .\REG.mem_26_14 (\REG.mem_26_14 ), 
            .\dc32_fifo_data_in[5] (\dc32_fifo_data_in[5] ), .\REG.mem_42_2 (\REG.mem_42_2 ), 
            .\REG.mem_43_2 (\REG.mem_43_2 ), .\REG.mem_41_2 (\REG.mem_41_2 ), 
            .\REG.mem_40_2 (\REG.mem_40_2 ), .\REG.mem_14_10 (\REG.mem_14_10 ), 
            .\REG.mem_15_10 (\REG.mem_15_10 ), .reset_all(reset_all), .\REG.mem_55_8 (\REG.mem_55_8 ), 
            .\REG.mem_13_10 (\REG.mem_13_10 ), .\REG.mem_12_10 (\REG.mem_12_10 ), 
            .\dc32_fifo_data_in[4] (\dc32_fifo_data_in[4] ), .\REG.mem_42_3 (\REG.mem_42_3 ), 
            .\REG.mem_43_3 (\REG.mem_43_3 ), .\REG.mem_41_3 (\REG.mem_41_3 ), 
            .\REG.mem_40_3 (\REG.mem_40_3 ), .\rd_grey_sync_r[0] (\rd_grey_sync_r[0] ), 
            .\dc32_fifo_data_in[3] (\dc32_fifo_data_in[3] ), .\REG.mem_58_8 (\REG.mem_58_8 ), 
            .DEBUG_5_c(DEBUG_5_c), .wr_grey_sync_r({wr_grey_sync_r}), .\REG.mem_48_5 (\REG.mem_48_5 ), 
            .\REG.mem_49_5 (\REG.mem_49_5 ), .\aempty_flag_impl.ae_flag_nxt_w (\aempty_flag_impl.ae_flag_nxt_w ), 
            .dc32_fifo_almost_empty(dc32_fifo_almost_empty), .\dc32_fifo_data_in[2] (\dc32_fifo_data_in[2] ), 
            .\REG.mem_55_11 (\REG.mem_55_11 ), .\REG.mem_50_5 (\REG.mem_50_5 ), 
            .\REG.mem_51_5 (\REG.mem_51_5 ), .\dc32_fifo_data_in[1] (\dc32_fifo_data_in[1] ), 
            .\REG.mem_55_5 (\REG.mem_55_5 ), .\REG.mem_63_4 (\REG.mem_63_4 ), 
            .\REG.mem_23_11 (\REG.mem_23_11 ), .\dc32_fifo_data_in[0] (\dc32_fifo_data_in[0] ), 
            .\REG.mem_10_12 (\REG.mem_10_12 ), .\REG.mem_11_12 (\REG.mem_11_12 ), 
            .\REG.mem_9_12 (\REG.mem_9_12 ), .\REG.mem_8_12 (\REG.mem_8_12 ), 
            .\REG.mem_38_11 (\REG.mem_38_11 ), .\REG.mem_39_11 (\REG.mem_39_11 ), 
            .\REG.mem_37_11 (\REG.mem_37_11 ), .\REG.mem_36_11 (\REG.mem_36_11 ), 
            .\REG.mem_14_12 (\REG.mem_14_12 ), .\REG.mem_15_12 (\REG.mem_15_12 ), 
            .\REG.mem_14_13 (\REG.mem_14_13 ), .\REG.mem_15_13 (\REG.mem_15_13 ), 
            .\REG.mem_6_12 (\REG.mem_6_12 ), .\REG.mem_7_12 (\REG.mem_7_12 ), 
            .\REG.mem_4_12 (\REG.mem_4_12 ), .\REG.mem_5_12 (\REG.mem_5_12 ), 
            .\REG.mem_13_13 (\REG.mem_13_13 ), .\REG.mem_12_13 (\REG.mem_12_13 ), 
            .\REG.mem_13_12 (\REG.mem_13_12 ), .\REG.mem_12_12 (\REG.mem_12_12 ), 
            .\REG.mem_23_15 (\REG.mem_23_15 ), .\REG.mem_18_12 (\REG.mem_18_12 ), 
            .\REG.mem_19_12 (\REG.mem_19_12 ), .\REG.mem_6_8 (\REG.mem_6_8 ), 
            .\REG.mem_7_8 (\REG.mem_7_8 ), .\REG.mem_17_12 (\REG.mem_17_12 ), 
            .\REG.mem_16_12 (\REG.mem_16_12 ), .\wr_addr_nxt_c[2] (\wr_addr_nxt_c[2] ), 
            .\REG.mem_26_0 (\REG.mem_26_0 ), .\REG.mem_42_10 (\REG.mem_42_10 ), 
            .\REG.mem_43_10 (\REG.mem_43_10 ), .\REG.mem_18_8 (\REG.mem_18_8 ), 
            .\REG.mem_19_8 (\REG.mem_19_8 ), .\REG.mem_14_15 (\REG.mem_14_15 ), 
            .\REG.mem_15_15 (\REG.mem_15_15 ), .\REG.mem_17_8 (\REG.mem_17_8 ), 
            .\REG.mem_16_8 (\REG.mem_16_8 ), .\REG.mem_41_10 (\REG.mem_41_10 ), 
            .\REG.mem_40_10 (\REG.mem_40_10 ), .n60(n60), .\REG.mem_18_13 (\REG.mem_18_13 ), 
            .\REG.mem_19_13 (\REG.mem_19_13 ), .\REG.mem_17_13 (\REG.mem_17_13 ), 
            .\REG.mem_16_13 (\REG.mem_16_13 ), .n28(n28), .\REG.mem_13_15 (\REG.mem_13_15 ), 
            .\REG.mem_12_15 (\REG.mem_12_15 ), .\REG.mem_26_3 (\REG.mem_26_3 ), 
            .\REG.mem_46_6 (\REG.mem_46_6 ), .\REG.mem_47_6 (\REG.mem_47_6 ), 
            .\REG.mem_45_6 (\REG.mem_45_6 ), .\REG.mem_44_6 (\REG.mem_44_6 ), 
            .\REG.mem_63_8 (\REG.mem_63_8 ), .\REG.mem_46_2 (\REG.mem_46_2 ), 
            .\REG.mem_47_2 (\REG.mem_47_2 ), .\REG.mem_45_2 (\REG.mem_45_2 ), 
            .\REG.mem_44_2 (\REG.mem_44_2 ), .\dc32_fifo_data_in[15] (\dc32_fifo_data_in[15] ), 
            .\dc32_fifo_data_in[14] (\dc32_fifo_data_in[14] ), .\REG.mem_6_7 (\REG.mem_6_7 ), 
            .\REG.mem_7_7 (\REG.mem_7_7 ), .\dc32_fifo_data_in[13] (\dc32_fifo_data_in[13] ), 
            .\REG.mem_46_11 (\REG.mem_46_11 ), .\REG.mem_47_11 (\REG.mem_47_11 ), 
            .\dc32_fifo_data_in[12] (\dc32_fifo_data_in[12] ), .\REG.mem_5_7 (\REG.mem_5_7 ), 
            .\REG.mem_4_7 (\REG.mem_4_7 ), .\dc32_fifo_data_in[11] (\dc32_fifo_data_in[11] ), 
            .\REG.mem_45_11 (\REG.mem_45_11 ), .\REG.mem_44_11 (\REG.mem_44_11 ), 
            .\REG.mem_23_13 (\REG.mem_23_13 ), .\REG.mem_58_5 (\REG.mem_58_5 ), 
            .\REG.mem_23_8 (\REG.mem_23_8 ), .\REG.mem_46_3 (\REG.mem_46_3 ), 
            .\REG.mem_47_3 (\REG.mem_47_3 ), .\REG.mem_10_7 (\REG.mem_10_7 ), 
            .\REG.mem_11_7 (\REG.mem_11_7 ), .\REG.mem_45_3 (\REG.mem_45_3 ), 
            .\REG.mem_44_3 (\REG.mem_44_3 ), .\REG.mem_8_2 (\REG.mem_8_2 ), 
            .\REG.mem_9_2 (\REG.mem_9_2 ), .\REG.mem_9_7 (\REG.mem_9_7 ), 
            .\REG.mem_8_7 (\REG.mem_8_7 ), .\REG.mem_31_14 (\REG.mem_31_14 ), 
            .\REG.mem_10_2 (\REG.mem_10_2 ), .\REG.mem_11_2 (\REG.mem_11_2 ), 
            .\REG.mem_58_13 (\REG.mem_58_13 ), .\REG.mem_26_8 (\REG.mem_26_8 ), 
            .\REG.mem_14_2 (\REG.mem_14_2 ), .\REG.mem_15_2 (\REG.mem_15_2 ), 
            .\REG.mem_12_2 (\REG.mem_12_2 ), .\REG.mem_13_2 (\REG.mem_13_2 ), 
            .\REG.mem_14_7 (\REG.mem_14_7 ), .\REG.mem_15_7 (\REG.mem_15_7 ), 
            .\REG.mem_13_7 (\REG.mem_13_7 ), .\REG.mem_12_7 (\REG.mem_12_7 ), 
            .\REG.mem_26_13 (\REG.mem_26_13 ), .\REG.mem_6_3 (\REG.mem_6_3 ), 
            .\REG.mem_7_3 (\REG.mem_7_3 ), .\REG.mem_5_3 (\REG.mem_5_3 ), 
            .\REG.mem_4_3 (\REG.mem_4_3 ), .\REG.mem_40_1 (\REG.mem_40_1 ), 
            .\REG.mem_41_1 (\REG.mem_41_1 ), .\REG.mem_14_5 (\REG.mem_14_5 ), 
            .\REG.mem_15_5 (\REG.mem_15_5 ), .\REG.mem_13_5 (\REG.mem_13_5 ), 
            .\REG.mem_12_5 (\REG.mem_12_5 ), .\REG.mem_42_1 (\REG.mem_42_1 ), 
            .\REG.mem_43_1 (\REG.mem_43_1 ), .\REG.mem_46_1 (\REG.mem_46_1 ), 
            .\REG.mem_47_1 (\REG.mem_47_1 ), .\REG.mem_44_1 (\REG.mem_44_1 ), 
            .\REG.mem_45_1 (\REG.mem_45_1 ), .\REG.mem_31_8 (\REG.mem_31_8 ), 
            .\REG.mem_26_10 (\REG.mem_26_10 ), .\REG.mem_18_2 (\REG.mem_18_2 ), 
            .\REG.mem_19_2 (\REG.mem_19_2 ), .\REG.mem_31_3 (\REG.mem_31_3 ), 
            .\REG.mem_17_2 (\REG.mem_17_2 ), .\REG.mem_16_2 (\REG.mem_16_2 ), 
            .n61(n61), .\REG.mem_63_13 (\REG.mem_63_13 ), .n34(n34), .n29(n29), 
            .\REG.mem_50_6 (\REG.mem_50_6 ), .\REG.mem_51_6 (\REG.mem_51_6 ), 
            .n58(n58), .\REG.mem_6_14 (\REG.mem_6_14 ), .\REG.mem_7_14 (\REG.mem_7_14 ), 
            .n26(n26), .\REG.mem_6_10 (\REG.mem_6_10 ), .\REG.mem_7_10 (\REG.mem_7_10 ), 
            .\REG.mem_4_10 (\REG.mem_4_10 ), .\REG.mem_5_10 (\REG.mem_5_10 ), 
            .\REG.mem_4_14 (\REG.mem_4_14 ), .\REG.mem_5_14 (\REG.mem_5_14 ), 
            .n5896(n5896), .VCC_net(VCC_net), .\fifo_data_out[6] (\fifo_data_out[6] ), 
            .n5893(n5893), .\fifo_data_out[5] (\fifo_data_out[5] ), .\REG.mem_16_10 (\REG.mem_16_10 ), 
            .\REG.mem_17_10 (\REG.mem_17_10 ), .\REG.mem_18_10 (\REG.mem_18_10 ), 
            .\REG.mem_19_10 (\REG.mem_19_10 ), .n11119(n11119), .\fifo_data_out[7] (\fifo_data_out[7] ), 
            .\REG.mem_18_7 (\REG.mem_18_7 ), .\REG.mem_19_7 (\REG.mem_19_7 ), 
            .n11139(n11139), .\fifo_data_out[3] (\fifo_data_out[3] ), .\REG.mem_17_7 (\REG.mem_17_7 ), 
            .\REG.mem_16_7 (\REG.mem_16_7 ), .\REG.mem_50_2 (\REG.mem_50_2 ), 
            .\REG.mem_51_2 (\REG.mem_51_2 ), .\REG.mem_46_0 (\REG.mem_46_0 ), 
            .\REG.mem_47_0 (\REG.mem_47_0 ), .\REG.mem_46_9 (\REG.mem_46_9 ), 
            .\REG.mem_47_9 (\REG.mem_47_9 ), .\REG.mem_45_9 (\REG.mem_45_9 ), 
            .\REG.mem_44_9 (\REG.mem_44_9 ), .\REG.mem_49_6 (\REG.mem_49_6 ), 
            .\REG.mem_48_6 (\REG.mem_48_6 ), .\REG.mem_49_2 (\REG.mem_49_2 ), 
            .\REG.mem_48_2 (\REG.mem_48_2 ), .n11097(n11097), .\fifo_data_out[8] (\fifo_data_out[8] ), 
            .n5854(n5854), .\fifo_data_out[0] (\fifo_data_out[0] ), .\REG.mem_5_8 (\REG.mem_5_8 ), 
            .\REG.mem_4_8 (\REG.mem_4_8 ), .\REG.mem_6_11 (\REG.mem_6_11 ), 
            .\REG.mem_7_11 (\REG.mem_7_11 ), .\REG.mem_58_1 (\REG.mem_58_1 ), 
            .\REG.mem_26_15 (\REG.mem_26_15 ), .n11095(n11095), .\fifo_data_out[9] (\fifo_data_out[9] ), 
            .\REG.mem_23_7 (\REG.mem_23_7 ), .n11143(n11143), .\fifo_data_out[1] (\fifo_data_out[1] ), 
            .n11141(n11141), .\fifo_data_out[2] (\fifo_data_out[2] ), .n11089(n11089), 
            .\fifo_data_out[10] (\fifo_data_out[10] ), .n11135(n11135), 
            .\fifo_data_out[11] (\fifo_data_out[11] ), .\REG.mem_50_3 (\REG.mem_50_3 ), 
            .\REG.mem_51_3 (\REG.mem_51_3 ), .\REG.mem_31_13 (\REG.mem_31_13 ), 
            .\REG.mem_49_3 (\REG.mem_49_3 ), .\REG.mem_48_3 (\REG.mem_48_3 ), 
            .\REG.mem_10_9 (\REG.mem_10_9 ), .\REG.mem_11_9 (\REG.mem_11_9 ), 
            .\REG.mem_9_9 (\REG.mem_9_9 ), .\REG.mem_8_9 (\REG.mem_8_9 ), 
            .\REG.mem_23_10 (\REG.mem_23_10 ), .\REG.mem_26_1 (\REG.mem_26_1 ), 
            .n47(n47), .n5789(n5789), .\REG.mem_63_15 (\REG.mem_63_15 ), 
            .n5788(n5788), .\REG.mem_63_14 (\REG.mem_63_14 ), .n5787(n5787), 
            .\REG.mem_31_11 (\REG.mem_31_11 ), .\REG.mem_5_11 (\REG.mem_5_11 ), 
            .\REG.mem_4_11 (\REG.mem_4_11 ), .\REG.mem_31_1 (\REG.mem_31_1 ), 
            .\REG.mem_23_12 (\REG.mem_23_12 ), .n5786(n5786), .\REG.mem_63_12 (\REG.mem_63_12 ), 
            .n5785(n5785), .\REG.mem_63_11 (\REG.mem_63_11 ), .n5784(n5784), 
            .\REG.mem_63_10 (\REG.mem_63_10 ), .n5783(n5783), .\REG.mem_63_9 (\REG.mem_63_9 ), 
            .\REG.mem_14_9 (\REG.mem_14_9 ), .\REG.mem_15_9 (\REG.mem_15_9 ), 
            .n5782(n5782), .n5781(n5781), .\REG.mem_63_7 (\REG.mem_63_7 ), 
            .n5780(n5780), .\REG.mem_63_6 (\REG.mem_63_6 ), .n5779(n5779), 
            .\REG.mem_63_5 (\REG.mem_63_5 ), .n5778(n5778), .n5777(n5777), 
            .\REG.mem_63_3 (\REG.mem_63_3 ), .n5776(n5776), .\REG.mem_63_2 (\REG.mem_63_2 ), 
            .n5775(n5775), .\REG.mem_63_1 (\REG.mem_63_1 ), .n11133(n11133), 
            .\fifo_data_out[12] (\fifo_data_out[12] ), .n5773(n5773), .\REG.mem_63_0 (\REG.mem_63_0 ), 
            .\REG.mem_13_9 (\REG.mem_13_9 ), .\REG.mem_12_9 (\REG.mem_12_9 ), 
            .\REG.mem_38_10 (\REG.mem_38_10 ), .\REG.mem_39_10 (\REG.mem_39_10 ), 
            .n15(n15), .\REG.mem_36_10 (\REG.mem_36_10 ), .\REG.mem_37_10 (\REG.mem_37_10 ), 
            .\REG.mem_8_1 (\REG.mem_8_1 ), .\REG.mem_9_1 (\REG.mem_9_1 ), 
            .\REG.mem_10_1 (\REG.mem_10_1 ), .\REG.mem_11_1 (\REG.mem_11_1 ), 
            .n11137(n11137), .\fifo_data_out[4] (\fifo_data_out[4] ), .\REG.mem_14_1 (\REG.mem_14_1 ), 
            .\REG.mem_15_1 (\REG.mem_15_1 ), .\REG.mem_12_1 (\REG.mem_12_1 ), 
            .\REG.mem_13_1 (\REG.mem_13_1 ), .\REG.mem_38_12 (\REG.mem_38_12 ), 
            .\REG.mem_39_12 (\REG.mem_39_12 ), .\REG.mem_36_12 (\REG.mem_36_12 ), 
            .\REG.mem_37_12 (\REG.mem_37_12 ), .\REG.mem_38_5 (\REG.mem_38_5 ), 
            .\REG.mem_39_5 (\REG.mem_39_5 ), .n5709(n5709), .rp_sync1_r({rp_sync1_r}), 
            .n5708(n5708), .n5707(n5707), .n5706(n5706), .n5705(n5705), 
            .\REG.mem_36_5 (\REG.mem_36_5 ), .\REG.mem_37_5 (\REG.mem_37_5 ), 
            .\REG.mem_48_12 (\REG.mem_48_12 ), .\REG.mem_49_12 (\REG.mem_49_12 ), 
            .\wr_addr_r[0] (\wr_addr_r[0] ), .\REG.mem_50_12 (\REG.mem_50_12 ), 
            .\REG.mem_51_12 (\REG.mem_51_12 ), .\REG.mem_55_12 (\REG.mem_55_12 ), 
            .\wr_addr_p1_w[6] (\wr_addr_p1_w[6] ), .n5704(n5704), .\rd_sig_diff0_w[1] (\rd_sig_diff0_w[1] ), 
            .n5686(n5686), .n5685(n5685), .n5684(n5684), .n5683(n5683), 
            .n5682(n5682), .\REG.mem_58_15 (\REG.mem_58_15 ), .n5681(n5681), 
            .\REG.mem_58_14 (\REG.mem_58_14 ), .n5680(n5680), .n5679(n5679), 
            .\REG.mem_58_12 (\REG.mem_58_12 ), .n5678(n5678), .\REG.mem_58_11 (\REG.mem_58_11 ), 
            .n5677(n5677), .\REG.mem_58_10 (\REG.mem_58_10 ), .n5676(n5676), 
            .\REG.mem_58_9 (\REG.mem_58_9 ), .n5675(n5675), .n5674(n5674), 
            .\REG.mem_58_7 (\REG.mem_58_7 ), .n5673(n5673), .\REG.mem_58_6 (\REG.mem_58_6 ), 
            .\REG.mem_26_7 (\REG.mem_26_7 ), .\rd_sig_diff0_w[0] (\rd_sig_diff0_w[0] ), 
            .n5672(n5672), .n5671(n5671), .n5670(n5670), .\REG.mem_58_3 (\REG.mem_58_3 ), 
            .n5669(n5669), .\REG.mem_58_2 (\REG.mem_58_2 ), .n5668(n5668), 
            .n5667(n5667), .\REG.mem_58_0 (\REG.mem_58_0 ), .n5666(n5666), 
            .n5665(n5665), .n5664(n5664), .n5662(n5662), .n5660(n5660), 
            .\rd_addr_r[6] (\rd_addr_r[6] ), .\REG.out_raw[15] (\REG.out_raw[15] ), 
            .\REG.out_raw[14] (\REG.out_raw[14] ), .\REG.out_raw[13] (\REG.out_raw[13] ), 
            .\REG.out_raw[12] (\REG.out_raw[12] ), .\REG.out_raw[11] (\REG.out_raw[11] ), 
            .\REG.out_raw[10] (\REG.out_raw[10] ), .\REG.out_raw[9] (\REG.out_raw[9] ), 
            .\REG.out_raw[8] (\REG.out_raw[8] ), .\REG.out_raw[7] (\REG.out_raw[7] ), 
            .\REG.out_raw[6] (\REG.out_raw[6] ), .\REG.out_raw[5] (\REG.out_raw[5] ), 
            .\REG.out_raw[4] (\REG.out_raw[4] ), .\REG.out_raw[3] (\REG.out_raw[3] ), 
            .\REG.out_raw[2] (\REG.out_raw[2] ), .\REG.out_raw[1] (\REG.out_raw[1] ), 
            .\REG.mem_31_7 (\REG.mem_31_7 ), .\REG.mem_42_11 (\REG.mem_42_11 ), 
            .\REG.mem_43_11 (\REG.mem_43_11 ), .\REG.mem_41_11 (\REG.mem_41_11 ), 
            .\REG.mem_40_11 (\REG.mem_40_11 ), .n2(n2), .\REG.mem_6_1 (\REG.mem_6_1 ), 
            .\REG.mem_7_1 (\REG.mem_7_1 ), .\REG.mem_4_1 (\REG.mem_4_1 ), 
            .\REG.mem_5_1 (\REG.mem_5_1 ), .\REG.mem_38_4 (\REG.mem_38_4 ), 
            .\REG.mem_39_4 (\REG.mem_39_4 ), .\REG.mem_16_1 (\REG.mem_16_1 ), 
            .\REG.mem_17_1 (\REG.mem_17_1 ), .\REG.mem_37_4 (\REG.mem_37_4 ), 
            .\REG.mem_36_4 (\REG.mem_36_4 ), .\REG.mem_55_2 (\REG.mem_55_2 ), 
            .\REG.mem_18_1 (\REG.mem_18_1 ), .\REG.mem_19_1 (\REG.mem_19_1 ), 
            .n5626(n5626), .\REG.mem_55_15 (\REG.mem_55_15 ), .\REG.mem_23_1 (\REG.mem_23_1 ), 
            .\REG.mem_31_10 (\REG.mem_31_10 ), .n5625(n5625), .\REG.mem_55_14 (\REG.mem_55_14 ), 
            .n5624(n5624), .\REG.mem_55_13 (\REG.mem_55_13 ), .n5623(n5623), 
            .n5622(n5622), .n5621(n5621), .\REG.mem_55_10 (\REG.mem_55_10 ), 
            .n5620(n5620), .\REG.mem_55_9 (\REG.mem_55_9 ), .n5619(n5619), 
            .n5618(n5618), .\REG.mem_55_7 (\REG.mem_55_7 ), .n5617(n5617), 
            .\REG.mem_55_6 (\REG.mem_55_6 ), .n5616(n5616), .n5615(n5615), 
            .\REG.mem_55_4 (\REG.mem_55_4 ), .n5614(n5614), .\REG.mem_55_3 (\REG.mem_55_3 ), 
            .n5613(n5613), .n5612(n5612), .\REG.mem_55_1 (\REG.mem_55_1 ), 
            .n11073(n11073), .\fifo_data_out[13] (\fifo_data_out[13] ), 
            .n5610(n5610), .\REG.mem_55_0 (\REG.mem_55_0 ), .n5609(n5609), 
            .wp_sync1_r({wp_sync1_r}), .n5608(n5608), .n5607(n5607), .n5606(n5606), 
            .n5605(n5605), .n5604(n5604), .n5603(n5603), .n5586(n5586), 
            .n5585(n5585), .n5584(n5584), .n5583(n5583), .n5582(n5582), 
            .n11071(n11071), .\fifo_data_out[14] (\fifo_data_out[14] ), 
            .\REG.mem_38_1 (\REG.mem_38_1 ), .\REG.mem_39_1 (\REG.mem_39_1 ), 
            .\REG.mem_36_1 (\REG.mem_36_1 ), .\REG.mem_37_1 (\REG.mem_37_1 ), 
            .\REG.mem_6_2 (\REG.mem_6_2 ), .\REG.mem_7_2 (\REG.mem_7_2 ), 
            .\REG.mem_5_2 (\REG.mem_5_2 ), .\REG.mem_4_2 (\REG.mem_4_2 ), 
            .n5548(n5548), .\REG.mem_51_15 (\REG.mem_51_15 ), .n5547(n5547), 
            .\REG.mem_51_14 (\REG.mem_51_14 ), .n5546(n5546), .\REG.mem_51_13 (\REG.mem_51_13 ), 
            .n5545(n5545), .n5544(n5544), .\REG.mem_51_11 (\REG.mem_51_11 ), 
            .n5543(n5543), .\REG.mem_51_10 (\REG.mem_51_10 ), .n5542(n5542), 
            .\REG.mem_51_9 (\REG.mem_51_9 ), .n5541(n5541), .\REG.mem_51_8 (\REG.mem_51_8 ), 
            .n5540(n5540), .\REG.mem_51_7 (\REG.mem_51_7 ), .n5539(n5539), 
            .n5538(n5538), .n5537(n5537), .\REG.mem_51_4 (\REG.mem_51_4 ), 
            .n5536(n5536), .n5535(n5535), .n5534(n5534), .\REG.mem_51_1 (\REG.mem_51_1 ), 
            .n5533(n5533), .\REG.mem_51_0 (\REG.mem_51_0 ), .n5532(n5532), 
            .\REG.mem_50_15 (\REG.mem_50_15 ), .\REG.mem_48_1 (\REG.mem_48_1 ), 
            .\REG.mem_49_1 (\REG.mem_49_1 ), .n5531(n5531), .\REG.mem_50_14 (\REG.mem_50_14 ), 
            .n5530(n5530), .\REG.mem_50_13 (\REG.mem_50_13 ), .n5529(n5529), 
            .n5528(n5528), .\REG.mem_50_11 (\REG.mem_50_11 ), .n5527(n5527), 
            .\REG.mem_50_10 (\REG.mem_50_10 ), .n5526(n5526), .\REG.mem_50_9 (\REG.mem_50_9 ), 
            .n5525(n5525), .\REG.mem_50_8 (\REG.mem_50_8 ), .n5524(n5524), 
            .\REG.mem_50_7 (\REG.mem_50_7 ), .n5523(n5523), .n5522(n5522), 
            .n5521(n5521), .\REG.mem_50_4 (\REG.mem_50_4 ), .n5520(n5520), 
            .n5519(n5519), .n5518(n5518), .\REG.mem_50_1 (\REG.mem_50_1 ), 
            .n5517(n5517), .\REG.mem_50_0 (\REG.mem_50_0 ), .n5516(n5516), 
            .\REG.mem_49_15 (\REG.mem_49_15 ), .n5515(n5515), .\REG.mem_49_14 (\REG.mem_49_14 ), 
            .\REG.mem_31_12 (\REG.mem_31_12 ), .\REG.mem_26_11 (\REG.mem_26_11 ), 
            .n5514(n5514), .\REG.mem_49_13 (\REG.mem_49_13 ), .n5513(n5513), 
            .n5512(n5512), .\REG.mem_49_11 (\REG.mem_49_11 ), .n5511(n5511), 
            .\REG.mem_49_10 (\REG.mem_49_10 ), .n5510(n5510), .\REG.mem_49_9 (\REG.mem_49_9 ), 
            .n5509(n5509), .\REG.mem_49_8 (\REG.mem_49_8 ), .n5508(n5508), 
            .\REG.mem_49_7 (\REG.mem_49_7 ), .n5507(n5507), .n5506(n5506), 
            .n5505(n5505), .\REG.mem_49_4 (\REG.mem_49_4 ), .n5504(n5504), 
            .n5503(n5503), .n5502(n5502), .n5501(n5501), .\REG.mem_49_0 (\REG.mem_49_0 ), 
            .\REG.mem_31_0 (\REG.mem_31_0 ), .\REG.mem_26_4 (\REG.mem_26_4 ), 
            .n5492(n5492), .\REG.mem_48_15 (\REG.mem_48_15 ), .n5491(n5491), 
            .n5490(n5490), .\REG.mem_48_14 (\REG.mem_48_14 ), .n5489(n5489), 
            .\REG.mem_48_13 (\REG.mem_48_13 ), .n5488(n5488), .n5487(n5487), 
            .\REG.mem_48_11 (\REG.mem_48_11 ), .n5486(n5486), .\REG.mem_48_10 (\REG.mem_48_10 ), 
            .n5485(n5485), .\REG.mem_48_9 (\REG.mem_48_9 ), .n5484(n5484), 
            .\REG.mem_48_8 (\REG.mem_48_8 ), .n5483(n5483), .\REG.mem_48_7 (\REG.mem_48_7 ), 
            .\REG.mem_46_10 (\REG.mem_46_10 ), .\REG.mem_47_10 (\REG.mem_47_10 ), 
            .n5482(n5482), .n5481(n5481), .n5480(n5480), .\REG.mem_48_4 (\REG.mem_48_4 ), 
            .n5479(n5479), .n5478(n5478), .n5477(n5477), .n5476(n5476), 
            .\REG.mem_48_0 (\REG.mem_48_0 ), .n5474(n5474), .n5472(n5472), 
            .\REG.mem_47_15 (\REG.mem_47_15 ), .n5471(n5471), .\REG.mem_47_14 (\REG.mem_47_14 ), 
            .n5470(n5470), .\REG.mem_47_13 (\REG.mem_47_13 ), .n5469(n5469), 
            .\REG.mem_47_12 (\REG.mem_47_12 ), .n5468(n5468), .n5467(n5467), 
            .\REG.mem_45_0 (\REG.mem_45_0 ), .\REG.mem_44_0 (\REG.mem_44_0 ), 
            .\REG.mem_45_10 (\REG.mem_45_10 ), .\REG.mem_44_10 (\REG.mem_44_10 ), 
            .n5466(n5466), .n5465(n5465), .\REG.mem_47_8 (\REG.mem_47_8 ), 
            .n5464(n5464), .\REG.mem_47_7 (\REG.mem_47_7 ), .n5463(n5463), 
            .n5462(n5462), .\REG.mem_47_5 (\REG.mem_47_5 ), .n5461(n5461), 
            .\REG.mem_47_4 (\REG.mem_47_4 ), .n5460(n5460), .n5459(n5459), 
            .n5458(n5458), .n5457(n5457), .n5456(n5456), .\REG.mem_46_15 (\REG.mem_46_15 ), 
            .n5455(n5455), .\REG.mem_46_14 (\REG.mem_46_14 ), .n5454(n5454), 
            .\REG.mem_46_13 (\REG.mem_46_13 ), .n5453(n5453), .\REG.mem_46_12 (\REG.mem_46_12 ), 
            .n5452(n5452), .n5451(n5451), .n5450(n5450), .n5449(n5449), 
            .\REG.mem_46_8 (\REG.mem_46_8 ), .n5448(n5448), .\REG.mem_46_7 (\REG.mem_46_7 ), 
            .n5447(n5447), .n5446(n5446), .\REG.mem_46_5 (\REG.mem_46_5 ), 
            .n5445(n5445), .\REG.mem_46_4 (\REG.mem_46_4 ), .n5444(n5444), 
            .n5443(n5443), .n5442(n5442), .n5441(n5441), .n5440(n5440), 
            .\REG.mem_45_15 (\REG.mem_45_15 ), .n5439(n5439), .\REG.mem_45_14 (\REG.mem_45_14 ), 
            .n5438(n5438), .\REG.mem_45_13 (\REG.mem_45_13 ), .n5437(n5437), 
            .\REG.mem_45_12 (\REG.mem_45_12 ), .n5436(n5436), .n5435(n5435), 
            .n5434(n5434), .\REG.mem_38_7 (\REG.mem_38_7 ), .\REG.mem_39_7 (\REG.mem_39_7 ), 
            .\REG.mem_37_7 (\REG.mem_37_7 ), .\REG.mem_36_7 (\REG.mem_36_7 ), 
            .n5433(n5433), .\REG.mem_45_8 (\REG.mem_45_8 ), .n5432(n5432), 
            .\REG.mem_45_7 (\REG.mem_45_7 ), .n5431(n5431), .n5430(n5430), 
            .\REG.mem_45_5 (\REG.mem_45_5 ), .n5429(n5429), .\REG.mem_45_4 (\REG.mem_45_4 ), 
            .n5428(n5428), .n5427(n5427), .n5426(n5426), .n5425(n5425), 
            .n5424(n5424), .\REG.mem_44_15 (\REG.mem_44_15 ), .n5423(n5423), 
            .\REG.mem_44_14 (\REG.mem_44_14 ), .n5422(n5422), .\REG.mem_44_13 (\REG.mem_44_13 ), 
            .n5421(n5421), .\REG.mem_44_12 (\REG.mem_44_12 ), .n5420(n5420), 
            .n5419(n5419), .\REG.mem_10_0 (\REG.mem_10_0 ), .\REG.mem_11_0 (\REG.mem_11_0 ), 
            .n5418(n5418), .\REG.mem_9_0 (\REG.mem_9_0 ), .\REG.mem_8_0 (\REG.mem_8_0 ), 
            .n5417(n5417), .\REG.mem_44_8 (\REG.mem_44_8 ), .n5416(n5416), 
            .\REG.mem_44_7 (\REG.mem_44_7 ), .n5415(n5415), .n5414(n5414), 
            .\REG.mem_44_5 (\REG.mem_44_5 ), .n5413(n5413), .\REG.mem_44_4 (\REG.mem_44_4 ), 
            .n5412(n5412), .n5411(n5411), .n5410(n5410), .n5409(n5409), 
            .n5408(n5408), .n5407(n5407), .\REG.mem_43_15 (\REG.mem_43_15 ), 
            .n5406(n5406), .\REG.mem_43_14 (\REG.mem_43_14 ), .n5405(n5405), 
            .\REG.mem_43_13 (\REG.mem_43_13 ), .n5404(n5404), .\REG.mem_43_12 (\REG.mem_43_12 ), 
            .n5403(n5403), .n5402(n5402), .\REG.mem_10_5 (\REG.mem_10_5 ), 
            .\REG.mem_11_5 (\REG.mem_11_5 ), .\REG.mem_9_5 (\REG.mem_9_5 ), 
            .\REG.mem_8_5 (\REG.mem_8_5 ), .\wr_addr_p1_w[0] (\wr_addr_p1_w[0] ), 
            .n5401(n5401), .\REG.mem_43_9 (\REG.mem_43_9 ), .n5400(n5400), 
            .\REG.mem_43_8 (\REG.mem_43_8 ), .n5399(n5399), .\REG.mem_43_7 (\REG.mem_43_7 ), 
            .n5398(n5398), .\REG.mem_43_6 (\REG.mem_43_6 ), .n5397(n5397), 
            .\REG.mem_43_5 (\REG.mem_43_5 ), .n5396(n5396), .\REG.mem_43_4 (\REG.mem_43_4 ), 
            .n5395(n5395), .n5394(n5394), .n5393(n5393), .n5392(n5392), 
            .\REG.mem_43_0 (\REG.mem_43_0 ), .n11069(n11069), .\fifo_data_out[15] (\fifo_data_out[15] ), 
            .n5390(n5390), .\REG.mem_42_15 (\REG.mem_42_15 ), .n5389(n5389), 
            .\REG.mem_42_14 (\REG.mem_42_14 ), .n5388(n5388), .\REG.mem_42_13 (\REG.mem_42_13 ), 
            .n5387(n5387), .\REG.mem_42_12 (\REG.mem_42_12 ), .n5386(n5386), 
            .\REG.mem_42_4 (\REG.mem_42_4 ), .\REG.mem_41_4 (\REG.mem_41_4 ), 
            .\REG.mem_40_4 (\REG.mem_40_4 ), .n5385(n5385), .n5384(n5384), 
            .\REG.mem_42_9 (\REG.mem_42_9 ), .n5383(n5383), .\REG.mem_42_8 (\REG.mem_42_8 ), 
            .n5382(n5382), .\REG.mem_42_7 (\REG.mem_42_7 ), .n5381(n5381), 
            .\REG.mem_42_6 (\REG.mem_42_6 ), .n5380(n5380), .\REG.mem_42_5 (\REG.mem_42_5 ), 
            .n5379(n5379), .n5378(n5378), .n5377(n5377), .n5376(n5376), 
            .n5375(n5375), .\REG.mem_42_0 (\REG.mem_42_0 ), .n5374(n5374), 
            .\REG.mem_41_15 (\REG.mem_41_15 ), .n5373(n5373), .\REG.mem_41_14 (\REG.mem_41_14 ), 
            .n5372(n5372), .\REG.mem_41_13 (\REG.mem_41_13 ), .n5371(n5371), 
            .\REG.mem_41_12 (\REG.mem_41_12 ), .n4667(n4667), .n5370(n5370), 
            .n5369(n5369), .n5368(n5368), .\REG.mem_41_9 (\REG.mem_41_9 ), 
            .n5367(n5367), .\REG.mem_41_8 (\REG.mem_41_8 ), .n5366(n5366), 
            .\REG.mem_41_7 (\REG.mem_41_7 ), .n5365(n5365), .\REG.mem_41_6 (\REG.mem_41_6 ), 
            .n5364(n5364), .\REG.mem_41_5 (\REG.mem_41_5 ), .n5363(n5363), 
            .n5362(n5362), .n5361(n5361), .n5360(n5360), .n5358(n5358), 
            .\REG.mem_41_0 (\REG.mem_41_0 ), .n5357(n5357), .\REG.mem_40_15 (\REG.mem_40_15 ), 
            .n5356(n5356), .\REG.mem_40_14 (\REG.mem_40_14 ), .n5355(n5355), 
            .\REG.mem_40_13 (\REG.mem_40_13 ), .n5354(n5354), .\REG.mem_40_12 (\REG.mem_40_12 ), 
            .\REG.mem_38_13 (\REG.mem_38_13 ), .\REG.mem_39_13 (\REG.mem_39_13 ), 
            .\REG.mem_37_13 (\REG.mem_37_13 ), .\REG.mem_36_13 (\REG.mem_36_13 ), 
            .n5353(n5353), .n5352(n5352), .n5351(n5351), .\REG.mem_40_9 (\REG.mem_40_9 ), 
            .n5350(n5350), .\REG.mem_40_8 (\REG.mem_40_8 ), .n5349(n5349), 
            .\REG.mem_40_7 (\REG.mem_40_7 ), .n5348(n5348), .\REG.mem_40_6 (\REG.mem_40_6 ), 
            .n5347(n5347), .\REG.mem_40_5 (\REG.mem_40_5 ), .n5346(n5346), 
            .n5345(n5345), .n5344(n5344), .n5343(n5343), .n5342(n5342), 
            .\REG.mem_40_0 (\REG.mem_40_0 ), .n5341(n5341), .\REG.mem_39_15 (\REG.mem_39_15 ), 
            .n5340(n5340), .\REG.mem_39_14 (\REG.mem_39_14 ), .n5339(n5339), 
            .\REG.mem_23_5 (\REG.mem_23_5 ), .\REG.mem_14_0 (\REG.mem_14_0 ), 
            .\REG.mem_15_0 (\REG.mem_15_0 ), .\REG.mem_13_0 (\REG.mem_13_0 ), 
            .\REG.mem_12_0 (\REG.mem_12_0 ), .n5338(n5338), .n5337(n5337), 
            .n5336(n5336), .n5335(n5335), .\REG.mem_39_9 (\REG.mem_39_9 ), 
            .n5334(n5334), .\REG.mem_39_8 (\REG.mem_39_8 ), .n5333(n5333), 
            .n5332(n5332), .\REG.mem_39_6 (\REG.mem_39_6 ), .n5331(n5331), 
            .n5330(n5330), .n5329(n5329), .\REG.mem_39_3 (\REG.mem_39_3 ), 
            .n5328(n5328), .\REG.mem_39_2 (\REG.mem_39_2 ), .n5327(n5327), 
            .n5326(n5326), .\REG.mem_39_0 (\REG.mem_39_0 ), .n5323(n5323), 
            .\REG.mem_38_15 (\REG.mem_38_15 ), .n5322(n5322), .\REG.mem_38_14 (\REG.mem_38_14 ), 
            .n5321(n5321), .n5320(n5320), .n5319(n5319), .n5318(n5318), 
            .n5317(n5317), .\REG.mem_38_9 (\REG.mem_38_9 ), .n5316(n5316), 
            .\REG.mem_38_8 (\REG.mem_38_8 ), .n5315(n5315), .n5314(n5314), 
            .\REG.mem_38_6 (\REG.mem_38_6 ), .n5313(n5313), .n5312(n5312), 
            .n5311(n5311), .\REG.mem_38_3 (\REG.mem_38_3 ), .n5310(n5310), 
            .\REG.mem_38_2 (\REG.mem_38_2 ), .n5309(n5309), .n5308(n5308), 
            .\REG.mem_38_0 (\REG.mem_38_0 ), .n5302(n5302), .\REG.mem_37_15 (\REG.mem_37_15 ), 
            .n5301(n5301), .\REG.mem_37_14 (\REG.mem_37_14 ), .n5300(n5300), 
            .n5299(n5299), .n5298(n5298), .n5297(n5297), .n5296(n5296), 
            .\REG.mem_37_9 (\REG.mem_37_9 ), .n5295(n5295), .\REG.mem_37_8 (\REG.mem_37_8 ), 
            .n5294(n5294), .n5293(n5293), .\REG.mem_37_6 (\REG.mem_37_6 ), 
            .n5292(n5292), .n5291(n5291), .n5290(n5290), .\REG.mem_37_3 (\REG.mem_37_3 ), 
            .n5289(n5289), .\REG.mem_37_2 (\REG.mem_37_2 ), .n5288(n5288), 
            .n5286(n5286), .\REG.mem_37_0 (\REG.mem_37_0 ), .n5285(n5285), 
            .\REG.mem_36_15 (\REG.mem_36_15 ), .n5284(n5284), .\REG.mem_36_14 (\REG.mem_36_14 ), 
            .n5283(n5283), .n5282(n5282), .n5281(n5281), .n5280(n5280), 
            .n5279(n5279), .\REG.mem_36_9 (\REG.mem_36_9 ), .n5278(n5278), 
            .\REG.mem_36_8 (\REG.mem_36_8 ), .n5277(n5277), .n5276(n5276), 
            .\REG.mem_36_6 (\REG.mem_36_6 ), .n5275(n5275), .n5274(n5274), 
            .n5273(n5273), .\REG.mem_36_3 (\REG.mem_36_3 ), .n5272(n5272), 
            .\REG.mem_36_2 (\REG.mem_36_2 ), .n5271(n5271), .n5270(n5270), 
            .\REG.mem_36_0 (\REG.mem_36_0 ), .\REG.mem_26_12 (\REG.mem_26_12 ), 
            .\REG.mem_10_3 (\REG.mem_10_3 ), .\REG.mem_11_3 (\REG.mem_11_3 ), 
            .n5202(n5202), .\REG.mem_31_15 (\REG.mem_31_15 ), .n5201(n5201), 
            .n5200(n5200), .n5199(n5199), .n5198(n5198), .n5197(n5197), 
            .n5196(n5196), .\REG.mem_31_9 (\REG.mem_31_9 ), .n5195(n5195), 
            .n5194(n5194), .n5193(n5193), .\REG.mem_31_6 (\REG.mem_31_6 ), 
            .n5192(n5192), .\REG.mem_31_5 (\REG.mem_31_5 ), .n5191(n5191), 
            .\REG.mem_31_4 (\REG.mem_31_4 ), .n5190(n5190), .n5189(n5189), 
            .\REG.mem_31_2 (\REG.mem_31_2 ), .\REG.mem_9_3 (\REG.mem_9_3 ), 
            .\REG.mem_8_3 (\REG.mem_8_3 ), .n5188(n5188), .n5187(n5187), 
            .\REG.mem_10_14 (\REG.mem_10_14 ), .\REG.mem_11_14 (\REG.mem_11_14 ), 
            .\REG.mem_9_14 (\REG.mem_9_14 ), .\REG.mem_8_14 (\REG.mem_8_14 ), 
            .\REG.mem_23_2 (\REG.mem_23_2 ), .n5121(n5121), .n5120(n5120), 
            .n5119(n5119), .n5118(n5118), .n5117(n5117), .n5116(n5116), 
            .n5115(n5115), .\REG.mem_26_9 (\REG.mem_26_9 ), .n5114(n5114), 
            .n5113(n5113), .n5112(n5112), .\REG.mem_26_6 (\REG.mem_26_6 ), 
            .n5111(n5111), .\REG.mem_26_5 (\REG.mem_26_5 ), .n5110(n5110), 
            .n5109(n5109), .n5108(n5108), .\REG.mem_26_2 (\REG.mem_26_2 ), 
            .n5107(n5107), .n5106(n5106), .n5073(n5073), .n5072(n5072), 
            .\REG.mem_23_14 (\REG.mem_23_14 ), .n5071(n5071), .n5070(n5070), 
            .n5069(n5069), .n5068(n5068), .n5067(n5067), .\REG.mem_23_9 (\REG.mem_23_9 ), 
            .n5066(n5066), .\rd_grey_sync_r[5] (\rd_grey_sync_r[5] ), .\rd_grey_sync_r[4] (\rd_grey_sync_r[4] ), 
            .\REG.mem_10_6 (\REG.mem_10_6 ), .\REG.mem_11_6 (\REG.mem_11_6 ), 
            .\rd_grey_sync_r[3] (\rd_grey_sync_r[3] ), .\rd_grey_sync_r[2] (\rd_grey_sync_r[2] ), 
            .\rd_grey_sync_r[1] (\rd_grey_sync_r[1] ), .n5065(n5065), .n5064(n5064), 
            .\REG.mem_23_6 (\REG.mem_23_6 ), .n5063(n5063), .n5062(n5062), 
            .\REG.mem_23_4 (\REG.mem_23_4 ), .n5061(n5061), .\REG.mem_23_3 (\REG.mem_23_3 ), 
            .n5060(n5060), .n5059(n5059), .n5058(n5058), .\REG.mem_23_0 (\REG.mem_23_0 ), 
            .\REG.mem_9_6 (\REG.mem_9_6 ), .\REG.mem_8_6 (\REG.mem_8_6 ), 
            .n5(n5), .\REG.mem_14_6 (\REG.mem_14_6 ), .\REG.mem_15_6 (\REG.mem_15_6 ), 
            .\REG.mem_13_6 (\REG.mem_13_6 ), .\REG.mem_12_6 (\REG.mem_12_6 ), 
            .n5006(n5006), .\REG.mem_19_15 (\REG.mem_19_15 ), .n5005(n5005), 
            .\REG.mem_19_14 (\REG.mem_19_14 ), .n5004(n5004), .n5003(n5003), 
            .n5002(n5002), .\REG.mem_19_11 (\REG.mem_19_11 ), .n5001(n5001), 
            .n5000(n5000), .\REG.mem_19_9 (\REG.mem_19_9 ), .n4999(n4999), 
            .n4998(n4998), .n4997(n4997), .\REG.mem_19_6 (\REG.mem_19_6 ), 
            .n4996(n4996), .\REG.mem_19_5 (\REG.mem_19_5 ), .n4995(n4995), 
            .\REG.mem_19_4 (\REG.mem_19_4 ), .n4994(n4994), .\REG.mem_19_3 (\REG.mem_19_3 ), 
            .n4993(n4993), .n4992(n4992), .n4991(n4991), .\REG.mem_19_0 (\REG.mem_19_0 ), 
            .n4990(n4990), .\REG.mem_18_15 (\REG.mem_18_15 ), .n4989(n4989), 
            .\REG.mem_18_14 (\REG.mem_18_14 ), .n4988(n4988), .n4987(n4987), 
            .n4986(n4986), .\REG.mem_18_11 (\REG.mem_18_11 ), .n4985(n4985), 
            .n4984(n4984), .\REG.mem_18_9 (\REG.mem_18_9 ), .n4983(n4983), 
            .n4982(n4982), .n4981(n4981), .\REG.mem_18_6 (\REG.mem_18_6 ), 
            .n4980(n4980), .\REG.mem_18_5 (\REG.mem_18_5 ), .n4979(n4979), 
            .\REG.mem_18_4 (\REG.mem_18_4 ), .n4978(n4978), .\REG.mem_18_3 (\REG.mem_18_3 ), 
            .n4977(n4977), .n4976(n4976), .n4975(n4975), .\REG.mem_18_0 (\REG.mem_18_0 ), 
            .n4974(n4974), .\REG.mem_17_15 (\REG.mem_17_15 ), .n4973(n4973), 
            .\REG.mem_17_14 (\REG.mem_17_14 ), .n4972(n4972), .n4971(n4971), 
            .n4970(n4970), .\REG.mem_17_11 (\REG.mem_17_11 ), .n4969(n4969), 
            .n4968(n4968), .\REG.mem_17_9 (\REG.mem_17_9 ), .n4967(n4967), 
            .n4966(n4966), .n4965(n4965), .\REG.mem_17_6 (\REG.mem_17_6 ), 
            .n4964(n4964), .\REG.mem_17_5 (\REG.mem_17_5 ), .n4963(n4963), 
            .\REG.mem_17_4 (\REG.mem_17_4 ), .n4962(n4962), .\REG.mem_17_3 (\REG.mem_17_3 ), 
            .n4961(n4961), .n4960(n4960), .n4958(n4958), .\REG.mem_17_0 (\REG.mem_17_0 ), 
            .n4957(n4957), .\REG.mem_16_15 (\REG.mem_16_15 ), .n4956(n4956), 
            .\REG.mem_16_14 (\REG.mem_16_14 ), .n4955(n4955), .n4954(n4954), 
            .n4953(n4953), .\REG.mem_16_11 (\REG.mem_16_11 ), .n4952(n4952), 
            .n51(n51), .n4951(n4951), .\REG.mem_16_9 (\REG.mem_16_9 ), 
            .n4950(n4950), .n4949(n4949), .n4948(n4948), .\REG.mem_16_6 (\REG.mem_16_6 ), 
            .n4947(n4947), .\REG.mem_16_5 (\REG.mem_16_5 ), .n4946(n4946), 
            .\REG.mem_16_4 (\REG.mem_16_4 ), .n4945(n4945), .\REG.mem_16_3 (\REG.mem_16_3 ), 
            .n4944(n4944), .n4943(n4943), .n4942(n4942), .\REG.mem_16_0 (\REG.mem_16_0 ), 
            .n4941(n4941), .n4940(n4940), .\REG.mem_15_14 (\REG.mem_15_14 ), 
            .n4939(n4939), .n4938(n4938), .n4937(n4937), .\REG.mem_15_11 (\REG.mem_15_11 ), 
            .\rd_addr_nxt_c_6__N_465[5] (\rd_addr_nxt_c_6__N_465[5] ), .n19(n19), 
            .n4936(n4936), .n4935(n4935), .get_next_word(get_next_word), 
            .\rd_addr_nxt_c_6__N_465[3] (\rd_addr_nxt_c_6__N_465[3] ), .n4934(n4934), 
            .n4933(n4933), .n4932(n4932), .n4931(n4931), .n4930(n4930), 
            .\REG.mem_15_4 (\REG.mem_15_4 ), .n4929(n4929), .\REG.mem_15_3 (\REG.mem_15_3 ), 
            .n4928(n4928), .n4927(n4927), .n4926(n4926), .n4925(n4925), 
            .n4924(n4924), .\REG.mem_14_14 (\REG.mem_14_14 ), .n4923(n4923), 
            .n4922(n4922), .n4921(n4921), .\REG.mem_14_11 (\REG.mem_14_11 ), 
            .n4920(n4920), .n4919(n4919), .n4918(n4918), .\rd_addr_nxt_c_6__N_465[1] (\rd_addr_nxt_c_6__N_465[1] ), 
            .\state_timeout_counter[3] (\state_timeout_counter[3] ), .n718(n718), 
            .n7(n7), .n14424(n14424), .n4917(n4917), .n4916(n4916), 
            .n4915(n4915), .n4914(n4914), .\REG.mem_14_4 (\REG.mem_14_4 ), 
            .n4913(n4913), .\REG.mem_14_3 (\REG.mem_14_3 ), .n4912(n4912), 
            .n4911(n4911), .n4910(n4910), .\REG.mem_6_15 (\REG.mem_6_15 ), 
            .\REG.mem_7_15 (\REG.mem_7_15 ), .\REG.mem_5_15 (\REG.mem_5_15 ), 
            .\REG.mem_4_15 (\REG.mem_4_15 ), .\REG.mem_10_15 (\REG.mem_10_15 ), 
            .\REG.mem_11_15 (\REG.mem_11_15 ), .\REG.mem_9_15 (\REG.mem_9_15 ), 
            .\REG.mem_8_15 (\REG.mem_8_15 ), .n50(n50), .n52(n52), .n20(n20), 
            .n18(n18), .n4909(n4909), .n4908(n4908), .\REG.mem_13_14 (\REG.mem_13_14 ), 
            .n4907(n4907), .n4906(n4906), .n4905(n4905), .\REG.mem_13_11 (\REG.mem_13_11 ), 
            .n4904(n4904), .n4903(n4903), .n4902(n4902), .n4901(n4901), 
            .n46(n46), .n4900(n4900), .n4899(n4899), .n14(n14), .\REG.mem_10_11 (\REG.mem_10_11 ), 
            .\REG.mem_11_11 (\REG.mem_11_11 ), .n4898(n4898), .\REG.mem_13_4 (\REG.mem_13_4 ), 
            .n4897(n4897), .\REG.mem_13_3 (\REG.mem_13_3 ), .\REG.mem_9_11 (\REG.mem_9_11 ), 
            .\REG.mem_8_11 (\REG.mem_8_11 ), .\REG.mem_12_14 (\REG.mem_12_14 ), 
            .\REG.mem_12_11 (\REG.mem_12_11 ), .n4896(n4896), .n4895(n4895), 
            .n4894(n4894), .n4893(n4893), .n4892(n4892), .n53(n53), 
            .n4891(n4891), .n4890(n4890), .n21(n21), .n4889(n4889), 
            .n4888(n4888), .n4887(n4887), .n4886(n4886), .n4885(n4885), 
            .n4884(n4884), .n4883(n4883), .n4882(n4882), .\REG.mem_12_4 (\REG.mem_12_4 ), 
            .n4881(n4881), .\REG.mem_12_3 (\REG.mem_12_3 ), .n4880(n4880), 
            .n4879(n4879), .n4878(n4878), .n4646(n4646), .n4644(n4644), 
            .n4639(n4639), .n4877(n4877), .n4876(n4876), .n4875(n4875), 
            .n4874(n4874), .n4873(n4873), .n4872(n4872), .n4871(n4871), 
            .n4870(n4870), .\REG.mem_11_8 (\REG.mem_11_8 ), .n4869(n4869), 
            .n4638(n4638), .n4868(n4868), .n4867(n4867), .n4866(n4866), 
            .\REG.mem_11_4 (\REG.mem_11_4 ), .n4865(n4865), .n4864(n4864), 
            .n4863(n4863), .n4862(n4862), .n4861(n4861), .n4860(n4860), 
            .n4859(n4859), .n54(n54), .n22(n22), .n39(n39), .n7_adj_3(n7_adj_4), 
            .n4858(n4858), .n4857(n4857), .n4856(n4856), .n4855(n4855), 
            .n4854(n4854), .\REG.mem_10_8 (\REG.mem_10_8 ), .n4853(n4853), 
            .n4852(n4852), .n4851(n4851), .n56(n56), .n24(n24), .n4850(n4850), 
            .\REG.mem_10_4 (\REG.mem_10_4 ), .n4849(n4849), .n4848(n4848), 
            .n4847(n4847), .n4846(n4846), .n4845(n4845), .n4844(n4844), 
            .n4843(n4843), .n4842(n4842), .n4841(n4841), .n4840(n4840), 
            .n4839(n4839), .\afull_flag_impl.af_flag_p_w_N_603[3] (\afull_flag_impl.af_flag_p_w_N_603[3] ), 
            .n4838(n4838), .\REG.mem_9_8 (\REG.mem_9_8 ), .n4837(n4837), 
            .n4836(n4836), .n4835(n4835), .n4834(n4834), .\REG.mem_9_4 (\REG.mem_9_4 ), 
            .n4833(n4833), .n4832(n4832), .n4831(n4831), .n4830(n4830), 
            .n4829(n4829), .n4828(n4828), .n4827(n4827), .n4826(n4826), 
            .n4825(n4825), .n4824(n4824), .n4823(n4823), .n4822(n4822), 
            .\REG.mem_8_8 (\REG.mem_8_8 ), .n4821(n4821), .n4820(n4820), 
            .n4819(n4819), .n4818(n4818), .\REG.mem_8_4 (\REG.mem_8_4 ), 
            .n4817(n4817), .n4816(n4816), .n4815(n4815), .n4814(n4814), 
            .n4813(n4813), .n4812(n4812), .n4811(n4811), .\REG.mem_7_13 (\REG.mem_7_13 ), 
            .n4810(n4810), .n4809(n4809), .n4808(n4808), .n4807(n4807), 
            .\REG.mem_7_9 (\REG.mem_7_9 ), .n4806(n4806), .n4805(n4805), 
            .n4804(n4804), .\REG.mem_7_6 (\REG.mem_7_6 ), .n4803(n4803), 
            .\REG.mem_7_5 (\REG.mem_7_5 ), .n4802(n4802), .\REG.mem_7_4 (\REG.mem_7_4 ), 
            .n4801(n4801), .n4800(n4800), .n4799(n4799), .n4798(n4798), 
            .\REG.mem_7_0 (\REG.mem_7_0 ), .n4797(n4797), .n4796(n4796), 
            .n4795(n4795), .\REG.mem_6_13 (\REG.mem_6_13 ), .n4794(n4794), 
            .n4793(n4793), .n4792(n4792), .n4791(n4791), .\REG.mem_6_9 (\REG.mem_6_9 ), 
            .n4790(n4790), .n4789(n4789), .n4788(n4788), .\REG.mem_6_6 (\REG.mem_6_6 ), 
            .n4787(n4787), .\REG.mem_6_5 (\REG.mem_6_5 ), .n4786(n4786), 
            .\REG.mem_6_4 (\REG.mem_6_4 ), .n4785(n4785), .n4784(n4784), 
            .n4783(n4783), .n4779(n4779), .\REG.mem_6_0 (\REG.mem_6_0 ), 
            .n4778(n4778), .n4777(n4777), .n4776(n4776), .\REG.mem_5_13 (\REG.mem_5_13 ), 
            .n4775(n4775), .n4774(n4774), .n4773(n4773), .n4772(n4772), 
            .\REG.mem_5_9 (\REG.mem_5_9 ), .n4771(n4771), .n4770(n4770), 
            .n4769(n4769), .\REG.mem_5_6 (\REG.mem_5_6 ), .n4768(n4768), 
            .\REG.mem_5_5 (\REG.mem_5_5 ), .n4767(n4767), .\REG.mem_5_4 (\REG.mem_5_4 ), 
            .n4766(n4766), .n4765(n4765), .n4764(n4764), .n4763(n4763), 
            .\REG.mem_5_0 (\REG.mem_5_0 ), .n4762(n4762), .n4761(n4761), 
            .n4760(n4760), .\REG.mem_4_13 (\REG.mem_4_13 ), .n4759(n4759), 
            .n4758(n4758), .n4757(n4757), .n4756(n4756), .\REG.mem_4_9 (\REG.mem_4_9 ), 
            .n4755(n4755), .n4754(n4754), .n4753(n4753), .\REG.mem_4_6 (\REG.mem_4_6 ), 
            .n4752(n4752), .\REG.mem_4_5 (\REG.mem_4_5 ), .n4751(n4751), 
            .\REG.mem_4_4 (\REG.mem_4_4 ), .n4750(n4750), .n4749(n4749), 
            .n4748(n4748), .n4747(n4747), .\REG.mem_4_0 (\REG.mem_4_0 ), 
            .n4612(n4612), .n57(n57), .n25(n25), .n42(n42), .n10(n10), 
            .n49(n49), .n17(n17), .n48(n48), .n16(n16), .n55(n55), 
            .n23(n23), .n59(n59), .n27(n27)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_dc_32_lut_gen.v(53[33] 72[34])
    
endmodule
//
// Verilog Description of module fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1
//

module fifo_dc_32_lut_gen2_ipgen_lscc_fifo_dc_renamed_due_excessive_length_1 (\REG.mem_58_4 , 
            GND_net, \REG.mem_14_8 , \REG.mem_15_8 , \dc32_fifo_data_in[10] , 
            \dc32_fifo_data_in[9] , DEBUG_6_c_c, \REG.mem_13_8 , \REG.mem_12_8 , 
            \dc32_fifo_data_in[8] , \REG.mem_10_10 , \REG.mem_11_10 , 
            \REG.mem_9_10 , \REG.mem_8_10 , t_rd_fifo_en_w, \REG.out_raw[0] , 
            SLM_CLK_c, \dc32_fifo_data_in[7] , \REG.mem_10_13 , \REG.mem_11_13 , 
            \REG.mem_9_13 , \REG.mem_8_13 , \dc32_fifo_data_in[6] , DEBUG_9_c, 
            n7596, \wr_addr_nxt_c[4] , \REG.mem_26_14 , \dc32_fifo_data_in[5] , 
            \REG.mem_42_2 , \REG.mem_43_2 , \REG.mem_41_2 , \REG.mem_40_2 , 
            \REG.mem_14_10 , \REG.mem_15_10 , reset_all, \REG.mem_55_8 , 
            \REG.mem_13_10 , \REG.mem_12_10 , \dc32_fifo_data_in[4] , 
            \REG.mem_42_3 , \REG.mem_43_3 , \REG.mem_41_3 , \REG.mem_40_3 , 
            \rd_grey_sync_r[0] , \dc32_fifo_data_in[3] , \REG.mem_58_8 , 
            DEBUG_5_c, wr_grey_sync_r, \REG.mem_48_5 , \REG.mem_49_5 , 
            \aempty_flag_impl.ae_flag_nxt_w , dc32_fifo_almost_empty, \dc32_fifo_data_in[2] , 
            \REG.mem_55_11 , \REG.mem_50_5 , \REG.mem_51_5 , \dc32_fifo_data_in[1] , 
            \REG.mem_55_5 , \REG.mem_63_4 , \REG.mem_23_11 , \dc32_fifo_data_in[0] , 
            \REG.mem_10_12 , \REG.mem_11_12 , \REG.mem_9_12 , \REG.mem_8_12 , 
            \REG.mem_38_11 , \REG.mem_39_11 , \REG.mem_37_11 , \REG.mem_36_11 , 
            \REG.mem_14_12 , \REG.mem_15_12 , \REG.mem_14_13 , \REG.mem_15_13 , 
            \REG.mem_6_12 , \REG.mem_7_12 , \REG.mem_4_12 , \REG.mem_5_12 , 
            \REG.mem_13_13 , \REG.mem_12_13 , \REG.mem_13_12 , \REG.mem_12_12 , 
            \REG.mem_23_15 , \REG.mem_18_12 , \REG.mem_19_12 , \REG.mem_6_8 , 
            \REG.mem_7_8 , \REG.mem_17_12 , \REG.mem_16_12 , \wr_addr_nxt_c[2] , 
            \REG.mem_26_0 , \REG.mem_42_10 , \REG.mem_43_10 , \REG.mem_18_8 , 
            \REG.mem_19_8 , \REG.mem_14_15 , \REG.mem_15_15 , \REG.mem_17_8 , 
            \REG.mem_16_8 , \REG.mem_41_10 , \REG.mem_40_10 , n60, \REG.mem_18_13 , 
            \REG.mem_19_13 , \REG.mem_17_13 , \REG.mem_16_13 , n28, 
            \REG.mem_13_15 , \REG.mem_12_15 , \REG.mem_26_3 , \REG.mem_46_6 , 
            \REG.mem_47_6 , \REG.mem_45_6 , \REG.mem_44_6 , \REG.mem_63_8 , 
            \REG.mem_46_2 , \REG.mem_47_2 , \REG.mem_45_2 , \REG.mem_44_2 , 
            \dc32_fifo_data_in[15] , \dc32_fifo_data_in[14] , \REG.mem_6_7 , 
            \REG.mem_7_7 , \dc32_fifo_data_in[13] , \REG.mem_46_11 , \REG.mem_47_11 , 
            \dc32_fifo_data_in[12] , \REG.mem_5_7 , \REG.mem_4_7 , \dc32_fifo_data_in[11] , 
            \REG.mem_45_11 , \REG.mem_44_11 , \REG.mem_23_13 , \REG.mem_58_5 , 
            \REG.mem_23_8 , \REG.mem_46_3 , \REG.mem_47_3 , \REG.mem_10_7 , 
            \REG.mem_11_7 , \REG.mem_45_3 , \REG.mem_44_3 , \REG.mem_8_2 , 
            \REG.mem_9_2 , \REG.mem_9_7 , \REG.mem_8_7 , \REG.mem_31_14 , 
            \REG.mem_10_2 , \REG.mem_11_2 , \REG.mem_58_13 , \REG.mem_26_8 , 
            \REG.mem_14_2 , \REG.mem_15_2 , \REG.mem_12_2 , \REG.mem_13_2 , 
            \REG.mem_14_7 , \REG.mem_15_7 , \REG.mem_13_7 , \REG.mem_12_7 , 
            \REG.mem_26_13 , \REG.mem_6_3 , \REG.mem_7_3 , \REG.mem_5_3 , 
            \REG.mem_4_3 , \REG.mem_40_1 , \REG.mem_41_1 , \REG.mem_14_5 , 
            \REG.mem_15_5 , \REG.mem_13_5 , \REG.mem_12_5 , \REG.mem_42_1 , 
            \REG.mem_43_1 , \REG.mem_46_1 , \REG.mem_47_1 , \REG.mem_44_1 , 
            \REG.mem_45_1 , \REG.mem_31_8 , \REG.mem_26_10 , \REG.mem_18_2 , 
            \REG.mem_19_2 , \REG.mem_31_3 , \REG.mem_17_2 , \REG.mem_16_2 , 
            n61, \REG.mem_63_13 , n34, n29, \REG.mem_50_6 , \REG.mem_51_6 , 
            n58, \REG.mem_6_14 , \REG.mem_7_14 , n26, \REG.mem_6_10 , 
            \REG.mem_7_10 , \REG.mem_4_10 , \REG.mem_5_10 , \REG.mem_4_14 , 
            \REG.mem_5_14 , n5896, VCC_net, \fifo_data_out[6] , n5893, 
            \fifo_data_out[5] , \REG.mem_16_10 , \REG.mem_17_10 , \REG.mem_18_10 , 
            \REG.mem_19_10 , n11119, \fifo_data_out[7] , \REG.mem_18_7 , 
            \REG.mem_19_7 , n11139, \fifo_data_out[3] , \REG.mem_17_7 , 
            \REG.mem_16_7 , \REG.mem_50_2 , \REG.mem_51_2 , \REG.mem_46_0 , 
            \REG.mem_47_0 , \REG.mem_46_9 , \REG.mem_47_9 , \REG.mem_45_9 , 
            \REG.mem_44_9 , \REG.mem_49_6 , \REG.mem_48_6 , \REG.mem_49_2 , 
            \REG.mem_48_2 , n11097, \fifo_data_out[8] , n5854, \fifo_data_out[0] , 
            \REG.mem_5_8 , \REG.mem_4_8 , \REG.mem_6_11 , \REG.mem_7_11 , 
            \REG.mem_58_1 , \REG.mem_26_15 , n11095, \fifo_data_out[9] , 
            \REG.mem_23_7 , n11143, \fifo_data_out[1] , n11141, \fifo_data_out[2] , 
            n11089, \fifo_data_out[10] , n11135, \fifo_data_out[11] , 
            \REG.mem_50_3 , \REG.mem_51_3 , \REG.mem_31_13 , \REG.mem_49_3 , 
            \REG.mem_48_3 , \REG.mem_10_9 , \REG.mem_11_9 , \REG.mem_9_9 , 
            \REG.mem_8_9 , \REG.mem_23_10 , \REG.mem_26_1 , n47, n5789, 
            \REG.mem_63_15 , n5788, \REG.mem_63_14 , n5787, \REG.mem_31_11 , 
            \REG.mem_5_11 , \REG.mem_4_11 , \REG.mem_31_1 , \REG.mem_23_12 , 
            n5786, \REG.mem_63_12 , n5785, \REG.mem_63_11 , n5784, 
            \REG.mem_63_10 , n5783, \REG.mem_63_9 , \REG.mem_14_9 , 
            \REG.mem_15_9 , n5782, n5781, \REG.mem_63_7 , n5780, \REG.mem_63_6 , 
            n5779, \REG.mem_63_5 , n5778, n5777, \REG.mem_63_3 , n5776, 
            \REG.mem_63_2 , n5775, \REG.mem_63_1 , n11133, \fifo_data_out[12] , 
            n5773, \REG.mem_63_0 , \REG.mem_13_9 , \REG.mem_12_9 , \REG.mem_38_10 , 
            \REG.mem_39_10 , n15, \REG.mem_36_10 , \REG.mem_37_10 , 
            \REG.mem_8_1 , \REG.mem_9_1 , \REG.mem_10_1 , \REG.mem_11_1 , 
            n11137, \fifo_data_out[4] , \REG.mem_14_1 , \REG.mem_15_1 , 
            \REG.mem_12_1 , \REG.mem_13_1 , \REG.mem_38_12 , \REG.mem_39_12 , 
            \REG.mem_36_12 , \REG.mem_37_12 , \REG.mem_38_5 , \REG.mem_39_5 , 
            n5709, rp_sync1_r, n5708, n5707, n5706, n5705, \REG.mem_36_5 , 
            \REG.mem_37_5 , \REG.mem_48_12 , \REG.mem_49_12 , \wr_addr_r[0] , 
            \REG.mem_50_12 , \REG.mem_51_12 , \REG.mem_55_12 , \wr_addr_p1_w[6] , 
            n5704, \rd_sig_diff0_w[1] , n5686, n5685, n5684, n5683, 
            n5682, \REG.mem_58_15 , n5681, \REG.mem_58_14 , n5680, 
            n5679, \REG.mem_58_12 , n5678, \REG.mem_58_11 , n5677, 
            \REG.mem_58_10 , n5676, \REG.mem_58_9 , n5675, n5674, 
            \REG.mem_58_7 , n5673, \REG.mem_58_6 , \REG.mem_26_7 , \rd_sig_diff0_w[0] , 
            n5672, n5671, n5670, \REG.mem_58_3 , n5669, \REG.mem_58_2 , 
            n5668, n5667, \REG.mem_58_0 , n5666, n5665, n5664, n5662, 
            n5660, \rd_addr_r[6] , \REG.out_raw[15] , \REG.out_raw[14] , 
            \REG.out_raw[13] , \REG.out_raw[12] , \REG.out_raw[11] , \REG.out_raw[10] , 
            \REG.out_raw[9] , \REG.out_raw[8] , \REG.out_raw[7] , \REG.out_raw[6] , 
            \REG.out_raw[5] , \REG.out_raw[4] , \REG.out_raw[3] , \REG.out_raw[2] , 
            \REG.out_raw[1] , \REG.mem_31_7 , \REG.mem_42_11 , \REG.mem_43_11 , 
            \REG.mem_41_11 , \REG.mem_40_11 , n2, \REG.mem_6_1 , \REG.mem_7_1 , 
            \REG.mem_4_1 , \REG.mem_5_1 , \REG.mem_38_4 , \REG.mem_39_4 , 
            \REG.mem_16_1 , \REG.mem_17_1 , \REG.mem_37_4 , \REG.mem_36_4 , 
            \REG.mem_55_2 , \REG.mem_18_1 , \REG.mem_19_1 , n5626, \REG.mem_55_15 , 
            \REG.mem_23_1 , \REG.mem_31_10 , n5625, \REG.mem_55_14 , 
            n5624, \REG.mem_55_13 , n5623, n5622, n5621, \REG.mem_55_10 , 
            n5620, \REG.mem_55_9 , n5619, n5618, \REG.mem_55_7 , n5617, 
            \REG.mem_55_6 , n5616, n5615, \REG.mem_55_4 , n5614, \REG.mem_55_3 , 
            n5613, n5612, \REG.mem_55_1 , n11073, \fifo_data_out[13] , 
            n5610, \REG.mem_55_0 , n5609, wp_sync1_r, n5608, n5607, 
            n5606, n5605, n5604, n5603, n5586, n5585, n5584, n5583, 
            n5582, n11071, \fifo_data_out[14] , \REG.mem_38_1 , \REG.mem_39_1 , 
            \REG.mem_36_1 , \REG.mem_37_1 , \REG.mem_6_2 , \REG.mem_7_2 , 
            \REG.mem_5_2 , \REG.mem_4_2 , n5548, \REG.mem_51_15 , n5547, 
            \REG.mem_51_14 , n5546, \REG.mem_51_13 , n5545, n5544, 
            \REG.mem_51_11 , n5543, \REG.mem_51_10 , n5542, \REG.mem_51_9 , 
            n5541, \REG.mem_51_8 , n5540, \REG.mem_51_7 , n5539, n5538, 
            n5537, \REG.mem_51_4 , n5536, n5535, n5534, \REG.mem_51_1 , 
            n5533, \REG.mem_51_0 , n5532, \REG.mem_50_15 , \REG.mem_48_1 , 
            \REG.mem_49_1 , n5531, \REG.mem_50_14 , n5530, \REG.mem_50_13 , 
            n5529, n5528, \REG.mem_50_11 , n5527, \REG.mem_50_10 , 
            n5526, \REG.mem_50_9 , n5525, \REG.mem_50_8 , n5524, \REG.mem_50_7 , 
            n5523, n5522, n5521, \REG.mem_50_4 , n5520, n5519, n5518, 
            \REG.mem_50_1 , n5517, \REG.mem_50_0 , n5516, \REG.mem_49_15 , 
            n5515, \REG.mem_49_14 , \REG.mem_31_12 , \REG.mem_26_11 , 
            n5514, \REG.mem_49_13 , n5513, n5512, \REG.mem_49_11 , 
            n5511, \REG.mem_49_10 , n5510, \REG.mem_49_9 , n5509, 
            \REG.mem_49_8 , n5508, \REG.mem_49_7 , n5507, n5506, n5505, 
            \REG.mem_49_4 , n5504, n5503, n5502, n5501, \REG.mem_49_0 , 
            \REG.mem_31_0 , \REG.mem_26_4 , n5492, \REG.mem_48_15 , 
            n5491, n5490, \REG.mem_48_14 , n5489, \REG.mem_48_13 , 
            n5488, n5487, \REG.mem_48_11 , n5486, \REG.mem_48_10 , 
            n5485, \REG.mem_48_9 , n5484, \REG.mem_48_8 , n5483, \REG.mem_48_7 , 
            \REG.mem_46_10 , \REG.mem_47_10 , n5482, n5481, n5480, 
            \REG.mem_48_4 , n5479, n5478, n5477, n5476, \REG.mem_48_0 , 
            n5474, n5472, \REG.mem_47_15 , n5471, \REG.mem_47_14 , 
            n5470, \REG.mem_47_13 , n5469, \REG.mem_47_12 , n5468, 
            n5467, \REG.mem_45_0 , \REG.mem_44_0 , \REG.mem_45_10 , 
            \REG.mem_44_10 , n5466, n5465, \REG.mem_47_8 , n5464, 
            \REG.mem_47_7 , n5463, n5462, \REG.mem_47_5 , n5461, \REG.mem_47_4 , 
            n5460, n5459, n5458, n5457, n5456, \REG.mem_46_15 , 
            n5455, \REG.mem_46_14 , n5454, \REG.mem_46_13 , n5453, 
            \REG.mem_46_12 , n5452, n5451, n5450, n5449, \REG.mem_46_8 , 
            n5448, \REG.mem_46_7 , n5447, n5446, \REG.mem_46_5 , n5445, 
            \REG.mem_46_4 , n5444, n5443, n5442, n5441, n5440, \REG.mem_45_15 , 
            n5439, \REG.mem_45_14 , n5438, \REG.mem_45_13 , n5437, 
            \REG.mem_45_12 , n5436, n5435, n5434, \REG.mem_38_7 , 
            \REG.mem_39_7 , \REG.mem_37_7 , \REG.mem_36_7 , n5433, \REG.mem_45_8 , 
            n5432, \REG.mem_45_7 , n5431, n5430, \REG.mem_45_5 , n5429, 
            \REG.mem_45_4 , n5428, n5427, n5426, n5425, n5424, \REG.mem_44_15 , 
            n5423, \REG.mem_44_14 , n5422, \REG.mem_44_13 , n5421, 
            \REG.mem_44_12 , n5420, n5419, \REG.mem_10_0 , \REG.mem_11_0 , 
            n5418, \REG.mem_9_0 , \REG.mem_8_0 , n5417, \REG.mem_44_8 , 
            n5416, \REG.mem_44_7 , n5415, n5414, \REG.mem_44_5 , n5413, 
            \REG.mem_44_4 , n5412, n5411, n5410, n5409, n5408, n5407, 
            \REG.mem_43_15 , n5406, \REG.mem_43_14 , n5405, \REG.mem_43_13 , 
            n5404, \REG.mem_43_12 , n5403, n5402, \REG.mem_10_5 , 
            \REG.mem_11_5 , \REG.mem_9_5 , \REG.mem_8_5 , \wr_addr_p1_w[0] , 
            n5401, \REG.mem_43_9 , n5400, \REG.mem_43_8 , n5399, \REG.mem_43_7 , 
            n5398, \REG.mem_43_6 , n5397, \REG.mem_43_5 , n5396, \REG.mem_43_4 , 
            n5395, n5394, n5393, n5392, \REG.mem_43_0 , n11069, 
            \fifo_data_out[15] , n5390, \REG.mem_42_15 , n5389, \REG.mem_42_14 , 
            n5388, \REG.mem_42_13 , n5387, \REG.mem_42_12 , n5386, 
            \REG.mem_42_4 , \REG.mem_41_4 , \REG.mem_40_4 , n5385, n5384, 
            \REG.mem_42_9 , n5383, \REG.mem_42_8 , n5382, \REG.mem_42_7 , 
            n5381, \REG.mem_42_6 , n5380, \REG.mem_42_5 , n5379, n5378, 
            n5377, n5376, n5375, \REG.mem_42_0 , n5374, \REG.mem_41_15 , 
            n5373, \REG.mem_41_14 , n5372, \REG.mem_41_13 , n5371, 
            \REG.mem_41_12 , n4667, n5370, n5369, n5368, \REG.mem_41_9 , 
            n5367, \REG.mem_41_8 , n5366, \REG.mem_41_7 , n5365, \REG.mem_41_6 , 
            n5364, \REG.mem_41_5 , n5363, n5362, n5361, n5360, n5358, 
            \REG.mem_41_0 , n5357, \REG.mem_40_15 , n5356, \REG.mem_40_14 , 
            n5355, \REG.mem_40_13 , n5354, \REG.mem_40_12 , \REG.mem_38_13 , 
            \REG.mem_39_13 , \REG.mem_37_13 , \REG.mem_36_13 , n5353, 
            n5352, n5351, \REG.mem_40_9 , n5350, \REG.mem_40_8 , n5349, 
            \REG.mem_40_7 , n5348, \REG.mem_40_6 , n5347, \REG.mem_40_5 , 
            n5346, n5345, n5344, n5343, n5342, \REG.mem_40_0 , n5341, 
            \REG.mem_39_15 , n5340, \REG.mem_39_14 , n5339, \REG.mem_23_5 , 
            \REG.mem_14_0 , \REG.mem_15_0 , \REG.mem_13_0 , \REG.mem_12_0 , 
            n5338, n5337, n5336, n5335, \REG.mem_39_9 , n5334, \REG.mem_39_8 , 
            n5333, n5332, \REG.mem_39_6 , n5331, n5330, n5329, \REG.mem_39_3 , 
            n5328, \REG.mem_39_2 , n5327, n5326, \REG.mem_39_0 , n5323, 
            \REG.mem_38_15 , n5322, \REG.mem_38_14 , n5321, n5320, 
            n5319, n5318, n5317, \REG.mem_38_9 , n5316, \REG.mem_38_8 , 
            n5315, n5314, \REG.mem_38_6 , n5313, n5312, n5311, \REG.mem_38_3 , 
            n5310, \REG.mem_38_2 , n5309, n5308, \REG.mem_38_0 , n5302, 
            \REG.mem_37_15 , n5301, \REG.mem_37_14 , n5300, n5299, 
            n5298, n5297, n5296, \REG.mem_37_9 , n5295, \REG.mem_37_8 , 
            n5294, n5293, \REG.mem_37_6 , n5292, n5291, n5290, \REG.mem_37_3 , 
            n5289, \REG.mem_37_2 , n5288, n5286, \REG.mem_37_0 , n5285, 
            \REG.mem_36_15 , n5284, \REG.mem_36_14 , n5283, n5282, 
            n5281, n5280, n5279, \REG.mem_36_9 , n5278, \REG.mem_36_8 , 
            n5277, n5276, \REG.mem_36_6 , n5275, n5274, n5273, \REG.mem_36_3 , 
            n5272, \REG.mem_36_2 , n5271, n5270, \REG.mem_36_0 , \REG.mem_26_12 , 
            \REG.mem_10_3 , \REG.mem_11_3 , n5202, \REG.mem_31_15 , 
            n5201, n5200, n5199, n5198, n5197, n5196, \REG.mem_31_9 , 
            n5195, n5194, n5193, \REG.mem_31_6 , n5192, \REG.mem_31_5 , 
            n5191, \REG.mem_31_4 , n5190, n5189, \REG.mem_31_2 , \REG.mem_9_3 , 
            \REG.mem_8_3 , n5188, n5187, \REG.mem_10_14 , \REG.mem_11_14 , 
            \REG.mem_9_14 , \REG.mem_8_14 , \REG.mem_23_2 , n5121, n5120, 
            n5119, n5118, n5117, n5116, n5115, \REG.mem_26_9 , n5114, 
            n5113, n5112, \REG.mem_26_6 , n5111, \REG.mem_26_5 , n5110, 
            n5109, n5108, \REG.mem_26_2 , n5107, n5106, n5073, n5072, 
            \REG.mem_23_14 , n5071, n5070, n5069, n5068, n5067, 
            \REG.mem_23_9 , n5066, \rd_grey_sync_r[5] , \rd_grey_sync_r[4] , 
            \REG.mem_10_6 , \REG.mem_11_6 , \rd_grey_sync_r[3] , \rd_grey_sync_r[2] , 
            \rd_grey_sync_r[1] , n5065, n5064, \REG.mem_23_6 , n5063, 
            n5062, \REG.mem_23_4 , n5061, \REG.mem_23_3 , n5060, n5059, 
            n5058, \REG.mem_23_0 , \REG.mem_9_6 , \REG.mem_8_6 , n5, 
            \REG.mem_14_6 , \REG.mem_15_6 , \REG.mem_13_6 , \REG.mem_12_6 , 
            n5006, \REG.mem_19_15 , n5005, \REG.mem_19_14 , n5004, 
            n5003, n5002, \REG.mem_19_11 , n5001, n5000, \REG.mem_19_9 , 
            n4999, n4998, n4997, \REG.mem_19_6 , n4996, \REG.mem_19_5 , 
            n4995, \REG.mem_19_4 , n4994, \REG.mem_19_3 , n4993, n4992, 
            n4991, \REG.mem_19_0 , n4990, \REG.mem_18_15 , n4989, 
            \REG.mem_18_14 , n4988, n4987, n4986, \REG.mem_18_11 , 
            n4985, n4984, \REG.mem_18_9 , n4983, n4982, n4981, \REG.mem_18_6 , 
            n4980, \REG.mem_18_5 , n4979, \REG.mem_18_4 , n4978, \REG.mem_18_3 , 
            n4977, n4976, n4975, \REG.mem_18_0 , n4974, \REG.mem_17_15 , 
            n4973, \REG.mem_17_14 , n4972, n4971, n4970, \REG.mem_17_11 , 
            n4969, n4968, \REG.mem_17_9 , n4967, n4966, n4965, \REG.mem_17_6 , 
            n4964, \REG.mem_17_5 , n4963, \REG.mem_17_4 , n4962, \REG.mem_17_3 , 
            n4961, n4960, n4958, \REG.mem_17_0 , n4957, \REG.mem_16_15 , 
            n4956, \REG.mem_16_14 , n4955, n4954, n4953, \REG.mem_16_11 , 
            n4952, n51, n4951, \REG.mem_16_9 , n4950, n4949, n4948, 
            \REG.mem_16_6 , n4947, \REG.mem_16_5 , n4946, \REG.mem_16_4 , 
            n4945, \REG.mem_16_3 , n4944, n4943, n4942, \REG.mem_16_0 , 
            n4941, n4940, \REG.mem_15_14 , n4939, n4938, n4937, 
            \REG.mem_15_11 , \rd_addr_nxt_c_6__N_465[5] , n19, n4936, 
            n4935, get_next_word, \rd_addr_nxt_c_6__N_465[3] , n4934, 
            n4933, n4932, n4931, n4930, \REG.mem_15_4 , n4929, \REG.mem_15_3 , 
            n4928, n4927, n4926, n4925, n4924, \REG.mem_14_14 , 
            n4923, n4922, n4921, \REG.mem_14_11 , n4920, n4919, 
            n4918, \rd_addr_nxt_c_6__N_465[1] , \state_timeout_counter[3] , 
            n718, n7, n14424, n4917, n4916, n4915, n4914, \REG.mem_14_4 , 
            n4913, \REG.mem_14_3 , n4912, n4911, n4910, \REG.mem_6_15 , 
            \REG.mem_7_15 , \REG.mem_5_15 , \REG.mem_4_15 , \REG.mem_10_15 , 
            \REG.mem_11_15 , \REG.mem_9_15 , \REG.mem_8_15 , n50, n52, 
            n20, n18, n4909, n4908, \REG.mem_13_14 , n4907, n4906, 
            n4905, \REG.mem_13_11 , n4904, n4903, n4902, n4901, 
            n46, n4900, n4899, n14, \REG.mem_10_11 , \REG.mem_11_11 , 
            n4898, \REG.mem_13_4 , n4897, \REG.mem_13_3 , \REG.mem_9_11 , 
            \REG.mem_8_11 , \REG.mem_12_14 , \REG.mem_12_11 , n4896, 
            n4895, n4894, n4893, n4892, n53, n4891, n4890, n21, 
            n4889, n4888, n4887, n4886, n4885, n4884, n4883, n4882, 
            \REG.mem_12_4 , n4881, \REG.mem_12_3 , n4880, n4879, n4878, 
            n4646, n4644, n4639, n4877, n4876, n4875, n4874, n4873, 
            n4872, n4871, n4870, \REG.mem_11_8 , n4869, n4638, n4868, 
            n4867, n4866, \REG.mem_11_4 , n4865, n4864, n4863, n4862, 
            n4861, n4860, n4859, n54, n22, n39, n7_adj_3, n4858, 
            n4857, n4856, n4855, n4854, \REG.mem_10_8 , n4853, n4852, 
            n4851, n56, n24, n4850, \REG.mem_10_4 , n4849, n4848, 
            n4847, n4846, n4845, n4844, n4843, n4842, n4841, n4840, 
            n4839, \afull_flag_impl.af_flag_p_w_N_603[3] , n4838, \REG.mem_9_8 , 
            n4837, n4836, n4835, n4834, \REG.mem_9_4 , n4833, n4832, 
            n4831, n4830, n4829, n4828, n4827, n4826, n4825, n4824, 
            n4823, n4822, \REG.mem_8_8 , n4821, n4820, n4819, n4818, 
            \REG.mem_8_4 , n4817, n4816, n4815, n4814, n4813, n4812, 
            n4811, \REG.mem_7_13 , n4810, n4809, n4808, n4807, \REG.mem_7_9 , 
            n4806, n4805, n4804, \REG.mem_7_6 , n4803, \REG.mem_7_5 , 
            n4802, \REG.mem_7_4 , n4801, n4800, n4799, n4798, \REG.mem_7_0 , 
            n4797, n4796, n4795, \REG.mem_6_13 , n4794, n4793, n4792, 
            n4791, \REG.mem_6_9 , n4790, n4789, n4788, \REG.mem_6_6 , 
            n4787, \REG.mem_6_5 , n4786, \REG.mem_6_4 , n4785, n4784, 
            n4783, n4779, \REG.mem_6_0 , n4778, n4777, n4776, \REG.mem_5_13 , 
            n4775, n4774, n4773, n4772, \REG.mem_5_9 , n4771, n4770, 
            n4769, \REG.mem_5_6 , n4768, \REG.mem_5_5 , n4767, \REG.mem_5_4 , 
            n4766, n4765, n4764, n4763, \REG.mem_5_0 , n4762, n4761, 
            n4760, \REG.mem_4_13 , n4759, n4758, n4757, n4756, \REG.mem_4_9 , 
            n4755, n4754, n4753, \REG.mem_4_6 , n4752, \REG.mem_4_5 , 
            n4751, \REG.mem_4_4 , n4750, n4749, n4748, n4747, \REG.mem_4_0 , 
            n4612, n57, n25, n42, n10, n49, n17, n48, n16, 
            n55, n23, n59, n27) /* synthesis syn_module_defined=1 */ ;
    output \REG.mem_58_4 ;
    input GND_net;
    output \REG.mem_14_8 ;
    output \REG.mem_15_8 ;
    input \dc32_fifo_data_in[10] ;
    input \dc32_fifo_data_in[9] ;
    input DEBUG_6_c_c;
    output \REG.mem_13_8 ;
    output \REG.mem_12_8 ;
    input \dc32_fifo_data_in[8] ;
    output \REG.mem_10_10 ;
    output \REG.mem_11_10 ;
    output \REG.mem_9_10 ;
    output \REG.mem_8_10 ;
    output t_rd_fifo_en_w;
    output \REG.out_raw[0] ;
    input SLM_CLK_c;
    input \dc32_fifo_data_in[7] ;
    output \REG.mem_10_13 ;
    output \REG.mem_11_13 ;
    output \REG.mem_9_13 ;
    output \REG.mem_8_13 ;
    input \dc32_fifo_data_in[6] ;
    output DEBUG_9_c;
    output n7596;
    output \wr_addr_nxt_c[4] ;
    output \REG.mem_26_14 ;
    input \dc32_fifo_data_in[5] ;
    output \REG.mem_42_2 ;
    output \REG.mem_43_2 ;
    output \REG.mem_41_2 ;
    output \REG.mem_40_2 ;
    output \REG.mem_14_10 ;
    output \REG.mem_15_10 ;
    input reset_all;
    output \REG.mem_55_8 ;
    output \REG.mem_13_10 ;
    output \REG.mem_12_10 ;
    input \dc32_fifo_data_in[4] ;
    output \REG.mem_42_3 ;
    output \REG.mem_43_3 ;
    output \REG.mem_41_3 ;
    output \REG.mem_40_3 ;
    output \rd_grey_sync_r[0] ;
    input \dc32_fifo_data_in[3] ;
    output \REG.mem_58_8 ;
    output DEBUG_5_c;
    output [6:0]wr_grey_sync_r;
    output \REG.mem_48_5 ;
    output \REG.mem_49_5 ;
    input \aempty_flag_impl.ae_flag_nxt_w ;
    output dc32_fifo_almost_empty;
    input \dc32_fifo_data_in[2] ;
    output \REG.mem_55_11 ;
    output \REG.mem_50_5 ;
    output \REG.mem_51_5 ;
    input \dc32_fifo_data_in[1] ;
    output \REG.mem_55_5 ;
    output \REG.mem_63_4 ;
    output \REG.mem_23_11 ;
    input \dc32_fifo_data_in[0] ;
    output \REG.mem_10_12 ;
    output \REG.mem_11_12 ;
    output \REG.mem_9_12 ;
    output \REG.mem_8_12 ;
    output \REG.mem_38_11 ;
    output \REG.mem_39_11 ;
    output \REG.mem_37_11 ;
    output \REG.mem_36_11 ;
    output \REG.mem_14_12 ;
    output \REG.mem_15_12 ;
    output \REG.mem_14_13 ;
    output \REG.mem_15_13 ;
    output \REG.mem_6_12 ;
    output \REG.mem_7_12 ;
    output \REG.mem_4_12 ;
    output \REG.mem_5_12 ;
    output \REG.mem_13_13 ;
    output \REG.mem_12_13 ;
    output \REG.mem_13_12 ;
    output \REG.mem_12_12 ;
    output \REG.mem_23_15 ;
    output \REG.mem_18_12 ;
    output \REG.mem_19_12 ;
    output \REG.mem_6_8 ;
    output \REG.mem_7_8 ;
    output \REG.mem_17_12 ;
    output \REG.mem_16_12 ;
    output \wr_addr_nxt_c[2] ;
    output \REG.mem_26_0 ;
    output \REG.mem_42_10 ;
    output \REG.mem_43_10 ;
    output \REG.mem_18_8 ;
    output \REG.mem_19_8 ;
    output \REG.mem_14_15 ;
    output \REG.mem_15_15 ;
    output \REG.mem_17_8 ;
    output \REG.mem_16_8 ;
    output \REG.mem_41_10 ;
    output \REG.mem_40_10 ;
    output n60;
    output \REG.mem_18_13 ;
    output \REG.mem_19_13 ;
    output \REG.mem_17_13 ;
    output \REG.mem_16_13 ;
    output n28;
    output \REG.mem_13_15 ;
    output \REG.mem_12_15 ;
    output \REG.mem_26_3 ;
    output \REG.mem_46_6 ;
    output \REG.mem_47_6 ;
    output \REG.mem_45_6 ;
    output \REG.mem_44_6 ;
    output \REG.mem_63_8 ;
    output \REG.mem_46_2 ;
    output \REG.mem_47_2 ;
    output \REG.mem_45_2 ;
    output \REG.mem_44_2 ;
    input \dc32_fifo_data_in[15] ;
    input \dc32_fifo_data_in[14] ;
    output \REG.mem_6_7 ;
    output \REG.mem_7_7 ;
    input \dc32_fifo_data_in[13] ;
    output \REG.mem_46_11 ;
    output \REG.mem_47_11 ;
    input \dc32_fifo_data_in[12] ;
    output \REG.mem_5_7 ;
    output \REG.mem_4_7 ;
    input \dc32_fifo_data_in[11] ;
    output \REG.mem_45_11 ;
    output \REG.mem_44_11 ;
    output \REG.mem_23_13 ;
    output \REG.mem_58_5 ;
    output \REG.mem_23_8 ;
    output \REG.mem_46_3 ;
    output \REG.mem_47_3 ;
    output \REG.mem_10_7 ;
    output \REG.mem_11_7 ;
    output \REG.mem_45_3 ;
    output \REG.mem_44_3 ;
    output \REG.mem_8_2 ;
    output \REG.mem_9_2 ;
    output \REG.mem_9_7 ;
    output \REG.mem_8_7 ;
    output \REG.mem_31_14 ;
    output \REG.mem_10_2 ;
    output \REG.mem_11_2 ;
    output \REG.mem_58_13 ;
    output \REG.mem_26_8 ;
    output \REG.mem_14_2 ;
    output \REG.mem_15_2 ;
    output \REG.mem_12_2 ;
    output \REG.mem_13_2 ;
    output \REG.mem_14_7 ;
    output \REG.mem_15_7 ;
    output \REG.mem_13_7 ;
    output \REG.mem_12_7 ;
    output \REG.mem_26_13 ;
    output \REG.mem_6_3 ;
    output \REG.mem_7_3 ;
    output \REG.mem_5_3 ;
    output \REG.mem_4_3 ;
    output \REG.mem_40_1 ;
    output \REG.mem_41_1 ;
    output \REG.mem_14_5 ;
    output \REG.mem_15_5 ;
    output \REG.mem_13_5 ;
    output \REG.mem_12_5 ;
    output \REG.mem_42_1 ;
    output \REG.mem_43_1 ;
    output \REG.mem_46_1 ;
    output \REG.mem_47_1 ;
    output \REG.mem_44_1 ;
    output \REG.mem_45_1 ;
    output \REG.mem_31_8 ;
    output \REG.mem_26_10 ;
    output \REG.mem_18_2 ;
    output \REG.mem_19_2 ;
    output \REG.mem_31_3 ;
    output \REG.mem_17_2 ;
    output \REG.mem_16_2 ;
    output n61;
    output \REG.mem_63_13 ;
    output n34;
    output n29;
    output \REG.mem_50_6 ;
    output \REG.mem_51_6 ;
    output n58;
    output \REG.mem_6_14 ;
    output \REG.mem_7_14 ;
    output n26;
    output \REG.mem_6_10 ;
    output \REG.mem_7_10 ;
    output \REG.mem_4_10 ;
    output \REG.mem_5_10 ;
    output \REG.mem_4_14 ;
    output \REG.mem_5_14 ;
    input n5896;
    input VCC_net;
    output \fifo_data_out[6] ;
    input n5893;
    output \fifo_data_out[5] ;
    output \REG.mem_16_10 ;
    output \REG.mem_17_10 ;
    output \REG.mem_18_10 ;
    output \REG.mem_19_10 ;
    input n11119;
    output \fifo_data_out[7] ;
    output \REG.mem_18_7 ;
    output \REG.mem_19_7 ;
    input n11139;
    output \fifo_data_out[3] ;
    output \REG.mem_17_7 ;
    output \REG.mem_16_7 ;
    output \REG.mem_50_2 ;
    output \REG.mem_51_2 ;
    output \REG.mem_46_0 ;
    output \REG.mem_47_0 ;
    output \REG.mem_46_9 ;
    output \REG.mem_47_9 ;
    output \REG.mem_45_9 ;
    output \REG.mem_44_9 ;
    output \REG.mem_49_6 ;
    output \REG.mem_48_6 ;
    output \REG.mem_49_2 ;
    output \REG.mem_48_2 ;
    input n11097;
    output \fifo_data_out[8] ;
    input n5854;
    output \fifo_data_out[0] ;
    output \REG.mem_5_8 ;
    output \REG.mem_4_8 ;
    output \REG.mem_6_11 ;
    output \REG.mem_7_11 ;
    output \REG.mem_58_1 ;
    output \REG.mem_26_15 ;
    input n11095;
    output \fifo_data_out[9] ;
    output \REG.mem_23_7 ;
    input n11143;
    output \fifo_data_out[1] ;
    input n11141;
    output \fifo_data_out[2] ;
    input n11089;
    output \fifo_data_out[10] ;
    input n11135;
    output \fifo_data_out[11] ;
    output \REG.mem_50_3 ;
    output \REG.mem_51_3 ;
    output \REG.mem_31_13 ;
    output \REG.mem_49_3 ;
    output \REG.mem_48_3 ;
    output \REG.mem_10_9 ;
    output \REG.mem_11_9 ;
    output \REG.mem_9_9 ;
    output \REG.mem_8_9 ;
    output \REG.mem_23_10 ;
    output \REG.mem_26_1 ;
    output n47;
    input n5789;
    output \REG.mem_63_15 ;
    input n5788;
    output \REG.mem_63_14 ;
    input n5787;
    output \REG.mem_31_11 ;
    output \REG.mem_5_11 ;
    output \REG.mem_4_11 ;
    output \REG.mem_31_1 ;
    output \REG.mem_23_12 ;
    input n5786;
    output \REG.mem_63_12 ;
    input n5785;
    output \REG.mem_63_11 ;
    input n5784;
    output \REG.mem_63_10 ;
    input n5783;
    output \REG.mem_63_9 ;
    output \REG.mem_14_9 ;
    output \REG.mem_15_9 ;
    input n5782;
    input n5781;
    output \REG.mem_63_7 ;
    input n5780;
    output \REG.mem_63_6 ;
    input n5779;
    output \REG.mem_63_5 ;
    input n5778;
    input n5777;
    output \REG.mem_63_3 ;
    input n5776;
    output \REG.mem_63_2 ;
    input n5775;
    output \REG.mem_63_1 ;
    input n11133;
    output \fifo_data_out[12] ;
    input n5773;
    output \REG.mem_63_0 ;
    output \REG.mem_13_9 ;
    output \REG.mem_12_9 ;
    output \REG.mem_38_10 ;
    output \REG.mem_39_10 ;
    output n15;
    output \REG.mem_36_10 ;
    output \REG.mem_37_10 ;
    output \REG.mem_8_1 ;
    output \REG.mem_9_1 ;
    output \REG.mem_10_1 ;
    output \REG.mem_11_1 ;
    input n11137;
    output \fifo_data_out[4] ;
    output \REG.mem_14_1 ;
    output \REG.mem_15_1 ;
    output \REG.mem_12_1 ;
    output \REG.mem_13_1 ;
    output \REG.mem_38_12 ;
    output \REG.mem_39_12 ;
    output \REG.mem_36_12 ;
    output \REG.mem_37_12 ;
    output \REG.mem_38_5 ;
    output \REG.mem_39_5 ;
    input n5709;
    output [6:0]rp_sync1_r;
    input n5708;
    input n5707;
    input n5706;
    input n5705;
    output \REG.mem_36_5 ;
    output \REG.mem_37_5 ;
    output \REG.mem_48_12 ;
    output \REG.mem_49_12 ;
    output \wr_addr_r[0] ;
    output \REG.mem_50_12 ;
    output \REG.mem_51_12 ;
    output \REG.mem_55_12 ;
    output \wr_addr_p1_w[6] ;
    input n5704;
    output \rd_sig_diff0_w[1] ;
    input n5686;
    input n5685;
    input n5684;
    input n5683;
    input n5682;
    output \REG.mem_58_15 ;
    input n5681;
    output \REG.mem_58_14 ;
    input n5680;
    input n5679;
    output \REG.mem_58_12 ;
    input n5678;
    output \REG.mem_58_11 ;
    input n5677;
    output \REG.mem_58_10 ;
    input n5676;
    output \REG.mem_58_9 ;
    input n5675;
    input n5674;
    output \REG.mem_58_7 ;
    input n5673;
    output \REG.mem_58_6 ;
    output \REG.mem_26_7 ;
    output \rd_sig_diff0_w[0] ;
    input n5672;
    input n5671;
    input n5670;
    output \REG.mem_58_3 ;
    input n5669;
    output \REG.mem_58_2 ;
    input n5668;
    input n5667;
    output \REG.mem_58_0 ;
    input n5666;
    input n5665;
    input n5664;
    input n5662;
    input n5660;
    output \rd_addr_r[6] ;
    output \REG.out_raw[15] ;
    output \REG.out_raw[14] ;
    output \REG.out_raw[13] ;
    output \REG.out_raw[12] ;
    output \REG.out_raw[11] ;
    output \REG.out_raw[10] ;
    output \REG.out_raw[9] ;
    output \REG.out_raw[8] ;
    output \REG.out_raw[7] ;
    output \REG.out_raw[6] ;
    output \REG.out_raw[5] ;
    output \REG.out_raw[4] ;
    output \REG.out_raw[3] ;
    output \REG.out_raw[2] ;
    output \REG.out_raw[1] ;
    output \REG.mem_31_7 ;
    output \REG.mem_42_11 ;
    output \REG.mem_43_11 ;
    output \REG.mem_41_11 ;
    output \REG.mem_40_11 ;
    output n2;
    output \REG.mem_6_1 ;
    output \REG.mem_7_1 ;
    output \REG.mem_4_1 ;
    output \REG.mem_5_1 ;
    output \REG.mem_38_4 ;
    output \REG.mem_39_4 ;
    output \REG.mem_16_1 ;
    output \REG.mem_17_1 ;
    output \REG.mem_37_4 ;
    output \REG.mem_36_4 ;
    output \REG.mem_55_2 ;
    output \REG.mem_18_1 ;
    output \REG.mem_19_1 ;
    input n5626;
    output \REG.mem_55_15 ;
    output \REG.mem_23_1 ;
    output \REG.mem_31_10 ;
    input n5625;
    output \REG.mem_55_14 ;
    input n5624;
    output \REG.mem_55_13 ;
    input n5623;
    input n5622;
    input n5621;
    output \REG.mem_55_10 ;
    input n5620;
    output \REG.mem_55_9 ;
    input n5619;
    input n5618;
    output \REG.mem_55_7 ;
    input n5617;
    output \REG.mem_55_6 ;
    input n5616;
    input n5615;
    output \REG.mem_55_4 ;
    input n5614;
    output \REG.mem_55_3 ;
    input n5613;
    input n5612;
    output \REG.mem_55_1 ;
    input n11073;
    output \fifo_data_out[13] ;
    input n5610;
    output \REG.mem_55_0 ;
    input n5609;
    output [6:0]wp_sync1_r;
    input n5608;
    input n5607;
    input n5606;
    input n5605;
    input n5604;
    input n5603;
    input n5586;
    input n5585;
    input n5584;
    input n5583;
    input n5582;
    input n11071;
    output \fifo_data_out[14] ;
    output \REG.mem_38_1 ;
    output \REG.mem_39_1 ;
    output \REG.mem_36_1 ;
    output \REG.mem_37_1 ;
    output \REG.mem_6_2 ;
    output \REG.mem_7_2 ;
    output \REG.mem_5_2 ;
    output \REG.mem_4_2 ;
    input n5548;
    output \REG.mem_51_15 ;
    input n5547;
    output \REG.mem_51_14 ;
    input n5546;
    output \REG.mem_51_13 ;
    input n5545;
    input n5544;
    output \REG.mem_51_11 ;
    input n5543;
    output \REG.mem_51_10 ;
    input n5542;
    output \REG.mem_51_9 ;
    input n5541;
    output \REG.mem_51_8 ;
    input n5540;
    output \REG.mem_51_7 ;
    input n5539;
    input n5538;
    input n5537;
    output \REG.mem_51_4 ;
    input n5536;
    input n5535;
    input n5534;
    output \REG.mem_51_1 ;
    input n5533;
    output \REG.mem_51_0 ;
    input n5532;
    output \REG.mem_50_15 ;
    output \REG.mem_48_1 ;
    output \REG.mem_49_1 ;
    input n5531;
    output \REG.mem_50_14 ;
    input n5530;
    output \REG.mem_50_13 ;
    input n5529;
    input n5528;
    output \REG.mem_50_11 ;
    input n5527;
    output \REG.mem_50_10 ;
    input n5526;
    output \REG.mem_50_9 ;
    input n5525;
    output \REG.mem_50_8 ;
    input n5524;
    output \REG.mem_50_7 ;
    input n5523;
    input n5522;
    input n5521;
    output \REG.mem_50_4 ;
    input n5520;
    input n5519;
    input n5518;
    output \REG.mem_50_1 ;
    input n5517;
    output \REG.mem_50_0 ;
    input n5516;
    output \REG.mem_49_15 ;
    input n5515;
    output \REG.mem_49_14 ;
    output \REG.mem_31_12 ;
    output \REG.mem_26_11 ;
    input n5514;
    output \REG.mem_49_13 ;
    input n5513;
    input n5512;
    output \REG.mem_49_11 ;
    input n5511;
    output \REG.mem_49_10 ;
    input n5510;
    output \REG.mem_49_9 ;
    input n5509;
    output \REG.mem_49_8 ;
    input n5508;
    output \REG.mem_49_7 ;
    input n5507;
    input n5506;
    input n5505;
    output \REG.mem_49_4 ;
    input n5504;
    input n5503;
    input n5502;
    input n5501;
    output \REG.mem_49_0 ;
    output \REG.mem_31_0 ;
    output \REG.mem_26_4 ;
    input n5492;
    output \REG.mem_48_15 ;
    input n5491;
    input n5490;
    output \REG.mem_48_14 ;
    input n5489;
    output \REG.mem_48_13 ;
    input n5488;
    input n5487;
    output \REG.mem_48_11 ;
    input n5486;
    output \REG.mem_48_10 ;
    input n5485;
    output \REG.mem_48_9 ;
    input n5484;
    output \REG.mem_48_8 ;
    input n5483;
    output \REG.mem_48_7 ;
    output \REG.mem_46_10 ;
    output \REG.mem_47_10 ;
    input n5482;
    input n5481;
    input n5480;
    output \REG.mem_48_4 ;
    input n5479;
    input n5478;
    input n5477;
    input n5476;
    output \REG.mem_48_0 ;
    input n5474;
    input n5472;
    output \REG.mem_47_15 ;
    input n5471;
    output \REG.mem_47_14 ;
    input n5470;
    output \REG.mem_47_13 ;
    input n5469;
    output \REG.mem_47_12 ;
    input n5468;
    input n5467;
    output \REG.mem_45_0 ;
    output \REG.mem_44_0 ;
    output \REG.mem_45_10 ;
    output \REG.mem_44_10 ;
    input n5466;
    input n5465;
    output \REG.mem_47_8 ;
    input n5464;
    output \REG.mem_47_7 ;
    input n5463;
    input n5462;
    output \REG.mem_47_5 ;
    input n5461;
    output \REG.mem_47_4 ;
    input n5460;
    input n5459;
    input n5458;
    input n5457;
    input n5456;
    output \REG.mem_46_15 ;
    input n5455;
    output \REG.mem_46_14 ;
    input n5454;
    output \REG.mem_46_13 ;
    input n5453;
    output \REG.mem_46_12 ;
    input n5452;
    input n5451;
    input n5450;
    input n5449;
    output \REG.mem_46_8 ;
    input n5448;
    output \REG.mem_46_7 ;
    input n5447;
    input n5446;
    output \REG.mem_46_5 ;
    input n5445;
    output \REG.mem_46_4 ;
    input n5444;
    input n5443;
    input n5442;
    input n5441;
    input n5440;
    output \REG.mem_45_15 ;
    input n5439;
    output \REG.mem_45_14 ;
    input n5438;
    output \REG.mem_45_13 ;
    input n5437;
    output \REG.mem_45_12 ;
    input n5436;
    input n5435;
    input n5434;
    output \REG.mem_38_7 ;
    output \REG.mem_39_7 ;
    output \REG.mem_37_7 ;
    output \REG.mem_36_7 ;
    input n5433;
    output \REG.mem_45_8 ;
    input n5432;
    output \REG.mem_45_7 ;
    input n5431;
    input n5430;
    output \REG.mem_45_5 ;
    input n5429;
    output \REG.mem_45_4 ;
    input n5428;
    input n5427;
    input n5426;
    input n5425;
    input n5424;
    output \REG.mem_44_15 ;
    input n5423;
    output \REG.mem_44_14 ;
    input n5422;
    output \REG.mem_44_13 ;
    input n5421;
    output \REG.mem_44_12 ;
    input n5420;
    input n5419;
    output \REG.mem_10_0 ;
    output \REG.mem_11_0 ;
    input n5418;
    output \REG.mem_9_0 ;
    output \REG.mem_8_0 ;
    input n5417;
    output \REG.mem_44_8 ;
    input n5416;
    output \REG.mem_44_7 ;
    input n5415;
    input n5414;
    output \REG.mem_44_5 ;
    input n5413;
    output \REG.mem_44_4 ;
    input n5412;
    input n5411;
    input n5410;
    input n5409;
    input n5408;
    input n5407;
    output \REG.mem_43_15 ;
    input n5406;
    output \REG.mem_43_14 ;
    input n5405;
    output \REG.mem_43_13 ;
    input n5404;
    output \REG.mem_43_12 ;
    input n5403;
    input n5402;
    output \REG.mem_10_5 ;
    output \REG.mem_11_5 ;
    output \REG.mem_9_5 ;
    output \REG.mem_8_5 ;
    output \wr_addr_p1_w[0] ;
    input n5401;
    output \REG.mem_43_9 ;
    input n5400;
    output \REG.mem_43_8 ;
    input n5399;
    output \REG.mem_43_7 ;
    input n5398;
    output \REG.mem_43_6 ;
    input n5397;
    output \REG.mem_43_5 ;
    input n5396;
    output \REG.mem_43_4 ;
    input n5395;
    input n5394;
    input n5393;
    input n5392;
    output \REG.mem_43_0 ;
    input n11069;
    output \fifo_data_out[15] ;
    input n5390;
    output \REG.mem_42_15 ;
    input n5389;
    output \REG.mem_42_14 ;
    input n5388;
    output \REG.mem_42_13 ;
    input n5387;
    output \REG.mem_42_12 ;
    input n5386;
    output \REG.mem_42_4 ;
    output \REG.mem_41_4 ;
    output \REG.mem_40_4 ;
    input n5385;
    input n5384;
    output \REG.mem_42_9 ;
    input n5383;
    output \REG.mem_42_8 ;
    input n5382;
    output \REG.mem_42_7 ;
    input n5381;
    output \REG.mem_42_6 ;
    input n5380;
    output \REG.mem_42_5 ;
    input n5379;
    input n5378;
    input n5377;
    input n5376;
    input n5375;
    output \REG.mem_42_0 ;
    input n5374;
    output \REG.mem_41_15 ;
    input n5373;
    output \REG.mem_41_14 ;
    input n5372;
    output \REG.mem_41_13 ;
    input n5371;
    output \REG.mem_41_12 ;
    input n4667;
    input n5370;
    input n5369;
    input n5368;
    output \REG.mem_41_9 ;
    input n5367;
    output \REG.mem_41_8 ;
    input n5366;
    output \REG.mem_41_7 ;
    input n5365;
    output \REG.mem_41_6 ;
    input n5364;
    output \REG.mem_41_5 ;
    input n5363;
    input n5362;
    input n5361;
    input n5360;
    input n5358;
    output \REG.mem_41_0 ;
    input n5357;
    output \REG.mem_40_15 ;
    input n5356;
    output \REG.mem_40_14 ;
    input n5355;
    output \REG.mem_40_13 ;
    input n5354;
    output \REG.mem_40_12 ;
    output \REG.mem_38_13 ;
    output \REG.mem_39_13 ;
    output \REG.mem_37_13 ;
    output \REG.mem_36_13 ;
    input n5353;
    input n5352;
    input n5351;
    output \REG.mem_40_9 ;
    input n5350;
    output \REG.mem_40_8 ;
    input n5349;
    output \REG.mem_40_7 ;
    input n5348;
    output \REG.mem_40_6 ;
    input n5347;
    output \REG.mem_40_5 ;
    input n5346;
    input n5345;
    input n5344;
    input n5343;
    input n5342;
    output \REG.mem_40_0 ;
    input n5341;
    output \REG.mem_39_15 ;
    input n5340;
    output \REG.mem_39_14 ;
    input n5339;
    output \REG.mem_23_5 ;
    output \REG.mem_14_0 ;
    output \REG.mem_15_0 ;
    output \REG.mem_13_0 ;
    output \REG.mem_12_0 ;
    input n5338;
    input n5337;
    input n5336;
    input n5335;
    output \REG.mem_39_9 ;
    input n5334;
    output \REG.mem_39_8 ;
    input n5333;
    input n5332;
    output \REG.mem_39_6 ;
    input n5331;
    input n5330;
    input n5329;
    output \REG.mem_39_3 ;
    input n5328;
    output \REG.mem_39_2 ;
    input n5327;
    input n5326;
    output \REG.mem_39_0 ;
    input n5323;
    output \REG.mem_38_15 ;
    input n5322;
    output \REG.mem_38_14 ;
    input n5321;
    input n5320;
    input n5319;
    input n5318;
    input n5317;
    output \REG.mem_38_9 ;
    input n5316;
    output \REG.mem_38_8 ;
    input n5315;
    input n5314;
    output \REG.mem_38_6 ;
    input n5313;
    input n5312;
    input n5311;
    output \REG.mem_38_3 ;
    input n5310;
    output \REG.mem_38_2 ;
    input n5309;
    input n5308;
    output \REG.mem_38_0 ;
    input n5302;
    output \REG.mem_37_15 ;
    input n5301;
    output \REG.mem_37_14 ;
    input n5300;
    input n5299;
    input n5298;
    input n5297;
    input n5296;
    output \REG.mem_37_9 ;
    input n5295;
    output \REG.mem_37_8 ;
    input n5294;
    input n5293;
    output \REG.mem_37_6 ;
    input n5292;
    input n5291;
    input n5290;
    output \REG.mem_37_3 ;
    input n5289;
    output \REG.mem_37_2 ;
    input n5288;
    input n5286;
    output \REG.mem_37_0 ;
    input n5285;
    output \REG.mem_36_15 ;
    input n5284;
    output \REG.mem_36_14 ;
    input n5283;
    input n5282;
    input n5281;
    input n5280;
    input n5279;
    output \REG.mem_36_9 ;
    input n5278;
    output \REG.mem_36_8 ;
    input n5277;
    input n5276;
    output \REG.mem_36_6 ;
    input n5275;
    input n5274;
    input n5273;
    output \REG.mem_36_3 ;
    input n5272;
    output \REG.mem_36_2 ;
    input n5271;
    input n5270;
    output \REG.mem_36_0 ;
    output \REG.mem_26_12 ;
    output \REG.mem_10_3 ;
    output \REG.mem_11_3 ;
    input n5202;
    output \REG.mem_31_15 ;
    input n5201;
    input n5200;
    input n5199;
    input n5198;
    input n5197;
    input n5196;
    output \REG.mem_31_9 ;
    input n5195;
    input n5194;
    input n5193;
    output \REG.mem_31_6 ;
    input n5192;
    output \REG.mem_31_5 ;
    input n5191;
    output \REG.mem_31_4 ;
    input n5190;
    input n5189;
    output \REG.mem_31_2 ;
    output \REG.mem_9_3 ;
    output \REG.mem_8_3 ;
    input n5188;
    input n5187;
    output \REG.mem_10_14 ;
    output \REG.mem_11_14 ;
    output \REG.mem_9_14 ;
    output \REG.mem_8_14 ;
    output \REG.mem_23_2 ;
    input n5121;
    input n5120;
    input n5119;
    input n5118;
    input n5117;
    input n5116;
    input n5115;
    output \REG.mem_26_9 ;
    input n5114;
    input n5113;
    input n5112;
    output \REG.mem_26_6 ;
    input n5111;
    output \REG.mem_26_5 ;
    input n5110;
    input n5109;
    input n5108;
    output \REG.mem_26_2 ;
    input n5107;
    input n5106;
    input n5073;
    input n5072;
    output \REG.mem_23_14 ;
    input n5071;
    input n5070;
    input n5069;
    input n5068;
    input n5067;
    output \REG.mem_23_9 ;
    input n5066;
    output \rd_grey_sync_r[5] ;
    output \rd_grey_sync_r[4] ;
    output \REG.mem_10_6 ;
    output \REG.mem_11_6 ;
    output \rd_grey_sync_r[3] ;
    output \rd_grey_sync_r[2] ;
    output \rd_grey_sync_r[1] ;
    input n5065;
    input n5064;
    output \REG.mem_23_6 ;
    input n5063;
    input n5062;
    output \REG.mem_23_4 ;
    input n5061;
    output \REG.mem_23_3 ;
    input n5060;
    input n5059;
    input n5058;
    output \REG.mem_23_0 ;
    output \REG.mem_9_6 ;
    output \REG.mem_8_6 ;
    output n5;
    output \REG.mem_14_6 ;
    output \REG.mem_15_6 ;
    output \REG.mem_13_6 ;
    output \REG.mem_12_6 ;
    input n5006;
    output \REG.mem_19_15 ;
    input n5005;
    output \REG.mem_19_14 ;
    input n5004;
    input n5003;
    input n5002;
    output \REG.mem_19_11 ;
    input n5001;
    input n5000;
    output \REG.mem_19_9 ;
    input n4999;
    input n4998;
    input n4997;
    output \REG.mem_19_6 ;
    input n4996;
    output \REG.mem_19_5 ;
    input n4995;
    output \REG.mem_19_4 ;
    input n4994;
    output \REG.mem_19_3 ;
    input n4993;
    input n4992;
    input n4991;
    output \REG.mem_19_0 ;
    input n4990;
    output \REG.mem_18_15 ;
    input n4989;
    output \REG.mem_18_14 ;
    input n4988;
    input n4987;
    input n4986;
    output \REG.mem_18_11 ;
    input n4985;
    input n4984;
    output \REG.mem_18_9 ;
    input n4983;
    input n4982;
    input n4981;
    output \REG.mem_18_6 ;
    input n4980;
    output \REG.mem_18_5 ;
    input n4979;
    output \REG.mem_18_4 ;
    input n4978;
    output \REG.mem_18_3 ;
    input n4977;
    input n4976;
    input n4975;
    output \REG.mem_18_0 ;
    input n4974;
    output \REG.mem_17_15 ;
    input n4973;
    output \REG.mem_17_14 ;
    input n4972;
    input n4971;
    input n4970;
    output \REG.mem_17_11 ;
    input n4969;
    input n4968;
    output \REG.mem_17_9 ;
    input n4967;
    input n4966;
    input n4965;
    output \REG.mem_17_6 ;
    input n4964;
    output \REG.mem_17_5 ;
    input n4963;
    output \REG.mem_17_4 ;
    input n4962;
    output \REG.mem_17_3 ;
    input n4961;
    input n4960;
    input n4958;
    output \REG.mem_17_0 ;
    input n4957;
    output \REG.mem_16_15 ;
    input n4956;
    output \REG.mem_16_14 ;
    input n4955;
    input n4954;
    input n4953;
    output \REG.mem_16_11 ;
    input n4952;
    output n51;
    input n4951;
    output \REG.mem_16_9 ;
    input n4950;
    input n4949;
    input n4948;
    output \REG.mem_16_6 ;
    input n4947;
    output \REG.mem_16_5 ;
    input n4946;
    output \REG.mem_16_4 ;
    input n4945;
    output \REG.mem_16_3 ;
    input n4944;
    input n4943;
    input n4942;
    output \REG.mem_16_0 ;
    input n4941;
    input n4940;
    output \REG.mem_15_14 ;
    input n4939;
    input n4938;
    input n4937;
    output \REG.mem_15_11 ;
    output \rd_addr_nxt_c_6__N_465[5] ;
    output n19;
    input n4936;
    input n4935;
    input get_next_word;
    output \rd_addr_nxt_c_6__N_465[3] ;
    input n4934;
    input n4933;
    input n4932;
    input n4931;
    input n4930;
    output \REG.mem_15_4 ;
    input n4929;
    output \REG.mem_15_3 ;
    input n4928;
    input n4927;
    input n4926;
    input n4925;
    input n4924;
    output \REG.mem_14_14 ;
    input n4923;
    input n4922;
    input n4921;
    output \REG.mem_14_11 ;
    input n4920;
    input n4919;
    input n4918;
    output \rd_addr_nxt_c_6__N_465[1] ;
    input \state_timeout_counter[3] ;
    input n718;
    input n7;
    output n14424;
    input n4917;
    input n4916;
    input n4915;
    input n4914;
    output \REG.mem_14_4 ;
    input n4913;
    output \REG.mem_14_3 ;
    input n4912;
    input n4911;
    input n4910;
    output \REG.mem_6_15 ;
    output \REG.mem_7_15 ;
    output \REG.mem_5_15 ;
    output \REG.mem_4_15 ;
    output \REG.mem_10_15 ;
    output \REG.mem_11_15 ;
    output \REG.mem_9_15 ;
    output \REG.mem_8_15 ;
    output n50;
    output n52;
    output n20;
    output n18;
    input n4909;
    input n4908;
    output \REG.mem_13_14 ;
    input n4907;
    input n4906;
    input n4905;
    output \REG.mem_13_11 ;
    input n4904;
    input n4903;
    input n4902;
    input n4901;
    output n46;
    input n4900;
    input n4899;
    output n14;
    output \REG.mem_10_11 ;
    output \REG.mem_11_11 ;
    input n4898;
    output \REG.mem_13_4 ;
    input n4897;
    output \REG.mem_13_3 ;
    output \REG.mem_9_11 ;
    output \REG.mem_8_11 ;
    output \REG.mem_12_14 ;
    output \REG.mem_12_11 ;
    input n4896;
    input n4895;
    input n4894;
    input n4893;
    input n4892;
    output n53;
    input n4891;
    input n4890;
    output n21;
    input n4889;
    input n4888;
    input n4887;
    input n4886;
    input n4885;
    input n4884;
    input n4883;
    input n4882;
    output \REG.mem_12_4 ;
    input n4881;
    output \REG.mem_12_3 ;
    input n4880;
    input n4879;
    input n4878;
    input n4646;
    input n4644;
    input n4639;
    input n4877;
    input n4876;
    input n4875;
    input n4874;
    input n4873;
    input n4872;
    input n4871;
    input n4870;
    output \REG.mem_11_8 ;
    input n4869;
    input n4638;
    input n4868;
    input n4867;
    input n4866;
    output \REG.mem_11_4 ;
    input n4865;
    input n4864;
    input n4863;
    input n4862;
    input n4861;
    input n4860;
    input n4859;
    output n54;
    output n22;
    output n39;
    output n7_adj_3;
    input n4858;
    input n4857;
    input n4856;
    input n4855;
    input n4854;
    output \REG.mem_10_8 ;
    input n4853;
    input n4852;
    input n4851;
    output n56;
    output n24;
    input n4850;
    output \REG.mem_10_4 ;
    input n4849;
    input n4848;
    input n4847;
    input n4846;
    input n4845;
    input n4844;
    input n4843;
    input n4842;
    input n4841;
    input n4840;
    input n4839;
    input \afull_flag_impl.af_flag_p_w_N_603[3] ;
    input n4838;
    output \REG.mem_9_8 ;
    input n4837;
    input n4836;
    input n4835;
    input n4834;
    output \REG.mem_9_4 ;
    input n4833;
    input n4832;
    input n4831;
    input n4830;
    input n4829;
    input n4828;
    input n4827;
    input n4826;
    input n4825;
    input n4824;
    input n4823;
    input n4822;
    output \REG.mem_8_8 ;
    input n4821;
    input n4820;
    input n4819;
    input n4818;
    output \REG.mem_8_4 ;
    input n4817;
    input n4816;
    input n4815;
    input n4814;
    input n4813;
    input n4812;
    input n4811;
    output \REG.mem_7_13 ;
    input n4810;
    input n4809;
    input n4808;
    input n4807;
    output \REG.mem_7_9 ;
    input n4806;
    input n4805;
    input n4804;
    output \REG.mem_7_6 ;
    input n4803;
    output \REG.mem_7_5 ;
    input n4802;
    output \REG.mem_7_4 ;
    input n4801;
    input n4800;
    input n4799;
    input n4798;
    output \REG.mem_7_0 ;
    input n4797;
    input n4796;
    input n4795;
    output \REG.mem_6_13 ;
    input n4794;
    input n4793;
    input n4792;
    input n4791;
    output \REG.mem_6_9 ;
    input n4790;
    input n4789;
    input n4788;
    output \REG.mem_6_6 ;
    input n4787;
    output \REG.mem_6_5 ;
    input n4786;
    output \REG.mem_6_4 ;
    input n4785;
    input n4784;
    input n4783;
    input n4779;
    output \REG.mem_6_0 ;
    input n4778;
    input n4777;
    input n4776;
    output \REG.mem_5_13 ;
    input n4775;
    input n4774;
    input n4773;
    input n4772;
    output \REG.mem_5_9 ;
    input n4771;
    input n4770;
    input n4769;
    output \REG.mem_5_6 ;
    input n4768;
    output \REG.mem_5_5 ;
    input n4767;
    output \REG.mem_5_4 ;
    input n4766;
    input n4765;
    input n4764;
    input n4763;
    output \REG.mem_5_0 ;
    input n4762;
    input n4761;
    input n4760;
    output \REG.mem_4_13 ;
    input n4759;
    input n4758;
    input n4757;
    input n4756;
    output \REG.mem_4_9 ;
    input n4755;
    input n4754;
    input n4753;
    output \REG.mem_4_6 ;
    input n4752;
    output \REG.mem_4_5 ;
    input n4751;
    output \REG.mem_4_4 ;
    input n4750;
    input n4749;
    input n4748;
    input n4747;
    output \REG.mem_4_0 ;
    input n4612;
    output n57;
    output n25;
    output n42;
    output n10;
    output n49;
    output n17;
    output n48;
    output n16;
    output n55;
    output n23;
    output n59;
    output n27;
    
    wire DEBUG_6_c_c /* synthesis is_clock=1, SET_AS_NETWORK=DEBUG_6_c_c */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [6:0]rd_addr_r;   // src/fifo_dc_32_lut_gen.v(217[29:38])
    
    wire n11830, n11831, n13490, \REG.mem_59_4 , n14198, \REG.mem_57_4 , 
        \REG.mem_56_4 , n12066, n12405, n12420, n12794;
    wire [6:0]rd_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(221[30:42])
    
    wire n10640, n14192, n11792, n11791, n13493, n10641, n10639, 
        n42_c;
    wire [6:0]wr_addr_r;   // src/fifo_dc_32_lut_gen.v(196[29:38])
    
    wire \REG.mem_34_10 , n5248, n47_c, \REG.mem_53_9 , n5574, n12387, 
        n12375;
    wire [31:0]\REG.out_raw_31__N_526 ;
    
    wire n11674, n11675, n13484, n4729, \REG.mem_3_4 , n11648, n11647, 
        n13487, n11667, n12327, n12339, n12902, n11530, n11531, 
        n14186, n11510, n11509, n14189, \REG.mem_53_8 , n5573, n14180, 
        n14183, n12165, n12168, n13478, \REG.mem_53_7 , n5572, n14174, 
        n12075, n12150, n12144, n12282, \REG.mem_53_6 , n5571;
    wire [6:0]wr_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(212[30:44])
    
    wire n10784, n12276, n12255, n11436, n11463;
    wire [6:0]wr_addr_p1_w;   // src/fifo_dc_32_lut_gen.v(200[30:42])
    
    wire n4728, \REG.mem_3_3 , \REG.mem_27_14 , n13472, \REG.mem_53_5 , 
        n5570, n4727, \REG.mem_3_2 , \REG.mem_25_14 , \REG.mem_24_14 , 
        n13475, n14168, \REG.mem_34_9 , n5247, n12078, n12195, n12198, 
        n13466, n12180, n12177, n12288, n14162, \afull_flag_impl.af_flag_nxt_w , 
        n4726, \REG.mem_3_1 , \REG.mem_54_8 , n13460, \REG.mem_34_8 , 
        n5246, n4725, \REG.mem_3_0 , \REG.mem_34_7 , n5245, \REG.mem_52_8 , 
        n11853, n14165, \REG.mem_53_4 , n5569, n13454, n12013, n12014, 
        n14156, n13457, \REG.mem_34_6 , n5244;
    wire [6:0]rd_grey_w;   // src/fifo_dc_32_lut_gen.v(224[38:47])
    
    wire \REG.mem_53_3 , n5568, \REG.mem_34_5 , n5243, \REG.mem_34_4 , 
        n5242, n11999, n11998, n12080, n12043, n12044, n14150, 
        \REG.mem_59_8 , n13448, empty_nxt_c_N_596, n12035, n12034, 
        n12083, \REG.mem_57_8 , \REG.mem_56_8 , n11862;
    wire [6:0]wr_grey_w;   // src/fifo_dc_32_lut_gen.v(203[38:47])
    
    wire \REG.mem_34_3 , n5241, n12295, \REG.mem_53_2 , n5567, \REG.mem_54_11 , 
        n14144, n4723, \REG.mem_2_15 , n4722, \REG.mem_2_14 , n12240, 
        n12246, n13442, n12296, \REG.mem_53_11 , \REG.mem_52_11 , 
        n14147, n12183, n12162, \REG.mem_53_1 , n5566, \REG.mem_54_5 , 
        n12305, \REG.mem_52_5 , n12304, \REG.mem_62_4 , n14138, \REG.mem_22_11 , 
        n13436, \REG.mem_61_4 , \REG.mem_60_4 , n12093, \REG.mem_53_0 , 
        n5565, \REG.mem_0_12 , \REG.mem_1_12 , n12292, \REG.mem_21_11 , 
        \REG.mem_20_11 , n13439, \REG.mem_2_12 , \REG.mem_3_12 , n12293, 
        n13430, n13433, n12016, n12017, n14132, n12008, n12007, 
        n12098, n13424, n13427, \REG.mem_35_4 , n13418, \REG.mem_33_4 , 
        \REG.mem_32_4 , n13421, n4721, \REG.mem_2_13 , n13412, n14126, 
        n12299, n12298, n12102, full_nxt_c_N_593, full_o, n13415, 
        n4720, n4719, \REG.mem_2_11 , \REG.mem_22_15 , n12788, n13406, 
        n12824, n10627;
    wire [6:0]rp_sync_w;   // src/fifo_dc_32_lut_gen.v(205[30:39])
    
    wire n10628, \REG.mem_2_2 , n14120, n12312, n4718, \REG.mem_2_10 , 
        n4717, \REG.mem_2_9 , n4716, \REG.mem_2_8 , \REG.mem_1_2 , 
        \REG.mem_0_2 , n14123, n4715, \REG.mem_2_7 , n4714, \REG.mem_2_6 , 
        n13679, n14114, \REG.mem_27_0 , n13400, \REG.mem_25_0 , \REG.mem_24_0 , 
        n13403, n13673, n14117, n13394, n4713, \REG.mem_2_5 , n14108, 
        n12896, n11691, n13397, n15_c, n4712, \REG.mem_2_4 , n14102, 
        n4711, \REG.mem_2_3 , n12108, n12899, \REG.mem_27_3 , n14096, 
        n4710, n13388, n12315, n4709, \REG.mem_2_1 , n4708, \REG.mem_2_0 , 
        \REG.mem_25_3 , \REG.mem_24_3 , n14099, \REG.mem_62_8 , n13382, 
        \REG.mem_61_8 , \REG.mem_60_8 , n11874, n13355, n11747, n13376, 
        \REG.mem_3_7 , n14090, n11744, n13349, n13379, \REG.mem_1_7 , 
        \REG.mem_0_7 , n12111, n11844, n13370, n4707, \REG.mem_0_0 , 
        n14084, n11838, n11835, n13373, n12114, n11722, n11723, 
        n13364, n45, \REG.mem_52_15 , n5564, n13685, n14078, n11720, 
        n11719, n13367, n4706, \REG.mem_0_1 , n12095, n12094, n14081, 
        n11701, n11702, n13358, n11699, n11698, n13361, \REG.mem_52_14 , 
        n5563, n14072, n4705, n65, \REG.mem_30_4 , n5175, \REG.mem_52_13 , 
        n5562, n12890, n11680, n11681, n13352, n13817, n13667, 
        n11513, n11678, n11677, \REG.mem_34_2 , n5240, n13331, n11534, 
        \REG.mem_52_12 , n5561, n12120, n11656, n11657, n13346, 
        n5560, n12893, \REG.mem_22_13 , n14066, n11654, n11653, 
        \REG.mem_52_10 , n5559, \REG.mem_21_13 , \REG.mem_20_13 , n12123, 
        n4704, \REG.mem_0_3 , \REG.mem_59_5 , n13340, \REG.mem_57_5 , 
        \REG.mem_56_5 , n13343, \REG.mem_52_9 , n5558, \REG.mem_22_8 , 
        n14060, \REG.mem_34_1 , n5239, n5557, n10638, \REG.mem_34_0 , 
        n5238, \REG.mem_21_8 , \REG.mem_20_8 , n11709, n11643, n11670, 
        n14054, n13097, n11577, n13334, n14048, n13337, n11806, 
        n12126, \REG.mem_52_7 , n5556, \REG.mem_30_14 , n13328, \REG.mem_52_6 , 
        n5555, n11807, \REG.mem_29_14 , \REG.mem_28_14 , \REG.mem_59_13 , 
        n13322, \REG.mem_27_8 , n14042, \REG.mem_57_13 , \REG.mem_56_13 , 
        n11858, n12228, n12237, n13316, n11857, \REG.mem_25_8 , 
        \REG.mem_24_8 , n11718, n12222, n12210, n12330, n14036, 
        n5554, n12129, n12517, n12518, n13310, n12506, n12505, 
        n13313, \REG.mem_27_13 , n14030, \REG.mem_25_13 , \REG.mem_24_13 , 
        n12138, n12130, n12131, n12818, n11646, n13304, n14024, 
        n12827, n13073, n11880, n11559, \REG.mem_52_4 , n5553, \REG.mem_21_15 , 
        \REG.mem_20_15 , n12791, \REG.mem_52_3 , n5552, \REG.mem_52_2 , 
        n5551, \REG.mem_52_1 , n5550, \REG.mem_52_0 , n5549, n13265, 
        n11627, n13298, n11621, n13259, n13301, n13853, n14021, 
        n12500, n12481, n12482, n13292, n13, n13517, n12875, n12511, 
        n11704, n14018, n11705, n11714, n12476, n12475, n13295, 
        n11713, \REG.mem_30_8 , n14012, n13286, \REG.mem_29_8 , \REG.mem_28_8 , 
        n11736, n5025, \REG.mem_27_10 , n14006, n12258, \REG.mem_25_10 , 
        \REG.mem_24_10 , n14009, \REG.mem_20_14 , n5024, n13280, \REG.mem_30_3 , 
        n14000, n13283, \REG.mem_0_10 , \REG.mem_1_10 , n11524, \REG.mem_3_10 , 
        n11525, \REG.mem_29_3 , \REG.mem_28_3 , n14003, \REG.mem_62_13 , 
        n13274, n5023, \REG.mem_20_12 , n5022, \REG.mem_61_13 , \REG.mem_60_13 , 
        \REG.mem_0_14 , \REG.mem_1_14 , n12184, n35, n12782, n11671, 
        n11672, n13994, n11660, n11659, n11584, n11585, n13268, 
        n36, \REG.mem_3_14 , n12185, n11579, n11578, n13271, n12191, 
        n5021, n11528, n11527, n12190, n11695, n11696, n13988, 
        n11684, n11683, \REG.mem_20_10 , n5020, \REG.mem_20_9 , n5019, 
        n11545, n5018, \REG.mem_20_7 , n5017, \REG.mem_20_6 , n5016, 
        n11546, n11548, n11549, n13262, \REG.mem_20_5 , n5015, n13982, 
        n4702, \REG.mem_0_4 , n13976, \REG.mem_20_4 , n5014, \REG.mem_20_3 , 
        n5013, n12812, \REG.mem_20_2 , n5012, \REG.mem_20_1 , n5011, 
        n12800, n13256, n12803, n12785, n13979, \REG.mem_20_0 , 
        n5010, \REG.mem_56_1 , \REG.mem_57_1 , n11725, n12884, n13970, 
        \REG.mem_59_1 , n11726, n11750, n12512, n13250, n5041, \REG.mem_27_15 , 
        n12776, \REG.mem_21_14 , n5040, \REG.mem_22_7 , n13964, \REG.mem_21_7 , 
        n12499, n13253, n5039, n13244, \REG.mem_30_13 , n13958, 
        \REG.mem_29_13 , \REG.mem_28_13 , n12153, n13247, \REG.mem_21_12 , 
        n5038, n13238, n12347, n13232, n13235, n13193, n13226, 
        n13163, n13229, n5037, n13637, n13601, n13946, n13649, 
        n13661, n13949, \REG.mem_21_10 , n5036, \REG.mem_21_9 , n5035, 
        n13220, \REG.mem_22_10 , n13223, \REG.mem_24_1 , \REG.mem_25_1 , 
        \REG.mem_27_1 , n13214, n13217, n5034, n26_adj_1146, \REG.mem_30_11 , 
        n13940, n12887, n5033, \REG.mem_30_1 , \REG.mem_28_1 , \REG.mem_29_1 , 
        \REG.mem_22_12 , n13208, \REG.mem_21_6 , n5032, n12354, \REG.mem_21_5 , 
        n5031, \REG.mem_21_4 , n5030, \REG.mem_21_3 , n5029, n13202, 
        n5772, \REG.mem_62_15 , n5771, \REG.mem_62_14 , n5770, n5769, 
        \REG.mem_62_12 , n5768, \REG.mem_62_11 , n5767, \REG.mem_62_10 , 
        n5766, \REG.mem_62_9 , n5765, \REG.mem_21_2 , n5028, n5764, 
        \REG.mem_62_7 , n13205, n5763, \REG.mem_62_6 , n5762, \REG.mem_62_5 , 
        n5761, n5760, \REG.mem_62_3 , \REG.mem_29_11 , \REG.mem_28_11 , 
        n13943, n5759, \REG.mem_62_2 , n5758, \REG.mem_62_1 , n5757, 
        \REG.mem_62_0 , \REG.mem_21_1 , n5027, \REG.mem_21_0 , n5026, 
        n49_c, n5057, \REG.mem_22_14 , n5056, n12355, n12356, n13196, 
        \REG.mem_32_10 , \REG.mem_33_10 , \REG.mem_35_10 , n5749, \REG.mem_61_15 , 
        n5748, \REG.mem_61_14 , n5747, n5746, \REG.mem_61_12 , n5745, 
        \REG.mem_61_11 , n5744, \REG.mem_61_10 , n5743, \REG.mem_61_9 , 
        n5742, n5741, \REG.mem_61_7 , n5740, \REG.mem_61_6 , n5739, 
        \REG.mem_61_5 , n5738, n5737, \REG.mem_61_3 , n5055, n5054, 
        n12332, n12331, n13199;
    wire [6:0]rp_sync2_r;   // src/fifo_dc_32_lut_gen.v(202[37:47])
    wire [6:0]n1;
    
    wire n5053, n11638, n11639, n13934, n5052, n11552, n11551, 
        n13937, \REG.mem_22_9 , n5051, n11741, \REG.mem_60_1 , \REG.mem_61_1 , 
        n11740, n12271, n12272, n13190, \REG.mem_35_8 , n13928, 
        n5736, \REG.mem_61_2 , n5735, n5734, \REG.mem_61_0 , n5726, 
        \REG.mem_60_15 , n5724, \REG.mem_60_14 , n5723, n5722, \REG.mem_60_12 , 
        n5721, \REG.mem_60_11 , n5050, n5049, \REG.mem_32_12 , \REG.mem_33_12 , 
        \REG.mem_34_12 , \REG.mem_35_12 , \REG.mem_22_6 , n5048, \REG.mem_33_8 , 
        \REG.mem_32_8 , n11760, n10637, n10626, n10625, n13901, 
        n5720, \REG.mem_60_10 , n5719, \REG.mem_60_9 , n5718, n5717, 
        \REG.mem_60_7 , n5716, \REG.mem_60_6 , n5715, \REG.mem_60_5 , 
        n5714, n5713, \REG.mem_60_3 , n5712, \REG.mem_60_2 , n5711, 
        n5710, \REG.mem_60_0 , n6;
    wire [6:0]wp_sync2_r;   // src/fifo_dc_32_lut_gen.v(223[37:47])
    wire [6:0]n1_adj_1173;
    
    wire n10624;
    wire [6:0]rd_sig_diff0_w;   // src/fifo_dc_32_lut_gen.v(233[30:44])
    
    wire \REG.mem_22_5 , n5047, \REG.mem_54_12 , n7_c;
    wire [6:0]wp_sync_w;   // src/fifo_dc_32_lut_gen.v(226[30:39])
    
    wire n10623, \REG.mem_22_4 , n5046, n10636, \REG.mem_53_12 , n10622, 
        n10635, n5703, \REG.mem_59_15 , n5702, \REG.mem_59_14 , n5701, 
        n5700, \REG.mem_59_12 , n5699, \REG.mem_59_11 , n5698, \REG.mem_59_10 , 
        n5697, \REG.mem_59_9 , n5696, n5695, \REG.mem_59_7 , n5694, 
        \REG.mem_59_6 , n5693, n5692, n5691, \REG.mem_59_3 , n5690, 
        \REG.mem_59_2 , n5689, \REG.mem_22_3 , n5045, n8, n10621, 
        n10620, n10634, n11576, n12248, n12247, n14255, n10619, 
        n5688, \REG.mem_59_0 , \REG.mem_22_2 , n5044, \REG.mem_27_7 , 
        n13922, \REG.mem_22_1 , n5043, \REG.mem_25_7 , \REG.mem_24_7 , 
        n10633, \REG.mem_1_1 , n5663, n5661, n5659, n5658, \REG.mem_57_15 , 
        n10632, n5657, \REG.mem_57_14 , n5656, n5655, \REG.mem_57_12 , 
        n5654, \REG.mem_57_11 , n5653, \REG.mem_57_10 , n5652, \REG.mem_57_9 , 
        n5651, n5650, \REG.mem_57_7 , n5649, \REG.mem_57_6 , n5648, 
        n5647, n5646, \REG.mem_57_3 , n5645, \REG.mem_57_2 , n5644, 
        n5643, \REG.mem_57_0 , n5642, \REG.mem_56_15 , n5641, \REG.mem_56_14 , 
        \REG.mem_30_7 , n13916, n13184, n13187, \REG.mem_29_7 , \REG.mem_28_7 , 
        \REG.mem_22_0 , n5042, n13178, n13181, \REG.mem_54_2 , n13910, 
        n13913, n5640, n5639, \REG.mem_56_12 , n5638, \REG.mem_56_11 , 
        n5637, \REG.mem_56_10 , n5636, \REG.mem_56_9 , n5635, n5634, 
        \REG.mem_56_7 , n5633, \REG.mem_56_6 , n5632, n5631, n5630, 
        \REG.mem_56_3 , n5629, \REG.mem_56_2 , n5628, n5627, \REG.mem_56_0 , 
        \REG.mem_34_13 , \REG.mem_35_13 , n13904, \REG.mem_33_13 , \REG.mem_32_13 , 
        n12174, n12911, n11495, n13172, n11492, n12863, n13175, 
        \REG.mem_30_10 , n13898, n12460, n12461, n13166, n12446, 
        n12445, n13169, n4604, \REG.mem_29_10 , \REG.mem_28_10 , n53_c, 
        \REG.mem_24_15 , n5089, n5088, n5602, \REG.mem_54_15 , n5601, 
        \REG.mem_54_14 , n5600, \REG.mem_54_13 , n5599, n5598, n5597, 
        \REG.mem_54_10 , n5596, \REG.mem_54_9 , n5595, n5594, \REG.mem_54_7 , 
        n5593, \REG.mem_54_6 , n5592, n5591, \REG.mem_54_4 , n5590, 
        \REG.mem_54_3 , n5589, n5588, \REG.mem_54_1 , n5587, \REG.mem_54_0 , 
        \REG.mem_32_1 , \REG.mem_33_1 , n13892, \REG.mem_35_1 , n5580, 
        \REG.mem_53_15 , n5579, \REG.mem_53_14 , n5578, \REG.mem_53_13 , 
        n5577, n5576, n5575, \REG.mem_53_10 , n11765, n5087, \REG.mem_24_12 , 
        n5086, n13886, \REG.mem_24_11 , n5085, n13115, n13019, n13160, 
        n5084, n13889, n12941, n12815, n10631, n12453, n12456, 
        n13154, \REG.mem_24_9 , n5083, \REG.mem_35_7 , n13880, n12953, 
        n13157, \REG.mem_33_7 , \REG.mem_32_7 , n5082, \REG.mem_30_12 , 
        n12878, \REG.mem_27_11 , n13874, n5081, \REG.mem_25_11 , n13877, 
        \REG.mem_30_0 , n13148, \REG.mem_29_0 , \REG.mem_28_0 , n13151, 
        \REG.mem_24_6 , n5080, \REG.mem_29_12 , \REG.mem_28_12 , n12881, 
        n4691, \REG.mem_0_5 , \REG.mem_27_4 , n13868, n4690, \REG.mem_1_13 , 
        n4689, \REG.mem_0_6 , n5493, \REG.mem_24_5 , n5079, \REG.mem_24_4 , 
        n5078, n4688, n4687, \REG.mem_0_8 , n5077, n11598, n11625, 
        n12806, n13142, \REG.mem_24_2 , n5076, \REG.mem_25_4 , n13871, 
        n5475, n5473, n5075, n5074, n55_c, \REG.mem_25_15 , n5105, 
        n13145, n5104, n5103, \REG.mem_25_12 , n5102, n4684, \REG.mem_0_9 , 
        n4683, n4682, \REG.mem_0_11 , n4681, n4680, \REG.mem_0_13 , 
        n4678, n13136, n11898, n4675, n5101, n13862, n5100, \REG.mem_25_9 , 
        n5099, n11811, n11820, n13130, n11784, n11901, n5098, 
        n13124, n13856, n13859, n5097, \REG.mem_25_6 , n5096, n11, 
        n13127, n13850, n13118, \REG.mem_25_5 , n5095, n13121, n5094, 
        n4671, \REG.mem_0_15 , n5093, \REG.mem_25_2 , n5092, n5091, 
        n13844, \genblk16.rd_prev_r , n4666, n5090, n13847, n59_c, 
        n5138, n4665, \REG.mem_1_6 , n5137, n10630, n11475, n13838, 
        n12189, n5136, \REG.mem_27_12 , n5135, n5134, n5133, \REG.mem_35_0 , 
        n13112, \REG.mem_33_0 , \REG.mem_32_0 , n13031, n12983, n12872, 
        n13106, \REG.mem_27_9 , n5132, n13109, n13832, n5131, n13835, 
        n13100, n5130, n12372, n13826, \REG.mem_27_6 , n5129, n5269, 
        \REG.mem_35_15 , n5268, \REG.mem_35_14 , n5267, n5266, n5265, 
        \REG.mem_35_11 , n5264, n5263, \REG.mem_35_9 , n5262, n5261, 
        n5260, \REG.mem_35_6 , n5259, \REG.mem_35_5 , n5258, n5257, 
        \REG.mem_35_3 , n5256, \REG.mem_35_2 , n5255, n5254, n5253, 
        \REG.mem_34_15 , \REG.mem_27_5 , n5128, n13820, n5127, n5252, 
        \REG.mem_34_14 , n5251, n5250, n5249, \REG.mem_34_11 , n13094, 
        n5126, \REG.mem_27_2 , n5125, n5124, n5235, \REG.mem_33_15 , 
        n5234, \REG.mem_33_14 , n5233, n5232, n5231, \REG.mem_33_11 , 
        n5230, n5229, \REG.mem_33_9 , n5228, n5227, n5226, \REG.mem_33_6 , 
        n5225, \REG.mem_33_5 , n5224, n5223, \REG.mem_33_3 , n5222, 
        \REG.mem_33_2 , n5221, full_max_w, n11447, n11384, n12, 
        n5123, n5220, n5219, \REG.mem_32_15 , n5218, \REG.mem_32_14 , 
        n5217, n5216, n5215, \REG.mem_32_11 , n5214, n5213, \REG.mem_32_9 , 
        n5212, n5211, n5210, \REG.mem_32_6 , n5209, \REG.mem_32_5 , 
        n5208, n5207, \REG.mem_32_3 , n5206, \REG.mem_32_2 , n5205, 
        n61_adj_1154, \REG.mem_28_15 , n5154, n11402, n13088, n5153, 
        n11420, n10629, n5203, n12527, n5152, n11400, n11481, 
        n5151, n5186, \REG.mem_30_15 , n5185, n5184, n5183, n5182, 
        n5181, n5180, \REG.mem_30_9 , n5179, n5178, n5177, \REG.mem_30_6 , 
        n5176, \REG.mem_30_5 , n5174, n5150, n5149, \REG.mem_28_9 , 
        n5148, n5147, n5146, n13814, \REG.mem_28_6 , n5145, \REG.mem_28_5 , 
        n5144, \REG.mem_28_4 , n5143, n13082, n5173, \REG.mem_30_2 , 
        n5142, n11841, n11913, n5172, n5171, n5170, \REG.mem_29_15 , 
        n5169, n5168, n5167, n5166, n5165, n5164, \REG.mem_29_9 , 
        n5163, n5162, n5161, \REG.mem_29_6 , n5160, \REG.mem_29_5 , 
        n5159, \REG.mem_29_4 , n5158, n5157, \REG.mem_29_2 , n13076, 
        n12051, n12042, n13808, \REG.mem_28_2 , n5141, \REG.mem_3_8 , 
        n13070, n5140, n5139, n5156, n63, n5155, n13802, n12204, 
        \REG.mem_1_8 , n11755, n11756, n13796, n13064, n11663, n11662, 
        n13799, n13067, n12520, n12521, n13784, n13787, n13058, 
        n12515, n12514, n13739, n12182, n13052, n13055, n11523, 
        n12809, n13778, n13046, n13781, n13049, \REG.mem_3_15 , 
        n13040, \REG.mem_1_15 , n13043, n13772, n13775, n13034;
    wire [6:0]wr_addr_nxt_c;   // src/fifo_dc_32_lut_gen.v(198[29:42])
    
    wire n13028, n13022, n13760, n12947, n14411, n11498, n13013, 
        n13025, n14261, n13016, n14303, n13754, n14231, n13757, 
        n13631, n13691, n12376, n12377, n13010, n12346, n12474, 
        n11634, n13004, n12459, n13007, n12998, n13001, n12_adj_1156, 
        n16_c, n13748, n13751, n12992, n12995, n13742, n13745, 
        n12986, n13736, n12989, n17_c, n4027, n11445, n11408, 
        rd_fifo_en_w, n11430, n12980, n12866, n12869, n13730, n12343, 
        n12344, n12860, n12341, n12340, n13733, n4025, n10_c, 
        n8_adj_1157, n12_adj_1158, n11483, n10760, n12974, n12977, 
        n12225, n12968, n13724, n4648, n13718, n12962, n12965, 
        n12956, n12959, n13712, \REG.mem_3_11 , n12950, \REG.mem_1_11 , 
        n12944, n12067, n12068, n13706, n12057, n12030, n12038, 
        n13565, n13709, n12938, n12932, n13700, n12935, n12926, 
        n12929, n12920, n12923, n12070, n12071, n13688, n12059, 
        n12058, n12914, n12917, n12382, n12383, n12908, n12362, 
        n12361, n44, n12854, n11983, n11984, n13682, n11972, n11971, 
        n4741, n4739, \REG.mem_3_13 , n4738, n4737, n4736, n4735, 
        \REG.mem_3_9 , n4734, n4733, n4732, \REG.mem_3_6 , n4731, 
        \REG.mem_3_5 , n4730, n12031, n12032, n13676, n12020, n12019, 
        n13607, n14408, n20_adj_1160, n11995, n11996, n13670, n11987, 
        n11986, n12779, n14402, n13664, n14396, n13658, n12830, 
        n14390, n13652, n14384, n13646, n14387, n12857, n14378, 
        n4647, n4645, n4643, n4642, n4641, n4640, \REG.mem_1_3 , 
        n12471, n4636, n14372, n13640, n13634, n14366, n12480, 
        n14360, n14363, n11572, n11573, n13628, n11543, n25_c, 
        n14354, n12486, n13622, n14348, n12006, n14342, n12003, 
        n13616, n13619, n14336, n13610, n12848, n12054, n12012, 
        n13604, n12851, n12466, n12467, n14330, n12464, n12463, 
        n11516, n14324, n13598, n40, n14207, n12498, n12833, n13592, 
        n14318, n11991, n14312, n4614, \REG.mem_1_0 , n9, n11976, 
        n13586, n7612, n13589, n13580, n4613, \REG.mem_1_4 , n14306, 
        n14300, n12842, n11501, n11500, n13574, n14294, n4610, 
        \REG.mem_1_9 , n13577, n14288, n13568, n12845, n11761, n11762, 
        n13562, n12025, n12026, n14282, n4608, \REG.mem_1_5 , n11732, 
        n11731, n11981, n11980, n12836, n11506, n11507, n14276, 
        n12509, n12508, n14270, n13550, n14273, n3_adj_1166, n7616, 
        n12839, n12089, n12088, n12821, n14264, n11555, n14258, 
        n11489, n12493, n12494, n14252, n12488, n12487, n14246, 
        n13532, n14240, n11788, n11789, n13526, n10642, n11786, 
        n11785, n13529, n11635, n11636, n14228, n11630, n14222, 
        n13520, n13514, n14216, n13508, n13502, n14210, n13505, 
        n14204, n12002, n11990, n11975, n6_adj_1172;
    
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11749 (.I0(rd_addr_r[1]), .I1(n11830), 
            .I2(n11831), .I3(rd_addr_r[2]), .O(n13490));
    defparam rd_addr_r_1__bdd_4_lut_11749.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12313 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_4 ), 
            .I2(\REG.mem_59_4 ), .I3(rd_addr_r[1]), .O(n14198));
    defparam rd_addr_r_0__bdd_4_lut_12313.LUT_INIT = 16'he4aa;
    SB_LUT4 n14198_bdd_4_lut (.I0(n14198), .I1(\REG.mem_57_4 ), .I2(\REG.mem_56_4 ), 
            .I3(rd_addr_r[1]), .O(n12066));
    defparam n14198_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11360 (.I0(rd_addr_r[4]), .I1(n12405), 
            .I2(n12420), .I3(rd_addr_r[5]), .O(n12794));
    defparam rd_addr_r_4__bdd_4_lut_11360.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_6__I_0_151_6_lut (.I0(GND_net), .I1(rd_addr_r[4]), 
            .I2(GND_net), .I3(n10640), .O(rd_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12308 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_8 ), 
            .I2(\REG.mem_15_8 ), .I3(rd_addr_r[1]), .O(n14192));
    defparam rd_addr_r_0__bdd_4_lut_12308.LUT_INIT = 16'he4aa;
    SB_LUT4 n13490_bdd_4_lut (.I0(n13490), .I1(n11792), .I2(n11791), .I3(rd_addr_r[2]), 
            .O(n13493));
    defparam n13490_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY rd_addr_r_6__I_0_151_6 (.CI(n10640), .I0(rd_addr_r[4]), .I1(GND_net), 
            .CO(n10641));
    SB_LUT4 rd_addr_r_6__I_0_151_5_lut (.I0(GND_net), .I1(rd_addr_r[3]), 
            .I2(GND_net), .I3(n10639), .O(rd_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4046_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_34_10 ), .O(n5248));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4046_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4372_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_53_9 ), .O(n5574));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4372_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12794_bdd_4_lut (.I0(n12794), .I1(n12387), .I2(n12375), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_526 [13]));
    defparam n12794_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11720 (.I0(rd_addr_r[1]), .I1(n11674), 
            .I2(n11675), .I3(rd_addr_r[2]), .O(n13484));
    defparam rd_addr_r_1__bdd_4_lut_11720.LUT_INIT = 16'he4aa;
    SB_DFF i338_339 (.Q(\REG.mem_3_4 ), .C(DEBUG_6_c_c), .D(n4729));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13484_bdd_4_lut (.I0(n13484), .I1(n11648), .I2(n11647), .I3(rd_addr_r[2]), 
            .O(n13487));
    defparam n13484_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14192_bdd_4_lut (.I0(n14192), .I1(\REG.mem_13_8 ), .I2(\REG.mem_12_8 ), 
            .I3(rd_addr_r[1]), .O(n11667));
    defparam n14192_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11266 (.I0(rd_addr_r[2]), .I1(n12327), 
            .I2(n12339), .I3(rd_addr_r[3]), .O(n12902));
    defparam rd_addr_r_2__bdd_4_lut_11266.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12353 (.I0(rd_addr_r[1]), .I1(n11530), 
            .I2(n11531), .I3(rd_addr_r[2]), .O(n14186));
    defparam rd_addr_r_1__bdd_4_lut_12353.LUT_INIT = 16'he4aa;
    SB_LUT4 n14186_bdd_4_lut (.I0(n14186), .I1(n11510), .I2(n11509), .I3(rd_addr_r[2]), 
            .O(n14189));
    defparam n14186_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4371_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_53_8 ), .O(n5573));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4371_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12303 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_10 ), 
            .I2(\REG.mem_11_10 ), .I3(rd_addr_r[1]), .O(n14180));
    defparam rd_addr_r_0__bdd_4_lut_12303.LUT_INIT = 16'he4aa;
    SB_LUT4 n14180_bdd_4_lut (.I0(n14180), .I1(\REG.mem_9_10 ), .I2(\REG.mem_8_10 ), 
            .I3(rd_addr_r[1]), .O(n14183));
    defparam n14180_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11794 (.I0(rd_addr_r[2]), .I1(n12165), 
            .I2(n12168), .I3(rd_addr_r[3]), .O(n13478));
    defparam rd_addr_r_2__bdd_4_lut_11794.LUT_INIT = 16'he4aa;
    SB_DFFE \REG.out_raw__i1  (.Q(\REG.out_raw[0] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [0]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 i4370_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_53_7 ), .O(n5572));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4370_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12293 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_13 ), 
            .I2(\REG.mem_11_13 ), .I3(rd_addr_r[1]), .O(n14174));
    defparam rd_addr_r_0__bdd_4_lut_12293.LUT_INIT = 16'he4aa;
    SB_LUT4 n14174_bdd_4_lut (.I0(n14174), .I1(\REG.mem_9_13 ), .I2(\REG.mem_8_13 ), 
            .I3(rd_addr_r[1]), .O(n12075));
    defparam n14174_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13478_bdd_4_lut (.I0(n13478), .I1(n12150), .I2(n12144), .I3(rd_addr_r[3]), 
            .O(n12282));
    defparam n13478_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4369_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_53_6 ), .O(n5571));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4369_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut (.I0(wr_sig_diff0_w[2]), .I1(wr_sig_diff0_w[1]), .I2(wr_sig_diff0_w[0]), 
            .I3(GND_net), .O(n10784));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 n12902_bdd_4_lut (.I0(n12902), .I1(n12276), .I2(n12255), .I3(rd_addr_r[3]), 
            .O(n12420));
    defparam n12902_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9815_4_lut (.I0(DEBUG_9_c), .I1(n11436), .I2(n10784), .I3(wr_sig_diff0_w[3]), 
            .O(n11463));
    defparam i9815_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 wr_addr_r_6__I_0_135_i5_3_lut (.I0(wr_addr_r[4]), .I1(wr_addr_p1_w[4]), 
            .I2(n7596), .I3(GND_net), .O(\wr_addr_nxt_c[4] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i5_3_lut.LUT_INIT = 16'hacac;
    SB_DFF i335_336 (.Q(\REG.mem_3_3 ), .C(DEBUG_6_c_c), .D(n4728));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11729 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_14 ), 
            .I2(\REG.mem_27_14 ), .I3(rd_addr_r[1]), .O(n13472));
    defparam rd_addr_r_0__bdd_4_lut_11729.LUT_INIT = 16'he4aa;
    SB_LUT4 i4368_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_53_5 ), .O(n5570));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4368_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i332_333 (.Q(\REG.mem_3_2 ), .C(DEBUG_6_c_c), .D(n4727));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13472_bdd_4_lut (.I0(n13472), .I1(\REG.mem_25_14 ), .I2(\REG.mem_24_14 ), 
            .I3(rd_addr_r[1]), .O(n13475));
    defparam n13472_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12288 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_2 ), 
            .I2(\REG.mem_43_2 ), .I3(rd_addr_r[1]), .O(n14168));
    defparam rd_addr_r_0__bdd_4_lut_12288.LUT_INIT = 16'he4aa;
    SB_LUT4 i4045_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_34_9 ), .O(n5247));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4045_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14168_bdd_4_lut (.I0(n14168), .I1(\REG.mem_41_2 ), .I2(\REG.mem_40_2 ), 
            .I3(rd_addr_r[1]), .O(n12078));
    defparam n14168_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11710 (.I0(rd_addr_r[2]), .I1(n12195), 
            .I2(n12198), .I3(rd_addr_r[3]), .O(n13466));
    defparam rd_addr_r_2__bdd_4_lut_11710.LUT_INIT = 16'he4aa;
    SB_LUT4 n13466_bdd_4_lut (.I0(n13466), .I1(n12180), .I2(n12177), .I3(rd_addr_r[3]), 
            .O(n12288));
    defparam n13466_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12283 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_10 ), 
            .I2(\REG.mem_15_10 ), .I3(rd_addr_r[1]), .O(n14162));
    defparam rd_addr_r_0__bdd_4_lut_12283.LUT_INIT = 16'he4aa;
    SB_DFFSR \afull_flag_impl.af_flag_ext_r_121  (.Q(DEBUG_9_c), .C(DEBUG_6_c_c), 
            .D(\afull_flag_impl.af_flag_nxt_w ), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(410[29] 422[32])
    SB_DFF i329_330 (.Q(\REG.mem_3_1 ), .C(DEBUG_6_c_c), .D(n4726));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11705 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_8 ), 
            .I2(\REG.mem_55_8 ), .I3(rd_addr_r[1]), .O(n13460));
    defparam rd_addr_r_0__bdd_4_lut_11705.LUT_INIT = 16'he4aa;
    SB_LUT4 i4044_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_34_8 ), .O(n5246));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4044_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i326_327 (.Q(\REG.mem_3_0 ), .C(DEBUG_6_c_c), .D(n4725));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4043_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_34_7 ), .O(n5245));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4043_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13460_bdd_4_lut (.I0(n13460), .I1(\REG.mem_53_8 ), .I2(\REG.mem_52_8 ), 
            .I3(rd_addr_r[1]), .O(n11853));
    defparam n13460_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14162_bdd_4_lut (.I0(n14162), .I1(\REG.mem_13_10 ), .I2(\REG.mem_12_10 ), 
            .I3(rd_addr_r[1]), .O(n14165));
    defparam n14162_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4367_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_53_4 ), .O(n5569));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4367_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11695 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_3 ), 
            .I2(\REG.mem_43_3 ), .I3(rd_addr_r[1]), .O(n13454));
    defparam rd_addr_r_0__bdd_4_lut_11695.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12298 (.I0(rd_addr_r[1]), .I1(n12013), 
            .I2(n12014), .I3(rd_addr_r[2]), .O(n14156));
    defparam rd_addr_r_1__bdd_4_lut_12298.LUT_INIT = 16'he4aa;
    SB_LUT4 n13454_bdd_4_lut (.I0(n13454), .I1(\REG.mem_41_3 ), .I2(\REG.mem_40_3 ), 
            .I3(rd_addr_r[1]), .O(n13457));
    defparam n13454_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4042_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_34_6 ), .O(n5244));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4042_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFSR rd_grey_sync_r__i0 (.Q(\rd_grey_sync_r[0] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[0]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 i4366_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_53_3 ), .O(n5568));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4366_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4041_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_34_5 ), .O(n5243));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4041_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4040_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_34_4 ), .O(n5242));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4040_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14156_bdd_4_lut (.I0(n14156), .I1(n11999), .I2(n11998), .I3(rd_addr_r[2]), 
            .O(n12080));
    defparam n14156_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12273 (.I0(rd_addr_r[1]), .I1(n12043), 
            .I2(n12044), .I3(rd_addr_r[2]), .O(n14150));
    defparam rd_addr_r_1__bdd_4_lut_12273.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11690 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_8 ), 
            .I2(\REG.mem_59_8 ), .I3(rd_addr_r[1]), .O(n13448));
    defparam rd_addr_r_0__bdd_4_lut_11690.LUT_INIT = 16'he4aa;
    SB_DFFSS empty_ext_r_124 (.Q(DEBUG_5_c), .C(SLM_CLK_c), .D(empty_nxt_c_N_596), 
            .S(reset_all));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_LUT4 n14150_bdd_4_lut (.I0(n14150), .I1(n12035), .I2(n12034), .I3(rd_addr_r[2]), 
            .O(n12083));
    defparam n14150_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13448_bdd_4_lut (.I0(n13448), .I1(\REG.mem_57_8 ), .I2(\REG.mem_56_8 ), 
            .I3(rd_addr_r[1]), .O(n11862));
    defparam n13448_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR wr_grey_sync_r__i0 (.Q(wr_grey_sync_r[0]), .C(DEBUG_6_c_c), 
            .D(wr_grey_w[0]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_LUT4 i4039_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_34_3 ), .O(n5241));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4039_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10646_3_lut (.I0(\REG.mem_48_5 ), .I1(\REG.mem_49_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12295));
    defparam i10646_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFS \aempty_flag_impl.ae_flag_ext_r_130  (.Q(dc32_fifo_almost_empty), 
            .C(SLM_CLK_c), .D(\aempty_flag_impl.ae_flag_nxt_w ), .S(reset_all));   // src/fifo_dc_32_lut_gen.v(669[37] 672[40])
    SB_LUT4 i4365_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_53_2 ), .O(n5567));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4365_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12278 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_11 ), 
            .I2(\REG.mem_55_11 ), .I3(rd_addr_r[1]), .O(n14144));
    defparam rd_addr_r_0__bdd_4_lut_12278.LUT_INIT = 16'he4aa;
    SB_DFF i275_276 (.Q(\REG.mem_2_15 ), .C(DEBUG_6_c_c), .D(n4723));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i272_273 (.Q(\REG.mem_2_14 ), .C(DEBUG_6_c_c), .D(n4722));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_4__bdd_4_lut_12188 (.I0(rd_addr_r[4]), .I1(n12240), 
            .I2(n12246), .I3(rd_addr_r[5]), .O(n13442));
    defparam rd_addr_r_4__bdd_4_lut_12188.LUT_INIT = 16'he4aa;
    SB_LUT4 i10647_3_lut (.I0(\REG.mem_50_5 ), .I1(\REG.mem_51_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12296));
    defparam i10647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n14144_bdd_4_lut (.I0(n14144), .I1(\REG.mem_53_11 ), .I2(\REG.mem_52_11 ), 
            .I3(rd_addr_r[1]), .O(n14147));
    defparam n14144_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13442_bdd_4_lut (.I0(n13442), .I1(n12183), .I2(n12162), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_526 [4]));
    defparam n13442_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4364_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_53_1 ), .O(n5566));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4364_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10656_3_lut (.I0(\REG.mem_54_5 ), .I1(\REG.mem_55_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12305));
    defparam i10656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10655_3_lut (.I0(\REG.mem_52_5 ), .I1(\REG.mem_53_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12304));
    defparam i10655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12263 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_4 ), 
            .I2(\REG.mem_63_4 ), .I3(rd_addr_r[1]), .O(n14138));
    defparam rd_addr_r_0__bdd_4_lut_12263.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11685 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_11 ), 
            .I2(\REG.mem_23_11 ), .I3(rd_addr_r[1]), .O(n13436));
    defparam rd_addr_r_0__bdd_4_lut_11685.LUT_INIT = 16'he4aa;
    SB_LUT4 n14138_bdd_4_lut (.I0(n14138), .I1(\REG.mem_61_4 ), .I2(\REG.mem_60_4 ), 
            .I3(rd_addr_r[1]), .O(n12093));
    defparam n14138_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4363_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_53_0 ), .O(n5565));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4363_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10643_3_lut (.I0(\REG.mem_0_12 ), .I1(\REG.mem_1_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12292));
    defparam i10643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13436_bdd_4_lut (.I0(n13436), .I1(\REG.mem_21_11 ), .I2(\REG.mem_20_11 ), 
            .I3(rd_addr_r[1]), .O(n13439));
    defparam n13436_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10644_3_lut (.I0(\REG.mem_2_12 ), .I1(\REG.mem_3_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12293));
    defparam i10644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11675 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_12 ), 
            .I2(\REG.mem_11_12 ), .I3(rd_addr_r[1]), .O(n13430));
    defparam rd_addr_r_0__bdd_4_lut_11675.LUT_INIT = 16'he4aa;
    SB_LUT4 n13430_bdd_4_lut (.I0(n13430), .I1(\REG.mem_9_12 ), .I2(\REG.mem_8_12 ), 
            .I3(rd_addr_r[1]), .O(n13433));
    defparam n13430_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12268 (.I0(rd_addr_r[1]), .I1(n12016), 
            .I2(n12017), .I3(rd_addr_r[2]), .O(n14132));
    defparam rd_addr_r_1__bdd_4_lut_12268.LUT_INIT = 16'he4aa;
    SB_LUT4 n14132_bdd_4_lut (.I0(n14132), .I1(n12008), .I2(n12007), .I3(rd_addr_r[2]), 
            .O(n12098));
    defparam n14132_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11670 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_11 ), 
            .I2(\REG.mem_39_11 ), .I3(rd_addr_r[1]), .O(n13424));
    defparam rd_addr_r_0__bdd_4_lut_11670.LUT_INIT = 16'he4aa;
    SB_LUT4 n13424_bdd_4_lut (.I0(n13424), .I1(\REG.mem_37_11 ), .I2(\REG.mem_36_11 ), 
            .I3(rd_addr_r[1]), .O(n13427));
    defparam n13424_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11665 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_4 ), 
            .I2(\REG.mem_35_4 ), .I3(rd_addr_r[1]), .O(n13418));
    defparam rd_addr_r_0__bdd_4_lut_11665.LUT_INIT = 16'he4aa;
    SB_LUT4 n13418_bdd_4_lut (.I0(n13418), .I1(\REG.mem_33_4 ), .I2(\REG.mem_32_4 ), 
            .I3(rd_addr_r[1]), .O(n13421));
    defparam n13418_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i269_270 (.Q(\REG.mem_2_13 ), .C(DEBUG_6_c_c), .D(n4721));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11660 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_12 ), 
            .I2(\REG.mem_15_12 ), .I3(rd_addr_r[1]), .O(n13412));
    defparam rd_addr_r_0__bdd_4_lut_11660.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12258 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_13 ), 
            .I2(\REG.mem_15_13 ), .I3(rd_addr_r[1]), .O(n14126));
    defparam rd_addr_r_0__bdd_4_lut_12258.LUT_INIT = 16'he4aa;
    SB_LUT4 i10650_3_lut (.I0(\REG.mem_6_12 ), .I1(\REG.mem_7_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12299));
    defparam i10650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10649_3_lut (.I0(\REG.mem_4_12 ), .I1(\REG.mem_5_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12298));
    defparam i10649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n14126_bdd_4_lut (.I0(n14126), .I1(\REG.mem_13_13 ), .I2(\REG.mem_12_13 ), 
            .I3(rd_addr_r[1]), .O(n12102));
    defparam n14126_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSR full_ext_r_117 (.Q(full_o), .C(DEBUG_6_c_c), .D(full_nxt_c_N_593), 
            .R(reset_all));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 n13412_bdd_4_lut (.I0(n13412), .I1(\REG.mem_13_12 ), .I2(\REG.mem_12_12 ), 
            .I3(rd_addr_r[1]), .O(n13415));
    defparam n13412_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i266_267 (.Q(\REG.mem_2_12 ), .C(DEBUG_6_c_c), .D(n4720));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i263_264 (.Q(\REG.mem_2_11 ), .C(DEBUG_6_c_c), .D(n4719));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11148 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_15 ), 
            .I2(\REG.mem_23_15 ), .I3(rd_addr_r[1]), .O(n12788));
    defparam rd_addr_r_0__bdd_4_lut_11148.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11655 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_12 ), 
            .I2(\REG.mem_19_12 ), .I3(rd_addr_r[1]), .O(n13406));
    defparam rd_addr_r_0__bdd_4_lut_11655.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11171 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_8 ), 
            .I2(\REG.mem_7_8 ), .I3(rd_addr_r[1]), .O(n12824));
    defparam rd_addr_r_0__bdd_4_lut_11171.LUT_INIT = 16'he4aa;
    SB_CARRY wr_addr_r_6__I_0_add_2_5 (.CI(n10627), .I0(wr_addr_r[3]), .I1(rp_sync_w[3]), 
            .CO(n10628));
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12248 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_2 ), 
            .I2(\REG.mem_3_2 ), .I3(rd_addr_r[1]), .O(n14120));
    defparam rd_addr_r_0__bdd_4_lut_12248.LUT_INIT = 16'he4aa;
    SB_LUT4 n13406_bdd_4_lut (.I0(n13406), .I1(\REG.mem_17_12 ), .I2(\REG.mem_16_12 ), 
            .I3(rd_addr_r[1]), .O(n12312));
    defparam n13406_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i260_261 (.Q(\REG.mem_2_10 ), .C(DEBUG_6_c_c), .D(n4718));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i257_258 (.Q(\REG.mem_2_9 ), .C(DEBUG_6_c_c), .D(n4717));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i254_255 (.Q(\REG.mem_2_8 ), .C(DEBUG_6_c_c), .D(n4716));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14120_bdd_4_lut (.I0(n14120), .I1(\REG.mem_1_2 ), .I2(\REG.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(n14123));
    defparam n14120_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_r_6__I_0_135_i3_3_lut (.I0(wr_addr_r[2]), .I1(wr_addr_p1_w[2]), 
            .I2(n7596), .I3(GND_net), .O(\wr_addr_nxt_c[2] ));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i3_3_lut.LUT_INIT = 16'hacac;
    SB_DFF i251_252 (.Q(\REG.mem_2_7 ), .C(DEBUG_6_c_c), .D(n4715));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i248_249 (.Q(\REG.mem_2_6 ), .C(DEBUG_6_c_c), .D(n4714));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12333 (.I0(rd_addr_r[3]), .I1(n13679), 
            .I2(n12083), .I3(rd_addr_r[4]), .O(n14114));
    defparam rd_addr_r_3__bdd_4_lut_12333.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11650 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_0 ), 
            .I2(\REG.mem_27_0 ), .I3(rd_addr_r[1]), .O(n13400));
    defparam rd_addr_r_0__bdd_4_lut_11650.LUT_INIT = 16'he4aa;
    SB_LUT4 n13400_bdd_4_lut (.I0(n13400), .I1(\REG.mem_25_0 ), .I2(\REG.mem_24_0 ), 
            .I3(rd_addr_r[1]), .O(n13403));
    defparam n13400_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14114_bdd_4_lut (.I0(n14114), .I1(n12080), .I2(n13673), .I3(rd_addr_r[4]), 
            .O(n14117));
    defparam n14114_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11645 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_10 ), 
            .I2(\REG.mem_43_10 ), .I3(rd_addr_r[1]), .O(n13394));
    defparam rd_addr_r_0__bdd_4_lut_11645.LUT_INIT = 16'he4aa;
    SB_DFF i245_246 (.Q(\REG.mem_2_5 ), .C(DEBUG_6_c_c), .D(n4713));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12243 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_8 ), 
            .I2(\REG.mem_19_8 ), .I3(rd_addr_r[1]), .O(n14108));
    defparam rd_addr_r_0__bdd_4_lut_12243.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11241 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_15 ), 
            .I2(\REG.mem_15_15 ), .I3(rd_addr_r[1]), .O(n12896));
    defparam rd_addr_r_0__bdd_4_lut_11241.LUT_INIT = 16'he4aa;
    SB_LUT4 n14108_bdd_4_lut (.I0(n14108), .I1(\REG.mem_17_8 ), .I2(\REG.mem_16_8 ), 
            .I3(rd_addr_r[1]), .O(n11691));
    defparam n14108_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13394_bdd_4_lut (.I0(n13394), .I1(\REG.mem_41_10 ), .I2(\REG.mem_40_10 ), 
            .I3(rd_addr_r[1]), .O(n13397));
    defparam n13394_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i80_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n60));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i80_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_DFF i242_243 (.Q(\REG.mem_2_4 ), .C(DEBUG_6_c_c), .D(n4712));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12233 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_13 ), 
            .I2(\REG.mem_19_13 ), .I3(rd_addr_r[1]), .O(n14102));
    defparam rd_addr_r_0__bdd_4_lut_12233.LUT_INIT = 16'he4aa;
    SB_DFF i239_240 (.Q(\REG.mem_2_3 ), .C(DEBUG_6_c_c), .D(n4711));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14102_bdd_4_lut (.I0(n14102), .I1(\REG.mem_17_13 ), .I2(\REG.mem_16_13 ), 
            .I3(rd_addr_r[1]), .O(n12108));
    defparam n14102_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i79_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n28));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i79_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 n12896_bdd_4_lut (.I0(n12896), .I1(\REG.mem_13_15 ), .I2(\REG.mem_12_15 ), 
            .I3(rd_addr_r[1]), .O(n12899));
    defparam n12896_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12228 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_3 ), 
            .I2(\REG.mem_27_3 ), .I3(rd_addr_r[1]), .O(n14096));
    defparam rd_addr_r_0__bdd_4_lut_12228.LUT_INIT = 16'he4aa;
    SB_DFF i236_237 (.Q(\REG.mem_2_2 ), .C(DEBUG_6_c_c), .D(n4710));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11640 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_6 ), 
            .I2(\REG.mem_47_6 ), .I3(rd_addr_r[1]), .O(n13388));
    defparam rd_addr_r_0__bdd_4_lut_11640.LUT_INIT = 16'he4aa;
    SB_LUT4 n13388_bdd_4_lut (.I0(n13388), .I1(\REG.mem_45_6 ), .I2(\REG.mem_44_6 ), 
            .I3(rd_addr_r[1]), .O(n12315));
    defparam n13388_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i233_234 (.Q(\REG.mem_2_1 ), .C(DEBUG_6_c_c), .D(n4709));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i230_231 (.Q(\REG.mem_2_0 ), .C(DEBUG_6_c_c), .D(n4708));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14096_bdd_4_lut (.I0(n14096), .I1(\REG.mem_25_3 ), .I2(\REG.mem_24_3 ), 
            .I3(rd_addr_r[1]), .O(n14099));
    defparam n14096_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11635 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_8 ), 
            .I2(\REG.mem_63_8 ), .I3(rd_addr_r[1]), .O(n13382));
    defparam rd_addr_r_0__bdd_4_lut_11635.LUT_INIT = 16'he4aa;
    SB_LUT4 n13382_bdd_4_lut (.I0(n13382), .I1(\REG.mem_61_8 ), .I2(\REG.mem_60_8 ), 
            .I3(rd_addr_r[1]), .O(n11874));
    defparam n13382_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11834 (.I0(rd_addr_r[3]), .I1(n13355), 
            .I2(n11747), .I3(rd_addr_r[4]), .O(n13376));
    defparam rd_addr_r_3__bdd_4_lut_11834.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12223 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_7 ), 
            .I2(\REG.mem_3_7 ), .I3(rd_addr_r[1]), .O(n14090));
    defparam rd_addr_r_0__bdd_4_lut_12223.LUT_INIT = 16'he4aa;
    SB_LUT4 n13376_bdd_4_lut (.I0(n13376), .I1(n11744), .I2(n13349), .I3(rd_addr_r[4]), 
            .O(n13379));
    defparam n13376_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14090_bdd_4_lut (.I0(n14090), .I1(\REG.mem_1_7 ), .I2(\REG.mem_0_7 ), 
            .I3(rd_addr_r[1]), .O(n12111));
    defparam n14090_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11700 (.I0(rd_addr_r[2]), .I1(n11844), 
            .I2(n12315), .I3(rd_addr_r[3]), .O(n13370));
    defparam rd_addr_r_2__bdd_4_lut_11700.LUT_INIT = 16'he4aa;
    SB_DFF i38_39 (.Q(\REG.mem_0_0 ), .C(DEBUG_6_c_c), .D(n4707));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12218 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_2 ), 
            .I2(\REG.mem_47_2 ), .I3(rd_addr_r[1]), .O(n14084));
    defparam rd_addr_r_0__bdd_4_lut_12218.LUT_INIT = 16'he4aa;
    SB_LUT4 n13370_bdd_4_lut (.I0(n13370), .I1(n11838), .I2(n11835), .I3(rd_addr_r[3]), 
            .O(n13373));
    defparam n13370_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14084_bdd_4_lut (.I0(n14084), .I1(\REG.mem_45_2 ), .I2(\REG.mem_44_2 ), 
            .I3(rd_addr_r[1]), .O(n12114));
    defparam n14084_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11715 (.I0(rd_addr_r[1]), .I1(n11722), 
            .I2(n11723), .I3(rd_addr_r[2]), .O(n13364));
    defparam rd_addr_r_1__bdd_4_lut_11715.LUT_INIT = 16'he4aa;
    SB_LUT4 i4362_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_52_15 ), .O(n5564));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4362_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12238 (.I0(rd_addr_r[3]), .I1(n13685), 
            .I2(n12098), .I3(rd_addr_r[4]), .O(n14078));
    defparam rd_addr_r_3__bdd_4_lut_12238.LUT_INIT = 16'he4aa;
    SB_LUT4 n13364_bdd_4_lut (.I0(n13364), .I1(n11720), .I2(n11719), .I3(rd_addr_r[2]), 
            .O(n13367));
    defparam n13364_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i41_42 (.Q(\REG.mem_0_1 ), .C(DEBUG_6_c_c), .D(n4706));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14078_bdd_4_lut (.I0(n14078), .I1(n12095), .I2(n12094), .I3(rd_addr_r[4]), 
            .O(n14081));
    defparam n14078_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11615 (.I0(rd_addr_r[1]), .I1(n11701), 
            .I2(n11702), .I3(rd_addr_r[2]), .O(n13358));
    defparam rd_addr_r_1__bdd_4_lut_11615.LUT_INIT = 16'he4aa;
    SB_LUT4 n13358_bdd_4_lut (.I0(n13358), .I1(n11699), .I2(n11698), .I3(rd_addr_r[2]), 
            .O(n13361));
    defparam n13358_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4361_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_52_14 ), .O(n5563));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4361_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12213 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_7 ), 
            .I2(\REG.mem_7_7 ), .I3(rd_addr_r[1]), .O(n14072));
    defparam rd_addr_r_0__bdd_4_lut_12213.LUT_INIT = 16'he4aa;
    SB_DFF i44_45 (.Q(\REG.mem_0_2 ), .C(DEBUG_6_c_c), .D(n4705));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3973_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_30_4 ), .O(n5175));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3973_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4360_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_52_13 ), .O(n5562));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4360_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11226 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_11 ), 
            .I2(\REG.mem_47_11 ), .I3(rd_addr_r[1]), .O(n12890));
    defparam rd_addr_r_0__bdd_4_lut_11226.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11610 (.I0(rd_addr_r[1]), .I1(n11680), 
            .I2(n11681), .I3(rd_addr_r[2]), .O(n13352));
    defparam rd_addr_r_1__bdd_4_lut_11610.LUT_INIT = 16'he4aa;
    SB_LUT4 i9864_3_lut (.I0(n13817), .I1(n13667), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11513));
    defparam i9864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13352_bdd_4_lut (.I0(n13352), .I1(n11678), .I2(n11677), .I3(rd_addr_r[2]), 
            .O(n13355));
    defparam n13352_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4038_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_34_2 ), .O(n5240));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4038_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9885_3_lut (.I0(n13475), .I1(n13331), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11534));
    defparam i9885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4359_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_52_12 ), .O(n5561));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4359_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14072_bdd_4_lut (.I0(n14072), .I1(\REG.mem_5_7 ), .I2(\REG.mem_4_7 ), 
            .I3(rd_addr_r[1]), .O(n12120));
    defparam n14072_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11605 (.I0(rd_addr_r[1]), .I1(n11656), 
            .I2(n11657), .I3(rd_addr_r[2]), .O(n13346));
    defparam rd_addr_r_1__bdd_4_lut_11605.LUT_INIT = 16'he4aa;
    SB_CARRY rd_addr_r_6__I_0_151_5 (.CI(n10639), .I0(rd_addr_r[3]), .I1(GND_net), 
            .CO(n10640));
    SB_LUT4 i4358_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_52_11 ), .O(n5560));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4358_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12890_bdd_4_lut (.I0(n12890), .I1(\REG.mem_45_11 ), .I2(\REG.mem_44_11 ), 
            .I3(rd_addr_r[1]), .O(n12893));
    defparam n12890_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12203 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_13 ), 
            .I2(\REG.mem_23_13 ), .I3(rd_addr_r[1]), .O(n14066));
    defparam rd_addr_r_0__bdd_4_lut_12203.LUT_INIT = 16'he4aa;
    SB_LUT4 n13346_bdd_4_lut (.I0(n13346), .I1(n11654), .I2(n11653), .I3(rd_addr_r[2]), 
            .O(n13349));
    defparam n13346_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4357_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_52_10 ), .O(n5559));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4357_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14066_bdd_4_lut (.I0(n14066), .I1(\REG.mem_21_13 ), .I2(\REG.mem_20_13 ), 
            .I3(rd_addr_r[1]), .O(n12123));
    defparam n14066_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i47_48 (.Q(\REG.mem_0_3 ), .C(DEBUG_6_c_c), .D(n4704));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11630 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_5 ), 
            .I2(\REG.mem_59_5 ), .I3(rd_addr_r[1]), .O(n13340));
    defparam rd_addr_r_0__bdd_4_lut_11630.LUT_INIT = 16'he4aa;
    SB_LUT4 n13340_bdd_4_lut (.I0(n13340), .I1(\REG.mem_57_5 ), .I2(\REG.mem_56_5 ), 
            .I3(rd_addr_r[1]), .O(n13343));
    defparam n13340_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4356_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_52_9 ), .O(n5558));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4356_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12198 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_8 ), 
            .I2(\REG.mem_23_8 ), .I3(rd_addr_r[1]), .O(n14060));
    defparam rd_addr_r_0__bdd_4_lut_12198.LUT_INIT = 16'he4aa;
    SB_LUT4 i4037_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_34_1 ), .O(n5239));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4037_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4355_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_52_8 ), .O(n5557));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4355_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_6__I_0_151_4_lut (.I0(GND_net), .I1(rd_addr_r[2]), 
            .I2(GND_net), .I3(n10638), .O(rd_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4036_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_34_0 ), .O(n5238));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4036_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14060_bdd_4_lut (.I0(n14060), .I1(\REG.mem_21_8 ), .I2(\REG.mem_20_8 ), 
            .I3(rd_addr_r[1]), .O(n11709));
    defparam n14060_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_12403 (.I0(rd_addr_r[4]), .I1(n11643), 
            .I2(n11670), .I3(rd_addr_r[5]), .O(n14054));
    defparam rd_addr_r_4__bdd_4_lut_12403.LUT_INIT = 16'he4aa;
    SB_LUT4 n14054_bdd_4_lut (.I0(n14054), .I1(n13097), .I2(n11577), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_526 [12]));
    defparam n14054_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY rd_addr_r_6__I_0_151_4 (.CI(n10638), .I0(rd_addr_r[2]), .I1(GND_net), 
            .CO(n10639));
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11595 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_3 ), 
            .I2(\REG.mem_47_3 ), .I3(rd_addr_r[1]), .O(n13334));
    defparam rd_addr_r_0__bdd_4_lut_11595.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12193 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_7 ), 
            .I2(\REG.mem_11_7 ), .I3(rd_addr_r[1]), .O(n14048));
    defparam rd_addr_r_0__bdd_4_lut_12193.LUT_INIT = 16'he4aa;
    SB_LUT4 n13334_bdd_4_lut (.I0(n13334), .I1(\REG.mem_45_3 ), .I2(\REG.mem_44_3 ), 
            .I3(rd_addr_r[1]), .O(n13337));
    defparam n13334_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10157_3_lut (.I0(\REG.mem_8_2 ), .I1(\REG.mem_9_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11806));
    defparam i10157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n14048_bdd_4_lut (.I0(n14048), .I1(\REG.mem_9_7 ), .I2(\REG.mem_8_7 ), 
            .I3(rd_addr_r[1]), .O(n12126));
    defparam n14048_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4354_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_52_7 ), .O(n5556));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4354_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11590 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_14 ), 
            .I2(\REG.mem_31_14 ), .I3(rd_addr_r[1]), .O(n13328));
    defparam rd_addr_r_0__bdd_4_lut_11590.LUT_INIT = 16'he4aa;
    SB_LUT4 i4353_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_52_6 ), .O(n5555));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4353_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10158_3_lut (.I0(\REG.mem_10_2 ), .I1(\REG.mem_11_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11807));
    defparam i10158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13328_bdd_4_lut (.I0(n13328), .I1(\REG.mem_29_14 ), .I2(\REG.mem_28_14 ), 
            .I3(rd_addr_r[1]), .O(n13331));
    defparam n13328_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11585 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_13 ), 
            .I2(\REG.mem_59_13 ), .I3(rd_addr_r[1]), .O(n13322));
    defparam rd_addr_r_0__bdd_4_lut_11585.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12183 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_8 ), 
            .I2(\REG.mem_27_8 ), .I3(rd_addr_r[1]), .O(n14042));
    defparam rd_addr_r_0__bdd_4_lut_12183.LUT_INIT = 16'he4aa;
    SB_LUT4 n13322_bdd_4_lut (.I0(n13322), .I1(\REG.mem_57_13 ), .I2(\REG.mem_56_13 ), 
            .I3(rd_addr_r[1]), .O(n12327));
    defparam n13322_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10209_3_lut (.I0(\REG.mem_14_2 ), .I1(\REG.mem_15_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11858));
    defparam i10209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11620 (.I0(rd_addr_r[2]), .I1(n12228), 
            .I2(n12237), .I3(rd_addr_r[3]), .O(n13316));
    defparam rd_addr_r_2__bdd_4_lut_11620.LUT_INIT = 16'he4aa;
    SB_LUT4 i10208_3_lut (.I0(\REG.mem_12_2 ), .I1(\REG.mem_13_2 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11857));
    defparam i10208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n14042_bdd_4_lut (.I0(n14042), .I1(\REG.mem_25_8 ), .I2(\REG.mem_24_8 ), 
            .I3(rd_addr_r[1]), .O(n11718));
    defparam n14042_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13316_bdd_4_lut (.I0(n13316), .I1(n12222), .I2(n12210), .I3(rd_addr_r[3]), 
            .O(n12330));
    defparam n13316_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12178 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_7 ), 
            .I2(\REG.mem_15_7 ), .I3(rd_addr_r[1]), .O(n14036));
    defparam rd_addr_r_0__bdd_4_lut_12178.LUT_INIT = 16'he4aa;
    SB_LUT4 i4352_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_52_5 ), .O(n5554));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4352_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14036_bdd_4_lut (.I0(n14036), .I1(\REG.mem_13_7 ), .I2(\REG.mem_12_7 ), 
            .I3(rd_addr_r[1]), .O(n12129));
    defparam n14036_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11600 (.I0(rd_addr_r[1]), .I1(n12517), 
            .I2(n12518), .I3(rd_addr_r[2]), .O(n13310));
    defparam rd_addr_r_1__bdd_4_lut_11600.LUT_INIT = 16'he4aa;
    SB_LUT4 n13310_bdd_4_lut (.I0(n13310), .I1(n12506), .I2(n12505), .I3(rd_addr_r[2]), 
            .O(n13313));
    defparam n13310_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12173 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_13 ), 
            .I2(\REG.mem_27_13 ), .I3(rd_addr_r[1]), .O(n14030));
    defparam rd_addr_r_0__bdd_4_lut_12173.LUT_INIT = 16'he4aa;
    SB_LUT4 n14030_bdd_4_lut (.I0(n14030), .I1(\REG.mem_25_13 ), .I2(\REG.mem_24_13 ), 
            .I3(rd_addr_r[1]), .O(n12138));
    defparam n14030_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11196 (.I0(rd_addr_r[1]), .I1(n12130), 
            .I2(n12131), .I3(rd_addr_r[2]), .O(n12818));
    defparam rd_addr_r_1__bdd_4_lut_11196.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11575 (.I0(rd_addr_r[2]), .I1(n11646), 
            .I2(n11667), .I3(rd_addr_r[3]), .O(n13304));
    defparam rd_addr_r_2__bdd_4_lut_11575.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12168 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_3 ), 
            .I2(\REG.mem_7_3 ), .I3(rd_addr_r[1]), .O(n14024));
    defparam rd_addr_r_0__bdd_4_lut_12168.LUT_INIT = 16'he4aa;
    SB_LUT4 n13304_bdd_4_lut (.I0(n13304), .I1(n12827), .I2(n13073), .I3(rd_addr_r[3]), 
            .O(n11880));
    defparam n13304_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14024_bdd_4_lut (.I0(n14024), .I1(\REG.mem_5_3 ), .I2(\REG.mem_4_3 ), 
            .I3(rd_addr_r[1]), .O(n11559));
    defparam n14024_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4351_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_52_4 ), .O(n5553));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4351_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12788_bdd_4_lut (.I0(n12788), .I1(\REG.mem_21_15 ), .I2(\REG.mem_20_15 ), 
            .I3(rd_addr_r[1]), .O(n12791));
    defparam n12788_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4350_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_52_3 ), .O(n5552));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4350_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4349_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_52_2 ), .O(n5551));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4349_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4348_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_52_1 ), .O(n5550));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4348_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4347_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_52_0 ), .O(n5549));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4347_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11625 (.I0(rd_addr_r[3]), .I1(n13265), 
            .I2(n11627), .I3(rd_addr_r[4]), .O(n13298));
    defparam rd_addr_r_3__bdd_4_lut_11625.LUT_INIT = 16'he4aa;
    SB_LUT4 n13298_bdd_4_lut (.I0(n13298), .I1(n11621), .I2(n13259), .I3(rd_addr_r[4]), 
            .O(n13301));
    defparam n13298_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10851_3_lut (.I0(n13853), .I1(n14021), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12500));
    defparam i10851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11570 (.I0(rd_addr_r[1]), .I1(n12481), 
            .I2(n12482), .I3(rd_addr_r[2]), .O(n13292));
    defparam rd_addr_r_1__bdd_4_lut_11570.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i45_2_lut_3_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n45));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i45_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i10862_3_lut (.I0(n13517), .I1(n12875), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12511));
    defparam i10862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10055_3_lut (.I0(\REG.mem_40_1 ), .I1(\REG.mem_41_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11704));
    defparam i10055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12163 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_5 ), 
            .I2(\REG.mem_15_5 ), .I3(rd_addr_r[1]), .O(n14018));
    defparam rd_addr_r_0__bdd_4_lut_12163.LUT_INIT = 16'he4aa;
    SB_LUT4 n14018_bdd_4_lut (.I0(n14018), .I1(\REG.mem_13_5 ), .I2(\REG.mem_12_5 ), 
            .I3(rd_addr_r[1]), .O(n14021));
    defparam n14018_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10056_3_lut (.I0(\REG.mem_42_1 ), .I1(\REG.mem_43_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11705));
    defparam i10056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10065_3_lut (.I0(\REG.mem_46_1 ), .I1(\REG.mem_47_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11714));
    defparam i10065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13292_bdd_4_lut (.I0(n13292), .I1(n12476), .I2(n12475), .I3(rd_addr_r[2]), 
            .O(n13295));
    defparam n13292_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10064_3_lut (.I0(\REG.mem_44_1 ), .I1(\REG.mem_45_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11713));
    defparam i10064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12158 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_8 ), 
            .I2(\REG.mem_31_8 ), .I3(rd_addr_r[1]), .O(n14012));
    defparam rd_addr_r_0__bdd_4_lut_12158.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11680 (.I0(rd_addr_r[4]), .I1(n12288), 
            .I2(n12330), .I3(rd_addr_r[5]), .O(n13286));
    defparam rd_addr_r_4__bdd_4_lut_11680.LUT_INIT = 16'he4aa;
    SB_LUT4 n14012_bdd_4_lut (.I0(n14012), .I1(\REG.mem_29_8 ), .I2(\REG.mem_28_8 ), 
            .I3(rd_addr_r[1]), .O(n11736));
    defparam n14012_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3823_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_20_15 ), .O(n5025));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3823_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12153 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_10 ), 
            .I2(\REG.mem_27_10 ), .I3(rd_addr_r[1]), .O(n14006));
    defparam rd_addr_r_0__bdd_4_lut_12153.LUT_INIT = 16'he4aa;
    SB_LUT4 n13286_bdd_4_lut (.I0(n13286), .I1(n12282), .I2(n12258), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_526 [7]));
    defparam n13286_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14006_bdd_4_lut (.I0(n14006), .I1(\REG.mem_25_10 ), .I2(\REG.mem_24_10 ), 
            .I3(rd_addr_r[1]), .O(n14009));
    defparam n14006_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3822_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_20_14 ), .O(n5024));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3822_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11580 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_2 ), 
            .I2(\REG.mem_19_2 ), .I3(rd_addr_r[1]), .O(n13280));
    defparam rd_addr_r_0__bdd_4_lut_11580.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12148 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_3 ), 
            .I2(\REG.mem_31_3 ), .I3(rd_addr_r[1]), .O(n14000));
    defparam rd_addr_r_0__bdd_4_lut_12148.LUT_INIT = 16'he4aa;
    SB_LUT4 n13280_bdd_4_lut (.I0(n13280), .I1(\REG.mem_17_2 ), .I2(\REG.mem_16_2 ), 
            .I3(rd_addr_r[1]), .O(n13283));
    defparam n13280_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9875_3_lut (.I0(\REG.mem_0_10 ), .I1(\REG.mem_1_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11524));
    defparam i9875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9876_3_lut (.I0(\REG.mem_2_10 ), .I1(\REG.mem_3_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11525));
    defparam i9876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n14000_bdd_4_lut (.I0(n14000), .I1(\REG.mem_29_3 ), .I2(\REG.mem_28_3 ), 
            .I3(rd_addr_r[1]), .O(n14003));
    defparam n14000_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i78_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n61));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i78_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11545 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_13 ), 
            .I2(\REG.mem_63_13 ), .I3(rd_addr_r[1]), .O(n13274));
    defparam rd_addr_r_0__bdd_4_lut_11545.LUT_INIT = 16'he4aa;
    SB_LUT4 i3821_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_20_13 ), .O(n5023));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3821_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3820_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_20_12 ), .O(n5022));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3820_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13274_bdd_4_lut (.I0(n13274), .I1(\REG.mem_61_13 ), .I2(\REG.mem_60_13 ), 
            .I3(rd_addr_r[1]), .O(n12339));
    defparam n13274_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10535_3_lut (.I0(\REG.mem_0_14 ), .I1(\REG.mem_1_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12184));
    defparam i10535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i132_2_lut_3_lut (.I0(n35), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n34));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i132_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i77_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n29));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i77_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11139 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_6 ), 
            .I2(\REG.mem_51_6 ), .I3(rd_addr_r[1]), .O(n12782));
    defparam rd_addr_r_0__bdd_4_lut_11139.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12253 (.I0(rd_addr_r[1]), .I1(n11671), 
            .I2(n11672), .I3(rd_addr_r[2]), .O(n13994));
    defparam rd_addr_r_1__bdd_4_lut_12253.LUT_INIT = 16'he4aa;
    SB_LUT4 n13994_bdd_4_lut (.I0(n13994), .I1(n11660), .I2(n11659), .I3(rd_addr_r[2]), 
            .O(n11744));
    defparam n13994_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11555 (.I0(rd_addr_r[1]), .I1(n11584), 
            .I2(n11585), .I3(rd_addr_r[2]), .O(n13268));
    defparam rd_addr_r_1__bdd_4_lut_11555.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i84_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n58));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i84_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i10536_3_lut (.I0(\REG.mem_2_14 ), .I1(\REG.mem_3_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12185));
    defparam i10536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13268_bdd_4_lut (.I0(n13268), .I1(n11579), .I2(n11578), .I3(rd_addr_r[2]), 
            .O(n13271));
    defparam n13268_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10542_3_lut (.I0(\REG.mem_6_14 ), .I1(\REG.mem_7_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12191));
    defparam i10542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3819_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_20_11 ), .O(n5021));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3819_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i83_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n26));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i83_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i9879_3_lut (.I0(\REG.mem_6_10 ), .I1(\REG.mem_7_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11528));
    defparam i9879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9878_3_lut (.I0(\REG.mem_4_10 ), .I1(\REG.mem_5_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11527));
    defparam i9878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10541_3_lut (.I0(\REG.mem_4_14 ), .I1(\REG.mem_5_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12190));
    defparam i10541_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE \REG.out_buffer__i6  (.Q(\fifo_data_out[6] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n5896));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFFE \REG.out_buffer__i5  (.Q(\fifo_data_out[5] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n5893));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12138 (.I0(rd_addr_r[1]), .I1(n11695), 
            .I2(n11696), .I3(rd_addr_r[2]), .O(n13988));
    defparam rd_addr_r_1__bdd_4_lut_12138.LUT_INIT = 16'he4aa;
    SB_LUT4 n13988_bdd_4_lut (.I0(n13988), .I1(n11684), .I2(n11683), .I3(rd_addr_r[2]), 
            .O(n11747));
    defparam n13988_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3818_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_20_10 ), .O(n5020));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3818_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3817_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_20_9 ), .O(n5019));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3817_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9896_3_lut (.I0(\REG.mem_16_10 ), .I1(\REG.mem_17_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11545));
    defparam i9896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3816_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_20_8 ), .O(n5018));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3816_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3815_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_20_7 ), .O(n5017));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3815_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3814_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_20_6 ), .O(n5016));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3814_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9897_3_lut (.I0(\REG.mem_18_10 ), .I1(\REG.mem_19_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11546));
    defparam i9897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11535 (.I0(rd_addr_r[1]), .I1(n11548), 
            .I2(n11549), .I3(rd_addr_r[2]), .O(n13262));
    defparam rd_addr_r_1__bdd_4_lut_11535.LUT_INIT = 16'he4aa;
    SB_LUT4 i3813_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_20_5 ), .O(n5015));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3813_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF \REG.out_buffer__i7  (.Q(\fifo_data_out[7] ), .C(SLM_CLK_c), 
           .D(n11119));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12143 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_7 ), 
            .I2(\REG.mem_19_7 ), .I3(rd_addr_r[1]), .O(n13982));
    defparam rd_addr_r_0__bdd_4_lut_12143.LUT_INIT = 16'he4aa;
    SB_DFF \REG.out_buffer__i3  (.Q(\fifo_data_out[3] ), .C(SLM_CLK_c), 
           .D(n11139));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 n13982_bdd_4_lut (.I0(n13982), .I1(\REG.mem_17_7 ), .I2(\REG.mem_16_7 ), 
            .I3(rd_addr_r[1]), .O(n12144));
    defparam n13982_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13262_bdd_4_lut (.I0(n13262), .I1(n11546), .I2(n11545), .I3(rd_addr_r[2]), 
            .O(n13265));
    defparam n13262_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i50_51 (.Q(\REG.mem_0_4 ), .C(DEBUG_6_c_c), .D(n4702));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12128 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_2 ), 
            .I2(\REG.mem_51_2 ), .I3(rd_addr_r[1]), .O(n13976));
    defparam rd_addr_r_0__bdd_4_lut_12128.LUT_INIT = 16'he4aa;
    SB_LUT4 i3812_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_20_4 ), .O(n5014));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3812_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3811_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_20_3 ), .O(n5013));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3811_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11166 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_0 ), 
            .I2(\REG.mem_47_0 ), .I3(rd_addr_r[1]), .O(n12812));
    defparam rd_addr_r_0__bdd_4_lut_11166.LUT_INIT = 16'he4aa;
    SB_LUT4 i3810_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_20_2 ), .O(n5012));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3810_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3809_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_20_1 ), .O(n5011));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3809_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11157 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_9 ), 
            .I2(\REG.mem_47_9 ), .I3(rd_addr_r[1]), .O(n12800));
    defparam rd_addr_r_0__bdd_4_lut_11157.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11530 (.I0(rd_addr_r[1]), .I1(n11527), 
            .I2(n11528), .I3(rd_addr_r[2]), .O(n13256));
    defparam rd_addr_r_1__bdd_4_lut_11530.LUT_INIT = 16'he4aa;
    SB_LUT4 n12800_bdd_4_lut (.I0(n12800), .I1(\REG.mem_45_9 ), .I2(\REG.mem_44_9 ), 
            .I3(rd_addr_r[1]), .O(n12803));
    defparam n12800_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12782_bdd_4_lut (.I0(n12782), .I1(\REG.mem_49_6 ), .I2(\REG.mem_48_6 ), 
            .I3(rd_addr_r[1]), .O(n12785));
    defparam n12782_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13976_bdd_4_lut (.I0(n13976), .I1(\REG.mem_49_2 ), .I2(\REG.mem_48_2 ), 
            .I3(rd_addr_r[1]), .O(n13979));
    defparam n13976_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF \REG.out_buffer__i8  (.Q(\fifo_data_out[8] ), .C(SLM_CLK_c), 
           .D(n11097));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 n13256_bdd_4_lut (.I0(n13256), .I1(n11525), .I2(n11524), .I3(rd_addr_r[2]), 
            .O(n13259));
    defparam n13256_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3808_3_lut_4_lut (.I0(n45), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_20_0 ), .O(n5010));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3808_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE \REG.out_buffer__i0  (.Q(\fifo_data_out[0] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n5854));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 n12824_bdd_4_lut (.I0(n12824), .I1(\REG.mem_5_8 ), .I2(\REG.mem_4_8 ), 
            .I3(rd_addr_r[1]), .O(n12827));
    defparam n12824_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10076_3_lut (.I0(\REG.mem_56_1 ), .I1(\REG.mem_57_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11725));
    defparam i10076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11221 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_11 ), 
            .I2(\REG.mem_7_11 ), .I3(rd_addr_r[1]), .O(n12884));
    defparam rd_addr_r_0__bdd_4_lut_11221.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12133 (.I0(rd_addr_r[1]), .I1(n11713), 
            .I2(n11714), .I3(rd_addr_r[2]), .O(n13970));
    defparam rd_addr_r_1__bdd_4_lut_12133.LUT_INIT = 16'he4aa;
    SB_LUT4 i10077_3_lut (.I0(\REG.mem_58_1 ), .I1(\REG.mem_59_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11726));
    defparam i10077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13970_bdd_4_lut (.I0(n13970), .I1(n11705), .I2(n11704), .I3(rd_addr_r[2]), 
            .O(n11750));
    defparam n13970_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11560 (.I0(rd_addr_r[3]), .I1(n12511), 
            .I2(n12512), .I3(rd_addr_r[4]), .O(n13250));
    defparam rd_addr_r_3__bdd_4_lut_11560.LUT_INIT = 16'he4aa;
    SB_LUT4 i3839_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_21_15 ), .O(n5041));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3839_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11134 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_15 ), 
            .I2(\REG.mem_27_15 ), .I3(rd_addr_r[1]), .O(n12776));
    defparam rd_addr_r_0__bdd_4_lut_11134.LUT_INIT = 16'he4aa;
    SB_DFF \REG.out_buffer__i9  (.Q(\fifo_data_out[9] ), .C(SLM_CLK_c), 
           .D(n11095));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 i3838_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_21_14 ), .O(n5040));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3838_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12123 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_7 ), 
            .I2(\REG.mem_23_7 ), .I3(rd_addr_r[1]), .O(n13964));
    defparam rd_addr_r_0__bdd_4_lut_12123.LUT_INIT = 16'he4aa;
    SB_LUT4 n13964_bdd_4_lut (.I0(n13964), .I1(\REG.mem_21_7 ), .I2(\REG.mem_20_7 ), 
            .I3(rd_addr_r[1]), .O(n12150));
    defparam n13964_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13250_bdd_4_lut (.I0(n13250), .I1(n12500), .I2(n12499), .I3(rd_addr_r[4]), 
            .O(n13253));
    defparam n13250_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3837_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_21_13 ), .O(n5039));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3837_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF \REG.out_buffer__i1  (.Q(\fifo_data_out[1] ), .C(SLM_CLK_c), 
           .D(n11143));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i2  (.Q(\fifo_data_out[2] ), .C(SLM_CLK_c), 
           .D(n11141));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i10  (.Q(\fifo_data_out[10] ), .C(SLM_CLK_c), 
           .D(n11089));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF \REG.out_buffer__i11  (.Q(\fifo_data_out[11] ), .C(SLM_CLK_c), 
           .D(n11135));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11540 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_3 ), 
            .I2(\REG.mem_51_3 ), .I3(rd_addr_r[1]), .O(n13244));
    defparam rd_addr_r_0__bdd_4_lut_11540.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12113 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_13 ), 
            .I2(\REG.mem_31_13 ), .I3(rd_addr_r[1]), .O(n13958));
    defparam rd_addr_r_0__bdd_4_lut_12113.LUT_INIT = 16'he4aa;
    SB_LUT4 n13958_bdd_4_lut (.I0(n13958), .I1(\REG.mem_29_13 ), .I2(\REG.mem_28_13 ), 
            .I3(rd_addr_r[1]), .O(n12153));
    defparam n13958_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13244_bdd_4_lut (.I0(n13244), .I1(\REG.mem_49_3 ), .I2(\REG.mem_48_3 ), 
            .I3(rd_addr_r[1]), .O(n13247));
    defparam n13244_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3836_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_21_12 ), .O(n5038));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3836_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11525 (.I0(rd_addr_r[1]), .I1(n11857), 
            .I2(n11858), .I3(rd_addr_r[2]), .O(n13238));
    defparam rd_addr_r_1__bdd_4_lut_11525.LUT_INIT = 16'he4aa;
    SB_LUT4 n13238_bdd_4_lut (.I0(n13238), .I1(n11807), .I2(n11806), .I3(rd_addr_r[2]), 
            .O(n12347));
    defparam n13238_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11515 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_9 ), 
            .I2(\REG.mem_11_9 ), .I3(rd_addr_r[1]), .O(n13232));
    defparam rd_addr_r_0__bdd_4_lut_11515.LUT_INIT = 16'he4aa;
    SB_LUT4 n13232_bdd_4_lut (.I0(n13232), .I1(\REG.mem_9_9 ), .I2(\REG.mem_8_9 ), 
            .I3(rd_addr_r[1]), .O(n13235));
    defparam n13232_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11520 (.I0(rd_addr_r[3]), .I1(n13193), 
            .I2(n11534), .I3(rd_addr_r[4]), .O(n13226));
    defparam rd_addr_r_3__bdd_4_lut_11520.LUT_INIT = 16'he4aa;
    SB_LUT4 n13226_bdd_4_lut (.I0(n13226), .I1(n11513), .I2(n13163), .I3(rd_addr_r[4]), 
            .O(n13229));
    defparam n13226_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3835_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_21_11 ), .O(n5037));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3835_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12413 (.I0(rd_addr_r[2]), .I1(n13637), 
            .I2(n13601), .I3(rd_addr_r[3]), .O(n13946));
    defparam rd_addr_r_2__bdd_4_lut_12413.LUT_INIT = 16'he4aa;
    SB_LUT4 n13946_bdd_4_lut (.I0(n13946), .I1(n13649), .I2(n13661), .I3(rd_addr_r[3]), 
            .O(n13949));
    defparam n13946_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3834_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_21_10 ), .O(n5036));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3834_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3833_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_21_9 ), .O(n5035));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3833_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11510 (.I0(rd_addr_r[1]), .I1(n12298), 
            .I2(n12299), .I3(rd_addr_r[2]), .O(n13220));
    defparam rd_addr_r_1__bdd_4_lut_11510.LUT_INIT = 16'he4aa;
    SB_LUT4 i9900_3_lut (.I0(\REG.mem_22_10 ), .I1(\REG.mem_23_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11549));
    defparam i9900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9899_3_lut (.I0(\REG.mem_20_10 ), .I1(\REG.mem_21_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11548));
    defparam i9899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13220_bdd_4_lut (.I0(n13220), .I1(n12293), .I2(n12292), .I3(rd_addr_r[2]), 
            .O(n13223));
    defparam n13220_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10034_3_lut (.I0(\REG.mem_24_1 ), .I1(\REG.mem_25_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11683));
    defparam i10034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10035_3_lut (.I0(\REG.mem_26_1 ), .I1(\REG.mem_27_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11684));
    defparam i10035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11495 (.I0(rd_addr_r[1]), .I1(n12304), 
            .I2(n12305), .I3(rd_addr_r[2]), .O(n13214));
    defparam rd_addr_r_1__bdd_4_lut_11495.LUT_INIT = 16'he4aa;
    SB_LUT4 n13214_bdd_4_lut (.I0(n13214), .I1(n12296), .I2(n12295), .I3(rd_addr_r[2]), 
            .O(n13217));
    defparam n13214_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3832_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_21_8 ), .O(n5034));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3832_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i106_2_lut_3_lut (.I0(n26_adj_1146), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n47));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i106_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i6131_6132 (.Q(\REG.mem_63_15 ), .C(DEBUG_6_c_c), .D(n5789));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6128_6129 (.Q(\REG.mem_63_14 ), .C(DEBUG_6_c_c), .D(n5788));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6125_6126 (.Q(\REG.mem_63_13 ), .C(DEBUG_6_c_c), .D(n5787));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12108 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_11 ), 
            .I2(\REG.mem_31_11 ), .I3(rd_addr_r[1]), .O(n13940));
    defparam rd_addr_r_0__bdd_4_lut_12108.LUT_INIT = 16'he4aa;
    SB_LUT4 n12884_bdd_4_lut (.I0(n12884), .I1(\REG.mem_5_11 ), .I2(\REG.mem_4_11 ), 
            .I3(rd_addr_r[1]), .O(n12887));
    defparam n12884_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3831_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_21_7 ), .O(n5033));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3831_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10047_3_lut (.I0(\REG.mem_30_1 ), .I1(\REG.mem_31_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11696));
    defparam i10047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10046_3_lut (.I0(\REG.mem_28_1 ), .I1(\REG.mem_29_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11695));
    defparam i10046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11505 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_12 ), 
            .I2(\REG.mem_23_12 ), .I3(rd_addr_r[1]), .O(n13208));
    defparam rd_addr_r_0__bdd_4_lut_11505.LUT_INIT = 16'he4aa;
    SB_LUT4 i3830_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_21_6 ), .O(n5032));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3830_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13208_bdd_4_lut (.I0(n13208), .I1(\REG.mem_21_12 ), .I2(\REG.mem_20_12 ), 
            .I3(rd_addr_r[1]), .O(n12354));
    defparam n13208_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3829_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_21_5 ), .O(n5031));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3829_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3828_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_21_4 ), .O(n5030));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3828_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i6122_6123 (.Q(\REG.mem_63_12 ), .C(DEBUG_6_c_c), .D(n5786));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6119_6120 (.Q(\REG.mem_63_11 ), .C(DEBUG_6_c_c), .D(n5785));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6116_6117 (.Q(\REG.mem_63_10 ), .C(DEBUG_6_c_c), .D(n5784));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3827_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_21_3 ), .O(n5029));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3827_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i6113_6114 (.Q(\REG.mem_63_9 ), .C(DEBUG_6_c_c), .D(n5783));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11485 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_9 ), 
            .I2(\REG.mem_15_9 ), .I3(rd_addr_r[1]), .O(n13202));
    defparam rd_addr_r_0__bdd_4_lut_11485.LUT_INIT = 16'he4aa;
    SB_DFF i6110_6111 (.Q(\REG.mem_63_8 ), .C(DEBUG_6_c_c), .D(n5782));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6107_6108 (.Q(\REG.mem_63_7 ), .C(DEBUG_6_c_c), .D(n5781));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6104_6105 (.Q(\REG.mem_63_6 ), .C(DEBUG_6_c_c), .D(n5780));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6101_6102 (.Q(\REG.mem_63_5 ), .C(DEBUG_6_c_c), .D(n5779));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6098_6099 (.Q(\REG.mem_63_4 ), .C(DEBUG_6_c_c), .D(n5778));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6095_6096 (.Q(\REG.mem_63_3 ), .C(DEBUG_6_c_c), .D(n5777));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6092_6093 (.Q(\REG.mem_63_2 ), .C(DEBUG_6_c_c), .D(n5776));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6089_6090 (.Q(\REG.mem_63_1 ), .C(DEBUG_6_c_c), .D(n5775));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF \REG.out_buffer__i12  (.Q(\fifo_data_out[12] ), .C(SLM_CLK_c), 
           .D(n11133));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF i6086_6087 (.Q(\REG.mem_63_0 ), .C(DEBUG_6_c_c), .D(n5773));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6035_6036 (.Q(\REG.mem_62_15 ), .C(DEBUG_6_c_c), .D(n5772));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6032_6033 (.Q(\REG.mem_62_14 ), .C(DEBUG_6_c_c), .D(n5771));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6029_6030 (.Q(\REG.mem_62_13 ), .C(DEBUG_6_c_c), .D(n5770));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6026_6027 (.Q(\REG.mem_62_12 ), .C(DEBUG_6_c_c), .D(n5769));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6023_6024 (.Q(\REG.mem_62_11 ), .C(DEBUG_6_c_c), .D(n5768));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6020_6021 (.Q(\REG.mem_62_10 ), .C(DEBUG_6_c_c), .D(n5767));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6017_6018 (.Q(\REG.mem_62_9 ), .C(DEBUG_6_c_c), .D(n5766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6014_6015 (.Q(\REG.mem_62_8 ), .C(DEBUG_6_c_c), .D(n5765));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3826_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_21_2 ), .O(n5028));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3826_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i6011_6012 (.Q(\REG.mem_62_7 ), .C(DEBUG_6_c_c), .D(n5764));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13202_bdd_4_lut (.I0(n13202), .I1(\REG.mem_13_9 ), .I2(\REG.mem_12_9 ), 
            .I3(rd_addr_r[1]), .O(n13205));
    defparam n13202_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i6008_6009 (.Q(\REG.mem_62_6 ), .C(DEBUG_6_c_c), .D(n5763));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6005_6006 (.Q(\REG.mem_62_5 ), .C(DEBUG_6_c_c), .D(n5762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i6002_6003 (.Q(\REG.mem_62_4 ), .C(DEBUG_6_c_c), .D(n5761));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5999_6000 (.Q(\REG.mem_62_3 ), .C(DEBUG_6_c_c), .D(n5760));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13940_bdd_4_lut (.I0(n13940), .I1(\REG.mem_29_11 ), .I2(\REG.mem_28_11 ), 
            .I3(rd_addr_r[1]), .O(n13943));
    defparam n13940_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5996_5997 (.Q(\REG.mem_62_2 ), .C(DEBUG_6_c_c), .D(n5759));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5993_5994 (.Q(\REG.mem_62_1 ), .C(DEBUG_6_c_c), .D(n5758));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5990_5991 (.Q(\REG.mem_62_0 ), .C(DEBUG_6_c_c), .D(n5757));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3825_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_21_1 ), .O(n5027));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3825_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3824_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_21_0 ), .O(n5026));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3824_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3855_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_22_15 ), .O(n5057));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3855_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3854_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_22_14 ), .O(n5056));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3854_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11490 (.I0(rd_addr_r[1]), .I1(n12355), 
            .I2(n12356), .I3(rd_addr_r[2]), .O(n13196));
    defparam rd_addr_r_1__bdd_4_lut_11490.LUT_INIT = 16'he4aa;
    SB_LUT4 i9929_3_lut (.I0(\REG.mem_32_10 ), .I1(\REG.mem_33_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11578));
    defparam i9929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9930_3_lut (.I0(\REG.mem_34_10 ), .I1(\REG.mem_35_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11579));
    defparam i9930_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5939_5940 (.Q(\REG.mem_61_15 ), .C(DEBUG_6_c_c), .D(n5749));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5936_5937 (.Q(\REG.mem_61_14 ), .C(DEBUG_6_c_c), .D(n5748));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5933_5934 (.Q(\REG.mem_61_13 ), .C(DEBUG_6_c_c), .D(n5747));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5930_5931 (.Q(\REG.mem_61_12 ), .C(DEBUG_6_c_c), .D(n5746));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5927_5928 (.Q(\REG.mem_61_11 ), .C(DEBUG_6_c_c), .D(n5745));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5924_5925 (.Q(\REG.mem_61_10 ), .C(DEBUG_6_c_c), .D(n5744));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5921_5922 (.Q(\REG.mem_61_9 ), .C(DEBUG_6_c_c), .D(n5743));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5918_5919 (.Q(\REG.mem_61_8 ), .C(DEBUG_6_c_c), .D(n5742));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5915_5916 (.Q(\REG.mem_61_7 ), .C(DEBUG_6_c_c), .D(n5741));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5912_5913 (.Q(\REG.mem_61_6 ), .C(DEBUG_6_c_c), .D(n5740));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5909_5910 (.Q(\REG.mem_61_5 ), .C(DEBUG_6_c_c), .D(n5739));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5906_5907 (.Q(\REG.mem_61_4 ), .C(DEBUG_6_c_c), .D(n5738));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5903_5904 (.Q(\REG.mem_61_3 ), .C(DEBUG_6_c_c), .D(n5737));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9936_3_lut (.I0(\REG.mem_38_10 ), .I1(\REG.mem_39_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11585));
    defparam i9936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3853_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_22_13 ), .O(n5055));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3853_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3852_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_22_12 ), .O(n5054));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3852_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13196_bdd_4_lut (.I0(n13196), .I1(n12332), .I2(n12331), .I3(rd_addr_r[2]), 
            .O(n13199));
    defparam n13196_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_r_6__I_0_inv_0_i7_1_lut (.I0(rp_sync2_r[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // src/fifo_dc_32_lut_gen.v(212[47:78])
    defparam wr_addr_r_6__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3851_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_22_11 ), .O(n5053));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3851_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i105_2_lut_3_lut (.I0(n26_adj_1146), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n15));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i105_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12118 (.I0(rd_addr_r[1]), .I1(n11638), 
            .I2(n11639), .I3(rd_addr_r[2]), .O(n13934));
    defparam rd_addr_r_1__bdd_4_lut_12118.LUT_INIT = 16'he4aa;
    SB_LUT4 i3850_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_22_10 ), .O(n5052));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3850_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9935_3_lut (.I0(\REG.mem_36_10 ), .I1(\REG.mem_37_10 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11584));
    defparam i9935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13934_bdd_4_lut (.I0(n13934), .I1(n11552), .I2(n11551), .I3(rd_addr_r[2]), 
            .O(n13937));
    defparam n13934_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3849_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_22_9 ), .O(n5051));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3849_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10010_3_lut (.I0(\REG.mem_8_1 ), .I1(\REG.mem_9_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11659));
    defparam i10010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10092_3_lut (.I0(\REG.mem_62_1 ), .I1(\REG.mem_63_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11741));
    defparam i10092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10091_3_lut (.I0(\REG.mem_60_1 ), .I1(\REG.mem_61_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11740));
    defparam i10091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11475 (.I0(rd_addr_r[1]), .I1(n12271), 
            .I2(n12272), .I3(rd_addr_r[2]), .O(n13190));
    defparam rd_addr_r_1__bdd_4_lut_11475.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12093 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_8 ), 
            .I2(\REG.mem_35_8 ), .I3(rd_addr_r[1]), .O(n13928));
    defparam rd_addr_r_0__bdd_4_lut_12093.LUT_INIT = 16'he4aa;
    SB_LUT4 i10011_3_lut (.I0(\REG.mem_10_1 ), .I1(\REG.mem_11_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11660));
    defparam i10011_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5900_5901 (.Q(\REG.mem_61_2 ), .C(DEBUG_6_c_c), .D(n5736));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5897_5898 (.Q(\REG.mem_61_1 ), .C(DEBUG_6_c_c), .D(n5735));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5894_5895 (.Q(\REG.mem_61_0 ), .C(DEBUG_6_c_c), .D(n5734));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5843_5844 (.Q(\REG.mem_60_15 ), .C(DEBUG_6_c_c), .D(n5726));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF \REG.out_buffer__i4  (.Q(\fifo_data_out[4] ), .C(SLM_CLK_c), 
           .D(n11137));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF i5840_5841 (.Q(\REG.mem_60_14 ), .C(DEBUG_6_c_c), .D(n5724));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5837_5838 (.Q(\REG.mem_60_13 ), .C(DEBUG_6_c_c), .D(n5723));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5834_5835 (.Q(\REG.mem_60_12 ), .C(DEBUG_6_c_c), .D(n5722));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5831_5832 (.Q(\REG.mem_60_11 ), .C(DEBUG_6_c_c), .D(n5721));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3848_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_22_8 ), .O(n5050));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3848_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10023_3_lut (.I0(\REG.mem_14_1 ), .I1(\REG.mem_15_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11672));
    defparam i10023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3847_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_22_7 ), .O(n5049));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3847_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10022_3_lut (.I0(\REG.mem_12_1 ), .I1(\REG.mem_13_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11671));
    defparam i10022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10826_3_lut (.I0(\REG.mem_32_12 ), .I1(\REG.mem_33_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12475));
    defparam i10826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10827_3_lut (.I0(\REG.mem_34_12 ), .I1(\REG.mem_35_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12476));
    defparam i10827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3846_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_22_6 ), .O(n5048));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3846_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10833_3_lut (.I0(\REG.mem_38_12 ), .I1(\REG.mem_39_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12482));
    defparam i10833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13928_bdd_4_lut (.I0(n13928), .I1(\REG.mem_33_8 ), .I2(\REG.mem_32_8 ), 
            .I3(rd_addr_r[1]), .O(n11760));
    defparam n13928_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_6__I_0_151_3_lut (.I0(GND_net), .I1(rd_addr_r[1]), 
            .I2(GND_net), .I3(n10637), .O(rd_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wr_addr_r_6__I_0_add_2_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(rp_sync_w[2]), .I3(n10626), .O(wr_sig_diff0_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10832_3_lut (.I0(\REG.mem_36_12 ), .I1(\REG.mem_37_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12481));
    defparam i10832_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY wr_addr_r_6__I_0_add_2_4 (.CI(n10626), .I0(wr_addr_r[2]), .I1(rp_sync_w[2]), 
            .CO(n10627));
    SB_CARRY rd_addr_r_6__I_0_151_3 (.CI(n10637), .I0(rd_addr_r[1]), .I1(GND_net), 
            .CO(n10638));
    SB_LUT4 wr_addr_r_6__I_0_add_2_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), 
            .I2(rp_sync_w[1]), .I3(n10625), .O(wr_sig_diff0_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9972_3_lut (.I0(n14183), .I1(n14165), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11621));
    defparam i9972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9978_3_lut (.I0(n14009), .I1(n13901), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11627));
    defparam i9978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10482_3_lut (.I0(\REG.mem_38_5 ), .I1(\REG.mem_39_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12131));
    defparam i10482_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5828_5829 (.Q(\REG.mem_60_10 ), .C(DEBUG_6_c_c), .D(n5720));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5825_5826 (.Q(\REG.mem_60_9 ), .C(DEBUG_6_c_c), .D(n5719));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5822_5823 (.Q(\REG.mem_60_8 ), .C(DEBUG_6_c_c), .D(n5718));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5819_5820 (.Q(\REG.mem_60_7 ), .C(DEBUG_6_c_c), .D(n5717));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5816_5817 (.Q(\REG.mem_60_6 ), .C(DEBUG_6_c_c), .D(n5716));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5813_5814 (.Q(\REG.mem_60_5 ), .C(DEBUG_6_c_c), .D(n5715));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5810_5811 (.Q(\REG.mem_60_4 ), .C(DEBUG_6_c_c), .D(n5714));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5807_5808 (.Q(\REG.mem_60_3 ), .C(DEBUG_6_c_c), .D(n5713));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5804_5805 (.Q(\REG.mem_60_2 ), .C(DEBUG_6_c_c), .D(n5712));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5801_5802 (.Q(\REG.mem_60_1 ), .C(DEBUG_6_c_c), .D(n5711));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5798_5799 (.Q(\REG.mem_60_0 ), .C(DEBUG_6_c_c), .D(n5710));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync1_r__i1 (.Q(rp_sync1_r[1]), .C(DEBUG_6_c_c), .D(n5709));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i2 (.Q(rp_sync1_r[2]), .C(DEBUG_6_c_c), .D(n5708));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i3 (.Q(rp_sync1_r[3]), .C(DEBUG_6_c_c), .D(n5707));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i4 (.Q(rp_sync1_r[4]), .C(DEBUG_6_c_c), .D(n5706));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync1_r__i5 (.Q(rp_sync1_r[5]), .C(DEBUG_6_c_c), .D(n5705));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_CARRY wr_addr_r_6__I_0_add_2_3 (.CI(n10625), .I0(wr_addr_r[1]), .I1(rp_sync_w[1]), 
            .CO(n10626));
    SB_LUT4 i10481_3_lut (.I0(\REG.mem_36_5 ), .I1(\REG.mem_37_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12130));
    defparam i10481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_6__I_0_151_2_lut (.I0(GND_net), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(VCC_net), .O(rd_addr_p1_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10856_3_lut (.I0(\REG.mem_48_12 ), .I1(\REG.mem_49_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12505));
    defparam i10856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_add_2_2_lut (.I0(GND_net), .I1(\wr_addr_r[0] ), 
            .I2(rp_sync_w[0]), .I3(VCC_net), .O(wr_sig_diff0_w[0])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wr_addr_r_6__I_0_add_2_2 (.CI(VCC_net), .I0(\wr_addr_r[0] ), 
            .I1(rp_sync_w[0]), .CO(n10625));
    SB_CARRY rd_addr_r_6__I_0_151_2 (.CI(VCC_net), .I0(rd_addr_r[0]), .I1(GND_net), 
            .CO(n10637));
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_8_lut (.I0(rd_sig_diff0_w[4]), .I1(wp_sync2_r[6]), 
            .I2(n1_adj_1173[6]), .I3(n10624), .O(n6)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i10857_3_lut (.I0(\REG.mem_50_12 ), .I1(\REG.mem_51_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12506));
    defparam i10857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3845_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_22_5 ), .O(n5047));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3845_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10869_3_lut (.I0(\REG.mem_54_12 ), .I1(\REG.mem_55_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12518));
    defparam i10869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_7_lut (.I0(rd_sig_diff0_w[2]), .I1(wp_sync_w[5]), 
            .I2(n1_adj_1173[5]), .I3(n10623), .O(n7_c)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i3844_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_22_4 ), .O(n5046));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3844_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wr_addr_r_6__I_0_141_8_lut (.I0(GND_net), .I1(wr_grey_sync_r[6]), 
            .I2(GND_net), .I3(n10636), .O(\wr_addr_p1_w[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_7 (.CI(n10623), .I0(wp_sync_w[5]), 
            .I1(n1_adj_1173[5]), .CO(n10624));
    SB_LUT4 i10868_3_lut (.I0(\REG.mem_52_12 ), .I1(\REG.mem_53_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12517));
    defparam i10868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_6_lut (.I0(GND_net), .I1(wp_sync_w[4]), 
            .I2(n1_adj_1173[4]), .I3(n10622), .O(rd_sig_diff0_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF rp_sync1_r__i6 (.Q(rp_sync1_r[6]), .C(DEBUG_6_c_c), .D(n5704));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_LUT4 wr_addr_r_6__I_0_141_7_lut (.I0(GND_net), .I1(wr_addr_r[5]), 
            .I2(GND_net), .I3(n10635), .O(wr_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF i5747_5748 (.Q(\REG.mem_59_15 ), .C(DEBUG_6_c_c), .D(n5703));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5744_5745 (.Q(\REG.mem_59_14 ), .C(DEBUG_6_c_c), .D(n5702));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5741_5742 (.Q(\REG.mem_59_13 ), .C(DEBUG_6_c_c), .D(n5701));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5738_5739 (.Q(\REG.mem_59_12 ), .C(DEBUG_6_c_c), .D(n5700));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5735_5736 (.Q(\REG.mem_59_11 ), .C(DEBUG_6_c_c), .D(n5699));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5732_5733 (.Q(\REG.mem_59_10 ), .C(DEBUG_6_c_c), .D(n5698));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5729_5730 (.Q(\REG.mem_59_9 ), .C(DEBUG_6_c_c), .D(n5697));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5726_5727 (.Q(\REG.mem_59_8 ), .C(DEBUG_6_c_c), .D(n5696));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5723_5724 (.Q(\REG.mem_59_7 ), .C(DEBUG_6_c_c), .D(n5695));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5720_5721 (.Q(\REG.mem_59_6 ), .C(DEBUG_6_c_c), .D(n5694));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5717_5718 (.Q(\REG.mem_59_5 ), .C(DEBUG_6_c_c), .D(n5693));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5714_5715 (.Q(\REG.mem_59_4 ), .C(DEBUG_6_c_c), .D(n5692));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5711_5712 (.Q(\REG.mem_59_3 ), .C(DEBUG_6_c_c), .D(n5691));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5708_5709 (.Q(\REG.mem_59_2 ), .C(DEBUG_6_c_c), .D(n5690));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5705_5706 (.Q(\REG.mem_59_1 ), .C(DEBUG_6_c_c), .D(n5689));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_6 (.CI(n10622), .I0(wp_sync_w[4]), 
            .I1(n1_adj_1173[4]), .CO(n10623));
    SB_LUT4 i3843_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_22_3 ), .O(n5045));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3843_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_5_lut (.I0(n6), .I1(wp_sync_w[3]), 
            .I2(n1_adj_1173[3]), .I3(n10621), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY wr_addr_r_6__I_0_141_7 (.CI(n10635), .I0(wr_addr_r[5]), .I1(GND_net), 
            .CO(n10636));
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_5 (.CI(n10621), .I0(wp_sync_w[3]), 
            .I1(n1_adj_1173[3]), .CO(n10622));
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_4_lut (.I0(GND_net), .I1(wp_sync_w[2]), 
            .I2(n1_adj_1173[2]), .I3(n10620), .O(rd_sig_diff0_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wr_addr_r_6__I_0_141_6_lut (.I0(GND_net), .I1(wr_addr_r[4]), 
            .I2(GND_net), .I3(n10634), .O(wr_addr_p1_w[4])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_4 (.CI(n10620), .I0(wp_sync_w[2]), 
            .I1(n1_adj_1173[2]), .CO(n10621));
    SB_LUT4 i9927_3_lut (.I0(n13433), .I1(n13415), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11576));
    defparam i9927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9928_3_lut (.I0(n13223), .I1(n11576), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n11577));
    defparam i9928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10021_3_lut (.I0(n13313), .I1(n14189), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n11670));
    defparam i10021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13190_bdd_4_lut (.I0(n13190), .I1(n12248), .I2(n12247), .I3(rd_addr_r[2]), 
            .O(n13193));
    defparam n13190_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9994_3_lut (.I0(n13295), .I1(n14255), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n11643));
    defparam i9994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_3_lut (.I0(GND_net), .I1(wp_sync_w[1]), 
            .I2(n1_adj_1173[1]), .I3(n10619), .O(\rd_sig_diff0_w[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF i5702_5703 (.Q(\REG.mem_59_0 ), .C(DEBUG_6_c_c), .D(n5688));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3842_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_22_2 ), .O(n5044));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3842_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF rp_sync2_r__i1 (.Q(rp_sync2_r[1]), .C(DEBUG_6_c_c), .D(n5686));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i2 (.Q(rp_sync2_r[2]), .C(DEBUG_6_c_c), .D(n5685));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i3 (.Q(rp_sync2_r[3]), .C(DEBUG_6_c_c), .D(n5684));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i4 (.Q(rp_sync2_r[4]), .C(DEBUG_6_c_c), .D(n5683));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i5651_5652 (.Q(\REG.mem_58_15 ), .C(DEBUG_6_c_c), .D(n5682));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5648_5649 (.Q(\REG.mem_58_14 ), .C(DEBUG_6_c_c), .D(n5681));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5645_5646 (.Q(\REG.mem_58_13 ), .C(DEBUG_6_c_c), .D(n5680));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5642_5643 (.Q(\REG.mem_58_12 ), .C(DEBUG_6_c_c), .D(n5679));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5639_5640 (.Q(\REG.mem_58_11 ), .C(DEBUG_6_c_c), .D(n5678));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5636_5637 (.Q(\REG.mem_58_10 ), .C(DEBUG_6_c_c), .D(n5677));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5633_5634 (.Q(\REG.mem_58_9 ), .C(DEBUG_6_c_c), .D(n5676));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5630_5631 (.Q(\REG.mem_58_8 ), .C(DEBUG_6_c_c), .D(n5675));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5627_5628 (.Q(\REG.mem_58_7 ), .C(DEBUG_6_c_c), .D(n5674));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5624_5625 (.Q(\REG.mem_58_6 ), .C(DEBUG_6_c_c), .D(n5673));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12083 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_7 ), 
            .I2(\REG.mem_27_7 ), .I3(rd_addr_r[1]), .O(n13922));
    defparam rd_addr_r_0__bdd_4_lut_12083.LUT_INIT = 16'he4aa;
    SB_LUT4 i3841_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_22_1 ), .O(n5043));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3841_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13922_bdd_4_lut (.I0(n13922), .I1(\REG.mem_25_7 ), .I2(\REG.mem_24_7 ), 
            .I3(rd_addr_r[1]), .O(n12165));
    defparam n13922_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY wr_addr_r_6__I_0_141_6 (.CI(n10634), .I0(wr_addr_r[4]), .I1(GND_net), 
            .CO(n10635));
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_3 (.CI(n10619), .I0(wp_sync_w[1]), 
            .I1(n1_adj_1173[1]), .CO(n10620));
    SB_LUT4 wp_sync2_r_6__I_0_149_add_2_2_lut (.I0(GND_net), .I1(wp_sync_w[0]), 
            .I2(n1_adj_1173[0]), .I3(VCC_net), .O(\rd_sig_diff0_w[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam wp_sync2_r_6__I_0_149_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 wr_addr_r_6__I_0_141_5_lut (.I0(GND_net), .I1(wr_addr_r[3]), 
            .I2(GND_net), .I3(n10633), .O(wr_addr_p1_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY wp_sync2_r_6__I_0_149_add_2_2 (.CI(VCC_net), .I0(wp_sync_w[0]), 
            .I1(n1_adj_1173[0]), .CO(n10619));
    SB_LUT4 i10004_3_lut (.I0(\REG.mem_0_1 ), .I1(\REG.mem_1_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11653));
    defparam i10004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10005_3_lut (.I0(\REG.mem_2_1 ), .I1(\REG.mem_3_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11654));
    defparam i10005_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5621_5622 (.Q(\REG.mem_58_5 ), .C(DEBUG_6_c_c), .D(n5672));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5618_5619 (.Q(\REG.mem_58_4 ), .C(DEBUG_6_c_c), .D(n5671));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5615_5616 (.Q(\REG.mem_58_3 ), .C(DEBUG_6_c_c), .D(n5670));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5612_5613 (.Q(\REG.mem_58_2 ), .C(DEBUG_6_c_c), .D(n5669));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5609_5610 (.Q(\REG.mem_58_1 ), .C(DEBUG_6_c_c), .D(n5668));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5606_5607 (.Q(\REG.mem_58_0 ), .C(DEBUG_6_c_c), .D(n5667));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync2_r__i5 (.Q(rp_sync2_r[5]), .C(DEBUG_6_c_c), .D(n5666));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rp_sync2_r__i6 (.Q(rp_sync2_r[6]), .C(DEBUG_6_c_c), .D(n5665));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(n5664));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .D(n5663));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i3 (.Q(rd_addr_r[3]), .C(SLM_CLK_c), .D(n5662));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i4 (.Q(rd_addr_r[4]), .C(SLM_CLK_c), .D(n5661));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i5 (.Q(rd_addr_r[5]), .C(SLM_CLK_c), .D(n5660));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF rd_addr_r__i6 (.Q(\rd_addr_r[6] ), .C(SLM_CLK_c), .D(n5659));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF i5555_5556 (.Q(\REG.mem_57_15 ), .C(DEBUG_6_c_c), .D(n5658));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFE \REG.out_raw__i16  (.Q(\REG.out_raw[15] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [15]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i15  (.Q(\REG.out_raw[14] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [14]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i14  (.Q(\REG.out_raw[13] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [13]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i13  (.Q(\REG.out_raw[12] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [12]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_CARRY wr_addr_r_6__I_0_141_5 (.CI(n10633), .I0(wr_addr_r[3]), .I1(GND_net), 
            .CO(n10634));
    SB_DFFE \REG.out_raw__i12  (.Q(\REG.out_raw[11] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [11]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i11  (.Q(\REG.out_raw[10] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [10]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i10  (.Q(\REG.out_raw[9] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [9]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i9  (.Q(\REG.out_raw[8] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [8]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i8  (.Q(\REG.out_raw[7] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [7]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i7  (.Q(\REG.out_raw[6] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [6]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_LUT4 wr_addr_r_6__I_0_141_4_lut (.I0(GND_net), .I1(wr_addr_r[2]), 
            .I2(GND_net), .I3(n10632), .O(wr_addr_p1_w[2])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \REG.out_raw__i6  (.Q(\REG.out_raw[5] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [5]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i5  (.Q(\REG.out_raw[4] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [4]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i4  (.Q(\REG.out_raw[3] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [3]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i3  (.Q(\REG.out_raw[2] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [2]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFFE \REG.out_raw__i2  (.Q(\REG.out_raw[1] ), .C(SLM_CLK_c), .E(t_rd_fifo_en_w), 
            .D(\REG.out_raw_31__N_526 [1]));   // src/fifo_dc_32_lut_gen.v(893[25] 899[28])
    SB_DFF i5552_5553 (.Q(\REG.mem_57_14 ), .C(DEBUG_6_c_c), .D(n5657));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5549_5550 (.Q(\REG.mem_57_13 ), .C(DEBUG_6_c_c), .D(n5656));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5546_5547 (.Q(\REG.mem_57_12 ), .C(DEBUG_6_c_c), .D(n5655));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5543_5544 (.Q(\REG.mem_57_11 ), .C(DEBUG_6_c_c), .D(n5654));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5540_5541 (.Q(\REG.mem_57_10 ), .C(DEBUG_6_c_c), .D(n5653));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5537_5538 (.Q(\REG.mem_57_9 ), .C(DEBUG_6_c_c), .D(n5652));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5534_5535 (.Q(\REG.mem_57_8 ), .C(DEBUG_6_c_c), .D(n5651));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5531_5532 (.Q(\REG.mem_57_7 ), .C(DEBUG_6_c_c), .D(n5650));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5528_5529 (.Q(\REG.mem_57_6 ), .C(DEBUG_6_c_c), .D(n5649));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5525_5526 (.Q(\REG.mem_57_5 ), .C(DEBUG_6_c_c), .D(n5648));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5522_5523 (.Q(\REG.mem_57_4 ), .C(DEBUG_6_c_c), .D(n5647));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5519_5520 (.Q(\REG.mem_57_3 ), .C(DEBUG_6_c_c), .D(n5646));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5516_5517 (.Q(\REG.mem_57_2 ), .C(DEBUG_6_c_c), .D(n5645));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5513_5514 (.Q(\REG.mem_57_1 ), .C(DEBUG_6_c_c), .D(n5644));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5510_5511 (.Q(\REG.mem_57_0 ), .C(DEBUG_6_c_c), .D(n5643));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5459_5460 (.Q(\REG.mem_56_15 ), .C(DEBUG_6_c_c), .D(n5642));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5456_5457 (.Q(\REG.mem_56_14 ), .C(DEBUG_6_c_c), .D(n5641));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12078 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_7 ), 
            .I2(\REG.mem_31_7 ), .I3(rd_addr_r[1]), .O(n13916));
    defparam rd_addr_r_0__bdd_4_lut_12078.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11480 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_11 ), 
            .I2(\REG.mem_43_11 ), .I3(rd_addr_r[1]), .O(n13184));
    defparam rd_addr_r_0__bdd_4_lut_11480.LUT_INIT = 16'he4aa;
    SB_LUT4 n13184_bdd_4_lut (.I0(n13184), .I1(\REG.mem_41_11 ), .I2(\REG.mem_40_11 ), 
            .I3(rd_addr_r[1]), .O(n13187));
    defparam n13184_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i131_2_lut_3_lut (.I0(n35), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n2));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i131_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i10008_3_lut (.I0(\REG.mem_6_1 ), .I1(\REG.mem_7_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11657));
    defparam i10008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13916_bdd_4_lut (.I0(n13916), .I1(\REG.mem_29_7 ), .I2(\REG.mem_28_7 ), 
            .I3(rd_addr_r[1]), .O(n12168));
    defparam n13916_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10007_3_lut (.I0(\REG.mem_4_1 ), .I1(\REG.mem_5_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11656));
    defparam i10007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3840_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_22_0 ), .O(n5042));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3840_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11465 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_4 ), 
            .I2(\REG.mem_39_4 ), .I3(rd_addr_r[1]), .O(n13178));
    defparam rd_addr_r_0__bdd_4_lut_11465.LUT_INIT = 16'he4aa;
    SB_LUT4 i10028_3_lut (.I0(\REG.mem_16_1 ), .I1(\REG.mem_17_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11677));
    defparam i10028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13178_bdd_4_lut (.I0(n13178), .I1(\REG.mem_37_4 ), .I2(\REG.mem_36_4 ), 
            .I3(rd_addr_r[1]), .O(n13181));
    defparam n13178_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12073 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_2 ), 
            .I2(\REG.mem_55_2 ), .I3(rd_addr_r[1]), .O(n13910));
    defparam rd_addr_r_0__bdd_4_lut_12073.LUT_INIT = 16'he4aa;
    SB_LUT4 n13910_bdd_4_lut (.I0(n13910), .I1(\REG.mem_53_2 ), .I2(\REG.mem_52_2 ), 
            .I3(rd_addr_r[1]), .O(n13913));
    defparam n13910_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i5453_5454 (.Q(\REG.mem_56_13 ), .C(DEBUG_6_c_c), .D(n5640));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10029_3_lut (.I0(\REG.mem_18_1 ), .I1(\REG.mem_19_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11678));
    defparam i10029_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i5450_5451 (.Q(\REG.mem_56_12 ), .C(DEBUG_6_c_c), .D(n5639));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5447_5448 (.Q(\REG.mem_56_11 ), .C(DEBUG_6_c_c), .D(n5638));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5444_5445 (.Q(\REG.mem_56_10 ), .C(DEBUG_6_c_c), .D(n5637));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5441_5442 (.Q(\REG.mem_56_9 ), .C(DEBUG_6_c_c), .D(n5636));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5438_5439 (.Q(\REG.mem_56_8 ), .C(DEBUG_6_c_c), .D(n5635));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5435_5436 (.Q(\REG.mem_56_7 ), .C(DEBUG_6_c_c), .D(n5634));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5432_5433 (.Q(\REG.mem_56_6 ), .C(DEBUG_6_c_c), .D(n5633));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5429_5430 (.Q(\REG.mem_56_5 ), .C(DEBUG_6_c_c), .D(n5632));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5426_5427 (.Q(\REG.mem_56_4 ), .C(DEBUG_6_c_c), .D(n5631));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5423_5424 (.Q(\REG.mem_56_3 ), .C(DEBUG_6_c_c), .D(n5630));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5420_5421 (.Q(\REG.mem_56_2 ), .C(DEBUG_6_c_c), .D(n5629));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5417_5418 (.Q(\REG.mem_56_1 ), .C(DEBUG_6_c_c), .D(n5628));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5414_5415 (.Q(\REG.mem_56_0 ), .C(DEBUG_6_c_c), .D(n5627));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5363_5364 (.Q(\REG.mem_55_15 ), .C(DEBUG_6_c_c), .D(n5626));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12068 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_13 ), 
            .I2(\REG.mem_35_13 ), .I3(rd_addr_r[1]), .O(n13904));
    defparam rd_addr_r_0__bdd_4_lut_12068.LUT_INIT = 16'he4aa;
    SB_LUT4 i10032_3_lut (.I0(\REG.mem_22_1 ), .I1(\REG.mem_23_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11681));
    defparam i10032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10031_3_lut (.I0(\REG.mem_20_1 ), .I1(\REG.mem_21_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11680));
    defparam i10031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13904_bdd_4_lut (.I0(n13904), .I1(\REG.mem_33_13 ), .I2(\REG.mem_32_13 ), 
            .I3(rd_addr_r[1]), .O(n12174));
    defparam n13904_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11500 (.I0(rd_addr_r[3]), .I1(n12911), 
            .I2(n11495), .I3(rd_addr_r[4]), .O(n13172));
    defparam rd_addr_r_3__bdd_4_lut_11500.LUT_INIT = 16'he4aa;
    SB_LUT4 n13172_bdd_4_lut (.I0(n13172), .I1(n11492), .I2(n12863), .I3(rd_addr_r[4]), 
            .O(n13175));
    defparam n13172_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12063 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_10 ), 
            .I2(\REG.mem_31_10 ), .I3(rd_addr_r[1]), .O(n13898));
    defparam rd_addr_r_0__bdd_4_lut_12063.LUT_INIT = 16'he4aa;
    SB_DFF i5360_5361 (.Q(\REG.mem_55_14 ), .C(DEBUG_6_c_c), .D(n5625));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5357_5358 (.Q(\REG.mem_55_13 ), .C(DEBUG_6_c_c), .D(n5624));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5354_5355 (.Q(\REG.mem_55_12 ), .C(DEBUG_6_c_c), .D(n5623));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5351_5352 (.Q(\REG.mem_55_11 ), .C(DEBUG_6_c_c), .D(n5622));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5348_5349 (.Q(\REG.mem_55_10 ), .C(DEBUG_6_c_c), .D(n5621));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5345_5346 (.Q(\REG.mem_55_9 ), .C(DEBUG_6_c_c), .D(n5620));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5342_5343 (.Q(\REG.mem_55_8 ), .C(DEBUG_6_c_c), .D(n5619));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5339_5340 (.Q(\REG.mem_55_7 ), .C(DEBUG_6_c_c), .D(n5618));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5336_5337 (.Q(\REG.mem_55_6 ), .C(DEBUG_6_c_c), .D(n5617));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5333_5334 (.Q(\REG.mem_55_5 ), .C(DEBUG_6_c_c), .D(n5616));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5330_5331 (.Q(\REG.mem_55_4 ), .C(DEBUG_6_c_c), .D(n5615));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5327_5328 (.Q(\REG.mem_55_3 ), .C(DEBUG_6_c_c), .D(n5614));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5324_5325 (.Q(\REG.mem_55_2 ), .C(DEBUG_6_c_c), .D(n5613));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5321_5322 (.Q(\REG.mem_55_1 ), .C(DEBUG_6_c_c), .D(n5612));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF \REG.out_buffer__i13  (.Q(\fifo_data_out[13] ), .C(SLM_CLK_c), 
           .D(n11073));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF i5318_5319 (.Q(\REG.mem_55_0 ), .C(DEBUG_6_c_c), .D(n5610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wp_sync1_r__i1 (.Q(wp_sync1_r[1]), .C(SLM_CLK_c), .D(n5609));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11470 (.I0(rd_addr_r[1]), .I1(n12460), 
            .I2(n12461), .I3(rd_addr_r[2]), .O(n13166));
    defparam rd_addr_r_1__bdd_4_lut_11470.LUT_INIT = 16'he4aa;
    SB_LUT4 n13166_bdd_4_lut (.I0(n13166), .I1(n12446), .I2(n12445), .I3(rd_addr_r[2]), 
            .O(n13169));
    defparam n13166_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i164_165 (.Q(\REG.mem_1_10 ), .C(DEBUG_6_c_c), .D(n4604));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wp_sync1_r__i2 (.Q(wp_sync1_r[2]), .C(SLM_CLK_c), .D(n5608));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 n13898_bdd_4_lut (.I0(n13898), .I1(\REG.mem_29_10 ), .I2(\REG.mem_28_10 ), 
            .I3(rd_addr_r[1]), .O(n13901));
    defparam n13898_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF wp_sync1_r__i3 (.Q(wp_sync1_r[3]), .C(SLM_CLK_c), .D(n5607));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 i3887_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_24_15 ), .O(n5089));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3887_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wp_sync1_r__i4 (.Q(wp_sync1_r[4]), .C(SLM_CLK_c), .D(n5606));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i5 (.Q(wp_sync1_r[5]), .C(SLM_CLK_c), .D(n5605));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync1_r__i6 (.Q(wp_sync1_r[6]), .C(SLM_CLK_c), .D(n5604));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 i3886_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_24_14 ), .O(n5088));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3886_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF wp_sync2_r__i1 (.Q(wp_sync2_r[1]), .C(SLM_CLK_c), .D(n5603));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i5267_5268 (.Q(\REG.mem_54_15 ), .C(DEBUG_6_c_c), .D(n5602));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5264_5265 (.Q(\REG.mem_54_14 ), .C(DEBUG_6_c_c), .D(n5601));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5261_5262 (.Q(\REG.mem_54_13 ), .C(DEBUG_6_c_c), .D(n5600));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5258_5259 (.Q(\REG.mem_54_12 ), .C(DEBUG_6_c_c), .D(n5599));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5255_5256 (.Q(\REG.mem_54_11 ), .C(DEBUG_6_c_c), .D(n5598));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5252_5253 (.Q(\REG.mem_54_10 ), .C(DEBUG_6_c_c), .D(n5597));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5249_5250 (.Q(\REG.mem_54_9 ), .C(DEBUG_6_c_c), .D(n5596));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5246_5247 (.Q(\REG.mem_54_8 ), .C(DEBUG_6_c_c), .D(n5595));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5243_5244 (.Q(\REG.mem_54_7 ), .C(DEBUG_6_c_c), .D(n5594));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5240_5241 (.Q(\REG.mem_54_6 ), .C(DEBUG_6_c_c), .D(n5593));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5237_5238 (.Q(\REG.mem_54_5 ), .C(DEBUG_6_c_c), .D(n5592));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5234_5235 (.Q(\REG.mem_54_4 ), .C(DEBUG_6_c_c), .D(n5591));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5231_5232 (.Q(\REG.mem_54_3 ), .C(DEBUG_6_c_c), .D(n5590));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5228_5229 (.Q(\REG.mem_54_2 ), .C(DEBUG_6_c_c), .D(n5589));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5225_5226 (.Q(\REG.mem_54_1 ), .C(DEBUG_6_c_c), .D(n5588));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5222_5223 (.Q(\REG.mem_54_0 ), .C(DEBUG_6_c_c), .D(n5587));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wp_sync2_r__i2 (.Q(wp_sync2_r[2]), .C(SLM_CLK_c), .D(n5586));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_LUT4 i10049_3_lut (.I0(\REG.mem_32_1 ), .I1(\REG.mem_33_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11698));
    defparam i10049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12088 (.I0(rd_addr_r[1]), .I1(n11740), 
            .I2(n11741), .I3(rd_addr_r[2]), .O(n13892));
    defparam rd_addr_r_1__bdd_4_lut_12088.LUT_INIT = 16'he4aa;
    SB_LUT4 i10050_3_lut (.I0(\REG.mem_34_1 ), .I1(\REG.mem_35_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11699));
    defparam i10050_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF wp_sync2_r__i3 (.Q(wp_sync2_r[3]), .C(SLM_CLK_c), .D(n5585));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i4 (.Q(wp_sync2_r[4]), .C(SLM_CLK_c), .D(n5584));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i5 (.Q(wp_sync2_r[5]), .C(SLM_CLK_c), .D(n5583));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF wp_sync2_r__i6 (.Q(wp_sync2_r[6]), .C(SLM_CLK_c), .D(n5582));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF \REG.out_buffer__i14  (.Q(\fifo_data_out[14] ), .C(SLM_CLK_c), 
           .D(n11071));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF i5171_5172 (.Q(\REG.mem_53_15 ), .C(DEBUG_6_c_c), .D(n5580));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5168_5169 (.Q(\REG.mem_53_14 ), .C(DEBUG_6_c_c), .D(n5579));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5165_5166 (.Q(\REG.mem_53_13 ), .C(DEBUG_6_c_c), .D(n5578));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5162_5163 (.Q(\REG.mem_53_12 ), .C(DEBUG_6_c_c), .D(n5577));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5159_5160 (.Q(\REG.mem_53_11 ), .C(DEBUG_6_c_c), .D(n5576));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5156_5157 (.Q(\REG.mem_53_10 ), .C(DEBUG_6_c_c), .D(n5575));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5153_5154 (.Q(\REG.mem_53_9 ), .C(DEBUG_6_c_c), .D(n5574));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5150_5151 (.Q(\REG.mem_53_8 ), .C(DEBUG_6_c_c), .D(n5573));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5147_5148 (.Q(\REG.mem_53_7 ), .C(DEBUG_6_c_c), .D(n5572));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5144_5145 (.Q(\REG.mem_53_6 ), .C(DEBUG_6_c_c), .D(n5571));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5141_5142 (.Q(\REG.mem_53_5 ), .C(DEBUG_6_c_c), .D(n5570));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13892_bdd_4_lut (.I0(n13892), .I1(n11726), .I2(n11725), .I3(rd_addr_r[2]), 
            .O(n11765));
    defparam n13892_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3885_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_24_13 ), .O(n5087));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3885_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10053_3_lut (.I0(\REG.mem_38_1 ), .I1(\REG.mem_39_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11702));
    defparam i10053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10052_3_lut (.I0(\REG.mem_36_1 ), .I1(\REG.mem_37_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11701));
    defparam i10052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3884_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_24_12 ), .O(n5086));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3884_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12058 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_2 ), 
            .I2(\REG.mem_7_2 ), .I3(rd_addr_r[1]), .O(n13886));
    defparam rd_addr_r_0__bdd_4_lut_12058.LUT_INIT = 16'he4aa;
    SB_LUT4 i3883_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_24_11 ), .O(n5085));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3883_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5138_5139 (.Q(\REG.mem_53_4 ), .C(DEBUG_6_c_c), .D(n5569));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5135_5136 (.Q(\REG.mem_53_3 ), .C(DEBUG_6_c_c), .D(n5568));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5132_5133 (.Q(\REG.mem_53_2 ), .C(DEBUG_6_c_c), .D(n5567));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5129_5130 (.Q(\REG.mem_53_1 ), .C(DEBUG_6_c_c), .D(n5566));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5126_5127 (.Q(\REG.mem_53_0 ), .C(DEBUG_6_c_c), .D(n5565));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5075_5076 (.Q(\REG.mem_52_15 ), .C(DEBUG_6_c_c), .D(n5564));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5072_5073 (.Q(\REG.mem_52_14 ), .C(DEBUG_6_c_c), .D(n5563));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5069_5070 (.Q(\REG.mem_52_13 ), .C(DEBUG_6_c_c), .D(n5562));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5066_5067 (.Q(\REG.mem_52_12 ), .C(DEBUG_6_c_c), .D(n5561));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5063_5064 (.Q(\REG.mem_52_11 ), .C(DEBUG_6_c_c), .D(n5560));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5060_5061 (.Q(\REG.mem_52_10 ), .C(DEBUG_6_c_c), .D(n5559));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5057_5058 (.Q(\REG.mem_52_9 ), .C(DEBUG_6_c_c), .D(n5558));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5054_5055 (.Q(\REG.mem_52_8 ), .C(DEBUG_6_c_c), .D(n5557));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5051_5052 (.Q(\REG.mem_52_7 ), .C(DEBUG_6_c_c), .D(n5556));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5048_5049 (.Q(\REG.mem_52_6 ), .C(DEBUG_6_c_c), .D(n5555));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5045_5046 (.Q(\REG.mem_52_5 ), .C(DEBUG_6_c_c), .D(n5554));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10445_3_lut (.I0(n13115), .I1(n13019), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12094));
    defparam i10445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11450 (.I0(rd_addr_r[1]), .I1(n12190), 
            .I2(n12191), .I3(rd_addr_r[2]), .O(n13160));
    defparam rd_addr_r_1__bdd_4_lut_11450.LUT_INIT = 16'he4aa;
    SB_LUT4 n13160_bdd_4_lut (.I0(n13160), .I1(n12185), .I2(n12184), .I3(rd_addr_r[2]), 
            .O(n13163));
    defparam n13160_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3882_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_24_10 ), .O(n5084));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3882_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13886_bdd_4_lut (.I0(n13886), .I1(\REG.mem_5_2 ), .I2(\REG.mem_4_2 ), 
            .I3(rd_addr_r[1]), .O(n13889));
    defparam n13886_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY wr_addr_r_6__I_0_141_4 (.CI(n10632), .I0(wr_addr_r[2]), .I1(GND_net), 
            .CO(n10633));
    SB_LUT4 i10446_3_lut (.I0(n12941), .I1(n12815), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12095));
    defparam i10446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wr_addr_r_6__I_0_141_3_lut (.I0(GND_net), .I1(wr_addr_r[1]), 
            .I2(GND_net), .I3(n10631), .O(wr_addr_p1_w[1])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11565 (.I0(rd_addr_r[2]), .I1(n12453), 
            .I2(n12456), .I3(rd_addr_r[3]), .O(n13154));
    defparam rd_addr_r_2__bdd_4_lut_11565.LUT_INIT = 16'he4aa;
    SB_DFF i5042_5043 (.Q(\REG.mem_52_4 ), .C(DEBUG_6_c_c), .D(n5553));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3881_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_24_9 ), .O(n5083));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3881_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i5039_5040 (.Q(\REG.mem_52_3 ), .C(DEBUG_6_c_c), .D(n5552));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5036_5037 (.Q(\REG.mem_52_2 ), .C(DEBUG_6_c_c), .D(n5551));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5033_5034 (.Q(\REG.mem_52_1 ), .C(DEBUG_6_c_c), .D(n5550));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i5030_5031 (.Q(\REG.mem_52_0 ), .C(DEBUG_6_c_c), .D(n5549));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4979_4980 (.Q(\REG.mem_51_15 ), .C(DEBUG_6_c_c), .D(n5548));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4976_4977 (.Q(\REG.mem_51_14 ), .C(DEBUG_6_c_c), .D(n5547));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4973_4974 (.Q(\REG.mem_51_13 ), .C(DEBUG_6_c_c), .D(n5546));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4970_4971 (.Q(\REG.mem_51_12 ), .C(DEBUG_6_c_c), .D(n5545));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4967_4968 (.Q(\REG.mem_51_11 ), .C(DEBUG_6_c_c), .D(n5544));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4964_4965 (.Q(\REG.mem_51_10 ), .C(DEBUG_6_c_c), .D(n5543));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4961_4962 (.Q(\REG.mem_51_9 ), .C(DEBUG_6_c_c), .D(n5542));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4958_4959 (.Q(\REG.mem_51_8 ), .C(DEBUG_6_c_c), .D(n5541));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4955_4956 (.Q(\REG.mem_51_7 ), .C(DEBUG_6_c_c), .D(n5540));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4952_4953 (.Q(\REG.mem_51_6 ), .C(DEBUG_6_c_c), .D(n5539));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4949_4950 (.Q(\REG.mem_51_5 ), .C(DEBUG_6_c_c), .D(n5538));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12048 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_7 ), 
            .I2(\REG.mem_35_7 ), .I3(rd_addr_r[1]), .O(n13880));
    defparam rd_addr_r_0__bdd_4_lut_12048.LUT_INIT = 16'he4aa;
    SB_LUT4 n13154_bdd_4_lut (.I0(n13154), .I1(n12887), .I2(n12953), .I3(rd_addr_r[3]), 
            .O(n13157));
    defparam n13154_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13880_bdd_4_lut (.I0(n13880), .I1(\REG.mem_33_7 ), .I2(\REG.mem_32_7 ), 
            .I3(rd_addr_r[1]), .O(n12177));
    defparam n13880_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4946_4947 (.Q(\REG.mem_51_4 ), .C(DEBUG_6_c_c), .D(n5537));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4943_4944 (.Q(\REG.mem_51_3 ), .C(DEBUG_6_c_c), .D(n5536));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4940_4941 (.Q(\REG.mem_51_2 ), .C(DEBUG_6_c_c), .D(n5535));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4937_4938 (.Q(\REG.mem_51_1 ), .C(DEBUG_6_c_c), .D(n5534));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4934_4935 (.Q(\REG.mem_51_0 ), .C(DEBUG_6_c_c), .D(n5533));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4883_4884 (.Q(\REG.mem_50_15 ), .C(DEBUG_6_c_c), .D(n5532));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10070_3_lut (.I0(\REG.mem_48_1 ), .I1(\REG.mem_49_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11719));
    defparam i10070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3880_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_24_8 ), .O(n5082));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3880_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4880_4881 (.Q(\REG.mem_50_14 ), .C(DEBUG_6_c_c), .D(n5531));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4877_4878 (.Q(\REG.mem_50_13 ), .C(DEBUG_6_c_c), .D(n5530));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4874_4875 (.Q(\REG.mem_50_12 ), .C(DEBUG_6_c_c), .D(n5529));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4871_4872 (.Q(\REG.mem_50_11 ), .C(DEBUG_6_c_c), .D(n5528));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4868_4869 (.Q(\REG.mem_50_10 ), .C(DEBUG_6_c_c), .D(n5527));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4865_4866 (.Q(\REG.mem_50_9 ), .C(DEBUG_6_c_c), .D(n5526));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4862_4863 (.Q(\REG.mem_50_8 ), .C(DEBUG_6_c_c), .D(n5525));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4859_4860 (.Q(\REG.mem_50_7 ), .C(DEBUG_6_c_c), .D(n5524));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4856_4857 (.Q(\REG.mem_50_6 ), .C(DEBUG_6_c_c), .D(n5523));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4853_4854 (.Q(\REG.mem_50_5 ), .C(DEBUG_6_c_c), .D(n5522));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4850_4851 (.Q(\REG.mem_50_4 ), .C(DEBUG_6_c_c), .D(n5521));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4847_4848 (.Q(\REG.mem_50_3 ), .C(DEBUG_6_c_c), .D(n5520));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4844_4845 (.Q(\REG.mem_50_2 ), .C(DEBUG_6_c_c), .D(n5519));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4841_4842 (.Q(\REG.mem_50_1 ), .C(DEBUG_6_c_c), .D(n5518));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4838_4839 (.Q(\REG.mem_50_0 ), .C(DEBUG_6_c_c), .D(n5517));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4787_4788 (.Q(\REG.mem_49_15 ), .C(DEBUG_6_c_c), .D(n5516));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4784_4785 (.Q(\REG.mem_49_14 ), .C(DEBUG_6_c_c), .D(n5515));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11216 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_12 ), 
            .I2(\REG.mem_31_12 ), .I3(rd_addr_r[1]), .O(n12878));
    defparam rd_addr_r_0__bdd_4_lut_11216.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12043 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_11 ), 
            .I2(\REG.mem_27_11 ), .I3(rd_addr_r[1]), .O(n13874));
    defparam rd_addr_r_0__bdd_4_lut_12043.LUT_INIT = 16'he4aa;
    SB_LUT4 i3879_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_24_7 ), .O(n5081));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3879_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13874_bdd_4_lut (.I0(n13874), .I1(\REG.mem_25_11 ), .I2(\REG.mem_24_11 ), 
            .I3(rd_addr_r[1]), .O(n13877));
    defparam n13874_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4781_4782 (.Q(\REG.mem_49_13 ), .C(DEBUG_6_c_c), .D(n5514));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4778_4779 (.Q(\REG.mem_49_12 ), .C(DEBUG_6_c_c), .D(n5513));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4775_4776 (.Q(\REG.mem_49_11 ), .C(DEBUG_6_c_c), .D(n5512));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4772_4773 (.Q(\REG.mem_49_10 ), .C(DEBUG_6_c_c), .D(n5511));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4769_4770 (.Q(\REG.mem_49_9 ), .C(DEBUG_6_c_c), .D(n5510));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4766_4767 (.Q(\REG.mem_49_8 ), .C(DEBUG_6_c_c), .D(n5509));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4763_4764 (.Q(\REG.mem_49_7 ), .C(DEBUG_6_c_c), .D(n5508));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4760_4761 (.Q(\REG.mem_49_6 ), .C(DEBUG_6_c_c), .D(n5507));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4757_4758 (.Q(\REG.mem_49_5 ), .C(DEBUG_6_c_c), .D(n5506));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4754_4755 (.Q(\REG.mem_49_4 ), .C(DEBUG_6_c_c), .D(n5505));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4751_4752 (.Q(\REG.mem_49_3 ), .C(DEBUG_6_c_c), .D(n5504));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4748_4749 (.Q(\REG.mem_49_2 ), .C(DEBUG_6_c_c), .D(n5503));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4745_4746 (.Q(\REG.mem_49_1 ), .C(DEBUG_6_c_c), .D(n5502));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4742_4743 (.Q(\REG.mem_49_0 ), .C(DEBUG_6_c_c), .D(n5501));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11460 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_0 ), 
            .I2(\REG.mem_31_0 ), .I3(rd_addr_r[1]), .O(n13148));
    defparam rd_addr_r_0__bdd_4_lut_11460.LUT_INIT = 16'he4aa;
    SB_LUT4 i10071_3_lut (.I0(\REG.mem_50_1 ), .I1(\REG.mem_51_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11720));
    defparam i10071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13148_bdd_4_lut (.I0(n13148), .I1(\REG.mem_29_0 ), .I2(\REG.mem_28_0 ), 
            .I3(rd_addr_r[1]), .O(n13151));
    defparam n13148_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3878_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_24_6 ), .O(n5080));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3878_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10074_3_lut (.I0(\REG.mem_54_1 ), .I1(\REG.mem_55_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11723));
    defparam i10074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12878_bdd_4_lut (.I0(n12878), .I1(\REG.mem_29_12 ), .I2(\REG.mem_28_12 ), 
            .I3(rd_addr_r[1]), .O(n12881));
    defparam n12878_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i53_54 (.Q(\REG.mem_0_5 ), .C(DEBUG_6_c_c), .D(n4691));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12038 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_4 ), 
            .I2(\REG.mem_27_4 ), .I3(rd_addr_r[1]), .O(n13868));
    defparam rd_addr_r_0__bdd_4_lut_12038.LUT_INIT = 16'he4aa;
    SB_DFF i173_174 (.Q(\REG.mem_1_13 ), .C(DEBUG_6_c_c), .D(n4690));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10073_3_lut (.I0(\REG.mem_52_1 ), .I1(\REG.mem_53_1 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11722));
    defparam i10073_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i56_57 (.Q(\REG.mem_0_6 ), .C(DEBUG_6_c_c), .D(n4689));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(DEBUG_6_c_c), .D(n5493));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i4691_4692 (.Q(\REG.mem_48_15 ), .C(DEBUG_6_c_c), .D(n5492));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(DEBUG_6_c_c), .D(n5491));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i4688_4689 (.Q(\REG.mem_48_14 ), .C(DEBUG_6_c_c), .D(n5490));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4685_4686 (.Q(\REG.mem_48_13 ), .C(DEBUG_6_c_c), .D(n5489));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4682_4683 (.Q(\REG.mem_48_12 ), .C(DEBUG_6_c_c), .D(n5488));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4679_4680 (.Q(\REG.mem_48_11 ), .C(DEBUG_6_c_c), .D(n5487));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4676_4677 (.Q(\REG.mem_48_10 ), .C(DEBUG_6_c_c), .D(n5486));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4673_4674 (.Q(\REG.mem_48_9 ), .C(DEBUG_6_c_c), .D(n5485));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4670_4671 (.Q(\REG.mem_48_8 ), .C(DEBUG_6_c_c), .D(n5484));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4667_4668 (.Q(\REG.mem_48_7 ), .C(DEBUG_6_c_c), .D(n5483));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3877_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_24_5 ), .O(n5079));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3877_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3876_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_24_4 ), .O(n5078));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3876_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i59_60 (.Q(\REG.mem_0_7 ), .C(DEBUG_6_c_c), .D(n4688));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i62_63 (.Q(\REG.mem_0_8 ), .C(DEBUG_6_c_c), .D(n4687));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3875_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_24_3 ), .O(n5077));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3875_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11231 (.I0(rd_addr_r[2]), .I1(n11598), 
            .I2(n11625), .I3(rd_addr_r[3]), .O(n12806));
    defparam rd_addr_r_2__bdd_4_lut_11231.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11435 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_10 ), 
            .I2(\REG.mem_47_10 ), .I3(rd_addr_r[1]), .O(n13142));
    defparam rd_addr_r_0__bdd_4_lut_11435.LUT_INIT = 16'he4aa;
    SB_DFF i4664_4665 (.Q(\REG.mem_48_6 ), .C(DEBUG_6_c_c), .D(n5482));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3874_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_24_2 ), .O(n5076));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3874_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13868_bdd_4_lut (.I0(n13868), .I1(\REG.mem_25_4 ), .I2(\REG.mem_24_4 ), 
            .I3(rd_addr_r[1]), .O(n13871));
    defparam n13868_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i4661_4662 (.Q(\REG.mem_48_5 ), .C(DEBUG_6_c_c), .D(n5481));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4658_4659 (.Q(\REG.mem_48_4 ), .C(DEBUG_6_c_c), .D(n5480));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4655_4656 (.Q(\REG.mem_48_3 ), .C(DEBUG_6_c_c), .D(n5479));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4652_4653 (.Q(\REG.mem_48_2 ), .C(DEBUG_6_c_c), .D(n5478));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4649_4650 (.Q(\REG.mem_48_1 ), .C(DEBUG_6_c_c), .D(n5477));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4646_4647 (.Q(\REG.mem_48_0 ), .C(DEBUG_6_c_c), .D(n5476));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wr_addr_r__i3 (.Q(wr_addr_r[3]), .C(DEBUG_6_c_c), .D(n5475));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i4 (.Q(wr_addr_r[4]), .C(DEBUG_6_c_c), .D(n5474));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF wr_addr_r__i5 (.Q(wr_addr_r[5]), .C(DEBUG_6_c_c), .D(n5473));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_DFF i4595_4596 (.Q(\REG.mem_47_15 ), .C(DEBUG_6_c_c), .D(n5472));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4592_4593 (.Q(\REG.mem_47_14 ), .C(DEBUG_6_c_c), .D(n5471));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4589_4590 (.Q(\REG.mem_47_13 ), .C(DEBUG_6_c_c), .D(n5470));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4586_4587 (.Q(\REG.mem_47_12 ), .C(DEBUG_6_c_c), .D(n5469));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4583_4584 (.Q(\REG.mem_47_11 ), .C(DEBUG_6_c_c), .D(n5468));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4580_4581 (.Q(\REG.mem_47_10 ), .C(DEBUG_6_c_c), .D(n5467));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12812_bdd_4_lut (.I0(n12812), .I1(\REG.mem_45_0 ), .I2(\REG.mem_44_0 ), 
            .I3(rd_addr_r[1]), .O(n12815));
    defparam n12812_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3873_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_24_1 ), .O(n5075));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3873_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3872_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_24_0 ), .O(n5074));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3872_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3903_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_25_15 ), .O(n5105));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3903_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13142_bdd_4_lut (.I0(n13142), .I1(\REG.mem_45_10 ), .I2(\REG.mem_44_10 ), 
            .I3(rd_addr_r[1]), .O(n13145));
    defparam n13142_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3902_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_25_14 ), .O(n5104));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3902_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3901_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_25_13 ), .O(n5103));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3901_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4577_4578 (.Q(\REG.mem_47_9 ), .C(DEBUG_6_c_c), .D(n5466));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4574_4575 (.Q(\REG.mem_47_8 ), .C(DEBUG_6_c_c), .D(n5465));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4571_4572 (.Q(\REG.mem_47_7 ), .C(DEBUG_6_c_c), .D(n5464));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4568_4569 (.Q(\REG.mem_47_6 ), .C(DEBUG_6_c_c), .D(n5463));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4565_4566 (.Q(\REG.mem_47_5 ), .C(DEBUG_6_c_c), .D(n5462));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4562_4563 (.Q(\REG.mem_47_4 ), .C(DEBUG_6_c_c), .D(n5461));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4559_4560 (.Q(\REG.mem_47_3 ), .C(DEBUG_6_c_c), .D(n5460));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4556_4557 (.Q(\REG.mem_47_2 ), .C(DEBUG_6_c_c), .D(n5459));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4553_4554 (.Q(\REG.mem_47_1 ), .C(DEBUG_6_c_c), .D(n5458));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4550_4551 (.Q(\REG.mem_47_0 ), .C(DEBUG_6_c_c), .D(n5457));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4499_4500 (.Q(\REG.mem_46_15 ), .C(DEBUG_6_c_c), .D(n5456));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4496_4497 (.Q(\REG.mem_46_14 ), .C(DEBUG_6_c_c), .D(n5455));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4493_4494 (.Q(\REG.mem_46_13 ), .C(DEBUG_6_c_c), .D(n5454));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4490_4491 (.Q(\REG.mem_46_12 ), .C(DEBUG_6_c_c), .D(n5453));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4487_4488 (.Q(\REG.mem_46_11 ), .C(DEBUG_6_c_c), .D(n5452));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4484_4485 (.Q(\REG.mem_46_10 ), .C(DEBUG_6_c_c), .D(n5451));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3900_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_25_12 ), .O(n5102));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3900_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i65_66 (.Q(\REG.mem_0_9 ), .C(DEBUG_6_c_c), .D(n4684));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i68_69 (.Q(\REG.mem_0_10 ), .C(DEBUG_6_c_c), .D(n4683));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10796_3_lut (.I0(\REG.mem_48_9 ), .I1(\REG.mem_49_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12445));
    defparam i10796_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i71_72 (.Q(\REG.mem_0_11 ), .C(DEBUG_6_c_c), .D(n4682));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i74_75 (.Q(\REG.mem_0_12 ), .C(DEBUG_6_c_c), .D(n4681));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10797_3_lut (.I0(\REG.mem_50_9 ), .I1(\REG.mem_51_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12446));
    defparam i10797_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i77_78 (.Q(\REG.mem_0_13 ), .C(DEBUG_6_c_c), .D(n4680));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i170_171 (.Q(\REG.mem_1_12 ), .C(DEBUG_6_c_c), .D(n4678));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11440 (.I0(rd_addr_r[2]), .I1(n11718), 
            .I2(n11736), .I3(rd_addr_r[3]), .O(n13136));
    defparam rd_addr_r_2__bdd_4_lut_11440.LUT_INIT = 16'he4aa;
    SB_LUT4 n13136_bdd_4_lut (.I0(n13136), .I1(n11709), .I2(n11691), .I3(rd_addr_r[3]), 
            .O(n11898));
    defparam n13136_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i80_81 (.Q(\REG.mem_0_14 ), .C(DEBUG_6_c_c), .D(n4675));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4481_4482 (.Q(\REG.mem_46_9 ), .C(DEBUG_6_c_c), .D(n5450));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4478_4479 (.Q(\REG.mem_46_8 ), .C(DEBUG_6_c_c), .D(n5449));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10812_3_lut (.I0(\REG.mem_54_9 ), .I1(\REG.mem_55_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12461));
    defparam i10812_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i4475_4476 (.Q(\REG.mem_46_7 ), .C(DEBUG_6_c_c), .D(n5448));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4472_4473 (.Q(\REG.mem_46_6 ), .C(DEBUG_6_c_c), .D(n5447));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4469_4470 (.Q(\REG.mem_46_5 ), .C(DEBUG_6_c_c), .D(n5446));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4466_4467 (.Q(\REG.mem_46_4 ), .C(DEBUG_6_c_c), .D(n5445));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4463_4464 (.Q(\REG.mem_46_3 ), .C(DEBUG_6_c_c), .D(n5444));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4460_4461 (.Q(\REG.mem_46_2 ), .C(DEBUG_6_c_c), .D(n5443));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4457_4458 (.Q(\REG.mem_46_1 ), .C(DEBUG_6_c_c), .D(n5442));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4454_4455 (.Q(\REG.mem_46_0 ), .C(DEBUG_6_c_c), .D(n5441));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4403_4404 (.Q(\REG.mem_45_15 ), .C(DEBUG_6_c_c), .D(n5440));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4400_4401 (.Q(\REG.mem_45_14 ), .C(DEBUG_6_c_c), .D(n5439));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4397_4398 (.Q(\REG.mem_45_13 ), .C(DEBUG_6_c_c), .D(n5438));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4394_4395 (.Q(\REG.mem_45_12 ), .C(DEBUG_6_c_c), .D(n5437));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4391_4392 (.Q(\REG.mem_45_11 ), .C(DEBUG_6_c_c), .D(n5436));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4388_4389 (.Q(\REG.mem_45_10 ), .C(DEBUG_6_c_c), .D(n5435));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10811_3_lut (.I0(\REG.mem_52_9 ), .I1(\REG.mem_53_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12460));
    defparam i10811_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i4385_4386 (.Q(\REG.mem_45_9 ), .C(DEBUG_6_c_c), .D(n5434));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3899_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_25_11 ), .O(n5101));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3899_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12033 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_7 ), 
            .I2(\REG.mem_39_7 ), .I3(rd_addr_r[1]), .O(n13862));
    defparam rd_addr_r_0__bdd_4_lut_12033.LUT_INIT = 16'he4aa;
    SB_LUT4 i3898_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_25_10 ), .O(n5100));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3898_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3897_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_25_9 ), .O(n5099));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3897_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11425 (.I0(rd_addr_r[2]), .I1(n11811), 
            .I2(n11820), .I3(rd_addr_r[3]), .O(n13130));
    defparam rd_addr_r_2__bdd_4_lut_11425.LUT_INIT = 16'he4aa;
    SB_LUT4 n13130_bdd_4_lut (.I0(n13130), .I1(n11784), .I2(n11760), .I3(rd_addr_r[3]), 
            .O(n11901));
    defparam n13130_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3896_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_25_8 ), .O(n5098));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3896_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13862_bdd_4_lut (.I0(n13862), .I1(\REG.mem_37_7 ), .I2(\REG.mem_36_7 ), 
            .I3(rd_addr_r[1]), .O(n12180));
    defparam n13862_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11430 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_3 ), 
            .I2(\REG.mem_55_3 ), .I3(rd_addr_r[1]), .O(n13124));
    defparam rd_addr_r_0__bdd_4_lut_11430.LUT_INIT = 16'he4aa;
    SB_DFF i4382_4383 (.Q(\REG.mem_45_8 ), .C(DEBUG_6_c_c), .D(n5433));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4379_4380 (.Q(\REG.mem_45_7 ), .C(DEBUG_6_c_c), .D(n5432));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4376_4377 (.Q(\REG.mem_45_6 ), .C(DEBUG_6_c_c), .D(n5431));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4373_4374 (.Q(\REG.mem_45_5 ), .C(DEBUG_6_c_c), .D(n5430));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4370_4371 (.Q(\REG.mem_45_4 ), .C(DEBUG_6_c_c), .D(n5429));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4367_4368 (.Q(\REG.mem_45_3 ), .C(DEBUG_6_c_c), .D(n5428));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4364_4365 (.Q(\REG.mem_45_2 ), .C(DEBUG_6_c_c), .D(n5427));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4361_4362 (.Q(\REG.mem_45_1 ), .C(DEBUG_6_c_c), .D(n5426));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4358_4359 (.Q(\REG.mem_45_0 ), .C(DEBUG_6_c_c), .D(n5425));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4307_4308 (.Q(\REG.mem_44_15 ), .C(DEBUG_6_c_c), .D(n5424));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4304_4305 (.Q(\REG.mem_44_14 ), .C(DEBUG_6_c_c), .D(n5423));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4301_4302 (.Q(\REG.mem_44_13 ), .C(DEBUG_6_c_c), .D(n5422));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4298_4299 (.Q(\REG.mem_44_12 ), .C(DEBUG_6_c_c), .D(n5421));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4295_4296 (.Q(\REG.mem_44_11 ), .C(DEBUG_6_c_c), .D(n5420));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4292_4293 (.Q(\REG.mem_44_10 ), .C(DEBUG_6_c_c), .D(n5419));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12028 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_0 ), 
            .I2(\REG.mem_11_0 ), .I3(rd_addr_r[1]), .O(n13856));
    defparam rd_addr_r_0__bdd_4_lut_12028.LUT_INIT = 16'he4aa;
    SB_DFF i4289_4290 (.Q(\REG.mem_44_9 ), .C(DEBUG_6_c_c), .D(n5418));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13856_bdd_4_lut (.I0(n13856), .I1(\REG.mem_9_0 ), .I2(\REG.mem_8_0 ), 
            .I3(rd_addr_r[1]), .O(n13859));
    defparam n13856_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3895_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_25_7 ), .O(n5097));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3895_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3894_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_25_6 ), .O(n5096));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3894_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i36_2_lut_3_lut (.I0(n11), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n36));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i36_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF i4286_4287 (.Q(\REG.mem_44_8 ), .C(DEBUG_6_c_c), .D(n5417));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4283_4284 (.Q(\REG.mem_44_7 ), .C(DEBUG_6_c_c), .D(n5416));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4280_4281 (.Q(\REG.mem_44_6 ), .C(DEBUG_6_c_c), .D(n5415));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4277_4278 (.Q(\REG.mem_44_5 ), .C(DEBUG_6_c_c), .D(n5414));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4274_4275 (.Q(\REG.mem_44_4 ), .C(DEBUG_6_c_c), .D(n5413));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4271_4272 (.Q(\REG.mem_44_3 ), .C(DEBUG_6_c_c), .D(n5412));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4268_4269 (.Q(\REG.mem_44_2 ), .C(DEBUG_6_c_c), .D(n5411));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4265_4266 (.Q(\REG.mem_44_1 ), .C(DEBUG_6_c_c), .D(n5410));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4262_4263 (.Q(\REG.mem_44_0 ), .C(DEBUG_6_c_c), .D(n5409));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wr_grey_sync_r__i6 (.Q(wr_grey_sync_r[6]), .C(DEBUG_6_c_c), .D(n5408));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF i4211_4212 (.Q(\REG.mem_43_15 ), .C(DEBUG_6_c_c), .D(n5407));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4208_4209 (.Q(\REG.mem_43_14 ), .C(DEBUG_6_c_c), .D(n5406));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4205_4206 (.Q(\REG.mem_43_13 ), .C(DEBUG_6_c_c), .D(n5405));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4202_4203 (.Q(\REG.mem_43_12 ), .C(DEBUG_6_c_c), .D(n5404));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4199_4200 (.Q(\REG.mem_43_11 ), .C(DEBUG_6_c_c), .D(n5403));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4196_4197 (.Q(\REG.mem_43_10 ), .C(DEBUG_6_c_c), .D(n5402));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13124_bdd_4_lut (.I0(n13124), .I1(\REG.mem_53_3 ), .I2(\REG.mem_52_3 ), 
            .I3(rd_addr_r[1]), .O(n13127));
    defparam n13124_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12023 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_5 ), 
            .I2(\REG.mem_11_5 ), .I3(rd_addr_r[1]), .O(n13850));
    defparam rd_addr_r_0__bdd_4_lut_12023.LUT_INIT = 16'he4aa;
    SB_LUT4 n13850_bdd_4_lut (.I0(n13850), .I1(\REG.mem_9_5 ), .I2(\REG.mem_8_5 ), 
            .I3(rd_addr_r[1]), .O(n13853));
    defparam n13850_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY wr_addr_r_6__I_0_141_3 (.CI(n10631), .I0(wr_addr_r[1]), .I1(GND_net), 
            .CO(n10632));
    SB_LUT4 wr_addr_r_6__I_0_141_2_lut (.I0(GND_net), .I1(\wr_addr_r[0] ), 
            .I2(GND_net), .I3(VCC_net), .O(\wr_addr_p1_w[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_141_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF i4193_4194 (.Q(\REG.mem_43_9 ), .C(DEBUG_6_c_c), .D(n5401));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4190_4191 (.Q(\REG.mem_43_8 ), .C(DEBUG_6_c_c), .D(n5400));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4187_4188 (.Q(\REG.mem_43_7 ), .C(DEBUG_6_c_c), .D(n5399));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4184_4185 (.Q(\REG.mem_43_6 ), .C(DEBUG_6_c_c), .D(n5398));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4181_4182 (.Q(\REG.mem_43_5 ), .C(DEBUG_6_c_c), .D(n5397));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4178_4179 (.Q(\REG.mem_43_4 ), .C(DEBUG_6_c_c), .D(n5396));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4175_4176 (.Q(\REG.mem_43_3 ), .C(DEBUG_6_c_c), .D(n5395));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4172_4173 (.Q(\REG.mem_43_2 ), .C(DEBUG_6_c_c), .D(n5394));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4169_4170 (.Q(\REG.mem_43_1 ), .C(DEBUG_6_c_c), .D(n5393));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4166_4167 (.Q(\REG.mem_43_0 ), .C(DEBUG_6_c_c), .D(n5392));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF \REG.out_buffer__i15  (.Q(\fifo_data_out[15] ), .C(SLM_CLK_c), 
           .D(n11069));   // src/fifo_dc_32_lut_gen.v(922[41] 933[44])
    SB_DFF i4115_4116 (.Q(\REG.mem_42_15 ), .C(DEBUG_6_c_c), .D(n5390));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4112_4113 (.Q(\REG.mem_42_14 ), .C(DEBUG_6_c_c), .D(n5389));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4109_4110 (.Q(\REG.mem_42_13 ), .C(DEBUG_6_c_c), .D(n5388));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4106_4107 (.Q(\REG.mem_42_12 ), .C(DEBUG_6_c_c), .D(n5387));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4103_4104 (.Q(\REG.mem_42_11 ), .C(DEBUG_6_c_c), .D(n5386));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11415 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_4 ), 
            .I2(\REG.mem_43_4 ), .I3(rd_addr_r[1]), .O(n13118));
    defparam rd_addr_r_0__bdd_4_lut_11415.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_r_6__I_0_135_i7_3_lut (.I0(wr_grey_sync_r[6]), .I1(\wr_addr_p1_w[6] ), 
            .I2(n7596), .I3(GND_net), .O(wr_grey_w[6]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3893_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_25_5 ), .O(n5095));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3893_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY wr_addr_r_6__I_0_141_2 (.CI(VCC_net), .I0(\wr_addr_r[0] ), 
            .I1(GND_net), .CO(n10631));
    SB_LUT4 n13118_bdd_4_lut (.I0(n13118), .I1(\REG.mem_41_4 ), .I2(\REG.mem_40_4 ), 
            .I3(rd_addr_r[1]), .O(n13121));
    defparam n13118_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3892_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_25_4 ), .O(n5094));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3892_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4100_4101 (.Q(\REG.mem_42_10 ), .C(DEBUG_6_c_c), .D(n5385));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4097_4098 (.Q(\REG.mem_42_9 ), .C(DEBUG_6_c_c), .D(n5384));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4094_4095 (.Q(\REG.mem_42_8 ), .C(DEBUG_6_c_c), .D(n5383));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4091_4092 (.Q(\REG.mem_42_7 ), .C(DEBUG_6_c_c), .D(n5382));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4088_4089 (.Q(\REG.mem_42_6 ), .C(DEBUG_6_c_c), .D(n5381));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4085_4086 (.Q(\REG.mem_42_5 ), .C(DEBUG_6_c_c), .D(n5380));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4082_4083 (.Q(\REG.mem_42_4 ), .C(DEBUG_6_c_c), .D(n5379));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4079_4080 (.Q(\REG.mem_42_3 ), .C(DEBUG_6_c_c), .D(n5378));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4076_4077 (.Q(\REG.mem_42_2 ), .C(DEBUG_6_c_c), .D(n5377));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4073_4074 (.Q(\REG.mem_42_1 ), .C(DEBUG_6_c_c), .D(n5376));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4070_4071 (.Q(\REG.mem_42_0 ), .C(DEBUG_6_c_c), .D(n5375));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4019_4020 (.Q(\REG.mem_41_15 ), .C(DEBUG_6_c_c), .D(n5374));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4016_4017 (.Q(\REG.mem_41_14 ), .C(DEBUG_6_c_c), .D(n5373));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4013_4014 (.Q(\REG.mem_41_13 ), .C(DEBUG_6_c_c), .D(n5372));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4010_4011 (.Q(\REG.mem_41_12 ), .C(DEBUG_6_c_c), .D(n5371));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i83_84 (.Q(\REG.mem_0_15 ), .C(DEBUG_6_c_c), .D(n4671));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3891_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_25_3 ), .O(n5093));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3891_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3890_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_25_2 ), .O(n5092));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3890_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3889_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_25_1 ), .O(n5091));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3889_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12208 (.I0(rd_addr_r[3]), .I1(n13367), 
            .I2(n11765), .I3(rd_addr_r[4]), .O(n13844));
    defparam rd_addr_r_3__bdd_4_lut_12208.LUT_INIT = 16'he4aa;
    SB_DFF \genblk16.rd_prev_r_132  (.Q(\genblk16.rd_prev_r ), .C(SLM_CLK_c), 
           .D(n4667));   // src/fifo_dc_32_lut_gen.v(751[29] 761[32])
    SB_DFF i137_138 (.Q(\REG.mem_1_1 ), .C(DEBUG_6_c_c), .D(n4666));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3888_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_25_0 ), .O(n5090));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3888_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13844_bdd_4_lut (.I0(n13844), .I1(n11750), .I2(n13361), .I3(rd_addr_r[4]), 
            .O(n13847));
    defparam n13844_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3936_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_27_15 ), .O(n5138));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3936_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i152_153 (.Q(\REG.mem_1_6 ), .C(DEBUG_6_c_c), .D(n4665));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i4007_4008 (.Q(\REG.mem_41_11 ), .C(DEBUG_6_c_c), .D(n5370));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i35_2_lut_3_lut (.I0(n11), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n35));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i35_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3935_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_27_14 ), .O(n5137));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3935_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i4004_4005 (.Q(\REG.mem_41_10 ), .C(DEBUG_6_c_c), .D(n5369));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_r_6__I_0_add_2_8_lut (.I0(n11475), .I1(wr_grey_sync_r[6]), 
            .I2(n1[6]), .I3(n10630), .O(\afull_flag_impl.af_flag_nxt_w )) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_DFF i4001_4002 (.Q(\REG.mem_41_9 ), .C(DEBUG_6_c_c), .D(n5368));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3998_3999 (.Q(\REG.mem_41_8 ), .C(DEBUG_6_c_c), .D(n5367));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3995_3996 (.Q(\REG.mem_41_7 ), .C(DEBUG_6_c_c), .D(n5366));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3992_3993 (.Q(\REG.mem_41_6 ), .C(DEBUG_6_c_c), .D(n5365));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3989_3990 (.Q(\REG.mem_41_5 ), .C(DEBUG_6_c_c), .D(n5364));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3986_3987 (.Q(\REG.mem_41_4 ), .C(DEBUG_6_c_c), .D(n5363));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3983_3984 (.Q(\REG.mem_41_3 ), .C(DEBUG_6_c_c), .D(n5362));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3980_3981 (.Q(\REG.mem_41_2 ), .C(DEBUG_6_c_c), .D(n5361));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3977_3978 (.Q(\REG.mem_41_1 ), .C(DEBUG_6_c_c), .D(n5360));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3974_3975 (.Q(\REG.mem_41_0 ), .C(DEBUG_6_c_c), .D(n5358));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3923_3924 (.Q(\REG.mem_40_15 ), .C(DEBUG_6_c_c), .D(n5357));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3920_3921 (.Q(\REG.mem_40_14 ), .C(DEBUG_6_c_c), .D(n5356));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3917_3918 (.Q(\REG.mem_40_13 ), .C(DEBUG_6_c_c), .D(n5355));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3914_3915 (.Q(\REG.mem_40_12 ), .C(DEBUG_6_c_c), .D(n5354));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12018 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_13 ), 
            .I2(\REG.mem_39_13 ), .I3(rd_addr_r[1]), .O(n13838));
    defparam rd_addr_r_0__bdd_4_lut_12018.LUT_INIT = 16'he4aa;
    SB_LUT4 n13838_bdd_4_lut (.I0(n13838), .I1(\REG.mem_37_13 ), .I2(\REG.mem_36_13 ), 
            .I3(rd_addr_r[1]), .O(n12189));
    defparam n13838_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3934_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_27_13 ), .O(n5136));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3934_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3933_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_27_12 ), .O(n5135));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3933_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3932_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_27_11 ), .O(n5134));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3932_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3931_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_27_10 ), .O(n5133));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3931_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11410 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_0 ), 
            .I2(\REG.mem_35_0 ), .I3(rd_addr_r[1]), .O(n13112));
    defparam rd_addr_r_0__bdd_4_lut_11410.LUT_INIT = 16'he4aa;
    SB_LUT4 i9843_3_lut (.I0(n13235), .I1(n13205), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11492));
    defparam i9843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13112_bdd_4_lut (.I0(n13112), .I1(\REG.mem_33_0 ), .I2(\REG.mem_32_0 ), 
            .I3(rd_addr_r[1]), .O(n13115));
    defparam n13112_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9846_3_lut (.I0(n13031), .I1(n12983), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11495));
    defparam i9846_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i3911_3912 (.Q(\REG.mem_40_11 ), .C(DEBUG_6_c_c), .D(n5353));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3908_3909 (.Q(\REG.mem_40_10 ), .C(DEBUG_6_c_c), .D(n5352));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3905_3906 (.Q(\REG.mem_40_9 ), .C(DEBUG_6_c_c), .D(n5351));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3902_3903 (.Q(\REG.mem_40_8 ), .C(DEBUG_6_c_c), .D(n5350));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3899_3900 (.Q(\REG.mem_40_7 ), .C(DEBUG_6_c_c), .D(n5349));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3896_3897 (.Q(\REG.mem_40_6 ), .C(DEBUG_6_c_c), .D(n5348));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3893_3894 (.Q(\REG.mem_40_5 ), .C(DEBUG_6_c_c), .D(n5347));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3890_3891 (.Q(\REG.mem_40_4 ), .C(DEBUG_6_c_c), .D(n5346));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3887_3888 (.Q(\REG.mem_40_3 ), .C(DEBUG_6_c_c), .D(n5345));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3884_3885 (.Q(\REG.mem_40_2 ), .C(DEBUG_6_c_c), .D(n5344));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3881_3882 (.Q(\REG.mem_40_1 ), .C(DEBUG_6_c_c), .D(n5343));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3878_3879 (.Q(\REG.mem_40_0 ), .C(DEBUG_6_c_c), .D(n5342));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3827_3828 (.Q(\REG.mem_39_15 ), .C(DEBUG_6_c_c), .D(n5341));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3824_3825 (.Q(\REG.mem_39_14 ), .C(DEBUG_6_c_c), .D(n5340));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3821_3822 (.Q(\REG.mem_39_13 ), .C(DEBUG_6_c_c), .D(n5339));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11211 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_5 ), 
            .I2(\REG.mem_23_5 ), .I3(rd_addr_r[1]), .O(n12872));
    defparam rd_addr_r_0__bdd_4_lut_11211.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11405 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_14 ), 
            .I2(\REG.mem_43_14 ), .I3(rd_addr_r[1]), .O(n13106));
    defparam rd_addr_r_0__bdd_4_lut_11405.LUT_INIT = 16'he4aa;
    SB_LUT4 i3930_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_27_9 ), .O(n5132));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3930_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13106_bdd_4_lut (.I0(n13106), .I1(\REG.mem_41_14 ), .I2(\REG.mem_40_14 ), 
            .I3(rd_addr_r[1]), .O(n13109));
    defparam n13106_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12008 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_0 ), 
            .I2(\REG.mem_15_0 ), .I3(rd_addr_r[1]), .O(n13832));
    defparam rd_addr_r_0__bdd_4_lut_12008.LUT_INIT = 16'he4aa;
    SB_LUT4 i3929_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_27_8 ), .O(n5131));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3929_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13832_bdd_4_lut (.I0(n13832), .I1(\REG.mem_13_0 ), .I2(\REG.mem_12_0 ), 
            .I3(rd_addr_r[1]), .O(n13835));
    defparam n13832_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i3818_3819 (.Q(\REG.mem_39_12 ), .C(DEBUG_6_c_c), .D(n5338));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3815_3816 (.Q(\REG.mem_39_11 ), .C(DEBUG_6_c_c), .D(n5337));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3812_3813 (.Q(\REG.mem_39_10 ), .C(DEBUG_6_c_c), .D(n5336));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3809_3810 (.Q(\REG.mem_39_9 ), .C(DEBUG_6_c_c), .D(n5335));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3806_3807 (.Q(\REG.mem_39_8 ), .C(DEBUG_6_c_c), .D(n5334));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3803_3804 (.Q(\REG.mem_39_7 ), .C(DEBUG_6_c_c), .D(n5333));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3800_3801 (.Q(\REG.mem_39_6 ), .C(DEBUG_6_c_c), .D(n5332));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3797_3798 (.Q(\REG.mem_39_5 ), .C(DEBUG_6_c_c), .D(n5331));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3794_3795 (.Q(\REG.mem_39_4 ), .C(DEBUG_6_c_c), .D(n5330));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3791_3792 (.Q(\REG.mem_39_3 ), .C(DEBUG_6_c_c), .D(n5329));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3788_3789 (.Q(\REG.mem_39_2 ), .C(DEBUG_6_c_c), .D(n5328));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3785_3786 (.Q(\REG.mem_39_1 ), .C(DEBUG_6_c_c), .D(n5327));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3782_3783 (.Q(\REG.mem_39_0 ), .C(DEBUG_6_c_c), .D(n5326));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3731_3732 (.Q(\REG.mem_38_15 ), .C(DEBUG_6_c_c), .D(n5323));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12872_bdd_4_lut (.I0(n12872), .I1(\REG.mem_21_5 ), .I2(\REG.mem_20_5 ), 
            .I3(rd_addr_r[1]), .O(n12875));
    defparam n12872_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i3728_3729 (.Q(\REG.mem_38_14 ), .C(DEBUG_6_c_c), .D(n5322));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFSR wr_grey_sync_r__i5 (.Q(wr_grey_sync_r[5]), .C(DEBUG_6_c_c), 
            .D(wr_grey_w[5]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFFSR wr_grey_sync_r__i4 (.Q(wr_grey_sync_r[4]), .C(DEBUG_6_c_c), 
            .D(wr_grey_w[4]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF i3725_3726 (.Q(\REG.mem_38_13 ), .C(DEBUG_6_c_c), .D(n5321));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFSR wr_grey_sync_r__i3 (.Q(wr_grey_sync_r[3]), .C(DEBUG_6_c_c), 
            .D(wr_grey_w[3]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF i3722_3723 (.Q(\REG.mem_38_12 ), .C(DEBUG_6_c_c), .D(n5320));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFSR wr_grey_sync_r__i2 (.Q(wr_grey_sync_r[2]), .C(DEBUG_6_c_c), 
            .D(wr_grey_w[2]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF i3719_3720 (.Q(\REG.mem_38_11 ), .C(DEBUG_6_c_c), .D(n5319));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFSR wr_grey_sync_r__i1 (.Q(wr_grey_sync_r[1]), .C(DEBUG_6_c_c), 
            .D(wr_grey_w[1]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(257[21] 267[24])
    SB_DFF i3716_3717 (.Q(\REG.mem_38_10 ), .C(DEBUG_6_c_c), .D(n5318));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3713_3714 (.Q(\REG.mem_38_9 ), .C(DEBUG_6_c_c), .D(n5317));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3710_3711 (.Q(\REG.mem_38_8 ), .C(DEBUG_6_c_c), .D(n5316));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3707_3708 (.Q(\REG.mem_38_7 ), .C(DEBUG_6_c_c), .D(n5315));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3704_3705 (.Q(\REG.mem_38_6 ), .C(DEBUG_6_c_c), .D(n5314));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3701_3702 (.Q(\REG.mem_38_5 ), .C(DEBUG_6_c_c), .D(n5313));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3698_3699 (.Q(\REG.mem_38_4 ), .C(DEBUG_6_c_c), .D(n5312));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3695_3696 (.Q(\REG.mem_38_3 ), .C(DEBUG_6_c_c), .D(n5311));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3692_3693 (.Q(\REG.mem_38_2 ), .C(DEBUG_6_c_c), .D(n5310));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3689_3690 (.Q(\REG.mem_38_1 ), .C(DEBUG_6_c_c), .D(n5309));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3686_3687 (.Q(\REG.mem_38_0 ), .C(DEBUG_6_c_c), .D(n5308));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3635_3636 (.Q(\REG.mem_37_15 ), .C(DEBUG_6_c_c), .D(n5302));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3632_3633 (.Q(\REG.mem_37_14 ), .C(DEBUG_6_c_c), .D(n5301));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3629_3630 (.Q(\REG.mem_37_13 ), .C(DEBUG_6_c_c), .D(n5300));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3626_3627 (.Q(\REG.mem_37_12 ), .C(DEBUG_6_c_c), .D(n5299));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3623_3624 (.Q(\REG.mem_37_11 ), .C(DEBUG_6_c_c), .D(n5298));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3620_3621 (.Q(\REG.mem_37_10 ), .C(DEBUG_6_c_c), .D(n5297));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3617_3618 (.Q(\REG.mem_37_9 ), .C(DEBUG_6_c_c), .D(n5296));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3614_3615 (.Q(\REG.mem_37_8 ), .C(DEBUG_6_c_c), .D(n5295));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3611_3612 (.Q(\REG.mem_37_7 ), .C(DEBUG_6_c_c), .D(n5294));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3608_3609 (.Q(\REG.mem_37_6 ), .C(DEBUG_6_c_c), .D(n5293));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3605_3606 (.Q(\REG.mem_37_5 ), .C(DEBUG_6_c_c), .D(n5292));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3602_3603 (.Q(\REG.mem_37_4 ), .C(DEBUG_6_c_c), .D(n5291));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3599_3600 (.Q(\REG.mem_37_3 ), .C(DEBUG_6_c_c), .D(n5290));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3596_3597 (.Q(\REG.mem_37_2 ), .C(DEBUG_6_c_c), .D(n5289));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3593_3594 (.Q(\REG.mem_37_1 ), .C(DEBUG_6_c_c), .D(n5288));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3590_3591 (.Q(\REG.mem_37_0 ), .C(DEBUG_6_c_c), .D(n5286));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3539_3540 (.Q(\REG.mem_36_15 ), .C(DEBUG_6_c_c), .D(n5285));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3536_3537 (.Q(\REG.mem_36_14 ), .C(DEBUG_6_c_c), .D(n5284));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3533_3534 (.Q(\REG.mem_36_13 ), .C(DEBUG_6_c_c), .D(n5283));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3530_3531 (.Q(\REG.mem_36_12 ), .C(DEBUG_6_c_c), .D(n5282));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3527_3528 (.Q(\REG.mem_36_11 ), .C(DEBUG_6_c_c), .D(n5281));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3524_3525 (.Q(\REG.mem_36_10 ), .C(DEBUG_6_c_c), .D(n5280));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3521_3522 (.Q(\REG.mem_36_9 ), .C(DEBUG_6_c_c), .D(n5279));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3518_3519 (.Q(\REG.mem_36_8 ), .C(DEBUG_6_c_c), .D(n5278));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3515_3516 (.Q(\REG.mem_36_7 ), .C(DEBUG_6_c_c), .D(n5277));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3512_3513 (.Q(\REG.mem_36_6 ), .C(DEBUG_6_c_c), .D(n5276));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3509_3510 (.Q(\REG.mem_36_5 ), .C(DEBUG_6_c_c), .D(n5275));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3506_3507 (.Q(\REG.mem_36_4 ), .C(DEBUG_6_c_c), .D(n5274));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3503_3504 (.Q(\REG.mem_36_3 ), .C(DEBUG_6_c_c), .D(n5273));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3500_3501 (.Q(\REG.mem_36_2 ), .C(DEBUG_6_c_c), .D(n5272));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3497_3498 (.Q(\REG.mem_36_1 ), .C(DEBUG_6_c_c), .D(n5271));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3494_3495 (.Q(\REG.mem_36_0 ), .C(DEBUG_6_c_c), .D(n5270));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11400 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_12 ), 
            .I2(\REG.mem_27_12 ), .I3(rd_addr_r[1]), .O(n13100));
    defparam rd_addr_r_0__bdd_4_lut_11400.LUT_INIT = 16'he4aa;
    SB_LUT4 i3928_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_27_7 ), .O(n5130));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3928_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13100_bdd_4_lut (.I0(n13100), .I1(\REG.mem_25_12 ), .I2(\REG.mem_24_12 ), 
            .I3(rd_addr_r[1]), .O(n12372));
    defparam n13100_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12003 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_7 ), 
            .I2(\REG.mem_43_7 ), .I3(rd_addr_r[1]), .O(n13826));
    defparam rd_addr_r_0__bdd_4_lut_12003.LUT_INIT = 16'he4aa;
    SB_LUT4 i3927_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_27_6 ), .O(n5129));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3927_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3443_3444 (.Q(\REG.mem_35_15 ), .C(DEBUG_6_c_c), .D(n5269));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13826_bdd_4_lut (.I0(n13826), .I1(\REG.mem_41_7 ), .I2(\REG.mem_40_7 ), 
            .I3(rd_addr_r[1]), .O(n12195));
    defparam n13826_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i3440_3441 (.Q(\REG.mem_35_14 ), .C(DEBUG_6_c_c), .D(n5268));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3437_3438 (.Q(\REG.mem_35_13 ), .C(DEBUG_6_c_c), .D(n5267));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3434_3435 (.Q(\REG.mem_35_12 ), .C(DEBUG_6_c_c), .D(n5266));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3431_3432 (.Q(\REG.mem_35_11 ), .C(DEBUG_6_c_c), .D(n5265));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3428_3429 (.Q(\REG.mem_35_10 ), .C(DEBUG_6_c_c), .D(n5264));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3425_3426 (.Q(\REG.mem_35_9 ), .C(DEBUG_6_c_c), .D(n5263));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3422_3423 (.Q(\REG.mem_35_8 ), .C(DEBUG_6_c_c), .D(n5262));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3419_3420 (.Q(\REG.mem_35_7 ), .C(DEBUG_6_c_c), .D(n5261));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3416_3417 (.Q(\REG.mem_35_6 ), .C(DEBUG_6_c_c), .D(n5260));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3413_3414 (.Q(\REG.mem_35_5 ), .C(DEBUG_6_c_c), .D(n5259));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3410_3411 (.Q(\REG.mem_35_4 ), .C(DEBUG_6_c_c), .D(n5258));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3407_3408 (.Q(\REG.mem_35_3 ), .C(DEBUG_6_c_c), .D(n5257));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3404_3405 (.Q(\REG.mem_35_2 ), .C(DEBUG_6_c_c), .D(n5256));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3401_3402 (.Q(\REG.mem_35_1 ), .C(DEBUG_6_c_c), .D(n5255));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3398_3399 (.Q(\REG.mem_35_0 ), .C(DEBUG_6_c_c), .D(n5254));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3347_3348 (.Q(\REG.mem_34_15 ), .C(DEBUG_6_c_c), .D(n5253));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3926_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_27_5 ), .O(n5128));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3926_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut (.I0(rp_sync2_r[3]), .I1(rp_sync_w[4]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11998 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_7 ), 
            .I2(\REG.mem_47_7 ), .I3(rd_addr_r[1]), .O(n13820));
    defparam rd_addr_r_0__bdd_4_lut_11998.LUT_INIT = 16'he4aa;
    SB_LUT4 rp_sync2_r_6__I_0_136_i1_2_lut (.I0(rp_sync2_r[5]), .I1(rp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(rp_sync_w[5]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam rp_sync2_r_6__I_0_136_i1_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 n13820_bdd_4_lut (.I0(n13820), .I1(\REG.mem_45_7 ), .I2(\REG.mem_44_7 ), 
            .I3(rd_addr_r[1]), .O(n12198));
    defparam n13820_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_45 (.I0(rp_sync2_r[1]), .I1(rp_sync_w[2]), .I2(GND_net), 
            .I3(GND_net), .O(rp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_adj_45.LUT_INIT = 16'h6666;
    SB_LUT4 i3925_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_27_4 ), .O(n5127));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3925_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3344_3345 (.Q(\REG.mem_34_14 ), .C(DEBUG_6_c_c), .D(n5252));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3341_3342 (.Q(\REG.mem_34_13 ), .C(DEBUG_6_c_c), .D(n5251));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3338_3339 (.Q(\REG.mem_34_12 ), .C(DEBUG_6_c_c), .D(n5250));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3335_3336 (.Q(\REG.mem_34_11 ), .C(DEBUG_6_c_c), .D(n5249));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3332_3333 (.Q(\REG.mem_34_10 ), .C(DEBUG_6_c_c), .D(n5248));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3329_3330 (.Q(\REG.mem_34_9 ), .C(DEBUG_6_c_c), .D(n5247));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3326_3327 (.Q(\REG.mem_34_8 ), .C(DEBUG_6_c_c), .D(n5246));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3323_3324 (.Q(\REG.mem_34_7 ), .C(DEBUG_6_c_c), .D(n5245));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3320_3321 (.Q(\REG.mem_34_6 ), .C(DEBUG_6_c_c), .D(n5244));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3317_3318 (.Q(\REG.mem_34_5 ), .C(DEBUG_6_c_c), .D(n5243));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3314_3315 (.Q(\REG.mem_34_4 ), .C(DEBUG_6_c_c), .D(n5242));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3311_3312 (.Q(\REG.mem_34_3 ), .C(DEBUG_6_c_c), .D(n5241));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3308_3309 (.Q(\REG.mem_34_2 ), .C(DEBUG_6_c_c), .D(n5240));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3305_3306 (.Q(\REG.mem_34_1 ), .C(DEBUG_6_c_c), .D(n5239));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3302_3303 (.Q(\REG.mem_34_0 ), .C(DEBUG_6_c_c), .D(n5238));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i2_3_lut_adj_46 (.I0(rp_sync2_r[5]), .I1(rp_sync2_r[4]), .I2(rp_sync2_r[6]), 
            .I3(GND_net), .O(rp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i2_3_lut_adj_46.LUT_INIT = 16'h6969;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11420 (.I0(rd_addr_r[2]), .I1(n12372), 
            .I2(n12881), .I3(rd_addr_r[3]), .O(n13094));
    defparam rd_addr_r_2__bdd_4_lut_11420.LUT_INIT = 16'he4aa;
    SB_LUT4 n13094_bdd_4_lut (.I0(n13094), .I1(n12354), .I2(n12312), .I3(rd_addr_r[3]), 
            .O(n13097));
    defparam n13094_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3924_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_27_3 ), .O(n5126));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3924_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3923_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_27_2 ), .O(n5125));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3923_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3922_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_27_1 ), .O(n5124));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3922_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3251_3252 (.Q(\REG.mem_33_15 ), .C(DEBUG_6_c_c), .D(n5235));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3248_3249 (.Q(\REG.mem_33_14 ), .C(DEBUG_6_c_c), .D(n5234));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3245_3246 (.Q(\REG.mem_33_13 ), .C(DEBUG_6_c_c), .D(n5233));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3242_3243 (.Q(\REG.mem_33_12 ), .C(DEBUG_6_c_c), .D(n5232));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3239_3240 (.Q(\REG.mem_33_11 ), .C(DEBUG_6_c_c), .D(n5231));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3236_3237 (.Q(\REG.mem_33_10 ), .C(DEBUG_6_c_c), .D(n5230));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3233_3234 (.Q(\REG.mem_33_9 ), .C(DEBUG_6_c_c), .D(n5229));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3230_3231 (.Q(\REG.mem_33_8 ), .C(DEBUG_6_c_c), .D(n5228));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3227_3228 (.Q(\REG.mem_33_7 ), .C(DEBUG_6_c_c), .D(n5227));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3224_3225 (.Q(\REG.mem_33_6 ), .C(DEBUG_6_c_c), .D(n5226));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3221_3222 (.Q(\REG.mem_33_5 ), .C(DEBUG_6_c_c), .D(n5225));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3218_3219 (.Q(\REG.mem_33_4 ), .C(DEBUG_6_c_c), .D(n5224));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3215_3216 (.Q(\REG.mem_33_3 ), .C(DEBUG_6_c_c), .D(n5223));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3212_3213 (.Q(\REG.mem_33_2 ), .C(DEBUG_6_c_c), .D(n5222));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3209_3210 (.Q(\REG.mem_33_1 ), .C(DEBUG_6_c_c), .D(n5221));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_p1_w_6__I_0_2_lut (.I0(\wr_addr_p1_w[6] ), .I1(rp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(full_max_w));   // src/fifo_dc_32_lut_gen.v(296[27:88])
    defparam wr_addr_p1_w_6__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9799_4_lut (.I0(wr_addr_p1_w[4]), .I1(wr_addr_p1_w[1]), .I2(rp_sync_w[4]), 
            .I3(rp_sync_w[1]), .O(n11447));
    defparam i9799_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i9736_4_lut (.I0(wr_addr_p1_w[5]), .I1(wr_addr_p1_w[3]), .I2(rp_sync_w[5]), 
            .I3(rp_sync_w[3]), .O(n11384));
    defparam i9736_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 i5_4_lut (.I0(\wr_addr_p1_w[0] ), .I1(n11447), .I2(full_max_w), 
            .I3(rp_sync_w[0]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h1020;
    SB_LUT4 i3921_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_27_0 ), .O(n5123));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3921_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i3206_3207 (.Q(\REG.mem_33_0 ), .C(DEBUG_6_c_c), .D(n5220));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3155_3156 (.Q(\REG.mem_32_15 ), .C(DEBUG_6_c_c), .D(n5219));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3152_3153 (.Q(\REG.mem_32_14 ), .C(DEBUG_6_c_c), .D(n5218));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3149_3150 (.Q(\REG.mem_32_13 ), .C(DEBUG_6_c_c), .D(n5217));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3146_3147 (.Q(\REG.mem_32_12 ), .C(DEBUG_6_c_c), .D(n5216));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3143_3144 (.Q(\REG.mem_32_11 ), .C(DEBUG_6_c_c), .D(n5215));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3140_3141 (.Q(\REG.mem_32_10 ), .C(DEBUG_6_c_c), .D(n5214));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3137_3138 (.Q(\REG.mem_32_9 ), .C(DEBUG_6_c_c), .D(n5213));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3134_3135 (.Q(\REG.mem_32_8 ), .C(DEBUG_6_c_c), .D(n5212));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3131_3132 (.Q(\REG.mem_32_7 ), .C(DEBUG_6_c_c), .D(n5211));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3128_3129 (.Q(\REG.mem_32_6 ), .C(DEBUG_6_c_c), .D(n5210));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3125_3126 (.Q(\REG.mem_32_5 ), .C(DEBUG_6_c_c), .D(n5209));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3122_3123 (.Q(\REG.mem_32_4 ), .C(DEBUG_6_c_c), .D(n5208));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3119_3120 (.Q(\REG.mem_32_3 ), .C(DEBUG_6_c_c), .D(n5207));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3116_3117 (.Q(\REG.mem_32_2 ), .C(DEBUG_6_c_c), .D(n5206));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3113_3114 (.Q(\REG.mem_32_1 ), .C(DEBUG_6_c_c), .D(n5205));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3952_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_28_15 ), .O(n5154));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3952_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9754_4_lut (.I0(wr_addr_r[5]), .I1(wr_addr_r[1]), .I2(rp_sync_w[5]), 
            .I3(rp_sync_w[1]), .O(n11402));
    defparam i9754_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11395 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_3 ), 
            .I2(\REG.mem_11_3 ), .I3(rd_addr_r[1]), .O(n13088));
    defparam rd_addr_r_0__bdd_4_lut_11395.LUT_INIT = 16'he4aa;
    SB_LUT4 i3951_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_28_14 ), .O(n5153));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3951_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9772_4_lut (.I0(wr_addr_r[2]), .I1(\wr_addr_r[0] ), .I2(rp_sync_w[2]), 
            .I3(rp_sync_w[0]), .O(n11420));
    defparam i9772_4_lut.LUT_INIT = 16'hedb7;
    SB_LUT4 wr_addr_r_6__I_0_add_2_7_lut (.I0(n11463), .I1(wr_addr_r[5]), 
            .I2(rp_sync_w[5]), .I3(n10629), .O(n11475)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_7_lut.LUT_INIT = 16'h8228;
    SB_DFF i3110_3111 (.Q(\REG.mem_32_0 ), .C(DEBUG_6_c_c), .D(n5203));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3059_3060 (.Q(\REG.mem_31_15 ), .C(DEBUG_6_c_c), .D(n5202));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3056_3057 (.Q(\REG.mem_31_14 ), .C(DEBUG_6_c_c), .D(n5201));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3053_3054 (.Q(\REG.mem_31_13 ), .C(DEBUG_6_c_c), .D(n5200));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3050_3051 (.Q(\REG.mem_31_12 ), .C(DEBUG_6_c_c), .D(n5199));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3047_3048 (.Q(\REG.mem_31_11 ), .C(DEBUG_6_c_c), .D(n5198));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3044_3045 (.Q(\REG.mem_31_10 ), .C(DEBUG_6_c_c), .D(n5197));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3041_3042 (.Q(\REG.mem_31_9 ), .C(DEBUG_6_c_c), .D(n5196));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3038_3039 (.Q(\REG.mem_31_8 ), .C(DEBUG_6_c_c), .D(n5195));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3035_3036 (.Q(\REG.mem_31_7 ), .C(DEBUG_6_c_c), .D(n5194));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3032_3033 (.Q(\REG.mem_31_6 ), .C(DEBUG_6_c_c), .D(n5193));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3029_3030 (.Q(\REG.mem_31_5 ), .C(DEBUG_6_c_c), .D(n5192));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3026_3027 (.Q(\REG.mem_31_4 ), .C(DEBUG_6_c_c), .D(n5191));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3023_3024 (.Q(\REG.mem_31_3 ), .C(DEBUG_6_c_c), .D(n5190));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3020_3021 (.Q(\REG.mem_31_2 ), .C(DEBUG_6_c_c), .D(n5189));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_6__I_0_add_2_7 (.CI(n10629), .I0(wr_addr_r[5]), .I1(rp_sync_w[5]), 
            .CO(n10630));
    SB_LUT4 i11017_4_lut (.I0(wr_addr_p1_w[2]), .I1(n12), .I2(n11384), 
            .I3(rp_sync_w[2]), .O(n12527));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam i11017_4_lut.LUT_INIT = 16'h0408;
    SB_LUT4 i3950_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_28_13 ), .O(n5152));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3950_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9832_3_lut (.I0(n11400), .I1(n11420), .I2(n11402), .I3(GND_net), 
            .O(n11481));
    defparam i9832_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 full_nxt_c_I_6_4_lut (.I0(n11481), .I1(n12527), .I2(n7596), 
            .I3(full_o), .O(full_nxt_c_N_593));   // src/fifo_dc_32_lut_gen.v(300[45:114])
    defparam full_nxt_c_I_6_4_lut.LUT_INIT = 16'h5c0c;
    SB_LUT4 i3949_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_28_12 ), .O(n5151));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3949_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13088_bdd_4_lut (.I0(n13088), .I1(\REG.mem_9_3 ), .I2(\REG.mem_8_3 ), 
            .I3(rd_addr_r[1]), .O(n11598));
    defparam n13088_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i3017_3018 (.Q(\REG.mem_31_1 ), .C(DEBUG_6_c_c), .D(n5188));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i3014_3015 (.Q(\REG.mem_31_0 ), .C(DEBUG_6_c_c), .D(n5187));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2963_2964 (.Q(\REG.mem_30_15 ), .C(DEBUG_6_c_c), .D(n5186));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2960_2961 (.Q(\REG.mem_30_14 ), .C(DEBUG_6_c_c), .D(n5185));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2957_2958 (.Q(\REG.mem_30_13 ), .C(DEBUG_6_c_c), .D(n5184));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2954_2955 (.Q(\REG.mem_30_12 ), .C(DEBUG_6_c_c), .D(n5183));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2951_2952 (.Q(\REG.mem_30_11 ), .C(DEBUG_6_c_c), .D(n5182));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2948_2949 (.Q(\REG.mem_30_10 ), .C(DEBUG_6_c_c), .D(n5181));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2945_2946 (.Q(\REG.mem_30_9 ), .C(DEBUG_6_c_c), .D(n5180));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2942_2943 (.Q(\REG.mem_30_8 ), .C(DEBUG_6_c_c), .D(n5179));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2939_2940 (.Q(\REG.mem_30_7 ), .C(DEBUG_6_c_c), .D(n5178));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2936_2937 (.Q(\REG.mem_30_6 ), .C(DEBUG_6_c_c), .D(n5177));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2933_2934 (.Q(\REG.mem_30_5 ), .C(DEBUG_6_c_c), .D(n5176));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2930_2931 (.Q(\REG.mem_30_4 ), .C(DEBUG_6_c_c), .D(n5175));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2927_2928 (.Q(\REG.mem_30_3 ), .C(DEBUG_6_c_c), .D(n5174));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3948_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_28_11 ), .O(n5150));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3948_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3947_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_28_10 ), .O(n5149));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3947_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3946_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_28_9 ), .O(n5148));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3946_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10358_3_lut (.I0(\REG.mem_56_0 ), .I1(\REG.mem_57_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12007));
    defparam i10358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3945_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_28_8 ), .O(n5147));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3945_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3944_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_28_7 ), .O(n5146));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3944_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11993 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_14 ), 
            .I2(\REG.mem_11_14 ), .I3(rd_addr_r[1]), .O(n13814));
    defparam rd_addr_r_0__bdd_4_lut_11993.LUT_INIT = 16'he4aa;
    SB_LUT4 i3943_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_28_6 ), .O(n5145));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3943_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10359_3_lut (.I0(\REG.mem_58_0 ), .I1(\REG.mem_59_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12008));
    defparam i10359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3942_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_28_5 ), .O(n5144));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3942_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3941_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_28_4 ), .O(n5143));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3941_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10368_3_lut (.I0(\REG.mem_62_0 ), .I1(\REG.mem_63_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12017));
    defparam i10368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11390 (.I0(rd_addr_r[2]), .I1(n11862), 
            .I2(n11874), .I3(rd_addr_r[3]), .O(n13082));
    defparam rd_addr_r_2__bdd_4_lut_11390.LUT_INIT = 16'he4aa;
    SB_DFF i2924_2925 (.Q(\REG.mem_30_2 ), .C(DEBUG_6_c_c), .D(n5173));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3940_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_28_3 ), .O(n5142));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3940_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13082_bdd_4_lut (.I0(n13082), .I1(n11853), .I2(n11841), .I3(rd_addr_r[3]), 
            .O(n11913));
    defparam n13082_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2921_2922 (.Q(\REG.mem_30_1 ), .C(DEBUG_6_c_c), .D(n5172));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13814_bdd_4_lut (.I0(n13814), .I1(\REG.mem_9_14 ), .I2(\REG.mem_8_14 ), 
            .I3(rd_addr_r[1]), .O(n13817));
    defparam n13814_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2918_2919 (.Q(\REG.mem_30_0 ), .C(DEBUG_6_c_c), .D(n5171));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2867_2868 (.Q(\REG.mem_29_15 ), .C(DEBUG_6_c_c), .D(n5170));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2864_2865 (.Q(\REG.mem_29_14 ), .C(DEBUG_6_c_c), .D(n5169));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2861_2862 (.Q(\REG.mem_29_13 ), .C(DEBUG_6_c_c), .D(n5168));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2858_2859 (.Q(\REG.mem_29_12 ), .C(DEBUG_6_c_c), .D(n5167));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2855_2856 (.Q(\REG.mem_29_11 ), .C(DEBUG_6_c_c), .D(n5166));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2852_2853 (.Q(\REG.mem_29_10 ), .C(DEBUG_6_c_c), .D(n5165));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2849_2850 (.Q(\REG.mem_29_9 ), .C(DEBUG_6_c_c), .D(n5164));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2846_2847 (.Q(\REG.mem_29_8 ), .C(DEBUG_6_c_c), .D(n5163));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2843_2844 (.Q(\REG.mem_29_7 ), .C(DEBUG_6_c_c), .D(n5162));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2840_2841 (.Q(\REG.mem_29_6 ), .C(DEBUG_6_c_c), .D(n5161));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2837_2838 (.Q(\REG.mem_29_5 ), .C(DEBUG_6_c_c), .D(n5160));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2834_2835 (.Q(\REG.mem_29_4 ), .C(DEBUG_6_c_c), .D(n5159));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2831_2832 (.Q(\REG.mem_29_3 ), .C(DEBUG_6_c_c), .D(n5158));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2828_2829 (.Q(\REG.mem_29_2 ), .C(DEBUG_6_c_c), .D(n5157));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10367_3_lut (.I0(\REG.mem_60_0 ), .I1(\REG.mem_61_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12016));
    defparam i10367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11380 (.I0(rd_addr_r[2]), .I1(n12075), 
            .I2(n12102), .I3(rd_addr_r[3]), .O(n13076));
    defparam rd_addr_r_2__bdd_4_lut_11380.LUT_INIT = 16'he4aa;
    SB_LUT4 n13076_bdd_4_lut (.I0(n13076), .I1(n12051), .I2(n12042), .I3(rd_addr_r[3]), 
            .O(n12375));
    defparam n13076_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11988 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_8 ), 
            .I2(\REG.mem_39_8 ), .I3(rd_addr_r[1]), .O(n13808));
    defparam rd_addr_r_0__bdd_4_lut_11988.LUT_INIT = 16'he4aa;
    SB_LUT4 i3939_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_28_2 ), .O(n5141));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3939_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13808_bdd_4_lut (.I0(n13808), .I1(\REG.mem_37_8 ), .I2(\REG.mem_36_8 ), 
            .I3(rd_addr_r[1]), .O(n11784));
    defparam n13808_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11385 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_8 ), 
            .I2(\REG.mem_3_8 ), .I3(rd_addr_r[1]), .O(n13070));
    defparam rd_addr_r_0__bdd_4_lut_11385.LUT_INIT = 16'he4aa;
    SB_LUT4 i3938_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_28_1 ), .O(n5140));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3938_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3937_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_28_0 ), .O(n5139));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3937_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i2825_2826 (.Q(\REG.mem_29_1 ), .C(DEBUG_6_c_c), .D(n5156));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3968_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_29_15 ), .O(n5170));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3968_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i2822_2823 (.Q(\REG.mem_29_0 ), .C(DEBUG_6_c_c), .D(n5155));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2771_2772 (.Q(\REG.mem_28_15 ), .C(DEBUG_6_c_c), .D(n5154));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2768_2769 (.Q(\REG.mem_28_14 ), .C(DEBUG_6_c_c), .D(n5153));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2765_2766 (.Q(\REG.mem_28_13 ), .C(DEBUG_6_c_c), .D(n5152));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2762_2763 (.Q(\REG.mem_28_12 ), .C(DEBUG_6_c_c), .D(n5151));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2759_2760 (.Q(\REG.mem_28_11 ), .C(DEBUG_6_c_c), .D(n5150));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2756_2757 (.Q(\REG.mem_28_10 ), .C(DEBUG_6_c_c), .D(n5149));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2753_2754 (.Q(\REG.mem_28_9 ), .C(DEBUG_6_c_c), .D(n5148));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2750_2751 (.Q(\REG.mem_28_8 ), .C(DEBUG_6_c_c), .D(n5147));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2747_2748 (.Q(\REG.mem_28_7 ), .C(DEBUG_6_c_c), .D(n5146));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2744_2745 (.Q(\REG.mem_28_6 ), .C(DEBUG_6_c_c), .D(n5145));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2741_2742 (.Q(\REG.mem_28_5 ), .C(DEBUG_6_c_c), .D(n5144));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2738_2739 (.Q(\REG.mem_28_4 ), .C(DEBUG_6_c_c), .D(n5143));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2735_2736 (.Q(\REG.mem_28_3 ), .C(DEBUG_6_c_c), .D(n5142));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2732_2733 (.Q(\REG.mem_28_2 ), .C(DEBUG_6_c_c), .D(n5141));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2729_2730 (.Q(\REG.mem_28_1 ), .C(DEBUG_6_c_c), .D(n5140));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11983 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_13 ), 
            .I2(\REG.mem_43_13 ), .I3(rd_addr_r[1]), .O(n13802));
    defparam rd_addr_r_0__bdd_4_lut_11983.LUT_INIT = 16'he4aa;
    SB_LUT4 n13802_bdd_4_lut (.I0(n13802), .I1(\REG.mem_41_13 ), .I2(\REG.mem_40_13 ), 
            .I3(rd_addr_r[1]), .O(n12204));
    defparam n13802_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13070_bdd_4_lut (.I0(n13070), .I1(\REG.mem_1_8 ), .I2(\REG.mem_0_8 ), 
            .I3(rd_addr_r[1]), .O(n13073));
    defparam n13070_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12053 (.I0(rd_addr_r[1]), .I1(n11755), 
            .I2(n11756), .I3(rd_addr_r[2]), .O(n13796));
    defparam rd_addr_r_1__bdd_4_lut_12053.LUT_INIT = 16'he4aa;
    SB_LUT4 i3967_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_29_14 ), .O(n5169));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3967_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i2726_2727 (.Q(\REG.mem_28_0 ), .C(DEBUG_6_c_c), .D(n5139));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11370 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_2 ), 
            .I2(\REG.mem_23_2 ), .I3(rd_addr_r[1]), .O(n13064));
    defparam rd_addr_r_0__bdd_4_lut_11370.LUT_INIT = 16'he4aa;
    SB_LUT4 n13796_bdd_4_lut (.I0(n13796), .I1(n11663), .I2(n11662), .I3(rd_addr_r[2]), 
            .O(n13799));
    defparam n13796_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i5_2_lut_4_lut (.I0(wr_addr_r[5]), .I1(wr_addr_p1_w[5]), 
            .I2(n7596), .I3(\wr_addr_nxt_c[4] ), .O(wr_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i5_2_lut_4_lut.LUT_INIT = 16'h53ac;
    SB_DFF i2675_2676 (.Q(\REG.mem_27_15 ), .C(DEBUG_6_c_c), .D(n5138));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2672_2673 (.Q(\REG.mem_27_14 ), .C(DEBUG_6_c_c), .D(n5137));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2669_2670 (.Q(\REG.mem_27_13 ), .C(DEBUG_6_c_c), .D(n5136));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2666_2667 (.Q(\REG.mem_27_12 ), .C(DEBUG_6_c_c), .D(n5135));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2663_2664 (.Q(\REG.mem_27_11 ), .C(DEBUG_6_c_c), .D(n5134));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2660_2661 (.Q(\REG.mem_27_10 ), .C(DEBUG_6_c_c), .D(n5133));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2657_2658 (.Q(\REG.mem_27_9 ), .C(DEBUG_6_c_c), .D(n5132));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2654_2655 (.Q(\REG.mem_27_8 ), .C(DEBUG_6_c_c), .D(n5131));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2651_2652 (.Q(\REG.mem_27_7 ), .C(DEBUG_6_c_c), .D(n5130));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2648_2649 (.Q(\REG.mem_27_6 ), .C(DEBUG_6_c_c), .D(n5129));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2645_2646 (.Q(\REG.mem_27_5 ), .C(DEBUG_6_c_c), .D(n5128));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2642_2643 (.Q(\REG.mem_27_4 ), .C(DEBUG_6_c_c), .D(n5127));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2639_2640 (.Q(\REG.mem_27_3 ), .C(DEBUG_6_c_c), .D(n5126));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2636_2637 (.Q(\REG.mem_27_2 ), .C(DEBUG_6_c_c), .D(n5125));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2633_2634 (.Q(\REG.mem_27_1 ), .C(DEBUG_6_c_c), .D(n5124));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2630_2631 (.Q(\REG.mem_27_0 ), .C(DEBUG_6_c_c), .D(n5123));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3966_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_29_13 ), .O(n5168));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3966_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i2579_2580 (.Q(\REG.mem_26_15 ), .C(DEBUG_6_c_c), .D(n5121));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3965_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_29_12 ), .O(n5167));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3965_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13064_bdd_4_lut (.I0(n13064), .I1(\REG.mem_21_2 ), .I2(\REG.mem_20_2 ), 
            .I3(rd_addr_r[1]), .O(n13067));
    defparam n13064_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3964_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_29_11 ), .O(n5166));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3964_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i2576_2577 (.Q(\REG.mem_26_14 ), .C(DEBUG_6_c_c), .D(n5120));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3963_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_29_10 ), .O(n5165));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3963_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i2573_2574 (.Q(\REG.mem_26_13 ), .C(DEBUG_6_c_c), .D(n5119));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2570_2571 (.Q(\REG.mem_26_12 ), .C(DEBUG_6_c_c), .D(n5118));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2567_2568 (.Q(\REG.mem_26_11 ), .C(DEBUG_6_c_c), .D(n5117));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2564_2565 (.Q(\REG.mem_26_10 ), .C(DEBUG_6_c_c), .D(n5116));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2561_2562 (.Q(\REG.mem_26_9 ), .C(DEBUG_6_c_c), .D(n5115));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2558_2559 (.Q(\REG.mem_26_8 ), .C(DEBUG_6_c_c), .D(n5114));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2555_2556 (.Q(\REG.mem_26_7 ), .C(DEBUG_6_c_c), .D(n5113));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2552_2553 (.Q(\REG.mem_26_6 ), .C(DEBUG_6_c_c), .D(n5112));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2549_2550 (.Q(\REG.mem_26_5 ), .C(DEBUG_6_c_c), .D(n5111));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2546_2547 (.Q(\REG.mem_26_4 ), .C(DEBUG_6_c_c), .D(n5110));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2543_2544 (.Q(\REG.mem_26_3 ), .C(DEBUG_6_c_c), .D(n5109));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2540_2541 (.Q(\REG.mem_26_2 ), .C(DEBUG_6_c_c), .D(n5108));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2537_2538 (.Q(\REG.mem_26_1 ), .C(DEBUG_6_c_c), .D(n5107));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2534_2535 (.Q(\REG.mem_26_0 ), .C(DEBUG_6_c_c), .D(n5106));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2483_2484 (.Q(\REG.mem_25_15 ), .C(DEBUG_6_c_c), .D(n5105));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2480_2481 (.Q(\REG.mem_25_14 ), .C(DEBUG_6_c_c), .D(n5104));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11973 (.I0(rd_addr_r[1]), .I1(n12520), 
            .I2(n12521), .I3(rd_addr_r[2]), .O(n13784));
    defparam rd_addr_r_1__bdd_4_lut_11973.LUT_INIT = 16'he4aa;
    SB_LUT4 i10513_3_lut (.I0(n13787), .I1(n13937), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n12162));
    defparam i10513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_11550 (.I0(rd_addr_r[4]), .I1(n11901), 
            .I2(n11913), .I3(rd_addr_r[5]), .O(n13058));
    defparam rd_addr_r_4__bdd_4_lut_11550.LUT_INIT = 16'he4aa;
    SB_LUT4 n13058_bdd_4_lut (.I0(n13058), .I1(n11898), .I2(n11880), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_526 [8]));
    defparam n13058_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13784_bdd_4_lut (.I0(n13784), .I1(n12515), .I2(n12514), .I3(rd_addr_r[2]), 
            .O(n13787));
    defparam n13784_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3962_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_29_9 ), .O(n5164));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3962_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10533_3_lut (.I0(n13871), .I1(n13739), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12182));
    defparam i10533_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2477_2478 (.Q(\REG.mem_25_13 ), .C(DEBUG_6_c_c), .D(n5103));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3961_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_29_8 ), .O(n5163));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3961_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10534_3_lut (.I0(n13799), .I1(n12182), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n12183));
    defparam i10534_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i2474_2475 (.Q(\REG.mem_25_12 ), .C(DEBUG_6_c_c), .D(n5102));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11365 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_3 ), 
            .I2(\REG.mem_59_3 ), .I3(rd_addr_r[1]), .O(n13052));
    defparam rd_addr_r_0__bdd_4_lut_11365.LUT_INIT = 16'he4aa;
    SB_DFF i2471_2472 (.Q(\REG.mem_25_11 ), .C(DEBUG_6_c_c), .D(n5101));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2468_2469 (.Q(\REG.mem_25_10 ), .C(DEBUG_6_c_c), .D(n5100));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2465_2466 (.Q(\REG.mem_25_9 ), .C(DEBUG_6_c_c), .D(n5099));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2462_2463 (.Q(\REG.mem_25_8 ), .C(DEBUG_6_c_c), .D(n5098));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2459_2460 (.Q(\REG.mem_25_7 ), .C(DEBUG_6_c_c), .D(n5097));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2456_2457 (.Q(\REG.mem_25_6 ), .C(DEBUG_6_c_c), .D(n5096));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2453_2454 (.Q(\REG.mem_25_5 ), .C(DEBUG_6_c_c), .D(n5095));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2450_2451 (.Q(\REG.mem_25_4 ), .C(DEBUG_6_c_c), .D(n5094));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2447_2448 (.Q(\REG.mem_25_3 ), .C(DEBUG_6_c_c), .D(n5093));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2444_2445 (.Q(\REG.mem_25_2 ), .C(DEBUG_6_c_c), .D(n5092));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2441_2442 (.Q(\REG.mem_25_1 ), .C(DEBUG_6_c_c), .D(n5091));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2438_2439 (.Q(\REG.mem_25_0 ), .C(DEBUG_6_c_c), .D(n5090));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2387_2388 (.Q(\REG.mem_24_15 ), .C(DEBUG_6_c_c), .D(n5089));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2384_2385 (.Q(\REG.mem_24_14 ), .C(DEBUG_6_c_c), .D(n5088));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13052_bdd_4_lut (.I0(n13052), .I1(\REG.mem_57_3 ), .I2(\REG.mem_56_3 ), 
            .I3(rd_addr_r[1]), .O(n13055));
    defparam n13052_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3960_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_29_7 ), .O(n5162));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3960_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i2381_2382 (.Q(\REG.mem_24_13 ), .C(DEBUG_6_c_c), .D(n5087));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3959_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_29_6 ), .O(n5161));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3959_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3958_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_29_5 ), .O(n5160));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3958_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3957_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_29_4 ), .O(n5159));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3957_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i2378_2379 (.Q(\REG.mem_24_12 ), .C(DEBUG_6_c_c), .D(n5086));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3956_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_29_3 ), .O(n5158));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3956_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3955_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_29_2 ), .O(n5157));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3955_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3954_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_29_1 ), .O(n5156));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3954_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i2375_2376 (.Q(\REG.mem_24_11 ), .C(DEBUG_6_c_c), .D(n5085));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2372_2373 (.Q(\REG.mem_24_10 ), .C(DEBUG_6_c_c), .D(n5084));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2369_2370 (.Q(\REG.mem_24_9 ), .C(DEBUG_6_c_c), .D(n5083));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2366_2367 (.Q(\REG.mem_24_8 ), .C(DEBUG_6_c_c), .D(n5082));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2363_2364 (.Q(\REG.mem_24_7 ), .C(DEBUG_6_c_c), .D(n5081));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2360_2361 (.Q(\REG.mem_24_6 ), .C(DEBUG_6_c_c), .D(n5080));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2357_2358 (.Q(\REG.mem_24_5 ), .C(DEBUG_6_c_c), .D(n5079));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2354_2355 (.Q(\REG.mem_24_4 ), .C(DEBUG_6_c_c), .D(n5078));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2351_2352 (.Q(\REG.mem_24_3 ), .C(DEBUG_6_c_c), .D(n5077));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2348_2349 (.Q(\REG.mem_24_2 ), .C(DEBUG_6_c_c), .D(n5076));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2345_2346 (.Q(\REG.mem_24_1 ), .C(DEBUG_6_c_c), .D(n5075));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2342_2343 (.Q(\REG.mem_24_0 ), .C(DEBUG_6_c_c), .D(n5074));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2291_2292 (.Q(\REG.mem_23_15 ), .C(DEBUG_6_c_c), .D(n5073));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2288_2289 (.Q(\REG.mem_23_14 ), .C(DEBUG_6_c_c), .D(n5072));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2285_2286 (.Q(\REG.mem_23_13 ), .C(DEBUG_6_c_c), .D(n5071));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2282_2283 (.Q(\REG.mem_23_12 ), .C(DEBUG_6_c_c), .D(n5070));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2279_2280 (.Q(\REG.mem_23_11 ), .C(DEBUG_6_c_c), .D(n5069));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2276_2277 (.Q(\REG.mem_23_10 ), .C(DEBUG_6_c_c), .D(n5068));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2273_2274 (.Q(\REG.mem_23_9 ), .C(DEBUG_6_c_c), .D(n5067));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12806_bdd_4_lut (.I0(n12806), .I1(n11559), .I2(n11523), .I3(rd_addr_r[3]), 
            .O(n12809));
    defparam n12806_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2270_2271 (.Q(\REG.mem_23_8 ), .C(DEBUG_6_c_c), .D(n5066));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFFSR rd_grey_sync_r__i5 (.Q(\rd_grey_sync_r[5] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[5]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_DFFSR rd_grey_sync_r__i4 (.Q(\rd_grey_sync_r[4] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[4]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 i3953_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_29_0 ), .O(n5155));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3953_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11978 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_6 ), 
            .I2(\REG.mem_11_6 ), .I3(rd_addr_r[1]), .O(n13778));
    defparam rd_addr_r_0__bdd_4_lut_11978.LUT_INIT = 16'he4aa;
    SB_DFFSR rd_grey_sync_r__i3 (.Q(\rd_grey_sync_r[3] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[3]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 i4570_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_62_15 ), .O(n5772));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4570_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFSR rd_grey_sync_r__i2 (.Q(\rd_grey_sync_r[2] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[2]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11355 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_14 ), 
            .I2(\REG.mem_47_14 ), .I3(rd_addr_r[1]), .O(n13046));
    defparam rd_addr_r_0__bdd_4_lut_11355.LUT_INIT = 16'he4aa;
    SB_DFFSR rd_grey_sync_r__i1 (.Q(\rd_grey_sync_r[1] ), .C(SLM_CLK_c), 
            .D(rd_grey_w[1]), .R(reset_all));   // src/fifo_dc_32_lut_gen.v(508[21] 518[24])
    SB_LUT4 EnabledDecoder_2_i42_2_lut (.I0(n26_adj_1146), .I1(wr_addr_r[4]), 
            .I2(GND_net), .I3(GND_net), .O(n42_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i42_2_lut.LUT_INIT = 16'h2222;
    SB_DFF i2267_2268 (.Q(\REG.mem_23_7 ), .C(DEBUG_6_c_c), .D(n5065));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4569_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_62_14 ), .O(n5771));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4569_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i2264_2265 (.Q(\REG.mem_23_6 ), .C(DEBUG_6_c_c), .D(n5064));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2261_2262 (.Q(\REG.mem_23_5 ), .C(DEBUG_6_c_c), .D(n5063));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2258_2259 (.Q(\REG.mem_23_4 ), .C(DEBUG_6_c_c), .D(n5062));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2255_2256 (.Q(\REG.mem_23_3 ), .C(DEBUG_6_c_c), .D(n5061));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2252_2253 (.Q(\REG.mem_23_2 ), .C(DEBUG_6_c_c), .D(n5060));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2249_2250 (.Q(\REG.mem_23_1 ), .C(DEBUG_6_c_c), .D(n5059));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2246_2247 (.Q(\REG.mem_23_0 ), .C(DEBUG_6_c_c), .D(n5058));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2195_2196 (.Q(\REG.mem_22_15 ), .C(DEBUG_6_c_c), .D(n5057));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2192_2193 (.Q(\REG.mem_22_14 ), .C(DEBUG_6_c_c), .D(n5056));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2189_2190 (.Q(\REG.mem_22_13 ), .C(DEBUG_6_c_c), .D(n5055));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2186_2187 (.Q(\REG.mem_22_12 ), .C(DEBUG_6_c_c), .D(n5054));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2183_2184 (.Q(\REG.mem_22_11 ), .C(DEBUG_6_c_c), .D(n5053));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2180_2181 (.Q(\REG.mem_22_10 ), .C(DEBUG_6_c_c), .D(n5052));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2177_2178 (.Q(\REG.mem_22_9 ), .C(DEBUG_6_c_c), .D(n5051));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2174_2175 (.Q(\REG.mem_22_8 ), .C(DEBUG_6_c_c), .D(n5050));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13778_bdd_4_lut (.I0(n13778), .I1(\REG.mem_9_6 ), .I2(\REG.mem_8_6 ), 
            .I3(rd_addr_r[1]), .O(n13781));
    defparam n13778_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13046_bdd_4_lut (.I0(n13046), .I1(\REG.mem_45_14 ), .I2(\REG.mem_44_14 ), 
            .I3(rd_addr_r[1]), .O(n13049));
    defparam n13046_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11350 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_15 ), 
            .I2(\REG.mem_3_15 ), .I3(rd_addr_r[1]), .O(n13040));
    defparam rd_addr_r_0__bdd_4_lut_11350.LUT_INIT = 16'he4aa;
    SB_LUT4 i4568_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_62_13 ), .O(n5770));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4568_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13040_bdd_4_lut (.I0(n13040), .I1(\REG.mem_1_15 ), .I2(\REG.mem_0_15 ), 
            .I3(rd_addr_r[1]), .O(n13043));
    defparam n13040_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4567_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_62_12 ), .O(n5769));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4567_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4566_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_62_11 ), .O(n5768));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4566_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_2_lut (.I0(n7_c), .I1(n8), .I2(GND_net), .I3(GND_net), 
            .O(n5));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11959 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_6 ), 
            .I2(\REG.mem_15_6 ), .I3(rd_addr_r[1]), .O(n13772));
    defparam rd_addr_r_0__bdd_4_lut_11959.LUT_INIT = 16'he4aa;
    SB_DFF i2171_2172 (.Q(\REG.mem_22_7 ), .C(DEBUG_6_c_c), .D(n5049));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13772_bdd_4_lut (.I0(n13772), .I1(\REG.mem_13_6 ), .I2(\REG.mem_12_6 ), 
            .I3(rd_addr_r[1]), .O(n13775));
    defparam n13772_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i2168_2169 (.Q(\REG.mem_22_6 ), .C(DEBUG_6_c_c), .D(n5048));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2165_2166 (.Q(\REG.mem_22_5 ), .C(DEBUG_6_c_c), .D(n5047));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2162_2163 (.Q(\REG.mem_22_4 ), .C(DEBUG_6_c_c), .D(n5046));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2159_2160 (.Q(\REG.mem_22_3 ), .C(DEBUG_6_c_c), .D(n5045));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2156_2157 (.Q(\REG.mem_22_2 ), .C(DEBUG_6_c_c), .D(n5044));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2153_2154 (.Q(\REG.mem_22_1 ), .C(DEBUG_6_c_c), .D(n5043));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2150_2151 (.Q(\REG.mem_22_0 ), .C(DEBUG_6_c_c), .D(n5042));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2099_2100 (.Q(\REG.mem_21_15 ), .C(DEBUG_6_c_c), .D(n5041));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2096_2097 (.Q(\REG.mem_21_14 ), .C(DEBUG_6_c_c), .D(n5040));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2093_2094 (.Q(\REG.mem_21_13 ), .C(DEBUG_6_c_c), .D(n5039));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2090_2091 (.Q(\REG.mem_21_12 ), .C(DEBUG_6_c_c), .D(n5038));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2087_2088 (.Q(\REG.mem_21_11 ), .C(DEBUG_6_c_c), .D(n5037));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2084_2085 (.Q(\REG.mem_21_10 ), .C(DEBUG_6_c_c), .D(n5036));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2081_2082 (.Q(\REG.mem_21_9 ), .C(DEBUG_6_c_c), .D(n5035));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2078_2079 (.Q(\REG.mem_21_8 ), .C(DEBUG_6_c_c), .D(n5034));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2075_2076 (.Q(\REG.mem_21_7 ), .C(DEBUG_6_c_c), .D(n5033));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2072_2073 (.Q(\REG.mem_21_6 ), .C(DEBUG_6_c_c), .D(n5032));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11375 (.I0(rd_addr_r[2]), .I1(n12138), 
            .I2(n12153), .I3(rd_addr_r[3]), .O(n13034));
    defparam rd_addr_r_2__bdd_4_lut_11375.LUT_INIT = 16'he4aa;
    SB_DFF i2069_2070 (.Q(\REG.mem_21_5 ), .C(DEBUG_6_c_c), .D(n5031));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2066_2067 (.Q(\REG.mem_21_4 ), .C(DEBUG_6_c_c), .D(n5030));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2063_2064 (.Q(\REG.mem_21_3 ), .C(DEBUG_6_c_c), .D(n5029));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2060_2061 (.Q(\REG.mem_21_2 ), .C(DEBUG_6_c_c), .D(n5028));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2057_2058 (.Q(\REG.mem_21_1 ), .C(DEBUG_6_c_c), .D(n5027));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2054_2055 (.Q(\REG.mem_21_0 ), .C(DEBUG_6_c_c), .D(n5026));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2003_2004 (.Q(\REG.mem_20_15 ), .C(DEBUG_6_c_c), .D(n5025));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i2000_2001 (.Q(\REG.mem_20_14 ), .C(DEBUG_6_c_c), .D(n5024));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1997_1998 (.Q(\REG.mem_20_13 ), .C(DEBUG_6_c_c), .D(n5023));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1994_1995 (.Q(\REG.mem_20_12 ), .C(DEBUG_6_c_c), .D(n5022));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1991_1992 (.Q(\REG.mem_20_11 ), .C(DEBUG_6_c_c), .D(n5021));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1988_1989 (.Q(\REG.mem_20_10 ), .C(DEBUG_6_c_c), .D(n5020));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1985_1986 (.Q(\REG.mem_20_9 ), .C(DEBUG_6_c_c), .D(n5019));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1982_1983 (.Q(\REG.mem_20_8 ), .C(DEBUG_6_c_c), .D(n5018));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1979_1980 (.Q(\REG.mem_20_7 ), .C(DEBUG_6_c_c), .D(n5017));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1976_1977 (.Q(\REG.mem_20_6 ), .C(DEBUG_6_c_c), .D(n5016));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1973_1974 (.Q(\REG.mem_20_5 ), .C(DEBUG_6_c_c), .D(n5015));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1970_1971 (.Q(\REG.mem_20_4 ), .C(DEBUG_6_c_c), .D(n5014));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1967_1968 (.Q(\REG.mem_20_3 ), .C(DEBUG_6_c_c), .D(n5013));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1964_1965 (.Q(\REG.mem_20_2 ), .C(DEBUG_6_c_c), .D(n5012));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1961_1962 (.Q(\REG.mem_20_1 ), .C(DEBUG_6_c_c), .D(n5011));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1958_1959 (.Q(\REG.mem_20_0 ), .C(DEBUG_6_c_c), .D(n5010));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13034_bdd_4_lut (.I0(n13034), .I1(n12123), .I2(n12108), .I3(rd_addr_r[3]), 
            .O(n12387));
    defparam n13034_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4565_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_62_10 ), .O(n5767));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4565_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1907_1908 (.Q(\REG.mem_19_15 ), .C(DEBUG_6_c_c), .D(n5006));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 wr_addr_r_6__I_0_135_i1_3_lut (.I0(\wr_addr_r[0] ), .I1(\wr_addr_p1_w[0] ), 
            .I2(n7596), .I3(GND_net), .O(wr_addr_nxt_c[0]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_r_6__I_0_135_i1_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4564_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_62_9 ), .O(n5766));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4564_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11345 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_9 ), 
            .I2(\REG.mem_27_9 ), .I3(rd_addr_r[1]), .O(n13028));
    defparam rd_addr_r_0__bdd_4_lut_11345.LUT_INIT = 16'he4aa;
    SB_LUT4 n13028_bdd_4_lut (.I0(n13028), .I1(\REG.mem_25_9 ), .I2(\REG.mem_24_9 ), 
            .I3(rd_addr_r[1]), .O(n13031));
    defparam n13028_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11335 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_10 ), 
            .I2(\REG.mem_51_10 ), .I3(rd_addr_r[1]), .O(n13022));
    defparam rd_addr_r_0__bdd_4_lut_11335.LUT_INIT = 16'he4aa;
    SB_LUT4 i10129_3_lut (.I0(n13379), .I1(n13847), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_526 [1]));
    defparam i10129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11954 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_7 ), 
            .I2(\REG.mem_51_7 ), .I3(rd_addr_r[1]), .O(n13760));
    defparam rd_addr_r_0__bdd_4_lut_11954.LUT_INIT = 16'he4aa;
    SB_LUT4 i9849_3_lut (.I0(n12947), .I1(n14411), .I2(rd_addr_r[4]), 
            .I3(GND_net), .O(n11498));
    defparam i9849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9850_3_lut (.I0(n13013), .I1(n11498), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_526 [2]));
    defparam i9850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4563_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_62_8 ), .O(n5765));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4563_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13022_bdd_4_lut (.I0(n13022), .I1(\REG.mem_49_10 ), .I2(\REG.mem_48_10 ), 
            .I3(rd_addr_r[1]), .O(n13025));
    defparam n13022_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9970_3_lut (.I0(n13253), .I1(n14261), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_526 [5]));
    defparam i9970_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1904_1905 (.Q(\REG.mem_19_14 ), .C(DEBUG_6_c_c), .D(n5005));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1901_1902 (.Q(\REG.mem_19_13 ), .C(DEBUG_6_c_c), .D(n5004));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1898_1899 (.Q(\REG.mem_19_12 ), .C(DEBUG_6_c_c), .D(n5003));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1895_1896 (.Q(\REG.mem_19_11 ), .C(DEBUG_6_c_c), .D(n5002));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1892_1893 (.Q(\REG.mem_19_10 ), .C(DEBUG_6_c_c), .D(n5001));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1889_1890 (.Q(\REG.mem_19_9 ), .C(DEBUG_6_c_c), .D(n5000));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1886_1887 (.Q(\REG.mem_19_8 ), .C(DEBUG_6_c_c), .D(n4999));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1883_1884 (.Q(\REG.mem_19_7 ), .C(DEBUG_6_c_c), .D(n4998));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1880_1881 (.Q(\REG.mem_19_6 ), .C(DEBUG_6_c_c), .D(n4997));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1877_1878 (.Q(\REG.mem_19_5 ), .C(DEBUG_6_c_c), .D(n4996));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1874_1875 (.Q(\REG.mem_19_4 ), .C(DEBUG_6_c_c), .D(n4995));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1871_1872 (.Q(\REG.mem_19_3 ), .C(DEBUG_6_c_c), .D(n4994));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1868_1869 (.Q(\REG.mem_19_2 ), .C(DEBUG_6_c_c), .D(n4993));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4562_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_62_7 ), .O(n5764));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4562_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11330 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_0 ), 
            .I2(\REG.mem_39_0 ), .I3(rd_addr_r[1]), .O(n13016));
    defparam rd_addr_r_0__bdd_4_lut_11330.LUT_INIT = 16'he4aa;
    SB_LUT4 n13760_bdd_4_lut (.I0(n13760), .I1(\REG.mem_49_7 ), .I2(\REG.mem_48_7 ), 
            .I3(rd_addr_r[1]), .O(n12210));
    defparam n13760_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4561_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_62_6 ), .O(n5763));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4561_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9871_3_lut (.I0(n13175), .I1(n14303), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_526 [9]));
    defparam i9871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4560_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_62_5 ), .O(n5762));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4560_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4559_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_62_4 ), .O(n5761));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4559_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4558_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_62_3 ), .O(n5760));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4558_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11944 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_11 ), 
            .I2(\REG.mem_35_11 ), .I3(rd_addr_r[1]), .O(n13754));
    defparam rd_addr_r_0__bdd_4_lut_11944.LUT_INIT = 16'he4aa;
    SB_DFF i1865_1866 (.Q(\REG.mem_19_1 ), .C(DEBUG_6_c_c), .D(n4992));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1862_1863 (.Q(\REG.mem_19_0 ), .C(DEBUG_6_c_c), .D(n4991));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1811_1812 (.Q(\REG.mem_18_15 ), .C(DEBUG_6_c_c), .D(n4990));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1808_1809 (.Q(\REG.mem_18_14 ), .C(DEBUG_6_c_c), .D(n4989));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1805_1806 (.Q(\REG.mem_18_13 ), .C(DEBUG_6_c_c), .D(n4988));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1802_1803 (.Q(\REG.mem_18_12 ), .C(DEBUG_6_c_c), .D(n4987));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1799_1800 (.Q(\REG.mem_18_11 ), .C(DEBUG_6_c_c), .D(n4986));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1796_1797 (.Q(\REG.mem_18_10 ), .C(DEBUG_6_c_c), .D(n4985));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1793_1794 (.Q(\REG.mem_18_9 ), .C(DEBUG_6_c_c), .D(n4984));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1790_1791 (.Q(\REG.mem_18_8 ), .C(DEBUG_6_c_c), .D(n4983));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1787_1788 (.Q(\REG.mem_18_7 ), .C(DEBUG_6_c_c), .D(n4982));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1784_1785 (.Q(\REG.mem_18_6 ), .C(DEBUG_6_c_c), .D(n4981));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1781_1782 (.Q(\REG.mem_18_5 ), .C(DEBUG_6_c_c), .D(n4980));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1778_1779 (.Q(\REG.mem_18_4 ), .C(DEBUG_6_c_c), .D(n4979));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1775_1776 (.Q(\REG.mem_18_3 ), .C(DEBUG_6_c_c), .D(n4978));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1772_1773 (.Q(\REG.mem_18_2 ), .C(DEBUG_6_c_c), .D(n4977));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1769_1770 (.Q(\REG.mem_18_1 ), .C(DEBUG_6_c_c), .D(n4976));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10003_3_lut (.I0(n13301), .I1(n14231), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_526 [10]));
    defparam i10003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13016_bdd_4_lut (.I0(n13016), .I1(\REG.mem_37_0 ), .I2(\REG.mem_36_0 ), 
            .I3(rd_addr_r[1]), .O(n13019));
    defparam n13016_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4557_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_62_2 ), .O(n5759));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4557_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1766_1767 (.Q(\REG.mem_18_0 ), .C(DEBUG_6_c_c), .D(n4975));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13754_bdd_4_lut (.I0(n13754), .I1(\REG.mem_33_11 ), .I2(\REG.mem_32_11 ), 
            .I3(rd_addr_r[1]), .O(n13757));
    defparam n13754_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1715_1716 (.Q(\REG.mem_17_15 ), .C(DEBUG_6_c_c), .D(n4974));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i9934_3_lut (.I0(n13229), .I1(n13631), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_526 [14]));
    defparam i9934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10456_3_lut (.I0(n13691), .I1(n14117), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_526 [15]));
    defparam i10456_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1712_1713 (.Q(\REG.mem_17_14 ), .C(DEBUG_6_c_c), .D(n4973));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11455 (.I0(rd_addr_r[3]), .I1(n12376), 
            .I2(n12377), .I3(rd_addr_r[4]), .O(n13010));
    defparam rd_addr_r_3__bdd_4_lut_11455.LUT_INIT = 16'he4aa;
    SB_LUT4 n13010_bdd_4_lut (.I0(n13010), .I1(n12347), .I2(n12346), .I3(rd_addr_r[4]), 
            .O(n13013));
    defparam n13010_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1709_1710 (.Q(\REG.mem_17_13 ), .C(DEBUG_6_c_c), .D(n4972));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11340 (.I0(rd_addr_r[2]), .I1(n12474), 
            .I2(n11634), .I3(rd_addr_r[3]), .O(n13004));
    defparam rd_addr_r_2__bdd_4_lut_11340.LUT_INIT = 16'he4aa;
    SB_LUT4 n13004_bdd_4_lut (.I0(n13004), .I1(n12459), .I2(n12785), .I3(rd_addr_r[3]), 
            .O(n13007));
    defparam n13004_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11325 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_3 ), 
            .I2(\REG.mem_63_3 ), .I3(rd_addr_r[1]), .O(n12998));
    defparam rd_addr_r_0__bdd_4_lut_11325.LUT_INIT = 16'he4aa;
    SB_DFF i1706_1707 (.Q(\REG.mem_17_12 ), .C(DEBUG_6_c_c), .D(n4971));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1703_1704 (.Q(\REG.mem_17_11 ), .C(DEBUG_6_c_c), .D(n4970));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1700_1701 (.Q(\REG.mem_17_10 ), .C(DEBUG_6_c_c), .D(n4969));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1697_1698 (.Q(\REG.mem_17_9 ), .C(DEBUG_6_c_c), .D(n4968));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1694_1695 (.Q(\REG.mem_17_8 ), .C(DEBUG_6_c_c), .D(n4967));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1691_1692 (.Q(\REG.mem_17_7 ), .C(DEBUG_6_c_c), .D(n4966));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1688_1689 (.Q(\REG.mem_17_6 ), .C(DEBUG_6_c_c), .D(n4965));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1685_1686 (.Q(\REG.mem_17_5 ), .C(DEBUG_6_c_c), .D(n4964));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1682_1683 (.Q(\REG.mem_17_4 ), .C(DEBUG_6_c_c), .D(n4963));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1679_1680 (.Q(\REG.mem_17_3 ), .C(DEBUG_6_c_c), .D(n4962));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1676_1677 (.Q(\REG.mem_17_2 ), .C(DEBUG_6_c_c), .D(n4961));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1673_1674 (.Q(\REG.mem_17_1 ), .C(DEBUG_6_c_c), .D(n4960));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1670_1671 (.Q(\REG.mem_17_0 ), .C(DEBUG_6_c_c), .D(n4958));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1619_1620 (.Q(\REG.mem_16_15 ), .C(DEBUG_6_c_c), .D(n4957));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1616_1617 (.Q(\REG.mem_16_14 ), .C(DEBUG_6_c_c), .D(n4956));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4556_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_62_1 ), .O(n5758));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4556_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10385_3_lut (.I0(\REG.mem_56_15 ), .I1(\REG.mem_57_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12034));
    defparam i10385_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1613_1614 (.Q(\REG.mem_16_13 ), .C(DEBUG_6_c_c), .D(n4955));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12998_bdd_4_lut (.I0(n12998), .I1(\REG.mem_61_3 ), .I2(\REG.mem_60_3 ), 
            .I3(rd_addr_r[1]), .O(n13001));
    defparam n12998_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4555_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_62_0 ), .O(n5757));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4555_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1610_1611 (.Q(\REG.mem_16_12 ), .C(DEBUG_6_c_c), .D(n4954));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i16_2_lut (.I0(n12_adj_1156), .I1(wr_addr_r[2]), 
            .I2(GND_net), .I3(GND_net), .O(n16_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i16_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11939 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_11 ), 
            .I2(\REG.mem_59_11 ), .I3(rd_addr_r[1]), .O(n13748));
    defparam rd_addr_r_0__bdd_4_lut_11939.LUT_INIT = 16'he4aa;
    SB_LUT4 n13748_bdd_4_lut (.I0(n13748), .I1(\REG.mem_57_11 ), .I2(\REG.mem_56_11 ), 
            .I3(rd_addr_r[1]), .O(n13751));
    defparam n13748_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1607_1608 (.Q(\REG.mem_16_11 ), .C(DEBUG_6_c_c), .D(n4953));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11311 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_4 ), 
            .I2(\REG.mem_47_4 ), .I3(rd_addr_r[1]), .O(n12992));
    defparam rd_addr_r_0__bdd_4_lut_11311.LUT_INIT = 16'he4aa;
    SB_LUT4 i10386_3_lut (.I0(\REG.mem_58_15 ), .I1(\REG.mem_59_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12035));
    defparam i10386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12992_bdd_4_lut (.I0(n12992), .I1(\REG.mem_45_4 ), .I2(\REG.mem_44_4 ), 
            .I3(rd_addr_r[1]), .O(n12995));
    defparam n12992_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11934 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_5 ), 
            .I2(\REG.mem_43_5 ), .I3(rd_addr_r[1]), .O(n13742));
    defparam rd_addr_r_0__bdd_4_lut_11934.LUT_INIT = 16'he4aa;
    SB_DFF i1604_1605 (.Q(\REG.mem_16_10 ), .C(DEBUG_6_c_c), .D(n4952));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13742_bdd_4_lut (.I0(n13742), .I1(\REG.mem_41_5 ), .I2(\REG.mem_40_5 ), 
            .I3(rd_addr_r[1]), .O(n13745));
    defparam n13742_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11306 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_5 ), 
            .I2(\REG.mem_63_5 ), .I3(rd_addr_r[1]), .O(n12986));
    defparam rd_addr_r_0__bdd_4_lut_11306.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11929 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_4 ), 
            .I2(\REG.mem_31_4 ), .I3(rd_addr_r[1]), .O(n13736));
    defparam rd_addr_r_0__bdd_4_lut_11929.LUT_INIT = 16'he4aa;
    SB_LUT4 n13736_bdd_4_lut (.I0(n13736), .I1(\REG.mem_29_4 ), .I2(\REG.mem_28_4 ), 
            .I3(rd_addr_r[1]), .O(n13739));
    defparam n13736_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12986_bdd_4_lut (.I0(n12986), .I1(\REG.mem_61_5 ), .I2(\REG.mem_60_5 ), 
            .I3(rd_addr_r[1]), .O(n12989));
    defparam n12986_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i98_2_lut_3_lut_4_lut (.I0(n17_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n51));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i98_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_adj_47 (.I0(wp_sync2_r[6]), .I1(wp_sync2_r[5]), .I2(GND_net), 
            .I3(GND_net), .O(n4027));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_47.LUT_INIT = 16'h6666;
    SB_DFF i1601_1602 (.Q(\REG.mem_16_9 ), .C(DEBUG_6_c_c), .D(n4951));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1598_1599 (.Q(\REG.mem_16_8 ), .C(DEBUG_6_c_c), .D(n4950));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1595_1596 (.Q(\REG.mem_16_7 ), .C(DEBUG_6_c_c), .D(n4949));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1592_1593 (.Q(\REG.mem_16_6 ), .C(DEBUG_6_c_c), .D(n4948));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1589_1590 (.Q(\REG.mem_16_5 ), .C(DEBUG_6_c_c), .D(n4947));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1586_1587 (.Q(\REG.mem_16_4 ), .C(DEBUG_6_c_c), .D(n4946));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i1_2_lut_adj_48 (.I0(wp_sync2_r[0]), .I1(wp_sync_w[1]), .I2(GND_net), 
            .I3(GND_net), .O(wp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_48.LUT_INIT = 16'h6666;
    SB_LUT4 i9797_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_r[4]), .I2(wp_sync_w[0]), 
            .I3(wp_sync_w[4]), .O(n11445));
    defparam i9797_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i9760_4_lut (.I0(rd_addr_r[5]), .I1(rd_addr_r[3]), .I2(n4027), 
            .I3(wp_sync_w[3]), .O(n11408));
    defparam i9760_4_lut.LUT_INIT = 16'h7bde;
    SB_DFF i1583_1584 (.Q(\REG.mem_16_3 ), .C(DEBUG_6_c_c), .D(n4945));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1580_1581 (.Q(\REG.mem_16_2 ), .C(DEBUG_6_c_c), .D(n4944));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1577_1578 (.Q(\REG.mem_16_1 ), .C(DEBUG_6_c_c), .D(n4943));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1574_1575 (.Q(\REG.mem_16_0 ), .C(DEBUG_6_c_c), .D(n4942));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1523_1524 (.Q(\REG.mem_15_15 ), .C(DEBUG_6_c_c), .D(n4941));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1520_1521 (.Q(\REG.mem_15_14 ), .C(DEBUG_6_c_c), .D(n4940));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1517_1518 (.Q(\REG.mem_15_13 ), .C(DEBUG_6_c_c), .D(n4939));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1514_1515 (.Q(\REG.mem_15_12 ), .C(DEBUG_6_c_c), .D(n4938));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1511_1512 (.Q(\REG.mem_15_11 ), .C(DEBUG_6_c_c), .D(n4937));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_6__I_0_i6_3_lut (.I0(rd_addr_r[5]), .I1(rd_addr_p1_w[5]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_465[5] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i97_2_lut_3_lut_4_lut (.I0(n17_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n19));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i97_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i9782_4_lut (.I0(rd_addr_r[1]), .I1(rd_addr_r[2]), .I2(wp_sync_w[1]), 
            .I3(wp_sync_w[2]), .O(n11430));
    defparam i9782_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11301 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_9 ), 
            .I2(\REG.mem_31_9 ), .I3(rd_addr_r[1]), .O(n12980));
    defparam rd_addr_r_0__bdd_4_lut_11301.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11206 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_14 ), 
            .I2(\REG.mem_55_14 ), .I3(rd_addr_r[1]), .O(n12866));
    defparam rd_addr_r_0__bdd_4_lut_11206.LUT_INIT = 16'he4aa;
    SB_LUT4 n12866_bdd_4_lut (.I0(n12866), .I1(\REG.mem_53_14 ), .I2(\REG.mem_52_14 ), 
            .I3(rd_addr_r[1]), .O(n12869));
    defparam n12866_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11924 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_2 ), 
            .I2(\REG.mem_59_2 ), .I3(rd_addr_r[1]), .O(n13730));
    defparam rd_addr_r_0__bdd_4_lut_11924.LUT_INIT = 16'he4aa;
    SB_DFF i1508_1509 (.Q(\REG.mem_15_10 ), .C(DEBUG_6_c_c), .D(n4936));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11236 (.I0(rd_addr_r[1]), .I1(n12343), 
            .I2(n12344), .I3(rd_addr_r[2]), .O(n12860));
    defparam rd_addr_r_1__bdd_4_lut_11236.LUT_INIT = 16'he4aa;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i6_2_lut_4_lut (.I0(wr_addr_r[5]), .I1(wr_addr_p1_w[5]), 
            .I2(n7596), .I3(wr_grey_w[6]), .O(wr_grey_w[5]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i6_2_lut_4_lut.LUT_INIT = 16'h53ac;
    SB_LUT4 n12860_bdd_4_lut (.I0(n12860), .I1(n12341), .I2(n12340), .I3(rd_addr_r[2]), 
            .O(n12863));
    defparam n12860_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4547_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_61_15 ), .O(n5749));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4547_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13730_bdd_4_lut (.I0(n13730), .I1(\REG.mem_57_2 ), .I2(\REG.mem_56_2 ), 
            .I3(rd_addr_r[1]), .O(n13733));
    defparam n13730_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12980_bdd_4_lut (.I0(n12980), .I1(\REG.mem_29_9 ), .I2(\REG.mem_28_9 ), 
            .I3(rd_addr_r[1]), .O(n12983));
    defparam n12980_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_49 (.I0(rd_addr_p1_w[4]), .I1(wp_sync_w[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4025));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_adj_49.LUT_INIT = 16'h6666;
    SB_LUT4 i4546_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_61_14 ), .O(n5748));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4546_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4545_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_61_13 ), .O(n5747));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4545_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4544_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_61_12 ), .O(n5746));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4544_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut (.I0(rd_addr_p1_w[5]), .I1(rd_addr_p1_w[3]), .I2(n4027), 
            .I3(wp_sync_w[3]), .O(n10_c));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_DFF i1505_1506 (.Q(\REG.mem_15_9 ), .C(DEBUG_6_c_c), .D(n4935));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i1_4_lut (.I0(wp_sync2_r[6]), .I1(rd_addr_p1_w[1]), .I2(rd_addr_p1_w[6]), 
            .I3(wp_sync_w[1]), .O(n8_adj_1157));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i1_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i4543_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_61_11 ), .O(n5745));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4543_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_4_lut_adj_50 (.I0(rd_addr_p1_w[0]), .I1(n10_c), .I2(n4025), 
            .I3(wp_sync_w[0]), .O(n12_adj_1158));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i5_4_lut_adj_50.LUT_INIT = 16'hfdfe;
    SB_LUT4 i9834_3_lut (.I0(n11430), .I1(n11408), .I2(n11445), .I3(GND_net), 
            .O(n11483));
    defparam i9834_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut (.I0(rd_addr_p1_w[2]), .I1(n12_adj_1158), .I2(n8_adj_1157), 
            .I3(wp_sync_w[2]), .O(n10760));   // src/fifo_dc_32_lut_gen.v(544[28:56])
    defparam i6_4_lut.LUT_INIT = 16'hfdfe;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11296 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_14 ), 
            .I2(\REG.mem_51_14 ), .I3(rd_addr_r[1]), .O(n12974));
    defparam rd_addr_r_0__bdd_4_lut_11296.LUT_INIT = 16'he4aa;
    SB_LUT4 i10968_4_lut (.I0(n10760), .I1(n11483), .I2(DEBUG_5_c), .I3(get_next_word), 
            .O(empty_nxt_c_N_596));   // src/fifo_dc_32_lut_gen.v(555[46:103])
    defparam i10968_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 n12974_bdd_4_lut (.I0(n12974), .I1(\REG.mem_49_14 ), .I2(\REG.mem_48_14 ), 
            .I3(rd_addr_r[1]), .O(n12977));
    defparam n12974_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_6__I_0_i4_3_lut (.I0(rd_addr_r[3]), .I1(rd_addr_p1_w[3]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_465[3] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11316 (.I0(rd_addr_r[2]), .I1(n12204), 
            .I2(n12225), .I3(rd_addr_r[3]), .O(n12968));
    defparam rd_addr_r_2__bdd_4_lut_11316.LUT_INIT = 16'he4aa;
    SB_DFF i1502_1503 (.Q(\REG.mem_15_8 ), .C(DEBUG_6_c_c), .D(n4934));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1499_1500 (.Q(\REG.mem_15_7 ), .C(DEBUG_6_c_c), .D(n4933));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1496_1497 (.Q(\REG.mem_15_6 ), .C(DEBUG_6_c_c), .D(n4932));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1493_1494 (.Q(\REG.mem_15_5 ), .C(DEBUG_6_c_c), .D(n4931));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1490_1491 (.Q(\REG.mem_15_4 ), .C(DEBUG_6_c_c), .D(n4930));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1487_1488 (.Q(\REG.mem_15_3 ), .C(DEBUG_6_c_c), .D(n4929));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1484_1485 (.Q(\REG.mem_15_2 ), .C(DEBUG_6_c_c), .D(n4928));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1481_1482 (.Q(\REG.mem_15_1 ), .C(DEBUG_6_c_c), .D(n4927));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11919 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_8 ), 
            .I2(\REG.mem_43_8 ), .I3(rd_addr_r[1]), .O(n13724));
    defparam rd_addr_r_0__bdd_4_lut_11919.LUT_INIT = 16'he4aa;
    SB_LUT4 i10395_3_lut (.I0(\REG.mem_62_15 ), .I1(\REG.mem_63_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12044));
    defparam i10395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12968_bdd_4_lut (.I0(n12968), .I1(n12189), .I2(n12174), .I3(rd_addr_r[3]), 
            .O(n12405));
    defparam n12968_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4542_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_61_10 ), .O(n5744));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4542_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i140_141 (.Q(\REG.mem_1_2 ), .C(DEBUG_6_c_c), .D(n4648));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13724_bdd_4_lut (.I0(n13724), .I1(\REG.mem_41_8 ), .I2(\REG.mem_40_8 ), 
            .I3(rd_addr_r[1]), .O(n11811));
    defparam n13724_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11914 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_7 ), 
            .I2(\REG.mem_55_7 ), .I3(rd_addr_r[1]), .O(n13718));
    defparam rd_addr_r_0__bdd_4_lut_11914.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11291 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_10 ), 
            .I2(\REG.mem_55_10 ), .I3(rd_addr_r[1]), .O(n12962));
    defparam rd_addr_r_0__bdd_4_lut_11291.LUT_INIT = 16'he4aa;
    SB_LUT4 i4541_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_61_9 ), .O(n5743));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4541_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4540_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_61_8 ), .O(n5742));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4540_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4539_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_61_7 ), .O(n5741));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4539_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10394_3_lut (.I0(\REG.mem_60_15 ), .I1(\REG.mem_61_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12043));
    defparam i10394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10349_3_lut (.I0(\REG.mem_40_15 ), .I1(\REG.mem_41_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11998));
    defparam i10349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n12962_bdd_4_lut (.I0(n12962), .I1(\REG.mem_53_10 ), .I2(\REG.mem_52_10 ), 
            .I3(rd_addr_r[1]), .O(n12965));
    defparam n12962_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4538_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_61_6 ), .O(n5740));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4538_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1478_1479 (.Q(\REG.mem_15_0 ), .C(DEBUG_6_c_c), .D(n4926));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11281 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_9 ), 
            .I2(\REG.mem_35_9 ), .I3(rd_addr_r[1]), .O(n12956));
    defparam rd_addr_r_0__bdd_4_lut_11281.LUT_INIT = 16'he4aa;
    SB_LUT4 n13718_bdd_4_lut (.I0(n13718), .I1(\REG.mem_53_7 ), .I2(\REG.mem_52_7 ), 
            .I3(rd_addr_r[1]), .O(n12222));
    defparam n13718_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12956_bdd_4_lut (.I0(n12956), .I1(\REG.mem_33_9 ), .I2(\REG.mem_32_9 ), 
            .I3(rd_addr_r[1]), .O(n12959));
    defparam n12956_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10350_3_lut (.I0(\REG.mem_42_15 ), .I1(\REG.mem_43_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11999));
    defparam i10350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4537_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_61_5 ), .O(n5739));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4537_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11909 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_13 ), 
            .I2(\REG.mem_47_13 ), .I3(rd_addr_r[1]), .O(n13712));
    defparam rd_addr_r_0__bdd_4_lut_11909.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11276 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_11 ), 
            .I2(\REG.mem_3_11 ), .I3(rd_addr_r[1]), .O(n12950));
    defparam rd_addr_r_0__bdd_4_lut_11276.LUT_INIT = 16'he4aa;
    SB_LUT4 n12950_bdd_4_lut (.I0(n12950), .I1(\REG.mem_1_11 ), .I2(\REG.mem_0_11 ), 
            .I3(rd_addr_r[1]), .O(n12953));
    defparam n12950_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4536_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_61_4 ), .O(n5738));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4536_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13712_bdd_4_lut (.I0(n13712), .I1(\REG.mem_45_13 ), .I2(\REG.mem_44_13 ), 
            .I3(rd_addr_r[1]), .O(n12225));
    defparam n13712_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1427_1428 (.Q(\REG.mem_14_15 ), .C(DEBUG_6_c_c), .D(n4925));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4535_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_61_3 ), .O(n5737));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4535_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1424_1425 (.Q(\REG.mem_14_14 ), .C(DEBUG_6_c_c), .D(n4924));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1421_1422 (.Q(\REG.mem_14_13 ), .C(DEBUG_6_c_c), .D(n4923));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1418_1419 (.Q(\REG.mem_14_12 ), .C(DEBUG_6_c_c), .D(n4922));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1415_1416 (.Q(\REG.mem_14_11 ), .C(DEBUG_6_c_c), .D(n4921));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1412_1413 (.Q(\REG.mem_14_10 ), .C(DEBUG_6_c_c), .D(n4920));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1409_1410 (.Q(\REG.mem_14_9 ), .C(DEBUG_6_c_c), .D(n4919));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1406_1407 (.Q(\REG.mem_14_8 ), .C(DEBUG_6_c_c), .D(n4918));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4534_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_61_2 ), .O(n5736));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4534_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11286 (.I0(rd_addr_r[2]), .I1(n12078), 
            .I2(n12114), .I3(rd_addr_r[3]), .O(n12944));
    defparam rd_addr_r_2__bdd_4_lut_11286.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12013 (.I0(rd_addr_r[3]), .I1(n12067), 
            .I2(n12068), .I3(rd_addr_r[4]), .O(n13706));
    defparam rd_addr_r_3__bdd_4_lut_12013.LUT_INIT = 16'he4aa;
    SB_LUT4 n12944_bdd_4_lut (.I0(n12944), .I1(n12057), .I2(n12030), .I3(rd_addr_r[3]), 
            .O(n12947));
    defparam n12944_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3972_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_30_3 ), .O(n5174));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3972_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13706_bdd_4_lut (.I0(n13706), .I1(n12038), .I2(n13565), .I3(rd_addr_r[4]), 
            .O(n13709));
    defparam n13706_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11271 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_0 ), 
            .I2(\REG.mem_43_0 ), .I3(rd_addr_r[1]), .O(n12938));
    defparam rd_addr_r_0__bdd_4_lut_11271.LUT_INIT = 16'he4aa;
    SB_LUT4 n12938_bdd_4_lut (.I0(n12938), .I1(\REG.mem_41_0 ), .I2(\REG.mem_40_0 ), 
            .I3(rd_addr_r[1]), .O(n12941));
    defparam n12938_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_6__I_0_i2_3_lut (.I0(rd_addr_r[1]), .I1(rd_addr_p1_w[1]), 
            .I2(rd_fifo_en_w), .I3(GND_net), .O(\rd_addr_nxt_c_6__N_465[1] ));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_r_6__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i1_1_lut (.I0(rd_addr_r[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1173[0]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11261 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_9 ), 
            .I2(\REG.mem_39_9 ), .I3(rd_addr_r[1]), .O(n12932));
    defparam rd_addr_r_0__bdd_4_lut_11261.LUT_INIT = 16'he4aa;
    SB_LUT4 i4271_2_lut_4_lut (.I0(wr_addr_r[5]), .I1(wr_addr_p1_w[5]), 
            .I2(n7596), .I3(reset_all), .O(n5473));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i4271_2_lut_4_lut.LUT_INIT = 16'h00ac;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11904 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_7 ), 
            .I2(\REG.mem_59_7 ), .I3(rd_addr_r[1]), .O(n13700));
    defparam rd_addr_r_0__bdd_4_lut_11904.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_51 (.I0(\state_timeout_counter[3] ), .I1(DEBUG_9_c), 
            .I2(n718), .I3(n7), .O(n14424));
    defparam i3_4_lut_adj_51.LUT_INIT = 16'h0040;
    SB_LUT4 i4533_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_61_1 ), .O(n5735));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4533_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13700_bdd_4_lut (.I0(n13700), .I1(\REG.mem_57_7 ), .I2(\REG.mem_56_7 ), 
            .I3(rd_addr_r[1]), .O(n12228));
    defparam n13700_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12932_bdd_4_lut (.I0(n12932), .I1(\REG.mem_37_9 ), .I2(\REG.mem_36_9 ), 
            .I3(rd_addr_r[1]), .O(n12935));
    defparam n12932_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4532_3_lut_4_lut (.I0(n63), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_61_0 ), .O(n5734));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4532_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1403_1404 (.Q(\REG.mem_14_7 ), .C(DEBUG_6_c_c), .D(n4917));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1400_1401 (.Q(\REG.mem_14_6 ), .C(DEBUG_6_c_c), .D(n4916));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1397_1398 (.Q(\REG.mem_14_5 ), .C(DEBUG_6_c_c), .D(n4915));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1394_1395 (.Q(\REG.mem_14_4 ), .C(DEBUG_6_c_c), .D(n4914));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1391_1392 (.Q(\REG.mem_14_3 ), .C(DEBUG_6_c_c), .D(n4913));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1388_1389 (.Q(\REG.mem_14_2 ), .C(DEBUG_6_c_c), .D(n4912));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1385_1386 (.Q(\REG.mem_14_1 ), .C(DEBUG_6_c_c), .D(n4911));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1382_1383 (.Q(\REG.mem_14_0 ), .C(DEBUG_6_c_c), .D(n4910));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11256 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_15 ), 
            .I2(\REG.mem_7_15 ), .I3(rd_addr_r[1]), .O(n12926));
    defparam rd_addr_r_0__bdd_4_lut_11256.LUT_INIT = 16'he4aa;
    SB_LUT4 n12926_bdd_4_lut (.I0(n12926), .I1(\REG.mem_5_15 ), .I2(\REG.mem_4_15 ), 
            .I3(rd_addr_r[1]), .O(n12929));
    defparam n12926_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11251 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_15 ), 
            .I2(\REG.mem_11_15 ), .I3(rd_addr_r[1]), .O(n12920));
    defparam rd_addr_r_0__bdd_4_lut_11251.LUT_INIT = 16'he4aa;
    SB_LUT4 n12920_bdd_4_lut (.I0(n12920), .I1(\REG.mem_9_15 ), .I2(\REG.mem_8_15 ), 
            .I3(rd_addr_r[1]), .O(n12923));
    defparam n12920_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11899 (.I0(rd_addr_r[3]), .I1(n12070), 
            .I2(n12071), .I3(rd_addr_r[4]), .O(n13688));
    defparam rd_addr_r_3__bdd_4_lut_11899.LUT_INIT = 16'he4aa;
    SB_LUT4 n13688_bdd_4_lut (.I0(n13688), .I1(n12059), .I2(n12058), .I3(rd_addr_r[4]), 
            .O(n13691));
    defparam n13688_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i100_2_lut_3_lut (.I0(n35), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n50));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i100_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11246 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_10 ), 
            .I2(\REG.mem_59_10 ), .I3(rd_addr_r[1]), .O(n12914));
    defparam rd_addr_r_0__bdd_4_lut_11246.LUT_INIT = 16'he4aa;
    SB_LUT4 n12914_bdd_4_lut (.I0(n12914), .I1(\REG.mem_57_10 ), .I2(\REG.mem_56_10 ), 
            .I3(rd_addr_r[1]), .O(n12917));
    defparam n12914_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11445 (.I0(rd_addr_r[1]), .I1(n12382), 
            .I2(n12383), .I3(rd_addr_r[2]), .O(n12908));
    defparam rd_addr_r_1__bdd_4_lut_11445.LUT_INIT = 16'he4aa;
    SB_LUT4 n12908_bdd_4_lut (.I0(n12908), .I1(n12362), .I2(n12361), .I3(rd_addr_r[2]), 
            .O(n12911));
    defparam n12908_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i96_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n52));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i96_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i95_2_lut_3_lut_4_lut (.I0(n15_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n20));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i95_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i3527_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_3_4 ), .O(n4729));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3527_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i99_2_lut_3_lut (.I0(n35), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n18));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i99_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i3526_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_3_3 ), .O(n4728));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3526_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11201 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_9 ), 
            .I2(\REG.mem_43_9 ), .I3(rd_addr_r[1]), .O(n12854));
    defparam rd_addr_r_0__bdd_4_lut_11201.LUT_INIT = 16'he4aa;
    SB_DFF i1331_1332 (.Q(\REG.mem_13_15 ), .C(DEBUG_6_c_c), .D(n4909));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3525_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_3_2 ), .O(n4727));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3525_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11964 (.I0(rd_addr_r[1]), .I1(n11983), 
            .I2(n11984), .I3(rd_addr_r[2]), .O(n13682));
    defparam rd_addr_r_1__bdd_4_lut_11964.LUT_INIT = 16'he4aa;
    SB_LUT4 i3524_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_3_1 ), .O(n4726));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3524_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3523_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_3_0 ), .O(n4725));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3523_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13682_bdd_4_lut (.I0(n13682), .I1(n11972), .I2(n11971), .I3(rd_addr_r[2]), 
            .O(n13685));
    defparam n13682_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1328_1329 (.Q(\REG.mem_13_14 ), .C(DEBUG_6_c_c), .D(n4908));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3539_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_3_15 ), .O(n4741));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3539_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3537_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_3_14 ), .O(n4739));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3537_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3536_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_3_13 ), .O(n4738));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3536_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3535_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_3_12 ), .O(n4737));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3535_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3534_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_3_11 ), .O(n4736));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3534_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3533_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_3_10 ), .O(n4735));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3533_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1325_1326 (.Q(\REG.mem_13_13 ), .C(DEBUG_6_c_c), .D(n4907));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1322_1323 (.Q(\REG.mem_13_12 ), .C(DEBUG_6_c_c), .D(n4906));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3532_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_3_9 ), .O(n4734));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3532_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1319_1320 (.Q(\REG.mem_13_11 ), .C(DEBUG_6_c_c), .D(n4905));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3531_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_3_8 ), .O(n4733));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3531_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1316_1317 (.Q(\REG.mem_13_10 ), .C(DEBUG_6_c_c), .D(n4904));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1313_1314 (.Q(\REG.mem_13_9 ), .C(DEBUG_6_c_c), .D(n4903));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3530_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_3_7 ), .O(n4732));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3530_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3529_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_3_6 ), .O(n4731));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3529_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3528_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_3_5 ), .O(n4730));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3528_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3984_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_30_15 ), .O(n5186));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3984_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1310_1311 (.Q(\REG.mem_13_8 ), .C(DEBUG_6_c_c), .D(n4902));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1307_1308 (.Q(\REG.mem_13_7 ), .C(DEBUG_6_c_c), .D(n4901));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11879 (.I0(rd_addr_r[1]), .I1(n12031), 
            .I2(n12032), .I3(rd_addr_r[2]), .O(n13676));
    defparam rd_addr_r_1__bdd_4_lut_11879.LUT_INIT = 16'he4aa;
    SB_LUT4 n13676_bdd_4_lut (.I0(n13676), .I1(n12020), .I2(n12019), .I3(rd_addr_r[2]), 
            .O(n13679));
    defparam n13676_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_2__bdd_4_lut (.I0(rd_addr_r[2]), .I1(n13733), .I2(n13607), 
            .I3(rd_addr_r[3]), .O(n14408));
    defparam rd_addr_r_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i108_2_lut_3_lut_4_lut (.I0(n20_adj_1160), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n46));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i108_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 n14408_bdd_4_lut (.I0(n14408), .I1(n13913), .I2(n13979), .I3(rd_addr_r[3]), 
            .O(n14411));
    defparam n14408_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1304_1305 (.Q(\REG.mem_13_6 ), .C(DEBUG_6_c_c), .D(n4900));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11874 (.I0(rd_addr_r[1]), .I1(n11995), 
            .I2(n11996), .I3(rd_addr_r[2]), .O(n13670));
    defparam rd_addr_r_1__bdd_4_lut_11874.LUT_INIT = 16'he4aa;
    SB_LUT4 i3983_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_30_14 ), .O(n5185));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3983_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1301_1302 (.Q(\REG.mem_13_5 ), .C(DEBUG_6_c_c), .D(n4899));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i107_2_lut_3_lut_4_lut (.I0(n20_adj_1160), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n14));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i107_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 n13670_bdd_4_lut (.I0(n13670), .I1(n11987), .I2(n11986), .I3(rd_addr_r[2]), 
            .O(n13673));
    defparam n13670_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n12776_bdd_4_lut (.I0(n12776), .I1(\REG.mem_25_15 ), .I2(\REG.mem_24_15 ), 
            .I3(rd_addr_r[1]), .O(n12779));
    defparam n12776_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\REG.mem_10_11 ), 
            .I2(\REG.mem_11_11 ), .I3(rd_addr_r[1]), .O(n14402));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF i1298_1299 (.Q(\REG.mem_13_4 ), .C(DEBUG_6_c_c), .D(n4898));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10365_3_lut (.I0(\REG.mem_46_15 ), .I1(\REG.mem_47_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12014));
    defparam i10365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10364_3_lut (.I0(\REG.mem_44_15 ), .I1(\REG.mem_45_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12013));
    defparam i10364_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1295_1296 (.Q(\REG.mem_13_3 ), .C(DEBUG_6_c_c), .D(n4897));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14402_bdd_4_lut (.I0(n14402), .I1(\REG.mem_9_11 ), .I2(\REG.mem_8_11 ), 
            .I3(rd_addr_r[1]), .O(n12453));
    defparam n14402_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4524_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_60_15 ), .O(n5726));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4524_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11894 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_14 ), 
            .I2(\REG.mem_15_14 ), .I3(rd_addr_r[1]), .O(n13664));
    defparam rd_addr_r_0__bdd_4_lut_11894.LUT_INIT = 16'he4aa;
    SB_LUT4 n13664_bdd_4_lut (.I0(n13664), .I1(\REG.mem_13_14 ), .I2(\REG.mem_12_14 ), 
            .I3(rd_addr_r[1]), .O(n13667));
    defparam n13664_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12478 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_11 ), 
            .I2(\REG.mem_15_11 ), .I3(rd_addr_r[1]), .O(n14396));
    defparam rd_addr_r_0__bdd_4_lut_12478.LUT_INIT = 16'he4aa;
    SB_LUT4 i4522_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_60_14 ), .O(n5724));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4522_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11864 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_6 ), 
            .I2(\REG.mem_19_6 ), .I3(rd_addr_r[1]), .O(n13658));
    defparam rd_addr_r_0__bdd_4_lut_11864.LUT_INIT = 16'he4aa;
    SB_LUT4 n13658_bdd_4_lut (.I0(n13658), .I1(\REG.mem_17_6 ), .I2(\REG.mem_16_6 ), 
            .I3(rd_addr_r[1]), .O(n13661));
    defparam n13658_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11176 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_15 ), 
            .I2(\REG.mem_19_15 ), .I3(rd_addr_r[1]), .O(n12830));
    defparam rd_addr_r_0__bdd_4_lut_11176.LUT_INIT = 16'he4aa;
    SB_LUT4 n14396_bdd_4_lut (.I0(n14396), .I1(\REG.mem_13_11 ), .I2(\REG.mem_12_11 ), 
            .I3(rd_addr_r[1]), .O(n12456));
    defparam n14396_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1292_1293 (.Q(\REG.mem_13_2 ), .C(DEBUG_6_c_c), .D(n4896));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4521_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_60_13 ), .O(n5723));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4521_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12473 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_6 ), 
            .I2(\REG.mem_55_6 ), .I3(rd_addr_r[1]), .O(n14390));
    defparam rd_addr_r_0__bdd_4_lut_12473.LUT_INIT = 16'he4aa;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i2_1_lut (.I0(rd_addr_r[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1173[1]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4520_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_60_12 ), .O(n5722));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4520_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11859 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_7 ), 
            .I2(\REG.mem_63_7 ), .I3(rd_addr_r[1]), .O(n13652));
    defparam rd_addr_r_0__bdd_4_lut_11859.LUT_INIT = 16'he4aa;
    SB_LUT4 i4519_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_60_11 ), .O(n5721));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4519_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14390_bdd_4_lut (.I0(n14390), .I1(\REG.mem_53_6 ), .I2(\REG.mem_52_6 ), 
            .I3(rd_addr_r[1]), .O(n12459));
    defparam n14390_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10598_3_lut (.I0(\REG.mem_16_14 ), .I1(\REG.mem_17_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12247));
    defparam i10598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10599_3_lut (.I0(\REG.mem_18_14 ), .I1(\REG.mem_19_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12248));
    defparam i10599_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i1289_1290 (.Q(\REG.mem_13_1 ), .C(DEBUG_6_c_c), .D(n4895));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1286_1287 (.Q(\REG.mem_13_0 ), .C(DEBUG_6_c_c), .D(n4894));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1235_1236 (.Q(\REG.mem_12_15 ), .C(DEBUG_6_c_c), .D(n4893));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4518_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_60_10 ), .O(n5720));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4518_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4517_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_60_9 ), .O(n5719));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4517_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4516_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_60_8 ), .O(n5718));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4516_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3982_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_30_13 ), .O(n5184));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3982_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4515_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_60_7 ), .O(n5717));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4515_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4514_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_60_6 ), .O(n5716));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4514_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4513_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_60_5 ), .O(n5715));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4513_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1232_1233 (.Q(\REG.mem_12_14 ), .C(DEBUG_6_c_c), .D(n4892));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4512_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_60_4 ), .O(n5714));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4512_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12468 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_15 ), 
            .I2(\REG.mem_31_15 ), .I3(rd_addr_r[1]), .O(n14384));
    defparam rd_addr_r_0__bdd_4_lut_12468.LUT_INIT = 16'he4aa;
    SB_LUT4 i4511_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_60_3 ), .O(n5713));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4511_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4510_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_60_2 ), .O(n5712));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4510_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4509_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_60_1 ), .O(n5711));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4509_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4508_3_lut_4_lut (.I0(n61_adj_1154), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_60_0 ), .O(n5710));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4508_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i61_2_lut_3_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n61_adj_1154));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i61_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n13652_bdd_4_lut (.I0(n13652), .I1(\REG.mem_61_7 ), .I2(\REG.mem_60_7 ), 
            .I3(rd_addr_r[1]), .O(n12237));
    defparam n13652_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i3_1_lut (.I0(rd_addr_r[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1173[2]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 EnabledDecoder_2_i94_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n53));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i94_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_DFF i1229_1230 (.Q(\REG.mem_12_13 ), .C(DEBUG_6_c_c), .D(n4891));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1226_1227 (.Q(\REG.mem_12_12 ), .C(DEBUG_6_c_c), .D(n4890));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11854 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_6 ), 
            .I2(\REG.mem_23_6 ), .I3(rd_addr_r[1]), .O(n13646));
    defparam rd_addr_r_0__bdd_4_lut_11854.LUT_INIT = 16'he4aa;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i4_1_lut (.I0(rd_addr_r[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1173[3]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 EnabledDecoder_2_i93_2_lut_3_lut_4_lut (.I0(n13), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n21));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i93_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_DFF i1223_1224 (.Q(\REG.mem_12_11 ), .C(DEBUG_6_c_c), .D(n4889));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13646_bdd_4_lut (.I0(n13646), .I1(\REG.mem_21_6 ), .I2(\REG.mem_20_6 ), 
            .I3(rd_addr_r[1]), .O(n13649));
    defparam n13646_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14384_bdd_4_lut (.I0(n14384), .I1(\REG.mem_29_15 ), .I2(\REG.mem_28_15 ), 
            .I3(rd_addr_r[1]), .O(n14387));
    defparam n14384_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1220_1221 (.Q(\REG.mem_12_10 ), .C(DEBUG_6_c_c), .D(n4888));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4501_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_59_15 ), .O(n5703));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4501_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4500_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_59_14 ), .O(n5702));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4500_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4499_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_59_13 ), .O(n5701));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4499_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4498_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_59_12 ), .O(n5700));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4498_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4497_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_59_11 ), .O(n5699));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4497_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4496_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_59_10 ), .O(n5698));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4496_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1217_1218 (.Q(\REG.mem_12_9 ), .C(DEBUG_6_c_c), .D(n4887));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12854_bdd_4_lut (.I0(n12854), .I1(\REG.mem_41_9 ), .I2(\REG.mem_40_9 ), 
            .I3(rd_addr_r[1]), .O(n12857));
    defparam n12854_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4067_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_35_15 ), .O(n5269));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4067_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1214_1215 (.Q(\REG.mem_12_8 ), .C(DEBUG_6_c_c), .D(n4886));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4495_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_59_9 ), .O(n5697));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4495_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4494_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_59_8 ), .O(n5696));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4494_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12463 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_11 ), 
            .I2(\REG.mem_19_11 ), .I3(rd_addr_r[1]), .O(n14378));
    defparam rd_addr_r_0__bdd_4_lut_12463.LUT_INIT = 16'he4aa;
    SB_LUT4 i4493_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_59_7 ), .O(n5695));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4493_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4492_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_59_6 ), .O(n5694));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4492_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1211_1212 (.Q(\REG.mem_12_7 ), .C(DEBUG_6_c_c), .D(n4885));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1208_1209 (.Q(\REG.mem_12_6 ), .C(DEBUG_6_c_c), .D(n4884));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1205_1206 (.Q(\REG.mem_12_5 ), .C(DEBUG_6_c_c), .D(n4883));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1202_1203 (.Q(\REG.mem_12_4 ), .C(DEBUG_6_c_c), .D(n4882));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1199_1200 (.Q(\REG.mem_12_3 ), .C(DEBUG_6_c_c), .D(n4881));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1196_1197 (.Q(\REG.mem_12_2 ), .C(DEBUG_6_c_c), .D(n4880));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1193_1194 (.Q(\REG.mem_12_1 ), .C(DEBUG_6_c_c), .D(n4879));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1190_1191 (.Q(\REG.mem_12_0 ), .C(DEBUG_6_c_c), .D(n4878));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i155_156 (.Q(\REG.mem_1_7 ), .C(DEBUG_6_c_c), .D(n4647));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wp_sync2_r__i0 (.Q(wp_sync2_r[0]), .C(SLM_CLK_c), .D(n4646));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i176_177 (.Q(\REG.mem_1_14 ), .C(DEBUG_6_c_c), .D(n4645));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF wp_sync1_r__i0 (.Q(wp_sync1_r[0]), .C(SLM_CLK_c), .D(n4644));   // src/fifo_dc_32_lut_gen.v(604[21] 616[24])
    SB_DFF i167_168 (.Q(\REG.mem_1_11 ), .C(DEBUG_6_c_c), .D(n4643));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n4642));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    SB_DFF i158_159 (.Q(\REG.mem_1_8 ), .C(DEBUG_6_c_c), .D(n4641));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i143_144 (.Q(\REG.mem_1_3 ), .C(DEBUG_6_c_c), .D(n4640));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync2_r__i0 (.Q(rp_sync2_r[0]), .C(DEBUG_6_c_c), .D(n4639));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i1139_1140 (.Q(\REG.mem_11_15 ), .C(DEBUG_6_c_c), .D(n4877));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4066_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_35_14 ), .O(n5268));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4066_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4491_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_59_5 ), .O(n5693));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4491_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4490_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_59_4 ), .O(n5692));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4490_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4065_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_35_13 ), .O(n5267));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4065_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3971_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_30_2 ), .O(n5173));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3971_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4489_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_59_3 ), .O(n5691));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4489_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4488_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_59_2 ), .O(n5690));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4488_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14378_bdd_4_lut (.I0(n14378), .I1(\REG.mem_17_11 ), .I2(\REG.mem_16_11 ), 
            .I3(rd_addr_r[1]), .O(n12471));
    defparam n14378_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4064_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_35_12 ), .O(n5266));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4064_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1136_1137 (.Q(\REG.mem_11_14 ), .C(DEBUG_6_c_c), .D(n4876));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1133_1134 (.Q(\REG.mem_11_13 ), .C(DEBUG_6_c_c), .D(n4875));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1130_1131 (.Q(\REG.mem_11_12 ), .C(DEBUG_6_c_c), .D(n4874));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1127_1128 (.Q(\REG.mem_11_11 ), .C(DEBUG_6_c_c), .D(n4873));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1124_1125 (.Q(\REG.mem_11_10 ), .C(DEBUG_6_c_c), .D(n4872));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1121_1122 (.Q(\REG.mem_11_9 ), .C(DEBUG_6_c_c), .D(n4871));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1118_1119 (.Q(\REG.mem_11_8 ), .C(DEBUG_6_c_c), .D(n4870));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1115_1116 (.Q(\REG.mem_11_7 ), .C(DEBUG_6_c_c), .D(n4869));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF rp_sync1_r__i0 (.Q(rp_sync1_r[0]), .C(DEBUG_6_c_c), .D(n4638));   // src/fifo_dc_32_lut_gen.v(354[21] 366[24])
    SB_DFF i179_180 (.Q(\REG.mem_1_15 ), .C(DEBUG_6_c_c), .D(n4636));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1112_1113 (.Q(\REG.mem_11_6 ), .C(DEBUG_6_c_c), .D(n4868));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12458 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_6 ), 
            .I2(\REG.mem_59_6 ), .I3(rd_addr_r[1]), .O(n14372));
    defparam rd_addr_r_0__bdd_4_lut_12458.LUT_INIT = 16'he4aa;
    SB_LUT4 i4063_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_35_11 ), .O(n5265));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4063_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4487_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_59_1 ), .O(n5689));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4487_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4486_3_lut_4_lut (.I0(n59_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_59_0 ), .O(n5688));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4486_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11849 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_8 ), 
            .I2(\REG.mem_47_8 ), .I3(rd_addr_r[1]), .O(n13640));
    defparam rd_addr_r_0__bdd_4_lut_11849.LUT_INIT = 16'he4aa;
    SB_LUT4 i4062_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_35_10 ), .O(n5264));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4062_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4061_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_35_9 ), .O(n5263));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4061_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1109_1110 (.Q(\REG.mem_11_5 ), .C(DEBUG_6_c_c), .D(n4867));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1106_1107 (.Q(\REG.mem_11_4 ), .C(DEBUG_6_c_c), .D(n4866));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1103_1104 (.Q(\REG.mem_11_3 ), .C(DEBUG_6_c_c), .D(n4865));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1100_1101 (.Q(\REG.mem_11_2 ), .C(DEBUG_6_c_c), .D(n4864));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1097_1098 (.Q(\REG.mem_11_1 ), .C(DEBUG_6_c_c), .D(n4863));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1094_1095 (.Q(\REG.mem_11_0 ), .C(DEBUG_6_c_c), .D(n4862));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1043_1044 (.Q(\REG.mem_10_15 ), .C(DEBUG_6_c_c), .D(n4861));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1040_1041 (.Q(\REG.mem_10_14 ), .C(DEBUG_6_c_c), .D(n4860));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1037_1038 (.Q(\REG.mem_10_13 ), .C(DEBUG_6_c_c), .D(n4859));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13640_bdd_4_lut (.I0(n13640), .I1(\REG.mem_45_8 ), .I2(\REG.mem_44_8 ), 
            .I3(rd_addr_r[1]), .O(n11820));
    defparam n13640_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n14372_bdd_4_lut (.I0(n14372), .I1(\REG.mem_57_6 ), .I2(\REG.mem_56_6 ), 
            .I3(rd_addr_r[1]), .O(n12474));
    defparam n14372_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i92_2_lut_3_lut_4_lut (.I0(n20_adj_1160), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n54));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i92_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i91_2_lut_3_lut_4_lut (.I0(n20_adj_1160), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n22));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i91_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11844 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_6 ), 
            .I2(\REG.mem_27_6 ), .I3(rd_addr_r[1]), .O(n13634));
    defparam rd_addr_r_0__bdd_4_lut_11844.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12483 (.I0(rd_addr_r[2]), .I1(n13877), 
            .I2(n13943), .I3(rd_addr_r[3]), .O(n14366));
    defparam rd_addr_r_2__bdd_4_lut_12483.LUT_INIT = 16'he4aa;
    SB_LUT4 n14366_bdd_4_lut (.I0(n14366), .I1(n13439), .I2(n12471), .I3(rd_addr_r[3]), 
            .O(n12480));
    defparam n14366_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4060_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_35_8 ), .O(n5262));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4060_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13634_bdd_4_lut (.I0(n13634), .I1(\REG.mem_25_6 ), .I2(\REG.mem_24_6 ), 
            .I3(rd_addr_r[1]), .O(n13637));
    defparam n13634_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3981_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_30_12 ), .O(n5183));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3981_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12453 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_2 ), 
            .I2(\REG.mem_31_2 ), .I3(rd_addr_r[1]), .O(n14360));
    defparam rd_addr_r_0__bdd_4_lut_12453.LUT_INIT = 16'he4aa;
    SB_LUT4 i4059_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_35_7 ), .O(n5261));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4059_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14360_bdd_4_lut (.I0(n14360), .I1(\REG.mem_29_2 ), .I2(\REG.mem_28_2 ), 
            .I3(rd_addr_r[1]), .O(n14363));
    defparam n14360_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4058_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_35_6 ), .O(n5260));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4058_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4057_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_35_5 ), .O(n5259));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4057_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_11884 (.I0(rd_addr_r[3]), .I1(n11572), 
            .I2(n11573), .I3(rd_addr_r[4]), .O(n13628));
    defparam rd_addr_r_3__bdd_4_lut_11884.LUT_INIT = 16'he4aa;
    SB_LUT4 n13628_bdd_4_lut (.I0(n13628), .I1(n11543), .I2(n13199), .I3(rd_addr_r[4]), 
            .O(n13631));
    defparam n13628_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4056_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_35_4 ), .O(n5258));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4056_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i122_2_lut_3_lut (.I0(n25_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n39));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i122_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12448 (.I0(rd_addr_r[2]), .I1(n13187), 
            .I2(n12893), .I3(rd_addr_r[3]), .O(n14354));
    defparam rd_addr_r_2__bdd_4_lut_12448.LUT_INIT = 16'he4aa;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i5_1_lut (.I0(rd_addr_r[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1173[4]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i6_1_lut (.I0(rd_addr_r[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1173[5]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 EnabledDecoder_2_i121_2_lut_3_lut (.I0(n25_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n7_adj_3));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i121_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3440_2_lut_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_p1_w[0]), 
            .I2(rd_fifo_en_w), .I3(reset_all), .O(n4642));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i3440_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i1_2_lut_4_lut (.I0(rd_addr_r[0]), .I1(rd_addr_p1_w[0]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_465[1] ), .O(rd_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i1_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4055_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_35_3 ), .O(n5257));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4055_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4054_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_35_2 ), .O(n5256));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4054_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wp_sync2_r_6__I_0_143_i1_2_lut (.I0(wp_sync2_r[5]), .I1(wp_sync2_r[6]), 
            .I2(GND_net), .I3(GND_net), .O(wp_sync_w[5]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam wp_sync2_r_6__I_0_143_i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n14354_bdd_4_lut (.I0(n14354), .I1(n13427), .I2(n13757), .I3(rd_addr_r[3]), 
            .O(n12486));
    defparam n14354_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1034_1035 (.Q(\REG.mem_10_12 ), .C(DEBUG_6_c_c), .D(n4858));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i1031_1032 (.Q(\REG.mem_10_11 ), .C(DEBUG_6_c_c), .D(n4857));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i2_2_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_465[1] ), .O(rd_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i2_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i3_2_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_465[3] ), .O(rd_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i3_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4053_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_35_1 ), .O(n5255));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4053_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4461_2_lut_4_lut (.I0(rd_addr_r[2]), .I1(rd_addr_p1_w[2]), 
            .I2(rd_fifo_en_w), .I3(reset_all), .O(n5663));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4461_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i4_2_lut_4_lut (.I0(rd_addr_r[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_465[3] ), .O(rd_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i4_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 wp_sync2_r_6__I_0_149_inv_0_i7_1_lut (.I0(\rd_addr_r[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_1173[6]));   // src/fifo_dc_32_lut_gen.v(233[47:78])
    defparam wp_sync2_r_6__I_0_149_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12098 (.I0(rd_addr_r[2]), .I1(n13121), 
            .I2(n12995), .I3(rd_addr_r[3]), .O(n13622));
    defparam rd_addr_r_2__bdd_4_lut_12098.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i5_2_lut_4_lut (.I0(rd_addr_r[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_465[5] ), .O(rd_grey_w[4]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i5_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4459_2_lut_4_lut (.I0(rd_addr_r[4]), .I1(rd_addr_p1_w[4]), 
            .I2(rd_fifo_en_w), .I3(reset_all), .O(n5661));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4459_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i4052_3_lut_4_lut (.I0(n44), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_35_0 ), .O(n5254));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4052_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1028_1029 (.Q(\REG.mem_10_10 ), .C(DEBUG_6_c_c), .D(n4856));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12443 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_4 ), 
            .I2(\REG.mem_51_4 ), .I3(rd_addr_r[1]), .O(n14348));
    defparam rd_addr_r_0__bdd_4_lut_12443.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_nxt_c_6__I_0_152_i6_2_lut_4_lut (.I0(\rd_addr_r[6] ), 
            .I1(rd_addr_p1_w[6]), .I2(rd_fifo_en_w), .I3(\rd_addr_nxt_c_6__N_465[5] ), 
            .O(rd_grey_w[5]));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam rd_addr_nxt_c_6__I_0_152_i6_2_lut_4_lut.LUT_INIT = 16'h35ca;
    SB_LUT4 i4457_2_lut_4_lut (.I0(\rd_addr_r[6] ), .I1(rd_addr_p1_w[6]), 
            .I2(rd_fifo_en_w), .I3(reset_all), .O(n5659));   // src/fifo_dc_32_lut_gen.v(550[59:99])
    defparam i4457_2_lut_4_lut.LUT_INIT = 16'h00ca;
    SB_LUT4 i3970_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_30_1 ), .O(n5172));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3970_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4456_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_57_15 ), .O(n5658));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4456_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4455_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_57_14 ), .O(n5657));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4455_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4454_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_57_13 ), .O(n5656));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4454_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13622_bdd_4_lut (.I0(n13622), .I1(n13181), .I2(n13421), .I3(rd_addr_r[3]), 
            .O(n12240));
    defparam n13622_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1025_1026 (.Q(\REG.mem_10_9 ), .C(DEBUG_6_c_c), .D(n4855));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4453_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_57_12 ), .O(n5655));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4453_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14348_bdd_4_lut (.I0(n14348), .I1(\REG.mem_49_4 ), .I2(\REG.mem_48_4 ), 
            .I3(rd_addr_r[1]), .O(n12006));
    defparam n14348_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4452_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_57_11 ), .O(n5654));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4452_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4451_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_57_10 ), .O(n5653));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4451_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4450_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_57_9 ), .O(n5652));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4450_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4449_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_57_8 ), .O(n5651));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4449_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_4__bdd_4_lut (.I0(rd_addr_r[4]), .I1(n13373), .I2(n13007), 
            .I3(rd_addr_r[5]), .O(n14342));
    defparam rd_addr_r_4__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i4448_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_57_7 ), .O(n5650));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4448_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4447_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_57_6 ), .O(n5649));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4447_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1022_1023 (.Q(\REG.mem_10_8 ), .C(DEBUG_6_c_c), .D(n4854));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14342_bdd_4_lut (.I0(n14342), .I1(n13949), .I2(n12003), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_526 [6]));
    defparam n14342_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4446_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_57_5 ), .O(n5648));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4446_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4445_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_57_4 ), .O(n5647));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4445_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1019_1020 (.Q(\REG.mem_10_7 ), .C(DEBUG_6_c_c), .D(n4853));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11839 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_11 ), 
            .I2(\REG.mem_63_11 ), .I3(rd_addr_r[1]), .O(n13616));
    defparam rd_addr_r_0__bdd_4_lut_11839.LUT_INIT = 16'he4aa;
    SB_LUT4 n13616_bdd_4_lut (.I0(n13616), .I1(\REG.mem_61_11 ), .I2(\REG.mem_60_11 ), 
            .I3(rd_addr_r[1]), .O(n13619));
    defparam n13616_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4444_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_57_3 ), .O(n5646));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4444_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12438 (.I0(rd_addr_r[2]), .I1(n13055), 
            .I2(n13001), .I3(rd_addr_r[3]), .O(n14336));
    defparam rd_addr_r_2__bdd_4_lut_12438.LUT_INIT = 16'he4aa;
    SB_LUT4 i4443_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_57_2 ), .O(n5645));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4443_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4442_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_57_1 ), .O(n5644));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4442_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i1016_1017 (.Q(\REG.mem_10_6 ), .C(DEBUG_6_c_c), .D(n4852));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4441_3_lut_4_lut (.I0(n55_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_57_0 ), .O(n5643));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4441_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11829 (.I0(rd_addr_r[2]), .I1(n12066), 
            .I2(n12093), .I3(rd_addr_r[3]), .O(n13610));
    defparam rd_addr_r_2__bdd_4_lut_11829.LUT_INIT = 16'he4aa;
    SB_DFF i1013_1014 (.Q(\REG.mem_10_5 ), .C(DEBUG_6_c_c), .D(n4851));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i88_2_lut_3_lut_4_lut (.I0(n16_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n56));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i88_2_lut_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 EnabledDecoder_2_i87_2_lut_3_lut_4_lut (.I0(n16_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n24));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i87_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i2_2_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(n7596), .I3(\wr_addr_nxt_c[2] ), .O(wr_grey_w[1]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i2_2_lut_4_lut.LUT_INIT = 16'h53ac;
    SB_LUT4 i4291_2_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(n7596), .I3(reset_all), .O(n5493));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i4291_2_lut_4_lut.LUT_INIT = 16'h00ac;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i1_2_lut_4_lut (.I0(wr_addr_r[1]), .I1(wr_addr_p1_w[1]), 
            .I2(n7596), .I3(wr_addr_nxt_c[0]), .O(wr_grey_w[0]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i1_2_lut_4_lut.LUT_INIT = 16'h53ac;
    SB_LUT4 i3521_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_2_15 ), .O(n4723));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3521_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1010_1011 (.Q(\REG.mem_10_4 ), .C(DEBUG_6_c_c), .D(n4850));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3520_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_2_14 ), .O(n4722));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3520_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3519_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_2_13 ), .O(n4721));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3519_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3518_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_2_12 ), .O(n4720));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3518_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3517_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_2_11 ), .O(n4719));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3517_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1007_1008 (.Q(\REG.mem_10_3 ), .C(DEBUG_6_c_c), .D(n4849));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11191 (.I0(rd_addr_r[0]), .I1(\REG.mem_26_2 ), 
            .I2(\REG.mem_27_2 ), .I3(rd_addr_r[1]), .O(n12848));
    defparam rd_addr_r_0__bdd_4_lut_11191.LUT_INIT = 16'he4aa;
    SB_LUT4 i3516_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_2_10 ), .O(n4718));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3516_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i1004_1005 (.Q(\REG.mem_10_2 ), .C(DEBUG_6_c_c), .D(n4848));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3515_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_2_9 ), .O(n4717));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3515_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n13610_bdd_4_lut (.I0(n13610), .I1(n12054), .I2(n12006), .I3(rd_addr_r[3]), 
            .O(n12246));
    defparam n13610_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3514_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_2_8 ), .O(n4716));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3514_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3513_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_2_7 ), .O(n4715));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3513_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14336_bdd_4_lut (.I0(n14336), .I1(n13127), .I2(n13247), .I3(rd_addr_r[3]), 
            .O(n12012));
    defparam n14336_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i1001_1002 (.Q(\REG.mem_10_1 ), .C(DEBUG_6_c_c), .D(n4847));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3512_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_2_6 ), .O(n4714));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3512_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3511_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_2_5 ), .O(n4713));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3511_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i998_999 (.Q(\REG.mem_10_0 ), .C(DEBUG_6_c_c), .D(n4846));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3980_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_30_11 ), .O(n5182));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3980_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11824 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_2 ), 
            .I2(\REG.mem_63_2 ), .I3(rd_addr_r[1]), .O(n13604));
    defparam rd_addr_r_0__bdd_4_lut_11824.LUT_INIT = 16'he4aa;
    SB_DFF i947_948 (.Q(\REG.mem_9_15 ), .C(DEBUG_6_c_c), .D(n4845));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n12848_bdd_4_lut (.I0(n12848), .I1(\REG.mem_25_2 ), .I2(\REG.mem_24_2 ), 
            .I3(rd_addr_r[1]), .O(n12851));
    defparam n12848_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i944_945 (.Q(\REG.mem_9_14 ), .C(DEBUG_6_c_c), .D(n4844));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13604_bdd_4_lut (.I0(n13604), .I1(\REG.mem_61_2 ), .I2(\REG.mem_60_2 ), 
            .I3(rd_addr_r[1]), .O(n13607));
    defparam n13604_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_1__bdd_4_lut (.I0(rd_addr_r[1]), .I1(n12466), .I2(n12467), 
            .I3(rd_addr_r[2]), .O(n14330));
    defparam rd_addr_r_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i3969_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_30_0 ), .O(n5171));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3969_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14330_bdd_4_lut (.I0(n14330), .I1(n12464), .I2(n12463), .I3(rd_addr_r[2]), 
            .O(n11516));
    defparam n14330_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i941_942 (.Q(\REG.mem_9_13 ), .C(DEBUG_6_c_c), .D(n4843));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3510_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_2_4 ), .O(n4712));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3510_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i938_939 (.Q(\REG.mem_9_12 ), .C(DEBUG_6_c_c), .D(n4842));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3509_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_2_3 ), .O(n4711));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3509_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_12423 (.I0(rd_addr_r[2]), .I1(n13751), 
            .I2(n13619), .I3(rd_addr_r[3]), .O(n14324));
    defparam rd_addr_r_2__bdd_4_lut_12423.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11814 (.I0(rd_addr_r[0]), .I1(\REG.mem_30_6 ), 
            .I2(\REG.mem_31_6 ), .I3(rd_addr_r[1]), .O(n13598));
    defparam rd_addr_r_0__bdd_4_lut_11814.LUT_INIT = 16'he4aa;
    SB_LUT4 n13598_bdd_4_lut (.I0(n13598), .I1(\REG.mem_29_6 ), .I2(\REG.mem_28_6 ), 
            .I3(rd_addr_r[1]), .O(n13601));
    defparam n13598_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_52 (.I0(DEBUG_5_c), .I1(get_next_word), .I2(GND_net), 
            .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(560[21] 576[24])
    defparam i1_2_lut_adj_52.LUT_INIT = 16'h4444;
    SB_LUT4 i3508_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_2_2 ), .O(n4710));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3508_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4033_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_33_15 ), .O(n5235));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4033_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3507_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_2_1 ), .O(n4709));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3507_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14324_bdd_4_lut (.I0(n14324), .I1(n14147), .I2(n14207), .I3(rd_addr_r[3]), 
            .O(n12498));
    defparam n14324_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i935_936 (.Q(\REG.mem_9_11 ), .C(DEBUG_6_c_c), .D(n4841));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i10468_3_lut (.I0(n13709), .I1(n14081), .I2(rd_addr_r[5]), 
            .I3(GND_net), .O(\REG.out_raw_31__N_526 [0]));
    defparam i10468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4032_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_33_14 ), .O(n5234));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4032_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n12830_bdd_4_lut (.I0(n12830), .I1(\REG.mem_17_15 ), .I2(\REG.mem_16_15 ), 
            .I3(rd_addr_r[1]), .O(n12833));
    defparam n12830_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i932_933 (.Q(\REG.mem_9_10 ), .C(DEBUG_6_c_c), .D(n4840));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i3506_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_2_0 ), .O(n4708));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3506_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11809 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_13 ), 
            .I2(\REG.mem_51_13 ), .I3(rd_addr_r[1]), .O(n13592));
    defparam rd_addr_r_0__bdd_4_lut_11809.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_12428 (.I0(rd_addr_r[4]), .I1(n12486), 
            .I2(n12498), .I3(rd_addr_r[5]), .O(n14318));
    defparam rd_addr_r_4__bdd_4_lut_12428.LUT_INIT = 16'he4aa;
    SB_LUT4 n13592_bdd_4_lut (.I0(n13592), .I1(\REG.mem_49_13 ), .I2(\REG.mem_48_13 ), 
            .I3(rd_addr_r[1]), .O(n12255));
    defparam n13592_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i929_930 (.Q(\REG.mem_9_9 ), .C(DEBUG_6_c_c), .D(n4839));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14318_bdd_4_lut (.I0(n14318), .I1(n12480), .I2(n13157), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_526 [11]));
    defparam n14318_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4031_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_33_13 ), .O(n5233));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4031_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9860_3_lut (.I0(\REG.mem_56_12 ), .I1(\REG.mem_57_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11509));
    defparam i9860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9861_3_lut (.I0(\REG.mem_58_12 ), .I1(\REG.mem_59_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11510));
    defparam i9861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_4__bdd_4_lut_12408 (.I0(rd_addr_r[4]), .I1(n11991), 
            .I2(n12012), .I3(rd_addr_r[5]), .O(n14312));
    defparam rd_addr_r_4__bdd_4_lut_12408.LUT_INIT = 16'he4aa;
    SB_LUT4 i9882_3_lut (.I0(\REG.mem_62_12 ), .I1(\REG.mem_63_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11531));
    defparam i9882_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF i134_135 (.Q(\REG.mem_1_0 ), .C(DEBUG_6_c_c), .D(n4614));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 EnabledDecoder_2_i25_2_lut_3_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n25_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i25_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i4030_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_33_12 ), .O(n5232));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4030_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9881_3_lut (.I0(\REG.mem_60_12 ), .I1(\REG.mem_61_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11530));
    defparam i9881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3979_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_30_10 ), .O(n5181));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3979_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14312_bdd_4_lut (.I0(n14312), .I1(n11976), .I2(n12809), .I3(rd_addr_r[5]), 
            .O(\REG.out_raw_31__N_526 [3]));
    defparam n14312_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i26_2_lut_3_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(GND_net), .O(n26_adj_1146));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i26_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11804 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_0 ), 
            .I2(\REG.mem_19_0 ), .I3(rd_addr_r[1]), .O(n13586));
    defparam rd_addr_r_0__bdd_4_lut_11804.LUT_INIT = 16'he4aa;
    SB_LUT4 i9998_3_lut (.I0(\REG.mem_16_3 ), .I1(\REG.mem_17_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11647));
    defparam i9998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9999_3_lut (.I0(\REG.mem_18_3 ), .I1(\REG.mem_19_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11648));
    defparam i9999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i13_2_lut_3_lut_4_lut (.I0(n7596), .I1(\wr_addr_r[0] ), 
            .I2(wr_addr_r[2]), .I3(wr_addr_r[1]), .O(n13));
    defparam EnabledDecoder_2_i13_2_lut_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i6433_2_lut_3_lut_4_lut (.I0(n7596), .I1(\wr_addr_r[0] ), .I2(wr_addr_r[2]), 
            .I3(wr_addr_r[1]), .O(n7612));
    defparam i6433_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4440_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_56_15 ), .O(n5642));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4440_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6417_2_lut (.I0(\afull_flag_impl.af_flag_p_w_N_603[3] ), .I1(full_o), 
            .I2(GND_net), .I3(GND_net), .O(n7596));
    defparam i6417_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i4439_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_56_14 ), .O(n5641));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4439_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n13586_bdd_4_lut (.I0(n13586), .I1(\REG.mem_17_0 ), .I2(\REG.mem_16_0 ), 
            .I3(rd_addr_r[1]), .O(n13589));
    defparam n13586_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4029_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_33_11 ), .O(n5231));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4029_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4438_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_56_13 ), .O(n5640));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4438_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_2__bdd_4_lut_11819 (.I0(rd_addr_r[2]), .I1(n12126), 
            .I2(n12129), .I3(rd_addr_r[3]), .O(n13580));
    defparam rd_addr_r_2__bdd_4_lut_11819.LUT_INIT = 16'he4aa;
    SB_LUT4 i4437_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_56_12 ), .O(n5639));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4437_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i146_147 (.Q(\REG.mem_1_4 ), .C(DEBUG_6_c_c), .D(n4613));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4436_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_56_11 ), .O(n5638));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4436_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12433 (.I0(rd_addr_r[0]), .I1(\REG.mem_14_3 ), 
            .I2(\REG.mem_15_3 ), .I3(rd_addr_r[1]), .O(n14306));
    defparam rd_addr_r_0__bdd_4_lut_12433.LUT_INIT = 16'he4aa;
    SB_LUT4 i4028_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_33_10 ), .O(n5230));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4028_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14306_bdd_4_lut (.I0(n14306), .I1(\REG.mem_13_3 ), .I2(\REG.mem_12_3 ), 
            .I3(rd_addr_r[1]), .O(n11625));
    defparam n14306_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n13580_bdd_4_lut (.I0(n13580), .I1(n12120), .I2(n12111), .I3(rd_addr_r[3]), 
            .O(n12258));
    defparam n13580_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4435_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_56_10 ), .O(n5637));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4435_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i926_927 (.Q(\REG.mem_9_8 ), .C(DEBUG_6_c_c), .D(n4838));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i923_924 (.Q(\REG.mem_9_7 ), .C(DEBUG_6_c_c), .D(n4837));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i920_921 (.Q(\REG.mem_9_6 ), .C(DEBUG_6_c_c), .D(n4836));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i917_918 (.Q(\REG.mem_9_5 ), .C(DEBUG_6_c_c), .D(n4835));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i914_915 (.Q(\REG.mem_9_4 ), .C(DEBUG_6_c_c), .D(n4834));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i911_912 (.Q(\REG.mem_9_3 ), .C(DEBUG_6_c_c), .D(n4833));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i908_909 (.Q(\REG.mem_9_2 ), .C(DEBUG_6_c_c), .D(n4832));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i905_906 (.Q(\REG.mem_9_1 ), .C(DEBUG_6_c_c), .D(n4831));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i902_903 (.Q(\REG.mem_9_0 ), .C(DEBUG_6_c_c), .D(n4830));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i851_852 (.Q(\REG.mem_8_15 ), .C(DEBUG_6_c_c), .D(n4829));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i848_849 (.Q(\REG.mem_8_14 ), .C(DEBUG_6_c_c), .D(n4828));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i845_846 (.Q(\REG.mem_8_13 ), .C(DEBUG_6_c_c), .D(n4827));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i842_843 (.Q(\REG.mem_8_12 ), .C(DEBUG_6_c_c), .D(n4826));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i839_840 (.Q(\REG.mem_8_11 ), .C(DEBUG_6_c_c), .D(n4825));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i836_837 (.Q(\REG.mem_8_10 ), .C(DEBUG_6_c_c), .D(n4824));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i833_834 (.Q(\REG.mem_8_9 ), .C(DEBUG_6_c_c), .D(n4823));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i830_831 (.Q(\REG.mem_8_8 ), .C(DEBUG_6_c_c), .D(n4822));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i827_828 (.Q(\REG.mem_8_7 ), .C(DEBUG_6_c_c), .D(n4821));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i824_825 (.Q(\REG.mem_8_6 ), .C(DEBUG_6_c_c), .D(n4820));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i821_822 (.Q(\REG.mem_8_5 ), .C(DEBUG_6_c_c), .D(n4819));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i818_819 (.Q(\REG.mem_8_4 ), .C(DEBUG_6_c_c), .D(n4818));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i815_816 (.Q(\REG.mem_8_3 ), .C(DEBUG_6_c_c), .D(n4817));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i812_813 (.Q(\REG.mem_8_2 ), .C(DEBUG_6_c_c), .D(n4816));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i809_810 (.Q(\REG.mem_8_1 ), .C(DEBUG_6_c_c), .D(n4815));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i806_807 (.Q(\REG.mem_8_0 ), .C(DEBUG_6_c_c), .D(n4814));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i755_756 (.Q(\REG.mem_7_15 ), .C(DEBUG_6_c_c), .D(n4813));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i752_753 (.Q(\REG.mem_7_14 ), .C(DEBUG_6_c_c), .D(n4812));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i749_750 (.Q(\REG.mem_7_13 ), .C(DEBUG_6_c_c), .D(n4811));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i746_747 (.Q(\REG.mem_7_12 ), .C(DEBUG_6_c_c), .D(n4810));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i743_744 (.Q(\REG.mem_7_11 ), .C(DEBUG_6_c_c), .D(n4809));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i740_741 (.Q(\REG.mem_7_10 ), .C(DEBUG_6_c_c), .D(n4808));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i737_738 (.Q(\REG.mem_7_9 ), .C(DEBUG_6_c_c), .D(n4807));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i734_735 (.Q(\REG.mem_7_8 ), .C(DEBUG_6_c_c), .D(n4806));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i731_732 (.Q(\REG.mem_7_7 ), .C(DEBUG_6_c_c), .D(n4805));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i728_729 (.Q(\REG.mem_7_6 ), .C(DEBUG_6_c_c), .D(n4804));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i725_726 (.Q(\REG.mem_7_5 ), .C(DEBUG_6_c_c), .D(n4803));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i722_723 (.Q(\REG.mem_7_4 ), .C(DEBUG_6_c_c), .D(n4802));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i719_720 (.Q(\REG.mem_7_3 ), .C(DEBUG_6_c_c), .D(n4801));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i716_717 (.Q(\REG.mem_7_2 ), .C(DEBUG_6_c_c), .D(n4800));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i713_714 (.Q(\REG.mem_7_1 ), .C(DEBUG_6_c_c), .D(n4799));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i710_711 (.Q(\REG.mem_7_0 ), .C(DEBUG_6_c_c), .D(n4798));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i659_660 (.Q(\REG.mem_6_15 ), .C(DEBUG_6_c_c), .D(n4797));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i656_657 (.Q(\REG.mem_6_14 ), .C(DEBUG_6_c_c), .D(n4796));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i653_654 (.Q(\REG.mem_6_13 ), .C(DEBUG_6_c_c), .D(n4795));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i650_651 (.Q(\REG.mem_6_12 ), .C(DEBUG_6_c_c), .D(n4794));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i647_648 (.Q(\REG.mem_6_11 ), .C(DEBUG_6_c_c), .D(n4793));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i644_645 (.Q(\REG.mem_6_10 ), .C(DEBUG_6_c_c), .D(n4792));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i641_642 (.Q(\REG.mem_6_9 ), .C(DEBUG_6_c_c), .D(n4791));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i638_639 (.Q(\REG.mem_6_8 ), .C(DEBUG_6_c_c), .D(n4790));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i635_636 (.Q(\REG.mem_6_7 ), .C(DEBUG_6_c_c), .D(n4789));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i632_633 (.Q(\REG.mem_6_6 ), .C(DEBUG_6_c_c), .D(n4788));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i629_630 (.Q(\REG.mem_6_5 ), .C(DEBUG_6_c_c), .D(n4787));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i626_627 (.Q(\REG.mem_6_4 ), .C(DEBUG_6_c_c), .D(n4786));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i623_624 (.Q(\REG.mem_6_3 ), .C(DEBUG_6_c_c), .D(n4785));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i620_621 (.Q(\REG.mem_6_2 ), .C(DEBUG_6_c_c), .D(n4784));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i617_618 (.Q(\REG.mem_6_1 ), .C(DEBUG_6_c_c), .D(n4783));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i614_615 (.Q(\REG.mem_6_0 ), .C(DEBUG_6_c_c), .D(n4779));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4434_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_56_9 ), .O(n5636));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4434_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4027_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_33_9 ), .O(n5229));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4027_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF i563_564 (.Q(\REG.mem_5_15 ), .C(DEBUG_6_c_c), .D(n4778));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i560_561 (.Q(\REG.mem_5_14 ), .C(DEBUG_6_c_c), .D(n4777));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i557_558 (.Q(\REG.mem_5_13 ), .C(DEBUG_6_c_c), .D(n4776));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i554_555 (.Q(\REG.mem_5_12 ), .C(DEBUG_6_c_c), .D(n4775));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i551_552 (.Q(\REG.mem_5_11 ), .C(DEBUG_6_c_c), .D(n4774));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i548_549 (.Q(\REG.mem_5_10 ), .C(DEBUG_6_c_c), .D(n4773));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i545_546 (.Q(\REG.mem_5_9 ), .C(DEBUG_6_c_c), .D(n4772));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i542_543 (.Q(\REG.mem_5_8 ), .C(DEBUG_6_c_c), .D(n4771));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i539_540 (.Q(\REG.mem_5_7 ), .C(DEBUG_6_c_c), .D(n4770));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i536_537 (.Q(\REG.mem_5_6 ), .C(DEBUG_6_c_c), .D(n4769));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i533_534 (.Q(\REG.mem_5_5 ), .C(DEBUG_6_c_c), .D(n4768));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i530_531 (.Q(\REG.mem_5_4 ), .C(DEBUG_6_c_c), .D(n4767));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i527_528 (.Q(\REG.mem_5_3 ), .C(DEBUG_6_c_c), .D(n4766));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i524_525 (.Q(\REG.mem_5_2 ), .C(DEBUG_6_c_c), .D(n4765));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i521_522 (.Q(\REG.mem_5_1 ), .C(DEBUG_6_c_c), .D(n4764));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i518_519 (.Q(\REG.mem_5_0 ), .C(DEBUG_6_c_c), .D(n4763));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i467_468 (.Q(\REG.mem_4_15 ), .C(DEBUG_6_c_c), .D(n4762));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i464_465 (.Q(\REG.mem_4_14 ), .C(DEBUG_6_c_c), .D(n4761));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i461_462 (.Q(\REG.mem_4_13 ), .C(DEBUG_6_c_c), .D(n4760));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i458_459 (.Q(\REG.mem_4_12 ), .C(DEBUG_6_c_c), .D(n4759));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i455_456 (.Q(\REG.mem_4_11 ), .C(DEBUG_6_c_c), .D(n4758));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i452_453 (.Q(\REG.mem_4_10 ), .C(DEBUG_6_c_c), .D(n4757));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i449_450 (.Q(\REG.mem_4_9 ), .C(DEBUG_6_c_c), .D(n4756));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i446_447 (.Q(\REG.mem_4_8 ), .C(DEBUG_6_c_c), .D(n4755));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i443_444 (.Q(\REG.mem_4_7 ), .C(DEBUG_6_c_c), .D(n4754));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i440_441 (.Q(\REG.mem_4_6 ), .C(DEBUG_6_c_c), .D(n4753));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i437_438 (.Q(\REG.mem_4_5 ), .C(DEBUG_6_c_c), .D(n4752));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i434_435 (.Q(\REG.mem_4_4 ), .C(DEBUG_6_c_c), .D(n4751));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i431_432 (.Q(\REG.mem_4_3 ), .C(DEBUG_6_c_c), .D(n4750));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i428_429 (.Q(\REG.mem_4_2 ), .C(DEBUG_6_c_c), .D(n4749));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i425_426 (.Q(\REG.mem_4_1 ), .C(DEBUG_6_c_c), .D(n4748));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i422_423 (.Q(\REG.mem_4_0 ), .C(DEBUG_6_c_c), .D(n4747));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4433_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_56_8 ), .O(n5635));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4433_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3978_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_30_9 ), .O(n5180));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3978_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 EnabledDecoder_2_i20_2_lut (.I0(n11), .I1(wr_addr_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_1160));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i20_2_lut.LUT_INIT = 16'h2222;
    SB_DFF wr_addr_r__i0 (.Q(\wr_addr_r[0] ), .C(DEBUG_6_c_c), .D(n4612));   // src/fifo_dc_32_lut_gen.v(310[21] 326[24])
    SB_LUT4 i4432_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_56_7 ), .O(n5634));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4432_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4431_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_56_6 ), .O(n5633));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4431_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4026_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_33_8 ), .O(n5228));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4026_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_3__bdd_4_lut (.I0(rd_addr_r[3]), .I1(n13169), .I2(n11516), 
            .I3(rd_addr_r[4]), .O(n14300));
    defparam rd_addr_r_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i4430_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_56_5 ), .O(n5632));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4430_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4429_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_56_4 ), .O(n5631));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4429_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4428_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_56_3 ), .O(n5630));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4428_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10026_3_lut (.I0(\REG.mem_22_3 ), .I1(\REG.mem_23_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11675));
    defparam i10026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10025_3_lut (.I0(\REG.mem_20_3 ), .I1(\REG.mem_21_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11674));
    defparam i10025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11186 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_10 ), 
            .I2(\REG.mem_63_10 ), .I3(rd_addr_r[1]), .O(n12842));
    defparam rd_addr_r_0__bdd_4_lut_11186.LUT_INIT = 16'he4aa;
    SB_LUT4 i4427_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_56_2 ), .O(n5629));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4427_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n14300_bdd_4_lut (.I0(n14300), .I1(n11501), .I2(n11500), .I3(rd_addr_r[4]), 
            .O(n14303));
    defparam n14300_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4426_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_56_1 ), .O(n5628));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4426_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4425_3_lut_4_lut (.I0(n53_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_56_0 ), .O(n5627));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4425_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11799 (.I0(rd_addr_r[0]), .I1(\REG.mem_46_5 ), 
            .I2(\REG.mem_47_5 ), .I3(rd_addr_r[1]), .O(n13574));
    defparam rd_addr_r_0__bdd_4_lut_11799.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12398 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_6 ), 
            .I2(\REG.mem_63_6 ), .I3(rd_addr_r[1]), .O(n14294));
    defparam rd_addr_r_0__bdd_4_lut_12398.LUT_INIT = 16'he4aa;
    SB_LUT4 n14294_bdd_4_lut (.I0(n14294), .I1(\REG.mem_61_6 ), .I2(\REG.mem_60_6 ), 
            .I3(rd_addr_r[1]), .O(n11634));
    defparam n14294_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF i161_162 (.Q(\REG.mem_1_9 ), .C(DEBUG_6_c_c), .D(n4610));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13574_bdd_4_lut (.I0(n13574), .I1(\REG.mem_45_5 ), .I2(\REG.mem_44_5 ), 
            .I3(rd_addr_r[1]), .O(n13577));
    defparam n13574_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12388 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_2 ), 
            .I2(\REG.mem_35_2 ), .I3(rd_addr_r[1]), .O(n14288));
    defparam rd_addr_r_0__bdd_4_lut_12388.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11789 (.I0(rd_addr_r[0]), .I1(\REG.mem_34_6 ), 
            .I2(\REG.mem_35_6 ), .I3(rd_addr_r[1]), .O(n13568));
    defparam rd_addr_r_0__bdd_4_lut_11789.LUT_INIT = 16'he4aa;
    SB_LUT4 n12842_bdd_4_lut (.I0(n12842), .I1(\REG.mem_61_10 ), .I2(\REG.mem_60_10 ), 
            .I3(rd_addr_r[1]), .O(n12845));
    defparam n12842_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10623_3_lut (.I0(\REG.mem_22_14 ), .I1(\REG.mem_23_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12272));
    defparam i10623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n13568_bdd_4_lut (.I0(n13568), .I1(\REG.mem_33_6 ), .I2(\REG.mem_32_6 ), 
            .I3(rd_addr_r[1]), .O(n11835));
    defparam n13568_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10622_3_lut (.I0(\REG.mem_20_14 ), .I1(\REG.mem_21_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12271));
    defparam i10622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n14288_bdd_4_lut (.I0(n14288), .I1(\REG.mem_33_2 ), .I2(\REG.mem_32_2 ), 
            .I3(rd_addr_r[1]), .O(n12030));
    defparam n14288_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9902_3_lut (.I0(\REG.mem_8_4 ), .I1(\REG.mem_9_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11551));
    defparam i9902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9903_3_lut (.I0(\REG.mem_10_4 ), .I1(\REG.mem_11_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11552));
    defparam i9903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9990_3_lut (.I0(\REG.mem_14_4 ), .I1(\REG.mem_15_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11639));
    defparam i9990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11869 (.I0(rd_addr_r[1]), .I1(n11761), 
            .I2(n11762), .I3(rd_addr_r[2]), .O(n13562));
    defparam rd_addr_r_1__bdd_4_lut_11869.LUT_INIT = 16'he4aa;
    SB_LUT4 i9989_3_lut (.I0(\REG.mem_12_4 ), .I1(\REG.mem_13_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11638));
    defparam i9989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i53_2_lut_3_lut (.I0(n7612), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[4]), .I3(GND_net), .O(n53_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i53_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 EnabledDecoder_2_i86_2_lut_3_lut_4_lut (.I0(n7612), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n57));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i86_2_lut_3_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12418 (.I0(rd_addr_r[1]), .I1(n12025), 
            .I2(n12026), .I3(rd_addr_r[2]), .O(n14282));
    defparam rd_addr_r_1__bdd_4_lut_12418.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i85_2_lut_3_lut_4_lut (.I0(n7612), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n25));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i85_2_lut_3_lut_4_lut.LUT_INIT = 16'h0040;
    SB_DFF i149_150 (.Q(\REG.mem_1_5 ), .C(DEBUG_6_c_c), .D(n4608));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n13562_bdd_4_lut (.I0(n13562), .I1(n11732), .I2(n11731), .I3(rd_addr_r[2]), 
            .O(n13565));
    defparam n13562_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10682_3_lut (.I0(\REG.mem_32_14 ), .I1(\REG.mem_33_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12331));
    defparam i10682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10683_3_lut (.I0(\REG.mem_34_14 ), .I1(\REG.mem_35_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12332));
    defparam i10683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3977_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_30_8 ), .O(n5179));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3977_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14282_bdd_4_lut (.I0(n14282), .I1(n11981), .I2(n11980), .I3(rd_addr_r[2]), 
            .O(n12512));
    defparam n14282_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11181 (.I0(rd_addr_r[0]), .I1(\REG.mem_58_14 ), 
            .I2(\REG.mem_59_14 ), .I3(rd_addr_r[1]), .O(n12836));
    defparam rd_addr_r_0__bdd_4_lut_11181.LUT_INIT = 16'he4aa;
    SB_LUT4 i4025_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_33_7 ), .O(n5227));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4025_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4024_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_33_6 ), .O(n5226));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4024_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i116_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n42));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i116_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 EnabledDecoder_2_i115_2_lut_3_lut (.I0(n36), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n10));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i115_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12378 (.I0(rd_addr_r[1]), .I1(n11506), 
            .I2(n11507), .I3(rd_addr_r[2]), .O(n14276));
    defparam rd_addr_r_1__bdd_4_lut_12378.LUT_INIT = 16'he4aa;
    SB_LUT4 n14276_bdd_4_lut (.I0(n14276), .I1(n12509), .I2(n12508), .I3(rd_addr_r[2]), 
            .O(n12499));
    defparam n14276_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12383 (.I0(rd_addr_r[0]), .I1(\REG.mem_62_14 ), 
            .I2(\REG.mem_63_14 ), .I3(rd_addr_r[1]), .O(n14270));
    defparam rd_addr_r_0__bdd_4_lut_12383.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11784 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_6 ), 
            .I2(\REG.mem_39_6 ), .I3(rd_addr_r[1]), .O(n13550));
    defparam rd_addr_r_0__bdd_4_lut_11784.LUT_INIT = 16'he4aa;
    SB_LUT4 n14270_bdd_4_lut (.I0(n14270), .I1(\REG.mem_61_14 ), .I2(\REG.mem_60_14 ), 
            .I3(rd_addr_r[1]), .O(n14273));
    defparam n14270_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 wr_addr_r_6__I_0_add_2_6_lut (.I0(n3_adj_1166), .I1(wr_addr_r[4]), 
            .I2(rp_sync_w[4]), .I3(n10628), .O(n11436)) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_6_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i4023_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_33_5 ), .O(n5225));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4023_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3469_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_0_15 ), .O(n4671));
    defparam i3469_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3473_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_0_14 ), .O(n4675));
    defparam i3473_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3478_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_0_13 ), .O(n4680));
    defparam i3478_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4022_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_33_4 ), .O(n5224));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4022_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4021_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_33_3 ), .O(n5223));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4021_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3479_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_0_12 ), .O(n4681));
    defparam i3479_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n13550_bdd_4_lut (.I0(n13550), .I1(\REG.mem_37_6 ), .I2(\REG.mem_36_6 ), 
            .I3(rd_addr_r[1]), .O(n11838));
    defparam n13550_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3480_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_0_11 ), .O(n4682));
    defparam i3480_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF i371_372 (.Q(\REG.mem_3_15 ), .C(DEBUG_6_c_c), .D(n4741));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_CARRY wr_addr_r_6__I_0_add_2_6 (.CI(n10628), .I0(wr_addr_r[4]), .I1(rp_sync_w[4]), 
            .CO(n10629));
    SB_LUT4 EnabledDecoder_2_i15_2_lut (.I0(n12_adj_1156), .I1(wr_addr_r[2]), 
            .I2(GND_net), .I3(GND_net), .O(n15_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i15_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3481_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_0_10 ), .O(n4683));
    defparam i3481_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n12836_bdd_4_lut (.I0(n12836), .I1(\REG.mem_57_14 ), .I2(\REG.mem_56_14 ), 
            .I3(rd_addr_r[1]), .O(n12839));
    defparam n12836_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4020_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_33_2 ), .O(n5222));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4020_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3482_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_0_9 ), .O(n4684));
    defparam i3482_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n12818_bdd_4_lut (.I0(n12818), .I1(n12089), .I2(n12088), .I3(rd_addr_r[2]), 
            .O(n12821));
    defparam n12818_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3485_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_0_8 ), .O(n4687));
    defparam i3485_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4019_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_33_1 ), .O(n5221));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4019_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3486_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_0_7 ), .O(n4688));
    defparam i3486_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3487_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_0_6 ), .O(n4689));
    defparam i3487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3489_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_0_5 ), .O(n4691));
    defparam i3489_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3500_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_0_4 ), .O(n4702));
    defparam i3500_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3502_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_0_3 ), .O(n4704));
    defparam i3502_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4018_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_33_0 ), .O(n5220));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4018_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12368 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_3 ), 
            .I2(\REG.mem_3_3 ), .I3(rd_addr_r[1]), .O(n14264));
    defparam rd_addr_r_0__bdd_4_lut_12368.LUT_INIT = 16'he4aa;
    SB_LUT4 i3503_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_0_2 ), .O(n4705));
    defparam i3503_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i3_2_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(n7596), .I3(\wr_addr_nxt_c[2] ), .O(wr_grey_w[2]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i3_2_lut_4_lut.LUT_INIT = 16'h53ac;
    SB_LUT4 n14264_bdd_4_lut (.I0(n14264), .I1(\REG.mem_1_3 ), .I2(\REG.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(n11523));
    defparam n14264_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3504_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_0_1 ), .O(n4706));
    defparam i3504_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 wr_addr_nxt_c_6__I_0_150_i4_2_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(n7596), .I3(\wr_addr_nxt_c[4] ), .O(wr_grey_w[3]));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam wr_addr_nxt_c_6__I_0_150_i4_2_lut_4_lut.LUT_INIT = 16'h53ac;
    SB_LUT4 i10142_3_lut (.I0(\REG.mem_32_3 ), .I1(\REG.mem_33_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11791));
    defparam i10142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3505_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_0_0 ), .O(n4707));
    defparam i3505_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4273_2_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_p1_w[3]), 
            .I2(n7596), .I3(reset_all), .O(n5475));   // src/fifo_dc_32_lut_gen.v(305[33:89])
    defparam i4273_2_lut_4_lut.LUT_INIT = 16'h00ac;
    SB_LUT4 i3402_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_1_10 ), .O(n4604));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3402_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12393 (.I0(rd_addr_r[3]), .I1(n13217), 
            .I2(n11555), .I3(rd_addr_r[4]), .O(n14258));
    defparam rd_addr_r_3__bdd_4_lut_12393.LUT_INIT = 16'he4aa;
    SB_LUT4 i3406_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_1_5 ), .O(n4608));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3406_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3464_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_1_1 ), .O(n4666));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3464_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10143_3_lut (.I0(\REG.mem_34_3 ), .I1(\REG.mem_35_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11792));
    defparam i10143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3443_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_1_14 ), .O(n4645));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3443_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3463_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_1_6 ), .O(n4665));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3463_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n14258_bdd_4_lut (.I0(n14258), .I1(n11489), .I2(n12821), .I3(rd_addr_r[4]), 
            .O(n14261));
    defparam n14258_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3411_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_1_4 ), .O(n4613));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3411_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4017_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_32_15 ), .O(n5219));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4017_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4016_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_32_14 ), .O(n5218));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4016_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10707_3_lut (.I0(\REG.mem_38_14 ), .I1(\REG.mem_39_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12356));
    defparam i10707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3438_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_1_3 ), .O(n4640));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3438_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10706_3_lut (.I0(\REG.mem_36_14 ), .I1(\REG.mem_37_14 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12355));
    defparam i10706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3446_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_1_2 ), .O(n4648));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3446_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i368_369 (.Q(\REG.mem_3_14 ), .C(DEBUG_6_c_c), .D(n4739));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i365_366 (.Q(\REG.mem_3_13 ), .C(DEBUG_6_c_c), .D(n4738));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_1__bdd_4_lut_12373 (.I0(rd_addr_r[1]), .I1(n12493), 
            .I2(n12494), .I3(rd_addr_r[2]), .O(n14252));
    defparam rd_addr_r_1__bdd_4_lut_12373.LUT_INIT = 16'he4aa;
    SB_DFF i362_363 (.Q(\REG.mem_3_12 ), .C(DEBUG_6_c_c), .D(n4737));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14252_bdd_4_lut (.I0(n14252), .I1(n12488), .I2(n12487), .I3(rd_addr_r[2]), 
            .O(n14255));
    defparam n14252_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3488_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_1_13 ), .O(n4690));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3488_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3412_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_1_0 ), .O(n4614));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3412_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i359_360 (.Q(\REG.mem_3_11 ), .C(DEBUG_6_c_c), .D(n4736));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i356_357 (.Q(\REG.mem_3_10 ), .C(DEBUG_6_c_c), .D(n4735));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i353_354 (.Q(\REG.mem_3_9 ), .C(DEBUG_6_c_c), .D(n4734));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 i4015_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_32_13 ), .O(n5217));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4015_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3434_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_1_15 ), .O(n4636));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3434_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3445_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_1_7 ), .O(n4647));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3445_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i350_351 (.Q(\REG.mem_3_8 ), .C(DEBUG_6_c_c), .D(n4733));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12363 (.I0(rd_addr_r[0]), .I1(\REG.mem_10_8 ), 
            .I2(\REG.mem_11_8 ), .I3(rd_addr_r[1]), .O(n14246));
    defparam rd_addr_r_0__bdd_4_lut_12363.LUT_INIT = 16'he4aa;
    SB_LUT4 i4014_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_32_12 ), .O(n5216));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4014_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11769 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_8 ), 
            .I2(\REG.mem_51_8 ), .I3(rd_addr_r[1]), .O(n13532));
    defparam rd_addr_r_0__bdd_4_lut_11769.LUT_INIT = 16'he4aa;
    SB_LUT4 n14246_bdd_4_lut (.I0(n14246), .I1(\REG.mem_9_8 ), .I2(\REG.mem_8_8 ), 
            .I3(rd_addr_r[1]), .O(n11646));
    defparam n14246_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3976_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_30_7 ), .O(n5178));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3976_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3476_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_1_12 ), .O(n4678));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3476_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3408_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_1_9 ), .O(n4610));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3408_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4013_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_32_11 ), .O(n5215));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4013_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n13532_bdd_4_lut (.I0(n13532), .I1(\REG.mem_49_8 ), .I2(\REG.mem_48_8 ), 
            .I3(rd_addr_r[1]), .O(n11841));
    defparam n13532_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4012_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_32_10 ), .O(n5214));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4012_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3439_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_1_8 ), .O(n4641));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3439_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3441_3_lut_4_lut (.I0(n40), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_1_11 ), .O(n4643));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3441_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF i347_348 (.Q(\REG.mem_3_7 ), .C(DEBUG_6_c_c), .D(n4732));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_DFF i344_345 (.Q(\REG.mem_3_6 ), .C(DEBUG_6_c_c), .D(n4731));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12348 (.I0(rd_addr_r[0]), .I1(\REG.mem_2_13 ), 
            .I2(\REG.mem_3_13 ), .I3(rd_addr_r[1]), .O(n14240));
    defparam rd_addr_r_0__bdd_4_lut_12348.LUT_INIT = 16'he4aa;
    SB_LUT4 i6437_2_lut_3_lut (.I0(n7612), .I1(wr_addr_r[3]), .I2(wr_addr_r[4]), 
            .I3(GND_net), .O(n7616));
    defparam i6437_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF i341_342 (.Q(\REG.mem_3_5 ), .C(DEBUG_6_c_c), .D(n4730));   // src/fifo_dc_32_lut_gen.v(878[78:81])
    SB_LUT4 n14240_bdd_4_lut (.I0(n14240), .I1(\REG.mem_1_13 ), .I2(\REG.mem_0_13 ), 
            .I3(rd_addr_r[1]), .O(n12042));
    defparam n14240_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i102_2_lut_3_lut_4_lut (.I0(n7612), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n49));
    defparam EnabledDecoder_2_i102_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 EnabledDecoder_2_i101_2_lut_3_lut_4_lut (.I0(n7612), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n17));
    defparam EnabledDecoder_2_i101_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 wr_addr_r_6__I_0_add_2_5_lut (.I0(GND_net), .I1(wr_addr_r[3]), 
            .I2(rp_sync_w[3]), .I3(n10627), .O(wr_sig_diff0_w[3])) /* synthesis syn_instantiated=1 */ ;
    defparam wr_addr_r_6__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3975_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_30_6 ), .O(n5177));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3975_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4011_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_32_9 ), .O(n5213));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4011_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 EnabledDecoder_2_i104_2_lut_3_lut_4_lut (.I0(n16_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n48));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i104_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 rd_addr_r_1__bdd_4_lut_11779 (.I0(rd_addr_r[1]), .I1(n11788), 
            .I2(n11789), .I3(rd_addr_r[2]), .O(n13526));
    defparam rd_addr_r_1__bdd_4_lut_11779.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_6__I_0_151_8_lut (.I0(GND_net), .I1(\rd_addr_r[6] ), 
            .I2(GND_net), .I3(n10642), .O(rd_addr_p1_w[6])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4010_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_32_8 ), .O(n5212));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4010_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n13526_bdd_4_lut (.I0(n13526), .I1(n11786), .I2(n11785), .I3(rd_addr_r[2]), 
            .O(n13529));
    defparam n13526_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_3__bdd_4_lut_12358 (.I0(rd_addr_r[3]), .I1(n11635), 
            .I2(n11636), .I3(rd_addr_r[4]), .O(n14228));
    defparam rd_addr_r_3__bdd_4_lut_12358.LUT_INIT = 16'he4aa;
    SB_LUT4 EnabledDecoder_2_i103_2_lut_3_lut_4_lut (.I0(n16_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n16));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i103_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 n14228_bdd_4_lut (.I0(n14228), .I1(n11630), .I2(n13271), .I3(rd_addr_r[4]), 
            .O(n14231));
    defparam n14228_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4009_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_32_7 ), .O(n5211));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4009_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 EnabledDecoder_2_i17_2_lut (.I0(n9), .I1(wr_addr_r[2]), .I2(GND_net), 
            .I3(GND_net), .O(n17_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i17_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 EnabledDecoder_2_i90_2_lut_3_lut (.I0(n25_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n55));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i90_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12343 (.I0(rd_addr_r[0]), .I1(\REG.mem_6_13 ), 
            .I2(\REG.mem_7_13 ), .I3(rd_addr_r[1]), .O(n14222));
    defparam rd_addr_r_0__bdd_4_lut_12343.LUT_INIT = 16'he4aa;
    SB_LUT4 n14222_bdd_4_lut (.I0(n14222), .I1(\REG.mem_5_13 ), .I2(\REG.mem_4_13 ), 
            .I3(rd_addr_r[1]), .O(n12051));
    defparam n14222_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11754 (.I0(rd_addr_r[0]), .I1(\REG.mem_42_6 ), 
            .I2(\REG.mem_43_6 ), .I3(rd_addr_r[1]), .O(n13520));
    defparam rd_addr_r_0__bdd_4_lut_11754.LUT_INIT = 16'he4aa;
    SB_LUT4 i4008_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_32_6 ), .O(n5210));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4008_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n13520_bdd_4_lut (.I0(n13520), .I1(\REG.mem_41_6 ), .I2(\REG.mem_40_6 ), 
            .I3(rd_addr_r[1]), .O(n11844));
    defparam n13520_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 EnabledDecoder_2_i89_2_lut_3_lut (.I0(n25_c), .I1(wr_addr_r[4]), 
            .I2(wr_addr_r[5]), .I3(GND_net), .O(n23));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i89_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11744 (.I0(rd_addr_r[0]), .I1(\REG.mem_18_5 ), 
            .I2(\REG.mem_19_5 ), .I3(rd_addr_r[1]), .O(n13514));
    defparam rd_addr_r_0__bdd_4_lut_11744.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12328 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_4 ), 
            .I2(\REG.mem_55_4 ), .I3(rd_addr_r[1]), .O(n14216));
    defparam rd_addr_r_0__bdd_4_lut_12328.LUT_INIT = 16'he4aa;
    SB_LUT4 n13514_bdd_4_lut (.I0(n13514), .I1(\REG.mem_17_5 ), .I2(\REG.mem_16_5 ), 
            .I3(rd_addr_r[1]), .O(n13517));
    defparam n13514_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_6__I_0_151_7_lut (.I0(GND_net), .I1(rd_addr_r[5]), 
            .I2(GND_net), .I3(n10641), .O(rd_addr_p1_w[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rd_addr_r_6__I_0_151_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n14216_bdd_4_lut (.I0(n14216), .I1(\REG.mem_53_4 ), .I2(\REG.mem_52_4 ), 
            .I3(rd_addr_r[1]), .O(n12054));
    defparam n14216_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11739 (.I0(rd_addr_r[0]), .I1(\REG.mem_54_13 ), 
            .I2(\REG.mem_55_13 ), .I3(rd_addr_r[1]), .O(n13508));
    defparam rd_addr_r_0__bdd_4_lut_11739.LUT_INIT = 16'he4aa;
    SB_LUT4 n13508_bdd_4_lut (.I0(n13508), .I1(\REG.mem_53_13 ), .I2(\REG.mem_52_13 ), 
            .I3(rd_addr_r[1]), .O(n12276));
    defparam n13508_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4400_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_54_15 ), .O(n5602));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4400_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4399_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_54_14 ), .O(n5601));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4399_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4007_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_32_5 ), .O(n5209));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4007_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11734 (.I0(rd_addr_r[0]), .I1(\REG.mem_22_0 ), 
            .I2(\REG.mem_23_0 ), .I3(rd_addr_r[1]), .O(n13502));
    defparam rd_addr_r_0__bdd_4_lut_11734.LUT_INIT = 16'he4aa;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12323 (.I0(rd_addr_r[0]), .I1(\REG.mem_38_2 ), 
            .I2(\REG.mem_39_2 ), .I3(rd_addr_r[1]), .O(n14210));
    defparam rd_addr_r_0__bdd_4_lut_12323.LUT_INIT = 16'he4aa;
    SB_LUT4 n13502_bdd_4_lut (.I0(n13502), .I1(\REG.mem_21_0 ), .I2(\REG.mem_20_0 ), 
            .I3(rd_addr_r[1]), .O(n13505));
    defparam n13502_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY rd_addr_r_6__I_0_151_7 (.CI(n10641), .I0(rd_addr_r[5]), .I1(GND_net), 
            .CO(n10642));
    SB_LUT4 n14210_bdd_4_lut (.I0(n14210), .I1(\REG.mem_37_2 ), .I2(\REG.mem_36_2 ), 
            .I3(rd_addr_r[1]), .O(n12057));
    defparam n14210_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4006_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_32_4 ), .O(n5208));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4006_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4398_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_54_13 ), .O(n5600));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4398_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4005_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_32_3 ), .O(n5207));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4005_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4397_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_54_12 ), .O(n5599));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4397_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4396_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_54_11 ), .O(n5598));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4396_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12318 (.I0(rd_addr_r[0]), .I1(\REG.mem_50_11 ), 
            .I2(\REG.mem_51_11 ), .I3(rd_addr_r[1]), .O(n14204));
    defparam rd_addr_r_0__bdd_4_lut_12318.LUT_INIT = 16'he4aa;
    SB_LUT4 i10182_3_lut (.I0(\REG.mem_38_3 ), .I1(\REG.mem_39_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11831));
    defparam i10182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4004_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_32_2 ), .O(n5206));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4004_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n14204_bdd_4_lut (.I0(n14204), .I1(\REG.mem_49_11 ), .I2(\REG.mem_48_11 ), 
            .I3(rd_addr_r[1]), .O(n14207));
    defparam n14204_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3974_3_lut_4_lut (.I0(n65), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_30_5 ), .O(n5176));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i3974_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10181_3_lut (.I0(\REG.mem_36_3 ), .I1(\REG.mem_37_3 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11830));
    defparam i10181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4395_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_54_10 ), .O(n5597));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4395_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10106_3_lut (.I0(\REG.mem_20_4 ), .I1(\REG.mem_21_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11755));
    defparam i10106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10107_3_lut (.I0(\REG.mem_22_4 ), .I1(\REG.mem_23_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11756));
    defparam i10107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10014_3_lut (.I0(\REG.mem_18_4 ), .I1(\REG.mem_19_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11663));
    defparam i10014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10013_3_lut (.I0(\REG.mem_16_4 ), .I1(\REG.mem_17_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11662));
    defparam i10013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4394_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[9] ), 
            .I3(\REG.mem_54_9 ), .O(n5596));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4394_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4393_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[8] ), 
            .I3(\REG.mem_54_8 ), .O(n5595));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4393_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4392_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[7] ), 
            .I3(\REG.mem_54_7 ), .O(n5594));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4392_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10871_3_lut (.I0(\REG.mem_4_4 ), .I1(\REG.mem_5_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12520));
    defparam i10871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10872_3_lut (.I0(\REG.mem_6_4 ), .I1(\REG.mem_7_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12521));
    defparam i10872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10866_3_lut (.I0(\REG.mem_2_4 ), .I1(\REG.mem_3_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12515));
    defparam i10866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10865_3_lut (.I0(\REG.mem_0_4 ), .I1(\REG.mem_1_4 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12514));
    defparam i10865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4391_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[6] ), 
            .I3(\REG.mem_54_6 ), .O(n5593));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4391_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4390_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[5] ), 
            .I3(\REG.mem_54_5 ), .O(n5592));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4390_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4389_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[4] ), 
            .I3(\REG.mem_54_4 ), .O(n5591));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4389_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4003_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_32_1 ), .O(n5205));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4003_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4388_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[3] ), 
            .I3(\REG.mem_54_3 ), .O(n5590));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4388_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(wp_sync2_r[3]), .I1(wp_sync2_r[4]), 
            .I2(wp_sync2_r[6]), .I3(wp_sync2_r[5]), .O(wp_sync_w[3]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 EnabledDecoder_2_i49_2_lut_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n49_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i49_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i4387_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[2] ), 
            .I3(\REG.mem_54_2 ), .O(n5589));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4387_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4001_3_lut_4_lut (.I0(n7616), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_32_0 ), .O(n5203));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4001_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4051_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_34_15 ), .O(n5253));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4051_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4386_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[1] ), 
            .I3(\REG.mem_54_1 ), .O(n5588));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4386_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4385_3_lut_4_lut (.I0(n49_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[0] ), 
            .I3(\REG.mem_54_0 ), .O(n5587));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4385_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i40_2_lut_3_lut_4_lut (.I0(n12_adj_1156), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n40));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i40_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i9_2_lut_3_lut_4_lut (.I0(\afull_flag_impl.af_flag_p_w_N_603[3] ), 
            .I1(full_o), .I2(\wr_addr_r[0] ), .I3(wr_addr_r[1]), .O(n9));
    defparam EnabledDecoder_2_i9_2_lut_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 rd_fifo_en_w_I_0_158_2_lut_3_lut (.I0(DEBUG_5_c), .I1(get_next_word), 
            .I2(\genblk16.rd_prev_r ), .I3(GND_net), .O(t_rd_fifo_en_w));   // src/fifo_dc_32_lut_gen.v(747[41:67])
    defparam rd_fifo_en_w_I_0_158_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_LUT4 EnabledDecoder_2_i55_2_lut_3_lut_4_lut (.I0(n12_adj_1156), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n55_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i55_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i59_2_lut_3_lut_4_lut (.I0(n11), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n59_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i59_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i4050_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_34_14 ), .O(n5252));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4050_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4049_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_34_13 ), .O(n5251));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4049_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4048_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_34_12 ), .O(n5250));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4048_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 EnabledDecoder_2_i11_2_lut_3_lut_4_lut (.I0(\afull_flag_impl.af_flag_p_w_N_603[3] ), 
            .I1(full_o), .I2(\wr_addr_r[0] ), .I3(wr_addr_r[1]), .O(n11));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 EnabledDecoder_2_i12_2_lut_3_lut_4_lut (.I0(\afull_flag_impl.af_flag_p_w_N_603[3] ), 
            .I1(full_o), .I2(\wr_addr_r[0] ), .I3(wr_addr_r[1]), .O(n12_adj_1156));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i12_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 EnabledDecoder_2_i44_2_lut_3_lut_4_lut (.I0(n11), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n44));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i44_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i82_2_lut_3_lut_4_lut (.I0(n17_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n59));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i82_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 EnabledDecoder_2_i63_2_lut_3_lut_4_lut (.I0(n12_adj_1156), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n63));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i63_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10727_3_lut (.I0(n13283), .I1(n13067), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12376));
    defparam i10727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10728_3_lut (.I0(n12851), .I1(n14363), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12377));
    defparam i10728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10697_3_lut (.I0(n14123), .I1(n13889), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12346));
    defparam i10697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i81_2_lut_3_lut_4_lut (.I0(n17_c), .I1(wr_addr_r[3]), 
            .I2(wr_addr_r[5]), .I3(wr_addr_r[4]), .O(n27));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i81_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut (.I0(wp_sync2_r[4]), .I1(wp_sync2_r[6]), .I2(wp_sync2_r[5]), 
            .I3(GND_net), .O(wp_sync_w[4]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i10694_3_lut (.I0(\REG.mem_4_9 ), .I1(\REG.mem_5_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12343));
    defparam i10694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10695_3_lut (.I0(\REG.mem_6_9 ), .I1(\REG.mem_7_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12344));
    defparam i10695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10692_3_lut (.I0(\REG.mem_2_9 ), .I1(\REG.mem_3_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12341));
    defparam i10692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10691_3_lut (.I0(\REG.mem_0_9 ), .I1(\REG.mem_1_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12340));
    defparam i10691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_53 (.I0(wp_sync2_r[2]), .I1(wp_sync2_r[3]), 
            .I2(wp_sync_w[4]), .I3(GND_net), .O(wp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_53.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_54 (.I0(wp_sync2_r[1]), .I1(wp_sync2_r[2]), 
            .I2(wp_sync_w[3]), .I3(GND_net), .O(wp_sync_w[1]));   // src/fifo_dc_32_lut_gen.v(539[38:77])
    defparam i1_2_lut_3_lut_adj_54.LUT_INIT = 16'h9696;
    SB_LUT4 i10418_3_lut (.I0(n13589), .I1(n13505), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12067));
    defparam i10418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10419_3_lut (.I0(n13403), .I1(n13151), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12068));
    defparam i10419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10389_3_lut (.I0(n13859), .I1(n13835), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12038));
    defparam i10389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10421_3_lut (.I0(n12833), .I1(n12791), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12070));
    defparam i10421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10422_3_lut (.I0(n12779), .I1(n14387), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12071));
    defparam i10422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10410_3_lut (.I0(n12923), .I1(n12899), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12059));
    defparam i10410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10409_3_lut (.I0(n13043), .I1(n12929), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12058));
    defparam i10409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10733_3_lut (.I0(\REG.mem_20_9 ), .I1(\REG.mem_21_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12382));
    defparam i10733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10734_3_lut (.I0(\REG.mem_22_9 ), .I1(\REG.mem_23_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12383));
    defparam i10734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10713_3_lut (.I0(\REG.mem_18_9 ), .I1(\REG.mem_19_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12362));
    defparam i10713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10712_3_lut (.I0(\REG.mem_16_9 ), .I1(\REG.mem_17_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12361));
    defparam i10712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i65_2_lut_3_lut_4_lut (.I0(n9), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n65));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i65_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10334_3_lut (.I0(\REG.mem_52_0 ), .I1(\REG.mem_53_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11983));
    defparam i10334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10335_3_lut (.I0(\REG.mem_54_0 ), .I1(\REG.mem_55_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11984));
    defparam i10335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10323_3_lut (.I0(\REG.mem_50_0 ), .I1(\REG.mem_51_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11972));
    defparam i10323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10322_3_lut (.I0(\REG.mem_48_0 ), .I1(\REG.mem_49_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11971));
    defparam i10322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10382_3_lut (.I0(\REG.mem_52_15 ), .I1(\REG.mem_53_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12031));
    defparam i10382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10383_3_lut (.I0(\REG.mem_54_15 ), .I1(\REG.mem_55_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12032));
    defparam i10383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10371_3_lut (.I0(\REG.mem_50_15 ), .I1(\REG.mem_51_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12020));
    defparam i10371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10370_3_lut (.I0(\REG.mem_48_15 ), .I1(\REG.mem_49_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12019));
    defparam i10370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10346_3_lut (.I0(\REG.mem_36_15 ), .I1(\REG.mem_37_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11995));
    defparam i10346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10347_3_lut (.I0(\REG.mem_38_15 ), .I1(\REG.mem_39_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11996));
    defparam i10347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10338_3_lut (.I0(\REG.mem_34_15 ), .I1(\REG.mem_35_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11987));
    defparam i10338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10337_3_lut (.I0(\REG.mem_32_15 ), .I1(\REG.mem_33_15 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11986));
    defparam i10337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4047_3_lut_4_lut (.I0(n42_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_34_11 ), .O(n5249));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4047_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9752_4_lut_4_lut (.I0(wr_addr_r[3]), .I1(wr_addr_r[4]), .I2(rp_sync2_r[3]), 
            .I3(rp_sync_w[4]), .O(n11400));
    defparam i9752_4_lut_4_lut.LUT_INIT = 16'hdeb7;
    SB_LUT4 i1_2_lut_3_lut_adj_55 (.I0(rp_sync2_r[0]), .I1(rp_sync2_r[1]), 
            .I2(rp_sync_w[2]), .I3(GND_net), .O(rp_sync_w[0]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_3_lut_adj_55.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_56 (.I0(rp_sync2_r[2]), .I1(rp_sync2_r[3]), 
            .I2(rp_sync_w[4]), .I3(GND_net), .O(rp_sync_w[2]));   // src/fifo_dc_32_lut_gen.v(288[38:77])
    defparam i1_2_lut_3_lut_adj_56.LUT_INIT = 16'h9696;
    SB_LUT4 i9923_3_lut (.I0(n12977), .I1(n12869), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11572));
    defparam i9923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9924_3_lut (.I0(n12839), .I1(n14273), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11573));
    defparam i9924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9894_3_lut (.I0(n13109), .I1(n13049), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11543));
    defparam i9894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10354_3_lut (.I0(n13529), .I1(n12002), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n12003));
    defparam i10354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10353_3_lut (.I0(n13781), .I1(n13775), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n12002));
    defparam i10353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10817_3_lut (.I0(\REG.mem_60_9 ), .I1(\REG.mem_61_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12466));
    defparam i10817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10818_3_lut (.I0(\REG.mem_62_9 ), .I1(\REG.mem_63_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12467));
    defparam i10818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10815_3_lut (.I0(\REG.mem_58_9 ), .I1(\REG.mem_59_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12464));
    defparam i10815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10814_3_lut (.I0(\REG.mem_56_9 ), .I1(\REG.mem_57_9 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12463));
    defparam i10814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10342_3_lut (.I0(n13493), .I1(n11990), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n11991));
    defparam i10342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10341_3_lut (.I0(n13457), .I1(n13337), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11990));
    defparam i10341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10327_3_lut (.I0(n13487), .I1(n11975), .I2(rd_addr_r[3]), 
            .I3(GND_net), .O(n11976));
    defparam i10327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10326_3_lut (.I0(n14099), .I1(n14003), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11975));
    defparam i10326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4378_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[15] ), 
            .I3(\REG.mem_53_15 ), .O(n5580));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4378_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4377_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[14] ), 
            .I3(\REG.mem_53_14 ), .O(n5579));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4377_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4376_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[13] ), 
            .I3(\REG.mem_53_13 ), .O(n5578));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4376_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4375_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[12] ), 
            .I3(\REG.mem_53_12 ), .O(n5577));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4375_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4374_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[11] ), 
            .I3(\REG.mem_53_11 ), .O(n5576));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4374_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4373_3_lut_4_lut (.I0(n47_c), .I1(wr_addr_r[5]), .I2(\dc32_fifo_data_in[10] ), 
            .I3(\REG.mem_53_10 ), .O(n5575));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam i4373_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i9852_3_lut (.I0(n12857), .I1(n12803), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11501));
    defparam i9852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9851_3_lut (.I0(n12959), .I1(n12935), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11500));
    defparam i9851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10112_3_lut (.I0(\REG.mem_4_0 ), .I1(\REG.mem_5_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11761));
    defparam i10112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10113_3_lut (.I0(\REG.mem_6_0 ), .I1(\REG.mem_7_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11762));
    defparam i10113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10376_3_lut (.I0(\REG.mem_28_5 ), .I1(\REG.mem_29_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12025));
    defparam i10376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10377_3_lut (.I0(\REG.mem_30_5 ), .I1(\REG.mem_31_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12026));
    defparam i10377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10083_3_lut (.I0(\REG.mem_2_0 ), .I1(\REG.mem_3_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11732));
    defparam i10083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10082_3_lut (.I0(\REG.mem_0_0 ), .I1(\REG.mem_1_0 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11731));
    defparam i10082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10332_3_lut (.I0(\REG.mem_26_5 ), .I1(\REG.mem_27_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11981));
    defparam i10332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10331_3_lut (.I0(\REG.mem_24_5 ), .I1(\REG.mem_25_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11980));
    defparam i10331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9857_3_lut (.I0(\REG.mem_4_5 ), .I1(\REG.mem_5_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11506));
    defparam i9857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9858_3_lut (.I0(\REG.mem_6_5 ), .I1(\REG.mem_7_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11507));
    defparam i9858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10860_3_lut (.I0(\REG.mem_2_5 ), .I1(\REG.mem_3_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12509));
    defparam i10860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10859_3_lut (.I0(\REG.mem_0_5 ), .I1(\REG.mem_1_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12508));
    defparam i10859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_57 (.I0(\afull_flag_impl.af_flag_p_w_N_603[3] ), 
            .I1(wr_sig_diff0_w[3]), .I2(n6_adj_1172), .I3(wr_sig_diff0_w[0]), 
            .O(n3_adj_1166));   // src/fifo_dc_32_lut_gen.v(403[38:87])
    defparam i1_4_lut_adj_57.LUT_INIT = 16'heccc;
    SB_LUT4 i2_2_lut (.I0(wr_sig_diff0_w[2]), .I1(wr_sig_diff0_w[1]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_1172));   // src/fifo_dc_32_lut_gen.v(403[38:87])
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10440_3_lut (.I0(\REG.mem_34_5 ), .I1(\REG.mem_35_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12089));
    defparam i10440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10439_3_lut (.I0(\REG.mem_32_5 ), .I1(\REG.mem_33_5 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12088));
    defparam i10439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9906_3_lut (.I0(n13343), .I1(n12989), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11555));
    defparam i9906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9840_3_lut (.I0(n13745), .I1(n13577), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11489));
    defparam i9840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10844_3_lut (.I0(\REG.mem_44_12 ), .I1(\REG.mem_45_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12493));
    defparam i10844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10845_3_lut (.I0(\REG.mem_46_12 ), .I1(\REG.mem_47_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12494));
    defparam i10845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10839_3_lut (.I0(\REG.mem_42_12 ), .I1(\REG.mem_43_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12488));
    defparam i10839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10838_3_lut (.I0(\REG.mem_40_12 ), .I1(\REG.mem_41_12 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n12487));
    defparam i10838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 EnabledDecoder_2_i47_2_lut_3_lut_4_lut (.I0(n12_adj_1156), .I1(wr_addr_r[2]), 
            .I2(wr_addr_r[3]), .I3(wr_addr_r[4]), .O(n47_c));   // src/fifo_dc_32_lut_gen.v(889[37:55])
    defparam EnabledDecoder_2_i47_2_lut_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i10139_3_lut (.I0(\REG.mem_4_6 ), .I1(\REG.mem_5_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11788));
    defparam i10139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10140_3_lut (.I0(\REG.mem_6_6 ), .I1(\REG.mem_7_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11789));
    defparam i10140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10137_3_lut (.I0(\REG.mem_2_6 ), .I1(\REG.mem_3_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11786));
    defparam i10137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10136_3_lut (.I0(\REG.mem_0_6 ), .I1(\REG.mem_1_6 ), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(n11785));
    defparam i10136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9986_3_lut (.I0(n13025), .I1(n12965), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11635));
    defparam i9986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9987_3_lut (.I0(n12917), .I1(n12845), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11636));
    defparam i9987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9981_3_lut (.I0(n13397), .I1(n13145), .I2(rd_addr_r[2]), 
            .I3(GND_net), .O(n11630));
    defparam i9981_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=20) 
//

module \uart_rx(CLKS_PER_BIT=20)  (SLM_CLK_c, r_Rx_Data, UART_RX_c, GND_net, 
            n4, n4_adj_1, n7455, n4_adj_2, n10847, debug_led3, n5869, 
            pc_data_rx, VCC_net, n5844, n5843, n5842, n5841, n5840, 
            n5839, n5838, n3997, n4002) /* synthesis syn_module_defined=1 */ ;
    input SLM_CLK_c;
    output r_Rx_Data;
    input UART_RX_c;
    input GND_net;
    output n4;
    output n4_adj_1;
    output n7455;
    output n4_adj_2;
    output n10847;
    output debug_led3;
    input n5869;
    output [7:0]pc_data_rx;
    input VCC_net;
    input n5844;
    input n5843;
    input n5842;
    input n5841;
    input n5840;
    input n5839;
    input n5838;
    output n3997;
    output n4002;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n3;
    wire [2:0]r_SM_Main;   // src/uart_rx.v(36[17:26])
    
    wire r_Rx_Data_R;
    wire [9:0]n45;
    
    wire n6490;
    wire [9:0]r_Clock_Count;   // src/uart_rx.v(32[17:30])
    
    wire n6481, n151, n5837;
    wire [2:0]r_Bit_Index;   // src/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main_2__N_732;
    
    wire n4140, n10927, n4081, n10901, n3_adj_1143, n55_adj_1144, 
        n145, n13, n125;
    wire [2:0]n340;
    
    wire n4470, n149, n8, n140, n6, n4_adj_1145, n6515, n6500, 
        n10711, n10710, n10709, n10708, n10707, n10706, n10705, 
        n10704, n10703;
    
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n3), .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(SLM_CLK_c), .D(r_Rx_Data_R));   // src/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Clock_Count_1111__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n6490), .D(n45[0]), .R(n6481));   // src/uart_rx.v(120[34:51])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(SLM_CLK_c), .D(UART_RX_c));   // src/uart_rx.v(41[10] 45[8])
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(n151), .I2(GND_net), .I3(GND_net), 
            .O(n5837));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_140_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // src/uart_rx.v(97[17:39])
    defparam equal_140_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_137_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // src/uart_rx.v(97[17:39])
    defparam equal_137_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i6277_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n7455));
    defparam i6277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main_2__N_732[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main[2]), .O(n4140));
    defparam i2_4_lut.LUT_INIT = 16'h0023;
    SB_LUT4 i12_3_lut (.I0(n4140), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n10927));   // src/uart_rx.v(36[17:26])
    defparam i12_3_lut.LUT_INIT = 16'h6464;
    SB_LUT4 equal_142_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // src/uart_rx.v(97[17:39])
    defparam equal_142_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[0]), .I1(n151), .I2(n4_adj_2), .I3(r_Bit_Index[0]), 
            .O(n10847));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_732[2]), 
            .I3(r_SM_Main[0]), .O(n4081));
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n4081), 
            .I3(debug_led3), .O(n10901));
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_DFF r_Rx_Byte_i0 (.Q(pc_data_rx[0]), .C(SLM_CLK_c), .D(n5869));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Rx_DV_52 (.Q(debug_led3), .C(SLM_CLK_c), .E(VCC_net), .D(n10901));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n10927));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(pc_data_rx[7]), .C(SLM_CLK_c), .D(n5844));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(pc_data_rx[6]), .C(SLM_CLK_c), .D(n5843));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(pc_data_rx[5]), .C(SLM_CLK_c), .D(n5842));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(pc_data_rx[4]), .C(SLM_CLK_c), .D(n5841));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(pc_data_rx[3]), .C(SLM_CLK_c), .D(n5840));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(pc_data_rx[2]), .C(SLM_CLK_c), .D(n5839));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(pc_data_rx[1]), .C(SLM_CLK_c), .D(n5838));   // src/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(n5837));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_2_lut_3_lut (.I0(r_SM_Main[0]), .I1(n151), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n3997));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_38 (.I0(r_SM_Main[0]), .I1(n151), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n4002));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_adj_38.LUT_INIT = 16'hbfbf;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n3_adj_1143), 
            .R(r_SM_Main[2]));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1111__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n6490), .D(n45[9]), .R(n6481));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1111__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n6490), .D(n45[8]), .R(n6481));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1111__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n6490), .D(n45[7]), .R(n6481));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1111__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n6490), .D(n45[6]), .R(n6481));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1111__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n6490), .D(n45[5]), .R(n6481));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1111__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n6490), .D(n45[4]), .R(n6481));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1111__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n6490), .D(n45[3]), .R(n6481));   // src/uart_rx.v(120[34:51])
    SB_LUT4 i1_2_lut_adj_39 (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_732[2]), 
            .I2(GND_net), .I3(GND_net), .O(n55_adj_1144));
    defparam i1_2_lut_adj_39.LUT_INIT = 16'h8888;
    SB_LUT4 i5323_4_lut (.I0(r_Rx_Data), .I1(n55_adj_1144), .I2(r_SM_Main[1]), 
            .I3(n145), .O(n3_adj_1143));   // src/uart_rx.v(36[17:26])
    defparam i5323_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main[0]), .I2(n13), .I3(GND_net), 
            .O(n125));   // src/uart_rx.v(30[17:26])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i11078_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[2]), .I2(n145), 
            .I3(r_SM_Main[1]), .O(n6490));
    defparam i11078_4_lut.LUT_INIT = 16'h3313;
    SB_DFFESR r_Clock_Count_1111__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n6490), .D(n45[2]), .R(n6481));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1111__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n6490), .D(n45[1]), .R(n6481));   // src/uart_rx.v(120[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(SLM_CLK_c), .E(n4140), 
            .D(n340[1]), .R(n4470));   // src/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(SLM_CLK_c), .E(n4140), 
            .D(n340[2]), .R(n4470));   // src/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1235_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n340[2]));   // src/uart_rx.v(49[10] 144[8])
    defparam i1235_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n149));   // src/uart_rx.v(49[10] 144[8])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i5281_4_lut_4_lut (.I0(r_SM_Main_2__N_732[2]), .I1(r_SM_Main[2]), 
            .I2(n125), .I3(r_SM_Main[1]), .O(n6481));   // src/uart_rx.v(49[10] 144[8])
    defparam i5281_4_lut_4_lut.LUT_INIT = 16'h2203;
    SB_LUT4 i1_2_lut_3_lut_adj_40 (.I0(r_SM_Main_2__N_732[2]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n151));   // src/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_adj_40.LUT_INIT = 16'h2020;
    SB_LUT4 i3_4_lut_adj_41 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), 
            .I2(r_Clock_Count[3]), .I3(r_Clock_Count[4]), .O(n8));
    defparam i3_4_lut_adj_41.LUT_INIT = 16'hffdf;
    SB_LUT4 i4_3_lut (.I0(n140), .I1(n8), .I2(r_Clock_Count[2]), .I3(GND_net), 
            .O(n13));
    defparam i4_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_42 (.I0(r_SM_Main[0]), .I1(n13), .I2(GND_net), 
            .I3(GND_net), .O(n145));   // src/uart_rx.v(36[17:26])
    defparam i1_2_lut_adj_42.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_43 (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // src/uart_rx.v(32[17:30])
    defparam i1_2_lut_adj_43.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[9]), 
            .I3(n6), .O(n140));   // src/uart_rx.v(32[17:30])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_44 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), 
            .I2(r_Clock_Count[1]), .I3(GND_net), .O(n4_adj_1145));   // src/uart_rx.v(118[17:47])
    defparam i1_3_lut_adj_44.LUT_INIT = 16'hecec;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[4]), .I1(n140), .I2(r_Clock_Count[3]), 
            .I3(n4_adj_1145), .O(r_SM_Main_2__N_732[2]));   // src/uart_rx.v(32[17:30])
    defparam i1_4_lut.LUT_INIT = 16'heeec;
    SB_LUT4 i5315_3_lut (.I0(n149), .I1(r_SM_Main[0]), .I2(r_SM_Main_2__N_732[2]), 
            .I3(GND_net), .O(n6515));   // src/uart_rx.v(36[17:26])
    defparam i5315_3_lut.LUT_INIT = 16'h2c2c;
    SB_LUT4 i5316_3_lut (.I0(n6500), .I1(n6515), .I2(r_SM_Main[1]), .I3(GND_net), 
            .O(n3));   // src/uart_rx.v(36[17:26])
    defparam i5316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_1111_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n10711), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1111_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1111_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n10710), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1111_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1111_add_4_10 (.CI(n10710), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n10711));
    SB_LUT4 r_Clock_Count_1111_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n10709), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1111_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1111_add_4_9 (.CI(n10709), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n10710));
    SB_LUT4 r_Clock_Count_1111_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n10708), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1111_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1111_add_4_8 (.CI(n10708), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n10709));
    SB_LUT4 r_Clock_Count_1111_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n10707), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1111_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1111_add_4_7 (.CI(n10707), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n10708));
    SB_LUT4 r_Clock_Count_1111_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n10706), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1111_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1111_add_4_6 (.CI(n10706), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n10707));
    SB_LUT4 r_Clock_Count_1111_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n10705), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1111_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1111_add_4_5 (.CI(n10705), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n10706));
    SB_LUT4 r_Clock_Count_1111_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n10704), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1111_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1111_add_4_4 (.CI(n10704), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n10705));
    SB_LUT4 r_Clock_Count_1111_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n10703), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1111_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1111_add_4_3 (.CI(n10703), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n10704));
    SB_LUT4 r_Clock_Count_1111_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1111_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1111_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n10703));
    SB_LUT4 i5300_4_lut_3_lut (.I0(r_SM_Main[0]), .I1(n13), .I2(r_Rx_Data), 
            .I3(GND_net), .O(n6500));   // src/uart_rx.v(30[17:26])
    defparam i5300_4_lut_3_lut.LUT_INIT = 16'h8d8d;
    SB_LUT4 i1228_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n340[1]));   // src/uart_rx.v(102[36:51])
    defparam i1228_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3268_3_lut (.I0(n4140), .I1(r_SM_Main[1]), .I2(n149), .I3(GND_net), 
            .O(n4470));   // src/uart_rx.v(49[10] 144[8])
    defparam i3268_3_lut.LUT_INIT = 16'ha2a2;
    
endmodule
//
// Verilog Description of module clock
//

module clock (GND_net, VCC_net, ICE_SYSCLK_c, pll_clk_unbuf) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    input ICE_SYSCLK_c;
    output pll_clk_unbuf;
    
    
    SB_PLL40_CORE pll_config (.REFERENCECLK(ICE_SYSCLK_c), .PLLOUTGLOBAL(pll_clk_unbuf), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=14, LSE_LCOL=7, LSE_RCOL=3, LSE_LLINE=222, LSE_RLINE=228 */ ;   // src/top.v(222[7] 228[3])
    defparam pll_config.FEEDBACK_PATH = "SIMPLE";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll_config.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll_config.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll_config.FDA_FEEDBACK = 0;
    defparam pll_config.FDA_RELATIVE = 0;
    defparam pll_config.PLLOUT_SELECT = "GENCLK";
    defparam pll_config.DIVR = 4'b0001;
    defparam pll_config.DIVF = 7'b1010010;
    defparam pll_config.DIVQ = 3'b100;
    defparam pll_config.FILTER_RANGE = 3'b001;
    defparam pll_config.ENABLE_ICEGATE = 1'b0;
    defparam pll_config.TEST_MODE = 1'b0;
    defparam pll_config.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module spi
//

module spi (\tx_data_byte[1] , \tx_shift_reg[0] , n1928, GND_net, \tx_data_byte[2] , 
            \tx_data_byte[3] , VCC_net, SEN_c_1, SLM_CLK_c, SOUT_c, 
            n4093, \rx_shift_reg[0] , \tx_data_byte[4] , \tx_data_byte[5] , 
            \tx_data_byte[6] , \tx_data_byte[7] , tx_addr_byte, n4070, 
            SDAT_c_15, multi_byte_spi_trans_flag_r, n11007, n5756, \rx_shift_reg[1] , 
            n5755, \rx_shift_reg[2] , n5754, \rx_shift_reg[3] , n5753, 
            \rx_shift_reg[4] , n5752, \rx_shift_reg[5] , n5751, \rx_shift_reg[6] , 
            n5750, \rx_shift_reg[7] , n5733, rx_buf_byte, n5732, n5731, 
            n5730, n5729, n5728, n5727, spi_rx_byte_ready, SCK_c_0, 
            spi_start_transfer_r, n4637, n3204) /* synthesis syn_module_defined=1 */ ;
    input \tx_data_byte[1] ;
    output \tx_shift_reg[0] ;
    output n1928;
    input GND_net;
    input \tx_data_byte[2] ;
    input \tx_data_byte[3] ;
    input VCC_net;
    output SEN_c_1;
    input SLM_CLK_c;
    input SOUT_c;
    output n4093;
    output \rx_shift_reg[0] ;
    input \tx_data_byte[4] ;
    input \tx_data_byte[5] ;
    input \tx_data_byte[6] ;
    input \tx_data_byte[7] ;
    input [7:0]tx_addr_byte;
    output n4070;
    output SDAT_c_15;
    input multi_byte_spi_trans_flag_r;
    input n11007;
    input n5756;
    output \rx_shift_reg[1] ;
    input n5755;
    output \rx_shift_reg[2] ;
    input n5754;
    output \rx_shift_reg[3] ;
    input n5753;
    output \rx_shift_reg[4] ;
    input n5752;
    output \rx_shift_reg[5] ;
    input n5751;
    output \rx_shift_reg[6] ;
    input n5750;
    output \rx_shift_reg[7] ;
    input n5733;
    output [7:0]rx_buf_byte;
    input n5732;
    input n5731;
    input n5730;
    input n5729;
    input n5728;
    input n5727;
    output spi_rx_byte_ready;
    output SCK_c_0;
    input spi_start_transfer_r;
    input n4637;
    output n3204;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [15:0]n1929;
    wire [15:0]tx_shift_reg;   // src/spi.v(70[12:24])
    
    wire n10698;
    wire [9:0]counter;   // src/spi.v(69[11:18])
    
    wire n10699;
    wire [9:0]n45;
    
    wire n10697;
    wire [2:0]n860;
    wire [3:0]state_3__N_905;
    
    wire n14414;
    wire [3:0]state;   // src/spi.v(71[11:16])
    
    wire n8, n12566, n12567, n4120, n10082, n10696, n10695, n10694, 
        n10090, n12605;
    wire [7:0]n315;
    wire [7:0]multi_byte_counter;   // src/spi.v(68[11:29])
    wire [7:0]n1985;
    
    wire n10659, n10658, n10657, n10656, n10655, n10654, n10653, 
        n11350, n11351, n11317, n2, n24, n16, n19, n11398, n10076, 
        n10081, n81, n12702, n12607, n19_adj_1139, n11345, n11346, 
        n11311, n4260, n2768, n4105, n6, n3, n4409, n3909, n14, 
        n9, n10, n14_adj_1140, n88, n10106, n14442, n12598, n4281, 
        n4455, n10702, n10701, n10700, n10119, n12586, n37, n21, 
        n12576, n3295, n11344, n12594;
    
    SB_LUT4 mux_946_i2_3_lut (.I0(\tx_data_byte[1] ), .I1(\tx_shift_reg[0] ), 
            .I2(n1928), .I3(GND_net), .O(n1929[1]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_946_i3_3_lut (.I0(\tx_data_byte[2] ), .I1(tx_shift_reg[1]), 
            .I2(n1928), .I3(GND_net), .O(n1929[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_946_i4_3_lut (.I0(\tx_data_byte[3] ), .I1(tx_shift_reg[2]), 
            .I2(n1928), .I3(GND_net), .O(n1929[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_1109_add_4_7 (.CI(n10698), .I0(VCC_net), .I1(counter[5]), 
            .CO(n10699));
    SB_LUT4 counter_1109_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[4]), 
            .I3(n10697), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1109_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF byte_recv_92_i2 (.Q(SEN_c_1), .C(SLM_CLK_c), .D(n860[1]));   // src/spi.v(88[9] 219[16])
    SB_DFFE rx_shift_reg_i0 (.Q(\rx_shift_reg[0] ), .C(SLM_CLK_c), .E(n4093), 
            .D(SOUT_c));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i0 (.Q(state[0]), .C(SLM_CLK_c), .E(n14414), .D(state_3__N_905[0]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 mux_946_i5_3_lut (.I0(\tx_data_byte[4] ), .I1(tx_shift_reg[3]), 
            .I2(n1928), .I3(GND_net), .O(n1929[4]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_946_i6_3_lut (.I0(\tx_data_byte[5] ), .I1(tx_shift_reg[4]), 
            .I2(n1928), .I3(GND_net), .O(n1929[5]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11041_4_lut (.I0(n8), .I1(state[1]), .I2(state[0]), .I3(state[2]), 
            .O(n12566));   // src/spi.v(88[9] 219[16])
    defparam i11041_4_lut.LUT_INIT = 16'hc08c;
    SB_LUT4 i1_4_lut (.I0(counter[4]), .I1(n12566), .I2(n12567), .I3(state[3]), 
            .O(n860[0]));   // src/spi.v(88[9] 219[16])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_CARRY counter_1109_add_4_6 (.CI(n10697), .I0(VCC_net), .I1(counter[4]), 
            .CO(n10698));
    SB_LUT4 mux_946_i7_3_lut (.I0(\tx_data_byte[6] ), .I1(tx_shift_reg[5]), 
            .I2(n1928), .I3(GND_net), .O(n1929[6]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR counter_1109__i0 (.Q(counter[0]), .C(SLM_CLK_c), .E(n4120), 
            .D(n45[0]), .R(n10082));   // src/spi.v(183[28:41])
    SB_LUT4 mux_946_i8_3_lut (.I0(\tx_data_byte[7] ), .I1(tx_shift_reg[6]), 
            .I2(n1928), .I3(GND_net), .O(n1929[7]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_946_i9_3_lut (.I0(tx_addr_byte[0]), .I1(tx_shift_reg[7]), 
            .I2(n1928), .I3(GND_net), .O(n1929[8]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_946_i10_3_lut (.I0(tx_addr_byte[1]), .I1(tx_shift_reg[8]), 
            .I2(n1928), .I3(GND_net), .O(n1929[9]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_946_i11_3_lut (.I0(tx_addr_byte[2]), .I1(tx_shift_reg[9]), 
            .I2(n1928), .I3(GND_net), .O(n1929[10]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_946_i12_3_lut (.I0(tx_addr_byte[3]), .I1(tx_shift_reg[10]), 
            .I2(n1928), .I3(GND_net), .O(n1929[11]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE tx_shift_reg_i0_i15 (.Q(SDAT_c_15), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[15]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 counter_1109_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[3]), 
            .I3(n10696), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1109_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1109_add_4_5 (.CI(n10696), .I0(VCC_net), .I1(counter[3]), 
            .CO(n10697));
    SB_LUT4 mux_946_i13_3_lut (.I0(tx_addr_byte[4]), .I1(tx_shift_reg[11]), 
            .I2(n1928), .I3(GND_net), .O(n1929[12]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_946_i14_3_lut (.I0(tx_addr_byte[5]), .I1(tx_shift_reg[12]), 
            .I2(n1928), .I3(GND_net), .O(n1929[13]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_946_i15_3_lut (.I0(tx_addr_byte[6]), .I1(tx_shift_reg[13]), 
            .I2(n1928), .I3(GND_net), .O(n1929[14]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_1109_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[2]), 
            .I3(n10695), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1109_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1109_add_4_4 (.CI(n10695), .I0(VCC_net), .I1(counter[2]), 
            .CO(n10696));
    SB_LUT4 counter_1109_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[1]), 
            .I3(n10694), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1109_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1109_add_4_3 (.CI(n10694), .I0(VCC_net), .I1(counter[1]), 
            .CO(n10695));
    SB_LUT4 i8576_4_lut_4_lut (.I0(state[3]), .I1(multi_byte_spi_trans_flag_r), 
            .I2(state[0]), .I3(state[2]), .O(n10090));   // src/spi.v(76[8] 221[4])
    defparam i8576_4_lut_4_lut.LUT_INIT = 16'ha0f4;
    SB_LUT4 i10988_3_lut_4_lut (.I0(state[3]), .I1(multi_byte_spi_trans_flag_r), 
            .I2(state[2]), .I3(state[0]), .O(n12605));   // src/spi.v(76[8] 221[4])
    defparam i10988_3_lut_4_lut.LUT_INIT = 16'h00f4;
    SB_DFFE tx_shift_reg_i0_i0 (.Q(\tx_shift_reg[0] ), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n11007));   // src/spi.v(76[8] 221[4])
    SB_LUT4 counter_1109_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1109_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1109_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n10694));
    SB_DFF rx_shift_reg_i1 (.Q(\rx_shift_reg[1] ), .C(SLM_CLK_c), .D(n5756));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i2 (.Q(\rx_shift_reg[2] ), .C(SLM_CLK_c), .D(n5755));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i3 (.Q(\rx_shift_reg[3] ), .C(SLM_CLK_c), .D(n5754));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i4 (.Q(\rx_shift_reg[4] ), .C(SLM_CLK_c), .D(n5753));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i5 (.Q(\rx_shift_reg[5] ), .C(SLM_CLK_c), .D(n5752));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i6 (.Q(\rx_shift_reg[6] ), .C(SLM_CLK_c), .D(n5751));   // src/spi.v(76[8] 221[4])
    SB_DFF rx_shift_reg_i7 (.Q(\rx_shift_reg[7] ), .C(SLM_CLK_c), .D(n5750));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i1 (.Q(rx_buf_byte[1]), .C(SLM_CLK_c), .D(n5733));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i2 (.Q(rx_buf_byte[2]), .C(SLM_CLK_c), .D(n5732));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i3 (.Q(rx_buf_byte[3]), .C(SLM_CLK_c), .D(n5731));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i4 (.Q(rx_buf_byte[4]), .C(SLM_CLK_c), .D(n5730));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i5 (.Q(rx_buf_byte[5]), .C(SLM_CLK_c), .D(n5729));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i6 (.Q(rx_buf_byte[6]), .C(SLM_CLK_c), .D(n5728));   // src/spi.v(76[8] 221[4])
    SB_DFF Rx_Recv_Byte_i7 (.Q(rx_buf_byte[7]), .C(SLM_CLK_c), .D(n5727));   // src/spi.v(76[8] 221[4])
    SB_LUT4 add_961_9_lut (.I0(GND_net), .I1(multi_byte_counter[7]), .I2(n1985[5]), 
            .I3(n10659), .O(n315[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_961_8_lut (.I0(GND_net), .I1(multi_byte_counter[6]), .I2(n1985[5]), 
            .I3(n10658), .O(n315[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_8 (.CI(n10658), .I0(multi_byte_counter[6]), .I1(n1985[5]), 
            .CO(n10659));
    SB_LUT4 add_961_7_lut (.I0(GND_net), .I1(multi_byte_counter[5]), .I2(n1985[5]), 
            .I3(n10657), .O(n315[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_7 (.CI(n10657), .I0(multi_byte_counter[5]), .I1(n1985[5]), 
            .CO(n10658));
    SB_LUT4 add_961_6_lut (.I0(GND_net), .I1(multi_byte_counter[4]), .I2(n1985[5]), 
            .I3(n10656), .O(n315[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_6 (.CI(n10656), .I0(multi_byte_counter[4]), .I1(n1985[5]), 
            .CO(n10657));
    SB_LUT4 add_961_5_lut (.I0(GND_net), .I1(multi_byte_counter[3]), .I2(n1985[5]), 
            .I3(n10655), .O(n315[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_5 (.CI(n10655), .I0(multi_byte_counter[3]), .I1(n1985[5]), 
            .CO(n10656));
    SB_LUT4 add_961_4_lut (.I0(GND_net), .I1(multi_byte_counter[2]), .I2(n1985[5]), 
            .I3(n10654), .O(n315[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_4 (.CI(n10654), .I0(multi_byte_counter[2]), .I1(n1985[5]), 
            .CO(n10655));
    SB_LUT4 add_961_3_lut (.I0(GND_net), .I1(multi_byte_counter[1]), .I2(n1985[5]), 
            .I3(n10653), .O(n315[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_961_3 (.CI(n10653), .I0(multi_byte_counter[1]), .I1(n1985[5]), 
            .CO(n10654));
    SB_LUT4 add_961_2_lut (.I0(GND_net), .I1(multi_byte_counter[0]), .I2(n1985[5]), 
            .I3(GND_net), .O(n315[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_961_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFE tx_shift_reg_i0_i14 (.Q(tx_shift_reg[14]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[14]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i13 (.Q(tx_shift_reg[13]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[13]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i12 (.Q(tx_shift_reg[12]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[12]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i11 (.Q(tx_shift_reg[11]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[11]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i10 (.Q(tx_shift_reg[10]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[10]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i9 (.Q(tx_shift_reg[9]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[9]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i8 (.Q(tx_shift_reg[8]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[8]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i7 (.Q(tx_shift_reg[7]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[7]));   // src/spi.v(76[8] 221[4])
    SB_DFF byte_recv_92_i3 (.Q(spi_rx_byte_ready), .C(SLM_CLK_c), .D(n860[2]));   // src/spi.v(88[9] 219[16])
    SB_DFFE tx_shift_reg_i0_i6 (.Q(tx_shift_reg[6]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[6]));   // src/spi.v(76[8] 221[4])
    SB_DFF byte_recv_92_i1 (.Q(SCK_c_0), .C(SLM_CLK_c), .D(n860[0]));   // src/spi.v(88[9] 219[16])
    SB_DFFE tx_shift_reg_i0_i5 (.Q(tx_shift_reg[5]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[5]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i4 (.Q(tx_shift_reg[4]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[4]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i3 (.Q(tx_shift_reg[3]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[3]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i2 (.Q(tx_shift_reg[2]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE tx_shift_reg_i0_i1 (.Q(tx_shift_reg[1]), .C(SLM_CLK_c), .E(n4070), 
            .D(n1929[1]));   // src/spi.v(76[8] 221[4])
    SB_CARRY add_961_2 (.CI(GND_net), .I0(multi_byte_counter[0]), .I1(n1985[5]), 
            .CO(n10653));
    SB_LUT4 i1_2_lut (.I0(state[3]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n11350));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_23 (.I0(counter[4]), .I1(n11351), .I2(n11317), 
            .I3(n2), .O(n1928));
    defparam i1_4_lut_adj_23.LUT_INIT = 16'h5040;
    SB_LUT4 i30_4_lut (.I0(spi_start_transfer_r), .I1(state[3]), .I2(state[1]), 
            .I3(state[0]), .O(n24));   // src/spi.v(88[9] 219[16])
    defparam i30_4_lut.LUT_INIT = 16'hcfc1;
    SB_LUT4 i1_4_lut_adj_24 (.I0(n11317), .I1(state[3]), .I2(counter[4]), 
            .I3(state[1]), .O(n16));   // src/spi.v(88[9] 219[16])
    defparam i1_4_lut_adj_24.LUT_INIT = 16'hf5c4;
    SB_LUT4 mux_946_i16_3_lut (.I0(tx_addr_byte[7]), .I1(tx_shift_reg[14]), 
            .I2(n1928), .I3(GND_net), .O(n1929[15]));   // src/spi.v(88[9] 219[16])
    defparam mux_946_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9750_3_lut (.I0(state[3]), .I1(state[2]), .I2(n19), .I3(GND_net), 
            .O(n11398));
    defparam i9750_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i8567_3_lut (.I0(n10076), .I1(n11398), .I2(state[0]), .I3(GND_net), 
            .O(n10081));   // src/spi.v(71[11:16])
    defparam i8567_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i8568_4_lut (.I0(n81), .I1(n10081), .I2(state[1]), .I3(state[0]), 
            .O(n10082));   // src/spi.v(71[11:16])
    defparam i8568_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i11053_2_lut (.I0(state[3]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n12702));   // src/spi.v(71[11:16])
    defparam i11053_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8614_4_lut (.I0(state[2]), .I1(n12607), .I2(state[1]), .I3(n12702), 
            .O(n4120));   // src/spi.v(71[11:16])
    defparam i8614_4_lut.LUT_INIT = 16'hc5c0;
    SB_DFFE state_i3 (.Q(state[3]), .C(SLM_CLK_c), .E(n19_adj_1139), .D(state_3__N_905[3]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i2 (.Q(state[2]), .C(SLM_CLK_c), .E(n11345), .D(state_3__N_905[2]));   // src/spi.v(76[8] 221[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(SLM_CLK_c), .E(n11346), .D(state_3__N_905[1]));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i1_2_lut_adj_25 (.I0(state[3]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n81));
    defparam i1_2_lut_adj_25.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut (.I0(state[3]), .I1(n19), .I2(state[1]), .I3(GND_net), 
            .O(n11311));
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i2_3_lut_adj_26 (.I0(n11311), .I1(state[0]), .I2(state[2]), 
            .I3(GND_net), .O(n4260));
    defparam i2_3_lut_adj_26.LUT_INIT = 16'hbfbf;
    SB_LUT4 i1584_2_lut (.I0(state[1]), .I1(state[2]), .I2(GND_net), .I3(GND_net), 
            .O(n2768));   // src/spi.v(88[9] 219[16])
    defparam i1584_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(n2768), .I1(state[3]), .I2(spi_start_transfer_r), 
            .I3(state[0]), .O(n4105));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(state[3]), .I1(n4105), .I2(n19), .I3(state[0]), 
            .O(n6));
    defparam i2_4_lut.LUT_INIT = 16'hcc4c;
    SB_LUT4 i3_4_lut (.I0(n2768), .I1(n6), .I2(n4260), .I3(state[3]), 
            .O(n14414));
    defparam i3_4_lut.LUT_INIT = 16'h40c0;
    SB_LUT4 i8618_4_lut (.I0(state[0]), .I1(n19), .I2(state[1]), .I3(multi_byte_spi_trans_flag_r), 
            .O(n3));   // src/spi.v(71[11:16])
    defparam i8618_4_lut.LUT_INIT = 16'h9095;
    SB_LUT4 i3238_3_lut (.I0(n3), .I1(state[0]), .I2(n81), .I3(GND_net), 
            .O(state_3__N_905[0]));   // src/spi.v(88[9] 219[16])
    defparam i3238_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i3_4_lut_adj_27 (.I0(counter[0]), .I1(counter[2]), .I2(counter[3]), 
            .I3(counter[1]), .O(n11317));
    defparam i3_4_lut_adj_27.LUT_INIT = 16'h8000;
    SB_LUT4 i11112_3_lut (.I0(counter[4]), .I1(n11317), .I2(n4409), .I3(GND_net), 
            .O(n4093));   // src/spi.v(88[9] 219[16])
    defparam i11112_3_lut.LUT_INIT = 16'h0808;
    SB_DFFESR counter_1109__i9 (.Q(counter[9]), .C(SLM_CLK_c), .E(n4120), 
            .D(n45[9]), .R(n10082));   // src/spi.v(183[28:41])
    SB_DFFESS counter_1109__i8 (.Q(counter[8]), .C(SLM_CLK_c), .E(n4120), 
            .D(n45[8]), .S(n10082));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1109__i7 (.Q(counter[7]), .C(SLM_CLK_c), .E(n4120), 
            .D(n45[7]), .R(n10082));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1109__i6 (.Q(counter[6]), .C(SLM_CLK_c), .E(n4120), 
            .D(n45[6]), .R(n10082));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1109__i5 (.Q(counter[5]), .C(SLM_CLK_c), .E(n4120), 
            .D(n45[5]), .R(n10082));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1109__i1 (.Q(counter[1]), .C(SLM_CLK_c), .E(n4120), 
            .D(n45[1]), .R(n10082));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1109__i2 (.Q(counter[2]), .C(SLM_CLK_c), .E(n4120), 
            .D(n45[2]), .R(n10082));   // src/spi.v(183[28:41])
    SB_DFFESR counter_1109__i3 (.Q(counter[3]), .C(SLM_CLK_c), .E(n4120), 
            .D(n45[3]), .R(n10082));   // src/spi.v(183[28:41])
    SB_DFF Rx_Recv_Byte_i0 (.Q(rx_buf_byte[0]), .C(SLM_CLK_c), .D(n4637));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i2_3_lut_adj_28 (.I0(counter[1]), .I1(counter[3]), .I2(counter[2]), 
            .I3(GND_net), .O(n3909));
    defparam i2_3_lut_adj_28.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(counter[5]), .I2(counter[8]), 
            .I3(counter[9]), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_29 (.I0(counter[4]), .I1(counter[7]), .I2(GND_net), 
            .I3(GND_net), .O(n9));
    defparam i1_2_lut_adj_29.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut (.I0(n9), .I1(n14), .I2(n3909), .I3(counter[0]), 
            .O(n19));
    defparam i7_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_2_lut (.I0(multi_byte_counter[2]), .I1(multi_byte_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // src/spi.v(208[21:52])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_30 (.I0(multi_byte_counter[3]), .I1(multi_byte_counter[1]), 
            .I2(multi_byte_counter[5]), .I3(multi_byte_counter[7]), .O(n14_adj_1140));   // src/spi.v(208[21:52])
    defparam i6_4_lut_adj_30.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_31 (.I0(multi_byte_counter[0]), .I1(n14_adj_1140), 
            .I2(n10), .I3(multi_byte_counter[6]), .O(n1985[5]));   // src/spi.v(208[21:52])
    defparam i7_4_lut_adj_31.LUT_INIT = 16'hfffd;
    SB_DFFESR counter_1109__i4 (.Q(counter[4]), .C(SLM_CLK_c), .E(n4120), 
            .D(n45[4]), .R(n10082));   // src/spi.v(183[28:41])
    SB_LUT4 i106_2_lut (.I0(state[2]), .I1(n19), .I2(GND_net), .I3(GND_net), 
            .O(n88));
    defparam i106_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i8592_4_lut (.I0(n1985[5]), .I1(n88), .I2(state[0]), .I3(state[3]), 
            .O(n10106));   // src/spi.v(71[11:16])
    defparam i8592_4_lut.LUT_INIT = 16'hf530;
    SB_LUT4 i1_rep_17_2_lut (.I0(state[3]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n14442));
    defparam i1_rep_17_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11039_3_lut (.I0(state[0]), .I1(state[2]), .I2(state[3]), 
            .I3(GND_net), .O(n12598));   // src/spi.v(71[11:16])
    defparam i11039_3_lut.LUT_INIT = 16'hcdcd;
    SB_LUT4 i1_4_lut_adj_32 (.I0(n12598), .I1(n14442), .I2(n10106), .I3(state[1]), 
            .O(n860[1]));
    defparam i1_4_lut_adj_32.LUT_INIT = 16'hfcee;
    SB_DFFESR multi_byte_counter_i0 (.Q(multi_byte_counter[0]), .C(SLM_CLK_c), 
            .E(n4281), .D(n315[0]), .R(n4455));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i1 (.Q(multi_byte_counter[1]), .C(SLM_CLK_c), 
            .E(n4281), .D(n315[1]), .R(n4455));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i2 (.Q(multi_byte_counter[2]), .C(SLM_CLK_c), 
            .E(n4281), .D(n315[2]), .R(n4455));   // src/spi.v(76[8] 221[4])
    SB_DFFESR multi_byte_counter_i3 (.Q(multi_byte_counter[3]), .C(SLM_CLK_c), 
            .E(n4281), .D(n315[3]), .R(n4455));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i11115_3_lut_4_lut (.I0(state[2]), .I1(state[0]), .I2(n24), 
            .I3(n16), .O(n4070));   // src/spi.v(88[9] 219[16])
    defparam i11115_3_lut_4_lut.LUT_INIT = 16'h000d;
    SB_DFFESR multi_byte_counter_i4 (.Q(multi_byte_counter[4]), .C(SLM_CLK_c), 
            .E(n4281), .D(n315[4]), .R(n4455));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i8562_4_lut_4_lut (.I0(state[2]), .I1(n1985[5]), .I2(n19), 
            .I3(state[3]), .O(n10076));   // src/spi.v(76[8] 221[4])
    defparam i8562_4_lut_4_lut.LUT_INIT = 16'h44af;
    SB_DFFESS multi_byte_counter_i5 (.Q(multi_byte_counter[5]), .C(SLM_CLK_c), 
            .E(n4281), .D(n315[5]), .S(n4455));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i11024_3_lut_4_lut (.I0(state[2]), .I1(n1985[5]), .I2(state[0]), 
            .I3(state[3]), .O(n12607));   // src/spi.v(76[8] 221[4])
    defparam i11024_3_lut_4_lut.LUT_INIT = 16'h04ff;
    SB_DFFESR multi_byte_counter_i6 (.Q(multi_byte_counter[6]), .C(SLM_CLK_c), 
            .E(n4281), .D(n315[6]), .R(n4455));   // src/spi.v(76[8] 221[4])
    SB_LUT4 i2_3_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(state[1]), 
            .I3(state[3]), .O(n2));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h00b0;
    SB_DFFESS multi_byte_counter_i7 (.Q(multi_byte_counter[7]), .C(SLM_CLK_c), 
            .E(n4281), .D(n315[7]), .S(n4455));   // src/spi.v(76[8] 221[4])
    SB_LUT4 counter_1109_add_4_11_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[9]), 
            .I3(n10702), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1109_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1109_add_4_10_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[8]), 
            .I3(n10701), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1109_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1109_add_4_10 (.CI(n10701), .I0(VCC_net), .I1(counter[8]), 
            .CO(n10702));
    SB_LUT4 counter_1109_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[7]), 
            .I3(n10700), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1109_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1109_add_4_9 (.CI(n10700), .I0(VCC_net), .I1(counter[7]), 
            .CO(n10701));
    SB_LUT4 counter_1109_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[6]), 
            .I3(n10699), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1109_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1109_add_4_8 (.CI(n10699), .I0(VCC_net), .I1(counter[6]), 
            .CO(n10700));
    SB_LUT4 counter_1109_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(counter[5]), 
            .I3(n10698), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1109_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut (.I0(n11311), .I1(state[0]), .I2(state[2]), 
            .I3(n4105), .O(n11345));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hba00;
    SB_LUT4 i8605_3_lut_3_lut (.I0(state[2]), .I1(state[3]), .I2(state[0]), 
            .I3(GND_net), .O(n10119));   // src/spi.v(71[11:16])
    defparam i8605_3_lut_3_lut.LUT_INIT = 16'h1a1a;
    SB_LUT4 i10998_2_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(state[2]), 
            .I3(GND_net), .O(n12586));   // src/spi.v(88[9] 219[16])
    defparam i10998_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mux_56_Mux_3_i15_4_lut (.I0(n12586), .I1(state[1]), .I2(state[3]), 
            .I3(n1985[5]), .O(state_3__N_905[3]));   // src/spi.v(88[9] 219[16])
    defparam mux_56_Mux_3_i15_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i11110_3_lut (.I0(state[3]), .I1(n37), .I2(state[2]), .I3(GND_net), 
            .O(n19_adj_1139));
    defparam i11110_3_lut.LUT_INIT = 16'h1313;
    SB_LUT4 i42_4_lut (.I0(n21), .I1(n12576), .I2(state[1]), .I3(state[0]), 
            .O(n37));
    defparam i42_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i44_4_lut (.I0(spi_start_transfer_r), .I1(n19), .I2(state[3]), 
            .I3(state[2]), .O(n21));
    defparam i44_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 i11009_4_lut (.I0(state[2]), .I1(state[0]), .I2(n19), .I3(state[3]), 
            .O(n12576));
    defparam i11009_4_lut.LUT_INIT = 16'hccd0;
    SB_LUT4 i2103_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n3295));   // src/spi.v(88[9] 219[16])
    defparam i2103_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_33 (.I0(n12605), .I1(n14442), .I2(n10119), .I3(state[1]), 
            .O(state_3__N_905[2]));
    defparam i1_4_lut_adj_33.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_3_lut (.I0(n4105), .I1(state[2]), .I2(n11311), .I3(GND_net), 
            .O(n11344));
    defparam i1_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i2026_4_lut_4_lut (.I0(state[0]), .I1(state[2]), .I2(state[1]), 
            .I3(state[3]), .O(n3204));   // src/spi.v(88[9] 219[16])
    defparam i2026_4_lut_4_lut.LUT_INIT = 16'hfdfb;
    SB_LUT4 i8583_4_lut (.I0(n10090), .I1(n12594), .I2(state[1]), .I3(state[3]), 
            .O(state_3__N_905[1]));   // src/spi.v(71[11:16])
    defparam i8583_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11033_3_lut (.I0(n19), .I1(state[0]), .I2(state[2]), .I3(GND_net), 
            .O(n12594));   // src/spi.v(71[11:16])
    defparam i11033_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i1_4_lut_adj_34 (.I0(state[3]), .I1(n11344), .I2(state[2]), 
            .I3(n3295), .O(n11346));
    defparam i1_4_lut_adj_34.LUT_INIT = 16'h444c;
    SB_LUT4 i2318_4_lut_4_lut (.I0(state[2]), .I1(state[0]), .I2(state[1]), 
            .I3(state[3]), .O(n4409));   // src/spi.v(88[9] 219[16])
    defparam i2318_4_lut_4_lut.LUT_INIT = 16'hfe2f;
    SB_LUT4 i2_3_lut_4_lut_adj_35 (.I0(state[3]), .I1(state[2]), .I2(state[1]), 
            .I3(state[0]), .O(n11351));
    defparam i2_3_lut_4_lut_adj_35.LUT_INIT = 16'h0002;
    SB_LUT4 i1_4_lut_adj_36 (.I0(state[1]), .I1(n11350), .I2(n11398), 
            .I3(state[0]), .O(n4281));
    defparam i1_4_lut_adj_36.LUT_INIT = 16'h0a88;
    SB_LUT4 i3253_2_lut (.I0(n4281), .I1(state[3]), .I2(GND_net), .I3(GND_net), 
            .O(n4455));   // src/spi.v(76[8] 221[4])
    defparam i3253_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_322_Mux_2_i15_4_lut_4_lut (.I0(state[0]), .I1(state[1]), 
            .I2(state[3]), .I3(state[2]), .O(n860[2]));   // src/spi.v(88[9] 219[16])
    defparam mux_322_Mux_2_i15_4_lut_4_lut.LUT_INIT = 16'h0240;
    SB_LUT4 i11020_2_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(n8), .O(n12567));   // src/spi.v(88[9] 219[16])
    defparam i11020_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_4_lut_adj_37 (.I0(counter[0]), .I1(counter[1]), .I2(counter[3]), 
            .I3(counter[2]), .O(n8));
    defparam i1_2_lut_4_lut_adj_37.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module \uart_tx(CLKS_PER_BIT=20) 
//

module \uart_tx(CLKS_PER_BIT=20)  (UART_TX_c, SLM_CLK_c, r_SM_Main, n4724, 
            r_Tx_Data, n5861, VCC_net, r_Bit_Index, n14415, \r_SM_Main_2__N_808[1] , 
            GND_net, n4133, \r_SM_Main_2__N_811[0] , n4632, n4631, 
            tx_uart_active_flag, n11319, n3710, n4746, n4745, n4744, 
            n4743, n4742, n4740, n11339) /* synthesis syn_module_defined=1 */ ;
    output UART_TX_c;
    input SLM_CLK_c;
    output [2:0]r_SM_Main;
    input n4724;
    output [7:0]r_Tx_Data;
    input n5861;
    input VCC_net;
    output [2:0]r_Bit_Index;
    input n14415;
    output \r_SM_Main_2__N_808[1] ;
    input GND_net;
    output n4133;
    input \r_SM_Main_2__N_811[0] ;
    input n4632;
    input n4631;
    output tx_uart_active_flag;
    output n11319;
    output n3710;
    input n4746;
    input n4745;
    input n4744;
    input n4743;
    input n4742;
    input n4740;
    output n11339;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    wire n3, n1, n2814, n3_adj_1138;
    wire [9:0]n45;
    wire [9:0]r_Clock_Count;   // src/uart_tx.v(32[16:29])
    
    wire n4577, n10720, n10719, n10718;
    wire [2:0]r_Bit_Index_c;   // src/uart_tx.v(33[16:27])
    
    wire n12139, n12140, n13790, n12134, n12133, o_Tx_Serial_N_840, 
        n10717, n10716, n10715, n4, n8, n7;
    wire [2:0]n312;
    
    wire n4468;
    wire [2:0]r_SM_Main_2__N_805;
    
    wire n2813, n10714, n10713, n10712;
    
    SB_DFFE o_Tx_Serial_44 (.Q(UART_TX_c), .C(SLM_CLK_c), .E(n1), .D(n3));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(SLM_CLK_c), .D(n2814), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(SLM_CLK_c), .D(n4724));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(SLM_CLK_c), .D(n3_adj_1138), 
            .R(r_SM_Main[2]));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Clock_Count_1113__i0 (.Q(r_Clock_Count[0]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[0]), .R(n4577));   // src/uart_tx.v(116[34:51])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n5861));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(SLM_CLK_c), .D(n14415));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i11085_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_808[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n4577));
    defparam i11085_4_lut.LUT_INIT = 16'h4445;
    SB_DFFESR r_Clock_Count_1113__i9 (.Q(r_Clock_Count[9]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[9]), .R(n4577));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1113__i8 (.Q(r_Clock_Count[8]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[8]), .R(n4577));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1113__i7 (.Q(r_Clock_Count[7]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[7]), .R(n4577));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1113__i6 (.Q(r_Clock_Count[6]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[6]), .R(n4577));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1113__i5 (.Q(r_Clock_Count[5]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[5]), .R(n4577));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1113__i4 (.Q(r_Clock_Count[4]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[4]), .R(n4577));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1113__i3 (.Q(r_Clock_Count[3]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[3]), .R(n4577));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1113__i2 (.Q(r_Clock_Count[2]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[2]), .R(n4577));   // src/uart_tx.v(116[34:51])
    SB_DFFESR r_Clock_Count_1113__i1 (.Q(r_Clock_Count[1]), .C(SLM_CLK_c), 
            .E(n1), .D(n45[1]), .R(n4577));   // src/uart_tx.v(116[34:51])
    SB_LUT4 r_Clock_Count_1113_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[9]), .I3(n10720), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1113_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1113_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n10719), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1113_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1113_add_4_10 (.CI(n10719), .I0(GND_net), .I1(r_Clock_Count[8]), 
            .CO(n10720));
    SB_LUT4 r_Clock_Count_1113_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n10718), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1113_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1113_add_4_9 (.CI(n10718), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n10719));
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index_c[1]), .I1(n12139), 
            .I2(n12140), .I3(r_Bit_Index_c[2]), .O(n13790));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n13790_bdd_4_lut (.I0(n13790), .I1(n12134), .I2(n12133), .I3(r_Bit_Index_c[2]), 
            .O(o_Tx_Serial_N_840));
    defparam n13790_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 r_Clock_Count_1113_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n10717), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1113_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1113_add_4_8 (.CI(n10717), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n10718));
    SB_LUT4 r_Clock_Count_1113_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n10716), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1113_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1113_add_4_7 (.CI(n10716), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n10717));
    SB_LUT4 r_Clock_Count_1113_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n10715), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1113_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n4));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[9]), .I2(GND_net), 
            .I3(GND_net), .O(n8));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[4]), 
            .I3(n4), .O(n7));
    defparam i1_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i5_4_lut (.I0(r_Clock_Count[5]), .I1(n7), .I2(r_Clock_Count[7]), 
            .I3(n8), .O(\r_SM_Main_2__N_808[1] ));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index_c[1]), .C(SLM_CLK_c), .E(n4133), 
            .D(n312[1]), .R(n4468));   // src/uart_tx.v(38[10] 141[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index_c[2]), .C(SLM_CLK_c), .E(n4133), 
            .D(n312[2]), .R(n4468));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i1627_3_lut (.I0(\r_SM_Main_2__N_811[0] ), .I1(r_SM_Main_2__N_805[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n2813));   // src/uart_tx.v(41[7] 140[14])
    defparam i1627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1628_3_lut (.I0(n2813), .I1(\r_SM_Main_2__N_808[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n2814));   // src/uart_tx.v(41[7] 140[14])
    defparam i1628_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(SLM_CLK_c), .D(n4632));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Active_46 (.Q(tx_uart_active_flag), .C(SLM_CLK_c), .D(n4631));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i1257_2_lut_3_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), 
            .I2(r_Bit_Index_c[2]), .I3(GND_net), .O(n312[2]));   // src/uart_tx.v(96[36:51])
    defparam i1257_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), 
            .I2(r_Bit_Index_c[2]), .I3(GND_net), .O(n11319));   // src/uart_tx.v(96[36:51])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_805[0]), .O(n4468));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_3_lut_4_lut_adj_22 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_808[1] ), .O(n4133));
    defparam i1_3_lut_4_lut_adj_22.LUT_INIT = 16'h1101;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_811[0] ), .O(n3710));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_SM_Main_2__I_0_55_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_840), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // src/uart_tx.v(41[7] 140[14])
    defparam r_SM_Main_2__I_0_55_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_CARRY r_Clock_Count_1113_add_4_6 (.CI(n10715), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n10716));
    SB_LUT4 r_Clock_Count_1113_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n10714), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1113_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1113_add_4_5 (.CI(n10714), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n10715));
    SB_LUT4 r_Clock_Count_1113_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n10713), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1113_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1113_add_4_4 (.CI(n10713), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n10714));
    SB_LUT4 r_Clock_Count_1113_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n10712), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1113_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1113_add_4_3 (.CI(n10712), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n10713));
    SB_LUT4 r_Clock_Count_1113_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1113_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1113_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n10712));
    SB_DFF r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(SLM_CLK_c), .D(n4746));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(SLM_CLK_c), .D(n4745));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(SLM_CLK_c), .D(n4744));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(SLM_CLK_c), .D(n4743));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(SLM_CLK_c), .D(n4742));   // src/uart_tx.v(38[10] 141[8])
    SB_DFF r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(SLM_CLK_c), .D(n4740));   // src/uart_tx.v(38[10] 141[8])
    SB_LUT4 i10490_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n12139));
    defparam i10490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10491_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n12140));
    defparam i10491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10485_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n12134));
    defparam i10485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10484_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n12133));
    defparam i10484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6427_2_lut_4_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), 
            .I2(r_Bit_Index_c[2]), .I3(\r_SM_Main_2__N_808[1] ), .O(r_SM_Main_2__N_805[0]));
    defparam i6427_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11046_4_lut_4_lut (.I0(\r_SM_Main_2__N_808[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_811[0] ), .O(n11339));
    defparam i11046_4_lut_4_lut.LUT_INIT = 16'h8380;
    SB_LUT4 i1250_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n312[1]));   // src/uart_tx.v(96[36:51])
    defparam i1250_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2305_2_lut_3_lut (.I0(\r_SM_Main_2__N_808[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_1138));
    defparam i2305_2_lut_3_lut.LUT_INIT = 16'h7878;
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word
//

module FIFO_Quad_Word (rd_fifo_en_w, \mem_LUT.data_raw_r[0] , SLM_CLK_c, 
            rd_addr_r, reset_all_w, wr_addr_r, n5905, VCC_net, \fifo_temp_output[7] , 
            \rd_addr_p1_w[2] , GND_net, n5902, \fifo_temp_output[6] , 
            n5899, \fifo_temp_output[5] , n5890, \fifo_temp_output[4] , 
            n5887, \fifo_temp_output[3] , n5884, \fifo_temp_output[2] , 
            n1, n5881, \fifo_temp_output[1] , n10921, is_tx_fifo_full_flag, 
            \wr_addr_p1_w[2] , n5857, \fifo_temp_output[0] , n10727, 
            \rd_addr_p1_w[1] , n4679, rx_buf_byte, n4670, n11324, 
            is_fifo_empty_flag, n4674, n4697, fifo_write_cmd, full_nxt_r, 
            n2207, \mem_LUT.data_raw_r[7] , \mem_LUT.data_raw_r[6] , \mem_LUT.data_raw_r[5] , 
            \mem_LUT.data_raw_r[4] , \mem_LUT.data_raw_r[3] , \mem_LUT.data_raw_r[2] , 
            \mem_LUT.data_raw_r[1] , n4700, fifo_read_cmd, n4249, empty_o_N_1116) /* synthesis syn_module_defined=1 */ ;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[0] ;
    input SLM_CLK_c;
    output [2:0]rd_addr_r;
    input reset_all_w;
    output [2:0]wr_addr_r;
    input n5905;
    input VCC_net;
    output \fifo_temp_output[7] ;
    output \rd_addr_p1_w[2] ;
    input GND_net;
    input n5902;
    output \fifo_temp_output[6] ;
    input n5899;
    output \fifo_temp_output[5] ;
    input n5890;
    output \fifo_temp_output[4] ;
    input n5887;
    output \fifo_temp_output[3] ;
    input n5884;
    output \fifo_temp_output[2] ;
    output n1;
    input n5881;
    output \fifo_temp_output[1] ;
    input n10921;
    output is_tx_fifo_full_flag;
    output \wr_addr_p1_w[2] ;
    input n5857;
    output \fifo_temp_output[0] ;
    output n10727;
    output \rd_addr_p1_w[1] ;
    input n4679;
    input [7:0]rx_buf_byte;
    input n4670;
    input n11324;
    output is_fifo_empty_flag;
    input n4674;
    input n4697;
    input fifo_write_cmd;
    output full_nxt_r;
    input n2207;
    output \mem_LUT.data_raw_r[7] ;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[3] ;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[1] ;
    input n4700;
    input fifo_read_cmd;
    output n4249;
    output empty_o_N_1116;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    
    FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2 lscc_fifo_inst (.rd_fifo_en_w(rd_fifo_en_w), 
            .\mem_LUT.data_raw_r[0] (\mem_LUT.data_raw_r[0] ), .SLM_CLK_c(SLM_CLK_c), 
            .rd_addr_r({rd_addr_r}), .reset_all_w(reset_all_w), .wr_addr_r({wr_addr_r}), 
            .n5905(n5905), .VCC_net(VCC_net), .\fifo_temp_output[7] (\fifo_temp_output[7] ), 
            .\rd_addr_p1_w[2] (\rd_addr_p1_w[2] ), .GND_net(GND_net), .n5902(n5902), 
            .\fifo_temp_output[6] (\fifo_temp_output[6] ), .n5899(n5899), 
            .\fifo_temp_output[5] (\fifo_temp_output[5] ), .n5890(n5890), 
            .\fifo_temp_output[4] (\fifo_temp_output[4] ), .n5887(n5887), 
            .\fifo_temp_output[3] (\fifo_temp_output[3] ), .n5884(n5884), 
            .\fifo_temp_output[2] (\fifo_temp_output[2] ), .n1(n1), .n5881(n5881), 
            .\fifo_temp_output[1] (\fifo_temp_output[1] ), .n10921(n10921), 
            .is_tx_fifo_full_flag(is_tx_fifo_full_flag), .\wr_addr_p1_w[2] (\wr_addr_p1_w[2] ), 
            .n5857(n5857), .\fifo_temp_output[0] (\fifo_temp_output[0] ), 
            .n10727(n10727), .\rd_addr_p1_w[1] (\rd_addr_p1_w[1] ), .n4679(n4679), 
            .rx_buf_byte({rx_buf_byte}), .n4670(n4670), .n11324(n11324), 
            .is_fifo_empty_flag(is_fifo_empty_flag), .n4674(n4674), .n4697(n4697), 
            .fifo_write_cmd(fifo_write_cmd), .full_nxt_r(full_nxt_r), .n2207(n2207), 
            .\mem_LUT.data_raw_r[7] (\mem_LUT.data_raw_r[7] ), .\mem_LUT.data_raw_r[6] (\mem_LUT.data_raw_r[6] ), 
            .\mem_LUT.data_raw_r[5] (\mem_LUT.data_raw_r[5] ), .\mem_LUT.data_raw_r[4] (\mem_LUT.data_raw_r[4] ), 
            .\mem_LUT.data_raw_r[3] (\mem_LUT.data_raw_r[3] ), .\mem_LUT.data_raw_r[2] (\mem_LUT.data_raw_r[2] ), 
            .\mem_LUT.data_raw_r[1] (\mem_LUT.data_raw_r[1] ), .n4700(n4700), 
            .fifo_read_cmd(fifo_read_cmd), .n4249(n4249), .empty_o_N_1116(empty_o_N_1116)) /* synthesis syn_module_defined=1 */ ;   // src/fifo_quad_word_mod.v(20[37:380])
    
endmodule
//
// Verilog Description of module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2
//

module FIFO_Quad_Word_ipgen_lscc_fifo_renamed_due_excessive_length_2 (rd_fifo_en_w, 
            \mem_LUT.data_raw_r[0] , SLM_CLK_c, rd_addr_r, reset_all_w, 
            wr_addr_r, n5905, VCC_net, \fifo_temp_output[7] , \rd_addr_p1_w[2] , 
            GND_net, n5902, \fifo_temp_output[6] , n5899, \fifo_temp_output[5] , 
            n5890, \fifo_temp_output[4] , n5887, \fifo_temp_output[3] , 
            n5884, \fifo_temp_output[2] , n1, n5881, \fifo_temp_output[1] , 
            n10921, is_tx_fifo_full_flag, \wr_addr_p1_w[2] , n5857, 
            \fifo_temp_output[0] , n10727, \rd_addr_p1_w[1] , n4679, 
            rx_buf_byte, n4670, n11324, is_fifo_empty_flag, n4674, 
            n4697, fifo_write_cmd, full_nxt_r, n2207, \mem_LUT.data_raw_r[7] , 
            \mem_LUT.data_raw_r[6] , \mem_LUT.data_raw_r[5] , \mem_LUT.data_raw_r[4] , 
            \mem_LUT.data_raw_r[3] , \mem_LUT.data_raw_r[2] , \mem_LUT.data_raw_r[1] , 
            n4700, fifo_read_cmd, n4249, empty_o_N_1116) /* synthesis syn_module_defined=1 */ ;
    output rd_fifo_en_w;
    output \mem_LUT.data_raw_r[0] ;
    input SLM_CLK_c;
    output [2:0]rd_addr_r;
    input reset_all_w;
    output [2:0]wr_addr_r;
    input n5905;
    input VCC_net;
    output \fifo_temp_output[7] ;
    output \rd_addr_p1_w[2] ;
    input GND_net;
    input n5902;
    output \fifo_temp_output[6] ;
    input n5899;
    output \fifo_temp_output[5] ;
    input n5890;
    output \fifo_temp_output[4] ;
    input n5887;
    output \fifo_temp_output[3] ;
    input n5884;
    output \fifo_temp_output[2] ;
    output n1;
    input n5881;
    output \fifo_temp_output[1] ;
    input n10921;
    output is_tx_fifo_full_flag;
    output \wr_addr_p1_w[2] ;
    input n5857;
    output \fifo_temp_output[0] ;
    output n10727;
    output \rd_addr_p1_w[1] ;
    input n4679;
    input [7:0]rx_buf_byte;
    input n4670;
    input n11324;
    output is_fifo_empty_flag;
    input n4674;
    input n4697;
    input fifo_write_cmd;
    output full_nxt_r;
    input n2207;
    output \mem_LUT.data_raw_r[7] ;
    output \mem_LUT.data_raw_r[6] ;
    output \mem_LUT.data_raw_r[5] ;
    output \mem_LUT.data_raw_r[4] ;
    output \mem_LUT.data_raw_r[3] ;
    output \mem_LUT.data_raw_r[2] ;
    output \mem_LUT.data_raw_r[1] ;
    input n4700;
    input fifo_read_cmd;
    output n4249;
    output empty_o_N_1116;
    
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [31:0]\mem_LUT.data_raw_r_31__N_1051 ;
    wire [2:0]n12;
    wire [2:0]n12_adj_1137;
    wire [2:0]wr_addr_p1_w;   // src/fifo_quad_word_mod.v(67[32:44])
    
    wire n3, \mem_LUT.mem_2_6 , \mem_LUT.mem_3_6 , n13952, n5821, 
        \mem_LUT.mem_3_7 , n5820, n5819, \mem_LUT.mem_3_5 , \mem_LUT.mem_1_6 , 
        \mem_LUT.mem_0_6 , n5818, \mem_LUT.mem_3_4 , n5817, \mem_LUT.mem_3_3 , 
        n5816, \mem_LUT.mem_3_2 , n5815, \mem_LUT.mem_3_1 , n5814, 
        \mem_LUT.mem_3_0 , n5813, \mem_LUT.mem_2_7 , n5812, n5811, 
        \mem_LUT.mem_2_5 , n5810, \mem_LUT.mem_2_4 , n5809, \mem_LUT.mem_2_3 , 
        n5808, \mem_LUT.mem_2_2 , n5807, \mem_LUT.mem_2_1 , n5806, 
        \mem_LUT.mem_2_0 , n5805, \mem_LUT.mem_1_7 , n5804, n5803, 
        \mem_LUT.mem_1_5 , n5802, \mem_LUT.mem_1_4 , n5801, \mem_LUT.mem_1_3 , 
        n5800, \mem_LUT.mem_1_2 , n5799, \mem_LUT.mem_1_1 , n5798, 
        \mem_LUT.mem_1_0 , n5797, \mem_LUT.mem_0_7 , n5796, n5795, 
        \mem_LUT.mem_0_5 , n5794, \mem_LUT.mem_0_4 , n5793, \mem_LUT.mem_0_3 , 
        n5792, \mem_LUT.mem_0_2 , n5791, \mem_LUT.mem_0_1 , n5790, 
        \mem_LUT.mem_0_0 , rd_fifo_en_prev_r, n3_adj_1136, n4, n13766, 
        n13694, n13556, n13544, n13538, n14234, n13496;
    
    SB_DFFE \mem_LUT.data_raw_r__i1  (.Q(\mem_LUT.data_raw_r[0] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1051 [0]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFSR rd_addr_r__i0 (.Q(rd_addr_r[0]), .C(SLM_CLK_c), .D(n12[0]), 
            .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFSR wr_addr_r__i0 (.Q(wr_addr_r[0]), .C(SLM_CLK_c), .D(n12_adj_1137[0]), 
            .R(reset_all_w));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFFE \mem_LUT.data_buff_r__i7  (.Q(\fifo_temp_output[7] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n5905));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 i1333_3_lut (.I0(rd_addr_r[2]), .I1(rd_addr_r[1]), .I2(rd_addr_r[0]), 
            .I3(GND_net), .O(\rd_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1333_3_lut.LUT_INIT = 16'h6a6a;
    SB_DFFE \mem_LUT.data_buff_r__i6  (.Q(\fifo_temp_output[6] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n5902));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_buff_r__i5  (.Q(\fifo_temp_output[5] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n5899));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_buff_r__i4  (.Q(\fifo_temp_output[4] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n5890));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_buff_r__i3  (.Q(\fifo_temp_output[3] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n5887));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE \mem_LUT.data_buff_r__i2  (.Q(\fifo_temp_output[2] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n5884));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 i1304_2_lut (.I0(wr_addr_r[1]), .I1(wr_addr_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(wr_addr_p1_w[1]));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam i1304_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 wr_addr_r_1__I_0_i1_2_lut (.I0(wr_addr_r[0]), .I1(rd_addr_r[0]), 
            .I2(GND_net), .I3(GND_net), .O(n1));   // src/fifo_quad_word_mod.v(115[26:58])
    defparam wr_addr_r_1__I_0_i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE \mem_LUT.data_buff_r__i1  (.Q(\fifo_temp_output[1] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n5881));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_DFFE full_r_84 (.Q(is_tx_fifo_full_flag), .C(SLM_CLK_c), .E(VCC_net), 
            .D(n10921));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i1311_3_lut (.I0(wr_addr_r[2]), .I1(wr_addr_r[1]), .I2(wr_addr_r[0]), 
            .I3(GND_net), .O(\wr_addr_p1_w[2] ));   // src/fifo_quad_word_mod.v(67[47:65])
    defparam i1311_3_lut.LUT_INIT = 16'h6a6a;
    SB_DFFE \mem_LUT.data_buff_r__i0  (.Q(\fifo_temp_output[0] ), .C(SLM_CLK_c), 
            .E(VCC_net), .D(n5857));   // src/fifo_quad_word_mod.v(473[37] 486[40])
    SB_LUT4 i2_4_lut (.I0(wr_addr_p1_w[1]), .I1(n1), .I2(rd_addr_r[1]), 
            .I3(n3), .O(n10727));
    defparam i2_4_lut.LUT_INIT = 16'h8400;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12338 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_6 ), 
            .I2(\mem_LUT.mem_3_6 ), .I3(rd_addr_r[1]), .O(n13952));
    defparam rd_addr_r_0__bdd_4_lut_12338.LUT_INIT = 16'he4aa;
    SB_DFF i347_348 (.Q(\mem_LUT.mem_3_7 ), .C(SLM_CLK_c), .D(n5821));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i344_345 (.Q(\mem_LUT.mem_3_6 ), .C(SLM_CLK_c), .D(n5820));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i341_342 (.Q(\mem_LUT.mem_3_5 ), .C(SLM_CLK_c), .D(n5819));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_LUT4 n13952_bdd_4_lut (.I0(n13952), .I1(\mem_LUT.mem_1_6 ), .I2(\mem_LUT.mem_0_6 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1051 [6]));
    defparam n13952_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1326_2_lut (.I0(rd_addr_r[1]), .I1(rd_addr_r[0]), .I2(GND_net), 
            .I3(GND_net), .O(\rd_addr_p1_w[1] ));   // src/fifo_quad_word_mod.v(71[47:65])
    defparam i1326_2_lut.LUT_INIT = 16'h6666;
    SB_DFF i338_339 (.Q(\mem_LUT.mem_3_4 ), .C(SLM_CLK_c), .D(n5818));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i335_336 (.Q(\mem_LUT.mem_3_3 ), .C(SLM_CLK_c), .D(n5817));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i332_333 (.Q(\mem_LUT.mem_3_2 ), .C(SLM_CLK_c), .D(n5816));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i329_330 (.Q(\mem_LUT.mem_3_1 ), .C(SLM_CLK_c), .D(n5815));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i326_327 (.Q(\mem_LUT.mem_3_0 ), .C(SLM_CLK_c), .D(n5814));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i251_252 (.Q(\mem_LUT.mem_2_7 ), .C(SLM_CLK_c), .D(n5813));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i248_249 (.Q(\mem_LUT.mem_2_6 ), .C(SLM_CLK_c), .D(n5812));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i245_246 (.Q(\mem_LUT.mem_2_5 ), .C(SLM_CLK_c), .D(n5811));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i242_243 (.Q(\mem_LUT.mem_2_4 ), .C(SLM_CLK_c), .D(n5810));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i239_240 (.Q(\mem_LUT.mem_2_3 ), .C(SLM_CLK_c), .D(n5809));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i236_237 (.Q(\mem_LUT.mem_2_2 ), .C(SLM_CLK_c), .D(n5808));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i233_234 (.Q(\mem_LUT.mem_2_1 ), .C(SLM_CLK_c), .D(n5807));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i230_231 (.Q(\mem_LUT.mem_2_0 ), .C(SLM_CLK_c), .D(n5806));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i155_156 (.Q(\mem_LUT.mem_1_7 ), .C(SLM_CLK_c), .D(n5805));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i152_153 (.Q(\mem_LUT.mem_1_6 ), .C(SLM_CLK_c), .D(n5804));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i149_150 (.Q(\mem_LUT.mem_1_5 ), .C(SLM_CLK_c), .D(n5803));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i146_147 (.Q(\mem_LUT.mem_1_4 ), .C(SLM_CLK_c), .D(n5802));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i143_144 (.Q(\mem_LUT.mem_1_3 ), .C(SLM_CLK_c), .D(n5801));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i140_141 (.Q(\mem_LUT.mem_1_2 ), .C(SLM_CLK_c), .D(n5800));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i137_138 (.Q(\mem_LUT.mem_1_1 ), .C(SLM_CLK_c), .D(n5799));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i134_135 (.Q(\mem_LUT.mem_1_0 ), .C(SLM_CLK_c), .D(n5798));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i59_60 (.Q(\mem_LUT.mem_0_7 ), .C(SLM_CLK_c), .D(n5797));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i56_57 (.Q(\mem_LUT.mem_0_6 ), .C(SLM_CLK_c), .D(n5796));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i53_54 (.Q(\mem_LUT.mem_0_5 ), .C(SLM_CLK_c), .D(n5795));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i50_51 (.Q(\mem_LUT.mem_0_4 ), .C(SLM_CLK_c), .D(n5794));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i47_48 (.Q(\mem_LUT.mem_0_3 ), .C(SLM_CLK_c), .D(n5793));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i44_45 (.Q(\mem_LUT.mem_0_2 ), .C(SLM_CLK_c), .D(n5792));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i41_42 (.Q(\mem_LUT.mem_0_1 ), .C(SLM_CLK_c), .D(n5791));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF i38_39 (.Q(\mem_LUT.mem_0_0 ), .C(SLM_CLK_c), .D(n5790));   // src/fifo_quad_word_mod.v(448[73:76])
    SB_DFF rd_fifo_en_prev_r_86 (.Q(rd_fifo_en_prev_r), .C(SLM_CLK_c), .D(n4679));   // src/fifo_quad_word_mod.v(353[29] 363[32])
    SB_LUT4 i4619_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_3_7 ), .O(n5821));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4619_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF rd_addr_r__i1 (.Q(rd_addr_r[1]), .C(SLM_CLK_c), .D(n4670));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF empty_r_85 (.Q(is_fifo_empty_flag), .C(SLM_CLK_c), .D(n11324));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_DFF rd_addr_r__i2 (.Q(rd_addr_r[2]), .C(SLM_CLK_c), .D(n4674));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i4618_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_3_6 ), .O(n5820));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4618_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4617_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_3_5 ), .O(n5819));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4617_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4616_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_3_4 ), .O(n5818));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4616_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4615_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_3_3 ), .O(n5817));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4615_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4614_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_3_2 ), .O(n5816));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4614_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4613_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_3_1 ), .O(n5815));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4613_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4612_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_3_0 ), .O(n5814));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4612_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF wr_addr_r__i1 (.Q(wr_addr_r[1]), .C(SLM_CLK_c), .D(n4697));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i4611_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_2_7 ), .O(n5813));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4611_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4610_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_2_6 ), .O(n5812));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4610_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4609_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_2_5 ), .O(n5811));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4609_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 wr_en_i_I_0_2_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(GND_net), .I3(GND_net), .O(full_nxt_r));   // src/fifo_quad_word_mod.v(103[21:60])
    defparam wr_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1516_2_lut (.I0(wr_addr_r[0]), .I1(n2207), .I2(GND_net), 
            .I3(GND_net), .O(n12_adj_1137[0]));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1516_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_12103 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_5 ), 
            .I2(\mem_LUT.mem_3_5 ), .I3(rd_addr_r[1]), .O(n13766));
    defparam rd_addr_r_0__bdd_4_lut_12103.LUT_INIT = 16'he4aa;
    SB_LUT4 n13766_bdd_4_lut (.I0(n13766), .I1(\mem_LUT.mem_1_5 ), .I2(\mem_LUT.mem_0_5 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1051 [5]));
    defparam n13766_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \mem_LUT.data_raw_r__i8  (.Q(\mem_LUT.data_raw_r[7] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1051 [7]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i7  (.Q(\mem_LUT.data_raw_r[6] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1051 [6]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i6  (.Q(\mem_LUT.data_raw_r[5] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1051 [5]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i5  (.Q(\mem_LUT.data_raw_r[4] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1051 [4]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i4  (.Q(\mem_LUT.data_raw_r[3] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1051 [3]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i3  (.Q(\mem_LUT.data_raw_r[2] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1051 [2]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFFE \mem_LUT.data_raw_r__i2  (.Q(\mem_LUT.data_raw_r[1] ), .C(SLM_CLK_c), 
            .E(rd_fifo_en_w), .D(\mem_LUT.data_raw_r_31__N_1051 [1]));   // src/fifo_quad_word_mod.v(461[21] 467[24])
    SB_DFF wr_addr_r__i2 (.Q(wr_addr_r[2]), .C(SLM_CLK_c), .D(n4700));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    SB_LUT4 i4608_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_2_4 ), .O(n5810));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4608_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4607_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_2_3 ), .O(n5809));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4607_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4606_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_2_2 ), .O(n5808));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4606_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4605_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_2_1 ), .O(n5807));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4605_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11949 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_4 ), 
            .I2(\mem_LUT.mem_3_4 ), .I3(rd_addr_r[1]), .O(n13694));
    defparam rd_addr_r_0__bdd_4_lut_11949.LUT_INIT = 16'he4aa;
    SB_LUT4 n13694_bdd_4_lut (.I0(n13694), .I1(\mem_LUT.mem_1_4 ), .I2(\mem_LUT.mem_0_4 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1051 [4]));
    defparam n13694_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4604_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_2_0 ), .O(n5806));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4604_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1518_2_lut_4_lut (.I0(rd_addr_r[0]), .I1(fifo_read_cmd), .I2(is_fifo_empty_flag), 
            .I3(reset_all_w), .O(n12[0]));   // src/fifo_quad_word_mod.v(145[21] 161[24])
    defparam i1518_2_lut_4_lut.LUT_INIT = 16'h55a6;
    SB_LUT4 i4603_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_1_7 ), .O(n5805));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4603_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4602_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_1_6 ), .O(n5804));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4602_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_en_i_I_0_2_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(GND_net), .I3(GND_net), .O(rd_fifo_en_w));   // src/fifo_quad_word_mod.v(62[29:51])
    defparam rd_en_i_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4601_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_1_5 ), .O(n5803));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4601_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4600_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_1_4 ), .O(n5802));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4600_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4599_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_1_3 ), .O(n5801));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4599_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4598_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_1_2 ), .O(n5800));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4598_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4597_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_1_1 ), .O(n5799));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4597_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4596_3_lut_4_lut (.I0(n3_adj_1136), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_1_0 ), .O(n5798));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4596_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4595_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[7]), 
            .I3(\mem_LUT.mem_0_7 ), .O(n5797));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4595_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4594_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[6]), 
            .I3(\mem_LUT.mem_0_6 ), .O(n5796));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4594_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4593_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[5]), 
            .I3(\mem_LUT.mem_0_5 ), .O(n5795));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4593_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4592_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[4]), 
            .I3(\mem_LUT.mem_0_4 ), .O(n5794));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4592_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4591_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[3]), 
            .I3(\mem_LUT.mem_0_3 ), .O(n5793));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4591_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4590_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[2]), 
            .I3(\mem_LUT.mem_0_2 ), .O(n5792));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4590_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4589_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[1]), 
            .I3(\mem_LUT.mem_0_1 ), .O(n5791));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4589_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4588_3_lut_4_lut (.I0(n4), .I1(wr_addr_r[1]), .I2(rx_buf_byte[0]), 
            .I3(\mem_LUT.mem_0_0 ), .O(n5790));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam i4588_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11889 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_3 ), 
            .I2(\mem_LUT.mem_3_3 ), .I3(rd_addr_r[1]), .O(n13556));
    defparam rd_addr_r_0__bdd_4_lut_11889.LUT_INIT = 16'he4aa;
    SB_LUT4 n13556_bdd_4_lut (.I0(n13556), .I1(\mem_LUT.mem_1_3 ), .I2(\mem_LUT.mem_0_3 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1051 [3]));
    defparam n13556_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11774 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_2 ), 
            .I2(\mem_LUT.mem_3_2 ), .I3(rd_addr_r[1]), .O(n13544));
    defparam rd_addr_r_0__bdd_4_lut_11774.LUT_INIT = 16'he4aa;
    SB_LUT4 n13544_bdd_4_lut (.I0(n13544), .I1(\mem_LUT.mem_1_2 ), .I2(\mem_LUT.mem_0_2 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1051 [2]));
    defparam n13544_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11764 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_1 ), 
            .I2(\mem_LUT.mem_3_1 ), .I3(rd_addr_r[1]), .O(n13538));
    defparam rd_addr_r_0__bdd_4_lut_11764.LUT_INIT = 16'he4aa;
    SB_LUT4 n13538_bdd_4_lut (.I0(n13538), .I1(\mem_LUT.mem_1_1 ), .I2(\mem_LUT.mem_0_1 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1051 [1]));
    defparam n13538_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_7 ), 
            .I2(\mem_LUT.mem_3_7 ), .I3(rd_addr_r[1]), .O(n14234));
    defparam rd_addr_r_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n14234_bdd_4_lut (.I0(n14234), .I1(\mem_LUT.mem_1_7 ), .I2(\mem_LUT.mem_0_7 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1051 [7]));
    defparam n14234_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 rd_addr_r_0__bdd_4_lut_11759 (.I0(rd_addr_r[0]), .I1(\mem_LUT.mem_2_0 ), 
            .I2(\mem_LUT.mem_3_0 ), .I3(rd_addr_r[1]), .O(n13496));
    defparam rd_addr_r_0__bdd_4_lut_11759.LUT_INIT = 16'he4aa;
    SB_LUT4 n13496_bdd_4_lut (.I0(n13496), .I1(\mem_LUT.mem_1_0 ), .I2(\mem_LUT.mem_0_0 ), 
            .I3(rd_addr_r[1]), .O(\mem_LUT.data_raw_r_31__N_1051 [0]));
    defparam n13496_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(rd_fifo_en_prev_r), .I1(fifo_read_cmd), 
            .I2(is_fifo_empty_flag), .I3(reset_all_w), .O(n4249));   // src/fifo_quad_word_mod.v(155[29] 160[32])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hffae;
    SB_LUT4 i3110_2_lut_3_lut (.I0(fifo_read_cmd), .I1(is_fifo_empty_flag), 
            .I2(reset_all_w), .I3(GND_net), .O(empty_o_N_1116));   // src/fifo_quad_word_mod.v(155[29] 160[32])
    defparam i3110_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 wr_addr_p1_w_2__I_0_i3_2_lut_4_lut (.I0(wr_addr_r[2]), .I1(wr_addr_r[1]), 
            .I2(wr_addr_r[0]), .I3(rd_addr_r[2]), .O(n3));   // src/fifo_quad_word_mod.v(107[37:64])
    defparam wr_addr_p1_w_2__I_0_i3_2_lut_4_lut.LUT_INIT = 16'h956a;
    SB_LUT4 EnabledDecoder_2_i3_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n3_adj_1136));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i3_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 EnabledDecoder_2_i4_2_lut_3_lut (.I0(fifo_write_cmd), .I1(is_tx_fifo_full_flag), 
            .I2(wr_addr_r[0]), .I3(GND_net), .O(n4));   // src/fifo_quad_word_mod.v(457[33:51])
    defparam EnabledDecoder_2_i4_2_lut_3_lut.LUT_INIT = 16'h0202;
    
endmodule
//
// Verilog Description of module usb3_if
//

module usb3_if (VCC_net, GND_net, \dc32_fifo_data_in[13] , DEBUG_6_c_c, 
            \dc32_fifo_data_in[12] , \dc32_fifo_data_in[11] , \dc32_fifo_data_in[10] , 
            \dc32_fifo_data_in[9] , \dc32_fifo_data_in[8] , \dc32_fifo_data_in[7] , 
            \dc32_fifo_data_in[6] , \dc32_fifo_data_in[5] , \dc32_fifo_data_in[4] , 
            DEBUG_3_c, \dc32_fifo_data_in[0] , buffer_switch_done, buffer_switch_done_latched, 
            SLM_CLK_c, reset_per_frame, FT_OE_c, \dc32_fifo_data_in[3] , 
            DEBUG_9_c, \dc32_fifo_data_in[2] , \dc32_fifo_data_in[1] , 
            DEBUG_2_c_c, \dc32_fifo_data_in[15] , DEBUG_5_c, FIFO_D15_c_15, 
            FIFO_D14_c_14, FIFO_D13_c_13, FIFO_D12_c_12, FIFO_D11_c_11, 
            FIFO_D10_c_10, FIFO_D9_c_9, FIFO_D8_c_8, FIFO_D7_c_7, FIFO_D6_c_6, 
            FIFO_D5_c_5, FIFO_D4_c_4, FIFO_D3_c_3, FIFO_D2_c_2, FIFO_D1_c_1, 
            \afull_flag_impl.af_flag_p_w_N_603[3] , \dc32_fifo_data_in[14] , 
            DEBUG_1_c_0_c) /* synthesis syn_module_defined=1 */ ;
    input VCC_net;
    input GND_net;
    output \dc32_fifo_data_in[13] ;
    input DEBUG_6_c_c;
    output \dc32_fifo_data_in[12] ;
    output \dc32_fifo_data_in[11] ;
    output \dc32_fifo_data_in[10] ;
    output \dc32_fifo_data_in[9] ;
    output \dc32_fifo_data_in[8] ;
    output \dc32_fifo_data_in[7] ;
    output \dc32_fifo_data_in[6] ;
    output \dc32_fifo_data_in[5] ;
    output \dc32_fifo_data_in[4] ;
    output DEBUG_3_c;
    output \dc32_fifo_data_in[0] ;
    input buffer_switch_done;
    output buffer_switch_done_latched;
    input SLM_CLK_c;
    input reset_per_frame;
    output FT_OE_c;
    output \dc32_fifo_data_in[3] ;
    input DEBUG_9_c;
    output \dc32_fifo_data_in[2] ;
    output \dc32_fifo_data_in[1] ;
    input DEBUG_2_c_c;
    output \dc32_fifo_data_in[15] ;
    input DEBUG_5_c;
    input FIFO_D15_c_15;
    input FIFO_D14_c_14;
    input FIFO_D13_c_13;
    input FIFO_D12_c_12;
    input FIFO_D11_c_11;
    input FIFO_D10_c_10;
    input FIFO_D9_c_9;
    input FIFO_D8_c_8;
    input FIFO_D7_c_7;
    input FIFO_D6_c_6;
    input FIFO_D5_c_5;
    input FIFO_D4_c_4;
    input FIFO_D3_c_3;
    input FIFO_D2_c_2;
    input FIFO_D1_c_1;
    output \afull_flag_impl.af_flag_p_w_N_603[3] ;
    output \dc32_fifo_data_in[14] ;
    input DEBUG_1_c_0_c;
    
    wire DEBUG_6_c_c /* synthesis is_clock=1, SET_AS_NETWORK=DEBUG_6_c_c */ ;   // src/top.v(84[12:20])
    wire SLM_CLK_c /* synthesis SET_AS_NETWORK=SLM_CLK_c, is_clock=1 */ ;   // src/top.v(29[12:19])
    wire [10:0]num_lines_clocked_out_10__N_368;
    wire [10:0]num_lines_clocked_out;   // src/usb3_if.v(67[12:33])
    
    wire n10665;
    wire [31:0]usb3_data_in_latched;   // src/usb3_if.v(63[12:32])
    wire [3:0]state_timeout_counter_3__N_379;
    
    wire n4061;
    wire [3:0]state_timeout_counter;   // src/usb3_if.v(68[11:32])
    
    wire n10666, FT_RD_N_387, reset_per_frame_latched, FT_OE_N_384, 
        n3684;
    wire [3:0]n134;
    wire [7:0]n547;
    
    wire n2798, n2912, n7505, n4403, n6904, n2760, n10664, n10663, 
        n2908, n10751, n4178, n10662, n10661, n10660, empty_o_N_599, 
        n5687, n7, n4, n21, n3686, n2744, n10750, n2754, n14425, 
        n4650, n7360, n3973, n10869, n18, n16, n20, n12582, 
        n10669, n10668, n10667, n2739, n534, n5, n10746, n2755;
    
    SB_LUT4 sub_113_add_2_8_lut (.I0(GND_net), .I1(num_lines_clocked_out[6]), 
            .I2(VCC_net), .I3(n10665), .O(num_lines_clocked_out_10__N_368[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFN dc32_fifo_data_in_i14 (.Q(\dc32_fifo_data_in[13] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[13]));   // src/usb3_if.v(159[8] 161[4])
    SB_DFFN dc32_fifo_data_in_i13 (.Q(\dc32_fifo_data_in[12] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[12]));   // src/usb3_if.v(159[8] 161[4])
    SB_DFFN dc32_fifo_data_in_i12 (.Q(\dc32_fifo_data_in[11] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[11]));   // src/usb3_if.v(159[8] 161[4])
    SB_DFFNE state_timeout_counter_i0_i0 (.Q(state_timeout_counter[0]), .C(DEBUG_6_c_c), 
            .E(n4061), .D(state_timeout_counter_3__N_379[0]));   // src/usb3_if.v(72[8] 146[4])
    SB_DFFN dc32_fifo_data_in_i11 (.Q(\dc32_fifo_data_in[10] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[10]));   // src/usb3_if.v(159[8] 161[4])
    SB_DFFN dc32_fifo_data_in_i10 (.Q(\dc32_fifo_data_in[9] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[9]));   // src/usb3_if.v(159[8] 161[4])
    SB_DFFN dc32_fifo_data_in_i9 (.Q(\dc32_fifo_data_in[8] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[8]));   // src/usb3_if.v(159[8] 161[4])
    SB_DFFN dc32_fifo_data_in_i8 (.Q(\dc32_fifo_data_in[7] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[7]));   // src/usb3_if.v(159[8] 161[4])
    SB_DFFN dc32_fifo_data_in_i7 (.Q(\dc32_fifo_data_in[6] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[6]));   // src/usb3_if.v(159[8] 161[4])
    SB_DFFN dc32_fifo_data_in_i6 (.Q(\dc32_fifo_data_in[5] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[5]));   // src/usb3_if.v(159[8] 161[4])
    SB_DFFN dc32_fifo_data_in_i5 (.Q(\dc32_fifo_data_in[4] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[4]));   // src/usb3_if.v(159[8] 161[4])
    SB_CARRY sub_113_add_2_8 (.CI(n10665), .I0(num_lines_clocked_out[6]), 
            .I1(VCC_net), .CO(n10666));
    SB_DFFNSS FT_RD_internal_75 (.Q(DEBUG_3_c), .C(DEBUG_6_c_c), .D(FT_RD_N_387), 
            .S(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_DFFN dc32_fifo_data_in_i1 (.Q(\dc32_fifo_data_in[0] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[0]));   // src/usb3_if.v(159[8] 161[4])
    SB_DFF buffer_switch_done_latched_81 (.Q(buffer_switch_done_latched), 
           .C(SLM_CLK_c), .D(buffer_switch_done));   // src/usb3_if.v(164[8] 173[4])
    SB_DFF reset_per_frame_latched_82 (.Q(reset_per_frame_latched), .C(SLM_CLK_c), 
           .D(reset_per_frame));   // src/usb3_if.v(164[8] 173[4])
    SB_DFFNSS FT_OE_internal_74 (.Q(FT_OE_c), .C(DEBUG_6_c_c), .D(FT_OE_N_384), 
            .S(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_DFFN dc32_fifo_data_in_i4 (.Q(\dc32_fifo_data_in[3] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[3]));   // src/usb3_if.v(159[8] 161[4])
    SB_LUT4 i1_2_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n3684));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1726_4_lut (.I0(n3684), .I1(n134[1]), .I2(n547[2]), .I3(n2798), 
            .O(n2912));   // src/usb3_if.v(80[9] 144[16])
    defparam i1726_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i1727_3_lut (.I0(n2912), .I1(DEBUG_9_c), .I2(n547[5]), .I3(GND_net), 
            .O(state_timeout_counter_3__N_379[1]));   // src/usb3_if.v(80[9] 144[16])
    defparam i1727_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFN dc32_fifo_data_in_i3 (.Q(\dc32_fifo_data_in[2] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[2]));   // src/usb3_if.v(159[8] 161[4])
    SB_LUT4 i5710_4_lut (.I0(n7505), .I1(n4403), .I2(n547[2]), .I3(n547[1]), 
            .O(n6904));   // src/usb3_if.v(80[9] 144[16])
    defparam i5710_4_lut.LUT_INIT = 16'h3530;
    SB_DFFN dc32_fifo_data_in_i2 (.Q(\dc32_fifo_data_in[1] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[1]));   // src/usb3_if.v(159[8] 161[4])
    SB_LUT4 i5713_4_lut (.I0(n6904), .I1(DEBUG_9_c), .I2(n547[5]), .I3(DEBUG_2_c_c), 
            .O(state_timeout_counter_3__N_379[2]));   // src/usb3_if.v(80[9] 144[16])
    defparam i5713_4_lut.LUT_INIT = 16'h3a0a;
    SB_DFFNSS state_FSM_i1 (.Q(n547[0]), .C(DEBUG_6_c_c), .D(n2760), .S(reset_per_frame_latched));   // src/usb3_if.v(80[9] 144[16])
    SB_LUT4 sub_113_add_2_7_lut (.I0(GND_net), .I1(num_lines_clocked_out[5]), 
            .I2(VCC_net), .I3(n10664), .O(num_lines_clocked_out_10__N_368[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_7 (.CI(n10664), .I0(num_lines_clocked_out[5]), 
            .I1(VCC_net), .CO(n10665));
    SB_LUT4 sub_113_add_2_6_lut (.I0(GND_net), .I1(num_lines_clocked_out[4]), 
            .I2(VCC_net), .I3(n10663), .O(num_lines_clocked_out_10__N_368[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFNESR state_timeout_counter_i0_i3 (.Q(state_timeout_counter[3]), 
            .C(DEBUG_6_c_c), .E(n4061), .D(n2908), .R(n10751));   // src/usb3_if.v(72[8] 146[4])
    SB_DFFNESR num_lines_clocked_out_i1 (.Q(num_lines_clocked_out[1]), .C(DEBUG_6_c_c), 
            .E(n4178), .D(num_lines_clocked_out_10__N_368[1]), .R(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_DFFNESR num_lines_clocked_out_i2 (.Q(num_lines_clocked_out[2]), .C(DEBUG_6_c_c), 
            .E(n4178), .D(num_lines_clocked_out_10__N_368[2]), .R(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_DFFNESR num_lines_clocked_out_i3 (.Q(num_lines_clocked_out[3]), .C(DEBUG_6_c_c), 
            .E(n4178), .D(num_lines_clocked_out_10__N_368[3]), .R(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_CARRY sub_113_add_2_6 (.CI(n10663), .I0(num_lines_clocked_out[4]), 
            .I1(VCC_net), .CO(n10664));
    SB_DFFNESS num_lines_clocked_out_i4 (.Q(num_lines_clocked_out[4]), .C(DEBUG_6_c_c), 
            .E(n4178), .D(num_lines_clocked_out_10__N_368[4]), .S(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_LUT4 sub_113_add_2_5_lut (.I0(GND_net), .I1(num_lines_clocked_out[3]), 
            .I2(VCC_net), .I3(n10662), .O(num_lines_clocked_out_10__N_368[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFNESR num_lines_clocked_out_i5 (.Q(num_lines_clocked_out[5]), .C(DEBUG_6_c_c), 
            .E(n4178), .D(num_lines_clocked_out_10__N_368[5]), .R(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_DFFNESR num_lines_clocked_out_i6 (.Q(num_lines_clocked_out[6]), .C(DEBUG_6_c_c), 
            .E(n4178), .D(num_lines_clocked_out_10__N_368[6]), .R(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_CARRY sub_113_add_2_5 (.CI(n10662), .I0(num_lines_clocked_out[3]), 
            .I1(VCC_net), .CO(n10663));
    SB_LUT4 sub_113_add_2_4_lut (.I0(GND_net), .I1(num_lines_clocked_out[2]), 
            .I2(VCC_net), .I3(n10661), .O(num_lines_clocked_out_10__N_368[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_4 (.CI(n10661), .I0(num_lines_clocked_out[2]), 
            .I1(VCC_net), .CO(n10662));
    SB_LUT4 sub_113_add_2_3_lut (.I0(GND_net), .I1(num_lines_clocked_out[1]), 
            .I2(VCC_net), .I3(n10660), .O(num_lines_clocked_out_10__N_368[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_3 (.CI(n10660), .I0(num_lines_clocked_out[1]), 
            .I1(VCC_net), .CO(n10661));
    SB_LUT4 sub_113_add_2_2_lut (.I0(GND_net), .I1(num_lines_clocked_out[0]), 
            .I2(empty_o_N_599), .I3(VCC_net), .O(num_lines_clocked_out_10__N_368[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_2 (.CI(VCC_net), .I0(num_lines_clocked_out[0]), 
            .I1(empty_o_N_599), .CO(n10660));
    SB_DFFN state_FSM_i5 (.Q(n547[4]), .C(DEBUG_6_c_c), .D(n5687));   // src/usb3_if.v(80[9] 144[16])
    SB_DFFN dc32_fifo_data_in_i16 (.Q(\dc32_fifo_data_in[15] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[15]));   // src/usb3_if.v(159[8] 161[4])
    SB_LUT4 i1_3_lut (.I0(n7), .I1(reset_per_frame_latched), .I2(n547[2]), 
            .I3(GND_net), .O(n4178));
    defparam i1_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 i1277_2_lut (.I0(state_timeout_counter[1]), .I1(state_timeout_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // src/usb3_if.v(126[42:69])
    defparam i1277_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mux_40_i4_4_lut (.I0(n21), .I1(n3686), .I2(n7), .I3(DEBUG_5_c), 
            .O(n134[3]));   // src/usb3_if.v(127[17] 142[20])
    defparam mux_40_i4_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i1722_4_lut (.I0(n3686), .I1(n134[3]), .I2(n547[2]), .I3(n2798), 
            .O(n2908));   // src/usb3_if.v(80[9] 144[16])
    defparam i1722_4_lut.LUT_INIT = 16'hc5c0;
    SB_DFFESR usb3_data_in_latched__i16 (.Q(usb3_data_in_latched[15]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D15_c_15), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i15 (.Q(usb3_data_in_latched[14]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D14_c_14), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i14 (.Q(usb3_data_in_latched[13]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D13_c_13), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i13 (.Q(usb3_data_in_latched[12]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D12_c_12), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i12 (.Q(usb3_data_in_latched[11]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D11_c_11), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i11 (.Q(usb3_data_in_latched[10]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D10_c_10), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i10 (.Q(usb3_data_in_latched[9]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D9_c_9), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i9 (.Q(usb3_data_in_latched[8]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D8_c_8), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i8 (.Q(usb3_data_in_latched[7]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D7_c_7), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i7 (.Q(usb3_data_in_latched[6]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D6_c_6), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i6 (.Q(usb3_data_in_latched[5]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D5_c_5), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i5 (.Q(usb3_data_in_latched[4]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D4_c_4), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i4 (.Q(usb3_data_in_latched[3]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D3_c_3), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i3 (.Q(usb3_data_in_latched[2]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D2_c_2), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFESR usb3_data_in_latched__i2 (.Q(usb3_data_in_latched[1]), .C(DEBUG_6_c_c), 
            .E(VCC_net), .D(FIFO_D1_c_1), .R(reset_per_frame_latched));   // src/usb3_if.v(149[8] 156[4])
    SB_DFFNE state_timeout_counter_i0_i2 (.Q(state_timeout_counter[2]), .C(DEBUG_6_c_c), 
            .E(n4061), .D(state_timeout_counter_3__N_379[2]));   // src/usb3_if.v(72[8] 146[4])
    SB_DFFNE state_timeout_counter_i0_i1 (.Q(state_timeout_counter[1]), .C(DEBUG_6_c_c), 
            .E(n4061), .D(state_timeout_counter_3__N_379[1]));   // src/usb3_if.v(72[8] 146[4])
    SB_DFFNSR state_FSM_i6 (.Q(n547[5]), .C(DEBUG_6_c_c), .D(n2744), .R(reset_per_frame_latched));   // src/usb3_if.v(80[9] 144[16])
    SB_DFFNSR state_FSM_i4 (.Q(n547[3]), .C(DEBUG_6_c_c), .D(n10750), 
            .R(reset_per_frame_latched));   // src/usb3_if.v(80[9] 144[16])
    SB_DFFNSR state_FSM_i3 (.Q(n547[2]), .C(DEBUG_6_c_c), .D(n2754), .R(reset_per_frame_latched));   // src/usb3_if.v(80[9] 144[16])
    SB_DFFNSR state_FSM_i2 (.Q(n547[1]), .C(DEBUG_6_c_c), .D(n14425), 
            .R(reset_per_frame_latched));   // src/usb3_if.v(80[9] 144[16])
    SB_DFF usb3_data_in_latched__i1 (.Q(usb3_data_in_latched[0]), .C(DEBUG_6_c_c), 
           .D(n4650));   // src/usb3_if.v(149[8] 156[4])
    SB_LUT4 i6327_2_lut_3_lut_4_lut (.I0(n7360), .I1(n7), .I2(n4), .I3(state_timeout_counter[2]), 
            .O(n7505));   // src/usb3_if.v(93[17] 100[20])
    defparam i6327_2_lut_3_lut_4_lut.LUT_INIT = 16'h0dd0;
    SB_LUT4 i2_3_lut (.I0(n7), .I1(n547[2]), .I2(DEBUG_5_c), .I3(GND_net), 
            .O(n3973));   // src/usb3_if.v(80[9] 144[16])
    defparam i2_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2_3_lut_adj_14 (.I0(buffer_switch_done_latched), .I1(DEBUG_2_c_c), 
            .I2(DEBUG_5_c), .I3(GND_net), .O(n10869));
    defparam i2_3_lut_adj_14.LUT_INIT = 16'hdfdf;
    SB_LUT4 i1576_4_lut (.I0(n10869), .I1(n21), .I2(n547[0]), .I3(n3973), 
            .O(n2760));   // src/usb3_if.v(80[9] 144[16])
    defparam i1576_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 i1_2_lut_adj_15 (.I0(reset_per_frame_latched), .I1(n547[3]), 
            .I2(GND_net), .I3(GND_net), .O(n5687));   // src/usb3_if.v(164[8] 173[4])
    defparam i1_2_lut_adj_15.LUT_INIT = 16'h4444;
    SB_DFFNESR num_lines_clocked_out_i7 (.Q(num_lines_clocked_out[7]), .C(DEBUG_6_c_c), 
            .E(n4178), .D(num_lines_clocked_out_10__N_368[7]), .R(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(n547[5]), .I1(n547[4]), .I2(n547[3]), 
            .I3(n7360), .O(FT_OE_N_384));
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'hab01;
    SB_DFFNESR num_lines_clocked_out_i8 (.Q(num_lines_clocked_out[8]), .C(DEBUG_6_c_c), 
            .E(n4178), .D(num_lines_clocked_out_10__N_368[8]), .R(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_DFFNESR num_lines_clocked_out_i9 (.Q(num_lines_clocked_out[9]), .C(DEBUG_6_c_c), 
            .E(n4178), .D(num_lines_clocked_out_10__N_368[9]), .R(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_DFFNESR num_lines_clocked_out_i10 (.Q(num_lines_clocked_out[10]), .C(DEBUG_6_c_c), 
            .E(n4178), .D(num_lines_clocked_out_10__N_368[10]), .R(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_LUT4 empty_o_I_0_1_lut (.I0(DEBUG_5_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(empty_o_N_599));   // src/fifo_dc_32_lut_gen.v(241[40:50])
    defparam empty_o_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_40_i3_3_lut_4_lut (.I0(state_timeout_counter[2]), .I1(n4), 
            .I2(n7), .I3(DEBUG_5_c), .O(n4403));
    defparam mux_40_i3_3_lut_4_lut.LUT_INIT = 16'h6f60;
    SB_DFFNESR num_lines_clocked_out_i0 (.Q(num_lines_clocked_out[0]), .C(DEBUG_6_c_c), 
            .E(n4178), .D(num_lines_clocked_out_10__N_368[0]), .R(reset_per_frame_latched));   // src/usb3_if.v(72[8] 146[4])
    SB_LUT4 i11082_3_lut (.I0(FT_OE_c), .I1(DEBUG_2_c_c), .I2(DEBUG_3_c), 
            .I3(GND_net), .O(\afull_flag_impl.af_flag_p_w_N_603[3] ));
    defparam i11082_3_lut.LUT_INIT = 16'h0101;
    SB_DFFN dc32_fifo_data_in_i15 (.Q(\dc32_fifo_data_in[14] ), .C(DEBUG_6_c_c), 
            .D(usb3_data_in_latched[14]));   // src/usb3_if.v(159[8] 161[4])
    SB_LUT4 i3_4_lut (.I0(state_timeout_counter[0]), .I1(state_timeout_counter[2]), 
            .I2(state_timeout_counter[1]), .I3(state_timeout_counter[3]), 
            .O(n7));   // src/usb3_if.v(127[21:49])
    defparam i3_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut (.I0(num_lines_clocked_out[7]), .I1(num_lines_clocked_out[2]), 
            .I2(num_lines_clocked_out[9]), .I3(num_lines_clocked_out[0]), 
            .O(n18));   // src/usb3_if.v(130[29:57])
    defparam i7_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i5_2_lut (.I0(num_lines_clocked_out[1]), .I1(num_lines_clocked_out[5]), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // src/usb3_if.v(130[29:57])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut (.I0(num_lines_clocked_out[6]), .I1(n18), .I2(num_lines_clocked_out[3]), 
            .I3(num_lines_clocked_out[10]), .O(n20));   // src/usb3_if.v(130[29:57])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(num_lines_clocked_out[4]), .I1(n20), .I2(n16), 
            .I3(num_lines_clocked_out[8]), .O(n21));   // src/usb3_if.v(130[29:57])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6182_2_lut (.I0(DEBUG_2_c_c), .I1(DEBUG_9_c), .I2(GND_net), 
            .I3(GND_net), .O(n7360));
    defparam i6182_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10966_2_lut (.I0(n547[1]), .I1(n547[2]), .I2(GND_net), .I3(GND_net), 
            .O(n12582));   // src/usb3_if.v(80[9] 144[16])
    defparam i10966_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(reset_per_frame_latched), .I1(n12582), .I2(n7360), 
            .I3(n547[5]), .O(n4061));   // src/usb3_if.v(164[8] 173[4])
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 sub_113_add_2_12_lut (.I0(GND_net), .I1(num_lines_clocked_out[10]), 
            .I2(VCC_net), .I3(n10669), .O(num_lines_clocked_out_10__N_368[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_113_add_2_11_lut (.I0(GND_net), .I1(num_lines_clocked_out[9]), 
            .I2(VCC_net), .I3(n10668), .O(num_lines_clocked_out_10__N_368[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_40_i1_4_lut (.I0(n21), .I1(state_timeout_counter[0]), .I2(n7), 
            .I3(DEBUG_5_c), .O(n134[0]));   // src/usb3_if.v(127[17] 142[20])
    defparam mux_40_i1_4_lut.LUT_INIT = 16'h3530;
    SB_CARRY sub_113_add_2_11 (.CI(n10668), .I0(num_lines_clocked_out[9]), 
            .I1(VCC_net), .CO(n10669));
    SB_LUT4 sub_113_add_2_10_lut (.I0(GND_net), .I1(num_lines_clocked_out[8]), 
            .I2(VCC_net), .I3(n10667), .O(num_lines_clocked_out_10__N_368[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_10 (.CI(n10667), .I0(num_lines_clocked_out[8]), 
            .I1(VCC_net), .CO(n10668));
    SB_LUT4 i1555_4_lut (.I0(state_timeout_counter[0]), .I1(n134[0]), .I2(n547[2]), 
            .I3(n2798), .O(n2739));   // src/usb3_if.v(80[9] 144[16])
    defparam i1555_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i1556_3_lut (.I0(n2739), .I1(DEBUG_9_c), .I2(n547[5]), .I3(GND_net), 
            .O(state_timeout_counter_3__N_379[0]));   // src/usb3_if.v(80[9] 144[16])
    defparam i1556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_113_add_2_9_lut (.I0(GND_net), .I1(num_lines_clocked_out[7]), 
            .I2(VCC_net), .I3(n10666), .O(num_lines_clocked_out_10__N_368[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_113_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_113_add_2_9 (.CI(n10666), .I0(num_lines_clocked_out[7]), 
            .I1(VCC_net), .CO(n10667));
    SB_LUT4 i1570_4_lut (.I0(n547[2]), .I1(DEBUG_9_c), .I2(n534), .I3(n547[5]), 
            .O(n2754));   // src/usb3_if.v(80[9] 144[16])
    defparam i1570_4_lut.LUT_INIT = 16'heca0;
    SB_LUT4 i3_4_lut_adj_16 (.I0(n5), .I1(n21), .I2(n10746), .I3(n3973), 
            .O(n14425));   // src/usb3_if.v(80[9] 144[16])
    defparam i3_4_lut_adj_16.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_17 (.I0(n2755), .I1(DEBUG_2_c_c), .I2(DEBUG_9_c), 
            .I3(n547[5]), .O(n5));   // src/usb3_if.v(80[9] 144[16])
    defparam i1_4_lut_adj_17.LUT_INIT = 16'haeaa;
    SB_LUT4 i3_4_lut_adj_18 (.I0(DEBUG_2_c_c), .I1(DEBUG_5_c), .I2(buffer_switch_done_latched), 
            .I3(n547[0]), .O(n10746));   // src/usb3_if.v(80[9] 144[16])
    defparam i3_4_lut_adj_18.LUT_INIT = 16'h4000;
    SB_LUT4 i1571_3_lut_4_lut (.I0(n547[1]), .I1(n7), .I2(DEBUG_2_c_c), 
            .I3(DEBUG_9_c), .O(n2755));   // src/usb3_if.v(80[9] 144[16])
    defparam i1571_3_lut_4_lut.LUT_INIT = 16'haaa8;
    SB_LUT4 i163_2_lut_2_lut (.I0(n7), .I1(DEBUG_5_c), .I2(GND_net), .I3(GND_net), 
            .O(n534));   // src/usb3_if.v(139[26] 141[24])
    defparam i163_2_lut_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut_4_lut (.I0(DEBUG_2_c_c), .I1(DEBUG_9_c), .I2(n7), 
            .I3(n547[1]), .O(n10750));   // src/usb3_if.v(80[9] 144[16])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_3_lut_4_lut (.I0(n547[5]), .I1(n547[4]), .I2(DEBUG_2_c_c), 
            .I3(DEBUG_9_c), .O(n2744));   // src/usb3_if.v(80[9] 144[16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hccce;
    SB_LUT4 i1_2_lut_3_lut_3_lut_4_lut (.I0(n547[5]), .I1(n547[4]), .I2(DEBUG_2_c_c), 
            .I3(DEBUG_9_c), .O(FT_RD_N_387));
    defparam i1_2_lut_3_lut_3_lut_4_lut.LUT_INIT = 16'hbbb1;
    SB_LUT4 i1_2_lut_adj_19 (.I0(reset_per_frame_latched), .I1(DEBUG_1_c_0_c), 
            .I2(GND_net), .I3(GND_net), .O(n4650));   // src/usb3_if.v(164[8] 173[4])
    defparam i1_2_lut_adj_19.LUT_INIT = 16'h4444;
    SB_LUT4 i1612_2_lut_3_lut_4_lut (.I0(DEBUG_2_c_c), .I1(DEBUG_9_c), .I2(n7), 
            .I3(n547[1]), .O(n2798));   // src/usb3_if.v(93[17] 100[20])
    defparam i1612_2_lut_3_lut_4_lut.LUT_INIT = 16'hf100;
    SB_LUT4 i2_3_lut_4_lut_adj_20 (.I0(n547[5]), .I1(DEBUG_2_c_c), .I2(DEBUG_9_c), 
            .I3(reset_per_frame_latched), .O(n10751));   // src/usb3_if.v(164[8] 173[4])
    defparam i2_3_lut_4_lut_adj_20.LUT_INIT = 16'h00a8;
    SB_LUT4 i1_3_lut_4_lut_adj_21 (.I0(state_timeout_counter[3]), .I1(state_timeout_counter[2]), 
            .I2(state_timeout_counter[1]), .I3(state_timeout_counter[0]), 
            .O(n3686));
    defparam i1_3_lut_4_lut_adj_21.LUT_INIT = 16'h5556;
    SB_LUT4 mux_40_i2_3_lut_4_lut (.I0(DEBUG_5_c), .I1(state_timeout_counter[1]), 
            .I2(state_timeout_counter[0]), .I3(n7), .O(n134[1]));   // src/usb3_if.v(127[17] 142[20])
    defparam mux_40_i2_3_lut_4_lut.LUT_INIT = 16'hc3aa;
    
endmodule

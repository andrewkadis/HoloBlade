-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Feb 27 2020 21:49:46

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    SOUT : in std_logic;
    SCK : out std_logic;
    FIFO_D31 : out std_logic;
    FIFO_D20 : out std_logic;
    FIFO_D13 : out std_logic;
    FIFO_D1 : out std_logic;
    FIFO_CLK : in std_logic;
    FIFO_BE2 : out std_logic;
    DATA15 : out std_logic;
    DATA4 : out std_logic;
    DATA23 : out std_logic;
    RST : out std_logic;
    FIFO_D4 : out std_logic;
    FIFO_D14 : out std_logic;
    UART_TX : out std_logic;
    DATA10 : out std_logic;
    DATA28 : out std_logic;
    DATA19 : out std_logic;
    SDAT : out std_logic;
    FT_SIWU : out std_logic;
    DATA0 : out std_logic;
    FT_WR : out std_logic;
    FIFO_D27 : out std_logic;
    FIFO_D10 : out std_logic;
    FIFO_D0 : in std_logic;
    FIFO_BE3 : out std_logic;
    DEBUG_0 : out std_logic;
    FIFO_D9 : out std_logic;
    DATA14 : out std_logic;
    UPDATE : out std_logic;
    RESET : out std_logic;
    FIFO_D21 : out std_logic;
    FIFO_D12 : out std_logic;
    FIFO_BE1 : out std_logic;
    DEBUG_6 : out std_logic;
    DATA5 : out std_logic;
    DATA24 : out std_logic;
    SEN : out std_logic;
    FIFO_D7 : out std_logic;
    FIFO_D15 : out std_logic;
    ICE_CREST : out std_logic;
    FIFO_D23 : out std_logic;
    DATA3 : out std_logic;
    DATA22 : out std_logic;
    DATA13 : out std_logic;
    INVERT : out std_logic;
    FT_RD : out std_logic;
    FIFO_D5 : out std_logic;
    FIFO_D24 : out std_logic;
    FIFO_D17 : out std_logic;
    DSR : out std_logic;
    DEBUG_3 : out std_logic;
    DATA29 : out std_logic;
    DATA18 : out std_logic;
    ICE_SYSCLK : in std_logic;
    ICE_CLK : out std_logic;
    DATA20 : out std_logic;
    DATA11 : out std_logic;
    DATA1 : out std_logic;
    VALID : out std_logic;
    SYNC : out std_logic;
    FIFO_D3 : out std_logic;
    FIFO_D26 : out std_logic;
    FIFO_D11 : out std_logic;
    DEBUG_1 : out std_logic;
    DATA8 : out std_logic;
    DATA31 : out std_logic;
    DATA27 : out std_logic;
    CTS : out std_logic;
    FIFO_D8 : out std_logic;
    FIFO_D18 : out std_logic;
    DEBUG_8 : out std_logic;
    DCD : out std_logic;
    DATA17 : out std_logic;
    SLM_CLK : out std_logic;
    DATA6 : out std_logic;
    DATA25 : out std_logic;
    ICE_CDONE : out std_logic;
    FIFO_D6 : out std_logic;
    FIFO_D29 : out std_logic;
    UART_RX : in std_logic;
    FIFO_D22 : out std_logic;
    FIFO_BE0 : out std_logic;
    DEBUG_5 : out std_logic;
    DATA12 : out std_logic;
    DTR : out std_logic;
    DATA21 : out std_logic;
    DATA2 : out std_logic;
    FIFO_D25 : out std_logic;
    FIFO_D2 : out std_logic;
    FIFO_D16 : out std_logic;
    DEBUG_2 : out std_logic;
    DATA9 : out std_logic;
    DATA30 : out std_logic;
    FT_TXE : in std_logic;
    FR_RXF : in std_logic;
    FIFO_D19 : out std_logic;
    DEBUG_9 : out std_logic;
    DATA16 : out std_logic;
    FT_OE : out std_logic;
    DATA7 : out std_logic;
    DATA26 : out std_logic;
    FIFO_D30 : out std_logic;
    FIFO_D28 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__13548\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \DEBUG_8_c_c\ : std_logic;
signal \ICE_SYSCLK_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DEBUG_9_c_c\ : std_logic;
signal \FT_OE_c\ : std_logic;
signal \FIFO_CLK_c\ : std_logic;
signal pll_clk_unbuf : std_logic;
signal \GB_BUFFER_pll_clk_unbuf_THRU_CO\ : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal fifo_temp_output_2 : std_logic;
signal \RESET_c\ : std_logic;
signal \n1819_cascade_\ : std_logic;
signal n1898 : std_logic;
signal \n1898_cascade_\ : std_logic;
signal n1819 : std_logic;
signal \pc_tx.n2550\ : std_logic;
signal \pc_tx.n2550_cascade_\ : std_logic;
signal \pc_tx.n1484\ : std_logic;
signal \pc_tx.r_Bit_Index_1\ : std_logic;
signal \pc_tx.r_Bit_Index_2\ : std_logic;
signal \pc_tx.n3385_cascade_\ : std_logic;
signal \pc_tx.n3323\ : std_logic;
signal \pc_tx.n3322\ : std_logic;
signal fifo_temp_output_0 : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal \mem_LUT_data_raw_r_2\ : std_logic;
signal \mem_LUT_mem_1_6\ : std_logic;
signal fifo_temp_output_3 : std_logic;
signal fifo_temp_output_4 : std_logic;
signal fifo_temp_output_5 : std_logic;
signal \mem_LUT_data_raw_r_6\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal \pc_tx.n3319\ : std_logic;
signal \reset_all_w_N_61_cascade_\ : std_logic;
signal \n2_adj_505_cascade_\ : std_logic;
signal \reset_all_w_N_61\ : std_logic;
signal reset_clk_counter_2 : std_logic;
signal reset_clk_counter_3 : std_logic;
signal reset_clk_counter_1 : std_logic;
signal reset_clk_counter_0 : std_logic;
signal \n4_cascade_\ : std_logic;
signal tx_uart_active_flag : std_logic;
signal \r_SM_Main_2_N_187_0\ : std_logic;
signal \pc_tx.o_Tx_Serial_N_216\ : std_logic;
signal \pc_tx.n3\ : std_logic;
signal \mem_LUT_data_raw_r_0\ : std_logic;
signal \mem_LUT_data_raw_r_5\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3397\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6\ : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal \mem_LUT_mem_1_0\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6\ : std_logic;
signal rd_fifo_en_prev_r : std_logic;
signal \n1795_cascade_\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3433\ : std_logic;
signal \mem_LUT_data_raw_r_4\ : std_logic;
signal fifo_temp_output_7 : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3403\ : std_logic;
signal \n32_cascade_\ : std_logic;
signal \n24_adj_510_cascade_\ : std_logic;
signal \mem_LUT_mem_3_4\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4\ : std_logic;
signal is_fifo_empty_flag : std_logic;
signal n4_adj_511 : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3409\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n4_cascade_\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0\ : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \r_Bit_Index_0_adj_498\ : std_logic;
signal \pc_tx.n3320\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5\ : std_logic;
signal \mem_LUT_mem_3_5\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3\ : std_logic;
signal \mem_LUT_mem_3_7\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2\ : std_logic;
signal fifo_temp_output_6 : std_logic;
signal n1636 : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2\ : std_logic;
signal \mem_LUT_mem_3_2\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3415\ : std_logic;
signal \mem_LUT_data_raw_r_7\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3391\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3\ : std_logic;
signal \mem_LUT_data_raw_r_3\ : std_logic;
signal \SDAT_c\ : std_logic;
signal \INVspi0.tx_shift_reg_i15C_net\ : std_logic;
signal \rd_addr_p1_w_2_cascade_\ : std_logic;
signal rd_fifo_en_w : std_logic;
signal \n3448_cascade_\ : std_logic;
signal rd_addr_p1_w_2 : std_logic;
signal n3289 : std_logic;
signal \mem_LUT_mem_3_1\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3427\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1\ : std_logic;
signal \mem_LUT_mem_1_1\ : std_logic;
signal \mem_LUT_mem_1_5\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n4\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7\ : std_logic;
signal n1795 : std_logic;
signal \mem_LUT_data_raw_r_1\ : std_logic;
signal fifo_temp_output_1 : std_logic;
signal \mem_LUT_mem_3_6\ : std_logic;
signal \mem_LUT_mem_3_3\ : std_logic;
signal \mem_LUT_mem_1_2\ : std_logic;
signal tx_addr_byte_7 : std_logic;
signal \mem_LUT_mem_1_3\ : std_logic;
signal \mem_LUT_mem_1_4\ : std_logic;
signal tx_addr_byte_4 : std_logic;
signal \spi0.n3176\ : std_logic;
signal tx_data_byte_3 : std_logic;
signal tx_addr_byte_3 : std_logic;
signal tx_shift_reg_11 : std_logic;
signal tx_shift_reg_10 : std_logic;
signal \INVspi0.tx_shift_reg_i12C_net\ : std_logic;
signal \r_SM_Main_0_adj_497\ : std_logic;
signal \r_SM_Main_1_adj_496\ : std_logic;
signal \r_SM_Main_2_adj_495\ : std_logic;
signal n2 : std_logic;
signal \n2_cascade_\ : std_logic;
signal \pc_tx.n2981_cascade_\ : std_logic;
signal \pc_tx.n2564_cascade_\ : std_logic;
signal \r_SM_Main_2_N_184_1\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0\ : std_logic;
signal \mem_LUT_mem_3_0\ : std_logic;
signal \tx_fifo.lscc_fifo_inst.n3421\ : std_logic;
signal \pc_tx.r_Clock_Count_0\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \pc_tx.r_Clock_Count_1\ : std_logic;
signal \pc_tx.n2929\ : std_logic;
signal \pc_tx.r_Clock_Count_2\ : std_logic;
signal \pc_tx.n2930\ : std_logic;
signal \pc_tx.r_Clock_Count_3\ : std_logic;
signal \pc_tx.n2931\ : std_logic;
signal \pc_tx.r_Clock_Count_4\ : std_logic;
signal \pc_tx.n2932\ : std_logic;
signal \pc_tx.r_Clock_Count_5\ : std_logic;
signal \pc_tx.n2933\ : std_logic;
signal \pc_tx.r_Clock_Count_6\ : std_logic;
signal \pc_tx.n2934\ : std_logic;
signal \pc_tx.r_Clock_Count_7\ : std_logic;
signal \pc_tx.n2935\ : std_logic;
signal \pc_tx.n2936\ : std_logic;
signal \pc_tx.r_Clock_Count_8\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \pc_tx.n2937\ : std_logic;
signal \pc_tx.r_Clock_Count_9\ : std_logic;
signal \pc_tx.n1\ : std_logic;
signal \pc_tx.n1919\ : std_logic;
signal n4_adj_494 : std_logic;
signal \mem_LUT_mem_1_7\ : std_logic;
signal \n3279_cascade_\ : std_logic;
signal \spi0.tx_shift_reg_14\ : std_logic;
signal tx_shift_reg_12 : std_logic;
signal tx_shift_reg_13 : std_logic;
signal \INVspi0.tx_shift_reg_i14C_net\ : std_logic;
signal tx_shift_reg_3 : std_logic;
signal tx_shift_reg_1 : std_logic;
signal tx_shift_reg_2 : std_logic;
signal tx_shift_reg_4 : std_logic;
signal \n1728_cascade_\ : std_logic;
signal tx_shift_reg_5 : std_logic;
signal tx_addr_byte_0 : std_logic;
signal tx_shift_reg_6 : std_logic;
signal tx_shift_reg_7 : std_logic;
signal n1728 : std_logic;
signal tx_shift_reg_8 : std_logic;
signal tx_shift_reg_9 : std_logic;
signal \INVspi0.tx_shift_reg_i6C_net\ : std_logic;
signal \DEBUG_5_c_c\ : std_logic;
signal rx_shift_reg_0 : std_logic;
signal \tx_fifo.lscc_fifo_inst.n2_cascade_\ : std_logic;
signal rd_addr_r_2 : std_logic;
signal wr_addr_p1_w_2 : std_logic;
signal \wr_addr_p1_w_2_cascade_\ : std_logic;
signal wr_addr_r_2 : std_logic;
signal rd_addr_r_0 : std_logic;
signal n1 : std_logic;
signal fifo_read_cmd : std_logic;
signal \n1_cascade_\ : std_logic;
signal rd_addr_r_1 : std_logic;
signal \n3275_cascade_\ : std_logic;
signal n2968 : std_logic;
signal \n15_adj_509_cascade_\ : std_logic;
signal is_tx_fifo_full_flag : std_logic;
signal fifo_write_cmd : std_logic;
signal wr_fifo_en_w : std_logic;
signal \wr_fifo_en_w_cascade_\ : std_logic;
signal wr_addr_r_0 : std_logic;
signal wr_addr_r_1 : std_logic;
signal tx_addr_byte_6 : std_logic;
signal tx_shift_reg_0 : std_logic;
signal \INVspi0.tx_shift_reg_i0C_net\ : std_logic;
signal \spi0.n890\ : std_logic;
signal \spi0.n3328_cascade_\ : std_logic;
signal \spi0.n1429_cascade_\ : std_logic;
signal \spi0.n3328\ : std_logic;
signal \spi0.n497\ : std_logic;
signal \spi0.n498\ : std_logic;
signal \n883_cascade_\ : std_logic;
signal \spi0.n2433\ : std_logic;
signal \spi0.n3337_cascade_\ : std_logic;
signal \spi0.n13\ : std_logic;
signal \spi0.n1429\ : std_logic;
signal \spi0.n13_cascade_\ : std_logic;
signal \spi0.state_next_2\ : std_logic;
signal \spi0.state_next_0_cascade_\ : std_logic;
signal \spi0.n4_cascade_\ : std_logic;
signal \spi0.CS_w\ : std_logic;
signal spi_busy_prev : std_logic;
signal spi_busy_falling_edge : std_logic;
signal tx_data_byte_0 : std_logic;
signal tx_addr_byte_5 : std_logic;
signal \spi0.n502\ : std_logic;
signal \spi0.state_next_2__N_311\ : std_logic;
signal \spi0.n487\ : std_logic;
signal \spi0.n488\ : std_logic;
signal \spi0.n489\ : std_logic;
signal \spi0.n490\ : std_logic;
signal \spi0.n491\ : std_logic;
signal rx_shift_reg_1 : std_logic;
signal \rx_shift_reg_15__N_319_cascade_\ : std_logic;
signal rx_buf_byte_0 : std_logic;
signal rx_buf_byte_1 : std_logic;
signal spi_busy : std_logic;
signal rx_buf_byte_6 : std_logic;
signal rx_buf_byte_3 : std_logic;
signal \spi0.n906\ : std_logic;
signal n883 : std_logic;
signal \spi0.n906_cascade_\ : std_logic;
signal \spi0.n492\ : std_logic;
signal \spi0.n493\ : std_logic;
signal \spi0.n494\ : std_logic;
signal \state_next_2__N_312\ : std_logic;
signal \spi0.n495\ : std_logic;
signal \spi0.state_next_2__N_310\ : std_logic;
signal \spi0.n4\ : std_logic;
signal \spi0.state_next_1\ : std_logic;
signal \spi0.n499\ : std_logic;
signal reset_all_w : std_logic;
signal state_reg_0 : std_logic;
signal state_reg_2 : std_logic;
signal state_reg_1 : std_logic;
signal \SEN_c\ : std_logic;
signal \DEBUG_6_c\ : std_logic;
signal tx_data_byte_4 : std_logic;
signal tx_data_byte_6 : std_logic;
signal start_transfer_prev : std_logic;
signal n5_adj_507 : std_logic;
signal start_transfer_edge : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \spi0.n2915\ : std_logic;
signal \spi0.n2916\ : std_logic;
signal \spi0.n2917\ : std_logic;
signal \spi0.n2918\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \spi0.n2919\ : std_logic;
signal \spi0.spi_clk_counter_1\ : std_logic;
signal \spi0.spi_clk_counter_5\ : std_logic;
signal \spi0.spi_clk_counter_0\ : std_logic;
signal \spi0.spi_clk_counter_2\ : std_logic;
signal \spi0.spi_clk_counter_3\ : std_logic;
signal \spi0.n10_cascade_\ : std_logic;
signal \spi0.spi_clk_counter_4\ : std_logic;
signal \spi0.n1896\ : std_logic;
signal tx_data_byte_1 : std_logic;
signal tx_addr_byte_1 : std_logic;
signal rx_shift_reg_2 : std_logic;
signal rx_buf_byte_7 : std_logic;
signal rx_buf_byte_4 : std_logic;
signal rx_buf_byte_2 : std_logic;
signal \rx_shift_reg_15__N_319\ : std_logic;
signal rx_buf_byte_5 : std_logic;
signal rx_shift_reg_3 : std_logic;
signal rx_shift_reg_4 : std_logic;
signal rx_shift_reg_7 : std_logic;
signal rx_shift_reg_8 : std_logic;
signal rx_shift_reg_5 : std_logic;
signal n3279 : std_logic;
signal rx_shift_reg_6 : std_logic;
signal \spi0.spi_clk\ : std_logic;
signal \pc_rx.n3291_cascade_\ : std_logic;
signal \pc_rx.n6\ : std_logic;
signal \pc_rx.n3260\ : std_logic;
signal \pc_rx.n3261_cascade_\ : std_logic;
signal \pc_rx.n2558_cascade_\ : std_logic;
signal \pc_rx.r_Clock_Count_0\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \pc_rx.r_Clock_Count_1\ : std_logic;
signal \pc_rx.n2920\ : std_logic;
signal \pc_rx.r_Clock_Count_2\ : std_logic;
signal \pc_rx.n2921\ : std_logic;
signal \pc_rx.r_Clock_Count_3\ : std_logic;
signal \pc_rx.n2922\ : std_logic;
signal \pc_rx.r_Clock_Count_4\ : std_logic;
signal \pc_rx.n2923\ : std_logic;
signal \pc_rx.r_Clock_Count_5\ : std_logic;
signal \pc_rx.n2924\ : std_logic;
signal \pc_rx.r_Clock_Count_6\ : std_logic;
signal \pc_rx.n2925\ : std_logic;
signal \pc_rx.r_Clock_Count_7\ : std_logic;
signal \pc_rx.n2926\ : std_logic;
signal \pc_rx.n2927\ : std_logic;
signal \pc_rx.r_Clock_Count_8\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \pc_rx.n2928\ : std_logic;
signal \pc_rx.r_Clock_Count_9\ : std_logic;
signal tx_data_byte_5 : std_logic;
signal tx_addr_byte_2 : std_logic;
signal tx_data_byte_2 : std_logic;
signal uart_rx_complete_prev : std_logic;
signal \n1764_cascade_\ : std_logic;
signal \DEBUG_1_c\ : std_logic;
signal \pc_rx.n3273_cascade_\ : std_logic;
signal \pc_rx.n1910\ : std_logic;
signal \pc_rx.n6_adj_492_cascade_\ : std_logic;
signal \pc_rx.n1815\ : std_logic;
signal \n1747_cascade_\ : std_logic;
signal pc_data_rx_6 : std_logic;
signal \n1754_cascade_\ : std_logic;
signal pc_data_rx_3 : std_logic;
signal n1747 : std_logic;
signal pc_data_rx_7 : std_logic;
signal tx_data_byte_7 : std_logic;
signal \pc_rx.n3271\ : std_logic;
signal \pc_rx.r_SM_Main_2_N_114_0\ : std_logic;
signal \pc_rx.n1_cascade_\ : std_logic;
signal \pc_rx.n2578\ : std_logic;
signal \pc_rx.n1715\ : std_logic;
signal n4_adj_504 : std_logic;
signal \n4_adj_504_cascade_\ : std_logic;
signal pc_data_rx_2 : std_logic;
signal \pc_rx.n3334_cascade_\ : std_logic;
signal \pc_rx.n1900\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal \r_SM_Main_2_N_108_2\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal n3293 : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \n3293_cascade_\ : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal n2540 : std_logic;
signal pc_data_rx_4 : std_logic;
signal n1750 : std_logic;
signal pc_data_rx_0 : std_logic;
signal n4_adj_506 : std_logic;
signal \n4_adj_506_cascade_\ : std_logic;
signal pc_data_rx_5 : std_logic;
signal \pc_rx.r_Bit_Index_2\ : std_logic;
signal \pc_rx.r_Bit_Index_1\ : std_logic;
signal n4_adj_500 : std_logic;
signal \n4_adj_500_cascade_\ : std_logic;
signal n1754 : std_logic;
signal pc_data_rx_1 : std_logic;
signal \r_Rx_Data\ : std_logic;
signal \DEBUG_2_c\ : std_logic;
signal uart_rx_complete_rising_edge : std_logic;
signal even_byte_flag : std_logic;
signal \UART_RX_c\ : std_logic;
signal \pc_rx.r_Rx_Data_R\ : std_logic;
signal n25 : std_logic;
signal \bfn_24_6_0_\ : std_logic;
signal n24 : std_logic;
signal n2938 : std_logic;
signal n23 : std_logic;
signal n2939 : std_logic;
signal n22 : std_logic;
signal n2940 : std_logic;
signal n21 : std_logic;
signal n2941 : std_logic;
signal n20 : std_logic;
signal n2942 : std_logic;
signal n19 : std_logic;
signal n2943 : std_logic;
signal n18 : std_logic;
signal n2944 : std_logic;
signal n2945 : std_logic;
signal n17 : std_logic;
signal \bfn_24_7_0_\ : std_logic;
signal n16 : std_logic;
signal n2946 : std_logic;
signal n15 : std_logic;
signal n2947 : std_logic;
signal n14 : std_logic;
signal n2948 : std_logic;
signal n13 : std_logic;
signal n2949 : std_logic;
signal n12 : std_logic;
signal n2950 : std_logic;
signal n11 : std_logic;
signal n2951 : std_logic;
signal n10 : std_logic;
signal n2952 : std_logic;
signal n2953 : std_logic;
signal n9 : std_logic;
signal \bfn_24_8_0_\ : std_logic;
signal n8_adj_501 : std_logic;
signal n2954 : std_logic;
signal n7 : std_logic;
signal n2955 : std_logic;
signal n6 : std_logic;
signal n2956 : std_logic;
signal n5 : std_logic;
signal n2957 : std_logic;
signal n4_adj_502 : std_logic;
signal n2958 : std_logic;
signal n3 : std_logic;
signal n2959 : std_logic;
signal n2_adj_503 : std_logic;
signal n2960 : std_logic;
signal n2961 : std_logic;
signal \bfn_24_9_0_\ : std_logic;
signal \DEBUG_0_c_24\ : std_logic;
signal \SLM_CLK_c\ : std_logic;
signal \GB_BUFFER_SLM_CLK_c_THRU_CO\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \FIFO_CLK_wire\ : std_logic;
signal \FIFO_BE1_wire\ : std_logic;
signal \VALID_wire\ : std_logic;
signal \FIFO_D14_wire\ : std_logic;
signal \DATA30_wire\ : std_logic;
signal \DEBUG_9_wire\ : std_logic;
signal \FIFO_D8_wire\ : std_logic;
signal \DATA7_wire\ : std_logic;
signal \DEBUG_1_wire\ : std_logic;
signal \DATA4_wire\ : std_logic;
signal \FIFO_D26_wire\ : std_logic;
signal \DATA24_wire\ : std_logic;
signal \DTR_wire\ : std_logic;
signal \DATA29_wire\ : std_logic;
signal \FIFO_D16_wire\ : std_logic;
signal \FT_SIWU_wire\ : std_logic;
signal \DEBUG_6_wire\ : std_logic;
signal \DATA17_wire\ : std_logic;
signal \DATA21_wire\ : std_logic;
signal \SYNC_wire\ : std_logic;
signal \SCK_wire\ : std_logic;
signal \UPDATE_wire\ : std_logic;
signal \DATA3_wire\ : std_logic;
signal \DATA18_wire\ : std_logic;
signal \DATA25_wire\ : std_logic;
signal \DEBUG_5_wire\ : std_logic;
signal \RESET_wire\ : std_logic;
signal \DATA22_wire\ : std_logic;
signal \DSR_wire\ : std_logic;
signal \FT_WR_wire\ : std_logic;
signal \DATA12_wire\ : std_logic;
signal \FIFO_D31_wire\ : std_logic;
signal \DATA11_wire\ : std_logic;
signal \DATA26_wire\ : std_logic;
signal \FT_RD_wire\ : std_logic;
signal \DATA1_wire\ : std_logic;
signal \DATA31_wire\ : std_logic;
signal \FIFO_D10_wire\ : std_logic;
signal \DATA5_wire\ : std_logic;
signal \INVERT_wire\ : std_logic;
signal \FIFO_D13_wire\ : std_logic;
signal \ICE_CREST_wire\ : std_logic;
signal \DEBUG_3_wire\ : std_logic;
signal \FIFO_D17_wire\ : std_logic;
signal \DATA8_wire\ : std_logic;
signal \FIFO_D27_wire\ : std_logic;
signal \FIFO_D1_wire\ : std_logic;
signal \DATA15_wire\ : std_logic;
signal \DATA20_wire\ : std_logic;
signal \SOUT_wire\ : std_logic;
signal \DATA16_wire\ : std_logic;
signal \DATA28_wire\ : std_logic;
signal \FIFO_D23_wire\ : std_logic;
signal \ICE_CLK_wire\ : std_logic;
signal \CTS_wire\ : std_logic;
signal \FR_RXF_wire\ : std_logic;
signal \SLM_CLK_wire\ : std_logic;
signal \FIFO_D20_wire\ : std_logic;
signal \FT_OE_wire\ : std_logic;
signal \FIFO_BE3_wire\ : std_logic;
signal \FIFO_D19_wire\ : std_logic;
signal \FIFO_D7_wire\ : std_logic;
signal \UART_RX_wire\ : std_logic;
signal \FIFO_D6_wire\ : std_logic;
signal \SDAT_wire\ : std_logic;
signal \FIFO_BE0_wire\ : std_logic;
signal \DATA19_wire\ : std_logic;
signal \FIFO_D28_wire\ : std_logic;
signal \DATA14_wire\ : std_logic;
signal \DATA10_wire\ : std_logic;
signal \DATA6_wire\ : std_logic;
signal \FIFO_BE2_wire\ : std_logic;
signal \FIFO_D11_wire\ : std_logic;
signal \FIFO_D3_wire\ : std_logic;
signal \RST_wire\ : std_logic;
signal \FIFO_D25_wire\ : std_logic;
signal \ICE_CDONE_wire\ : std_logic;
signal \SEN_wire\ : std_logic;
signal \DCD_wire\ : std_logic;
signal \FIFO_D9_wire\ : std_logic;
signal \DATA9_wire\ : std_logic;
signal \FIFO_D12_wire\ : std_logic;
signal \DATA27_wire\ : std_logic;
signal \DEBUG_0_wire\ : std_logic;
signal \DATA2_wire\ : std_logic;
signal \FIFO_D24_wire\ : std_logic;
signal \FIFO_D2_wire\ : std_logic;
signal \FIFO_D22_wire\ : std_logic;
signal \UART_TX_wire\ : std_logic;
signal \FIFO_D29_wire\ : std_logic;
signal \FIFO_D21_wire\ : std_logic;
signal \DEBUG_8_wire\ : std_logic;
signal \FIFO_D15_wire\ : std_logic;
signal \DEBUG_2_wire\ : std_logic;
signal \DATA13_wire\ : std_logic;
signal \FIFO_D5_wire\ : std_logic;
signal \FIFO_D4_wire\ : std_logic;
signal \FIFO_D18_wire\ : std_logic;
signal \DATA23_wire\ : std_logic;
signal \FIFO_D0_wire\ : std_logic;
signal \ICE_SYSCLK_wire\ : std_logic;
signal \FIFO_D30_wire\ : std_logic;
signal \DATA0_wire\ : std_logic;
signal \clock_inst.pll_config_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \FIFO_CLK_wire\ <= FIFO_CLK;
    FIFO_BE1 <= \FIFO_BE1_wire\;
    VALID <= \VALID_wire\;
    FIFO_D14 <= \FIFO_D14_wire\;
    DATA30 <= \DATA30_wire\;
    DEBUG_9 <= \DEBUG_9_wire\;
    FIFO_D8 <= \FIFO_D8_wire\;
    DATA7 <= \DATA7_wire\;
    DEBUG_1 <= \DEBUG_1_wire\;
    DATA4 <= \DATA4_wire\;
    FIFO_D26 <= \FIFO_D26_wire\;
    DATA24 <= \DATA24_wire\;
    DTR <= \DTR_wire\;
    DATA29 <= \DATA29_wire\;
    FIFO_D16 <= \FIFO_D16_wire\;
    FT_SIWU <= \FT_SIWU_wire\;
    DEBUG_6 <= \DEBUG_6_wire\;
    DATA17 <= \DATA17_wire\;
    DATA21 <= \DATA21_wire\;
    SYNC <= \SYNC_wire\;
    SCK <= \SCK_wire\;
    UPDATE <= \UPDATE_wire\;
    DATA3 <= \DATA3_wire\;
    DATA18 <= \DATA18_wire\;
    DATA25 <= \DATA25_wire\;
    DEBUG_5 <= \DEBUG_5_wire\;
    RESET <= \RESET_wire\;
    DATA22 <= \DATA22_wire\;
    DSR <= \DSR_wire\;
    FT_WR <= \FT_WR_wire\;
    DATA12 <= \DATA12_wire\;
    FIFO_D31 <= \FIFO_D31_wire\;
    DATA11 <= \DATA11_wire\;
    DATA26 <= \DATA26_wire\;
    FT_RD <= \FT_RD_wire\;
    DATA1 <= \DATA1_wire\;
    DATA31 <= \DATA31_wire\;
    FIFO_D10 <= \FIFO_D10_wire\;
    DATA5 <= \DATA5_wire\;
    INVERT <= \INVERT_wire\;
    FIFO_D13 <= \FIFO_D13_wire\;
    ICE_CREST <= \ICE_CREST_wire\;
    DEBUG_3 <= \DEBUG_3_wire\;
    FIFO_D17 <= \FIFO_D17_wire\;
    DATA8 <= \DATA8_wire\;
    FIFO_D27 <= \FIFO_D27_wire\;
    FIFO_D1 <= \FIFO_D1_wire\;
    DATA15 <= \DATA15_wire\;
    DATA20 <= \DATA20_wire\;
    \SOUT_wire\ <= SOUT;
    DATA16 <= \DATA16_wire\;
    DATA28 <= \DATA28_wire\;
    FIFO_D23 <= \FIFO_D23_wire\;
    ICE_CLK <= \ICE_CLK_wire\;
    CTS <= \CTS_wire\;
    \FR_RXF_wire\ <= FR_RXF;
    SLM_CLK <= \SLM_CLK_wire\;
    FIFO_D20 <= \FIFO_D20_wire\;
    FT_OE <= \FT_OE_wire\;
    FIFO_BE3 <= \FIFO_BE3_wire\;
    FIFO_D19 <= \FIFO_D19_wire\;
    FIFO_D7 <= \FIFO_D7_wire\;
    \UART_RX_wire\ <= UART_RX;
    FIFO_D6 <= \FIFO_D6_wire\;
    SDAT <= \SDAT_wire\;
    FIFO_BE0 <= \FIFO_BE0_wire\;
    DATA19 <= \DATA19_wire\;
    FIFO_D28 <= \FIFO_D28_wire\;
    DATA14 <= \DATA14_wire\;
    DATA10 <= \DATA10_wire\;
    DATA6 <= \DATA6_wire\;
    FIFO_BE2 <= \FIFO_BE2_wire\;
    FIFO_D11 <= \FIFO_D11_wire\;
    FIFO_D3 <= \FIFO_D3_wire\;
    RST <= \RST_wire\;
    FIFO_D25 <= \FIFO_D25_wire\;
    ICE_CDONE <= \ICE_CDONE_wire\;
    SEN <= \SEN_wire\;
    DCD <= \DCD_wire\;
    FIFO_D9 <= \FIFO_D9_wire\;
    DATA9 <= \DATA9_wire\;
    FIFO_D12 <= \FIFO_D12_wire\;
    DATA27 <= \DATA27_wire\;
    DEBUG_0 <= \DEBUG_0_wire\;
    DATA2 <= \DATA2_wire\;
    FIFO_D24 <= \FIFO_D24_wire\;
    FIFO_D2 <= \FIFO_D2_wire\;
    FIFO_D22 <= \FIFO_D22_wire\;
    UART_TX <= \UART_TX_wire\;
    FIFO_D29 <= \FIFO_D29_wire\;
    FIFO_D21 <= \FIFO_D21_wire\;
    DEBUG_8 <= \DEBUG_8_wire\;
    FIFO_D15 <= \FIFO_D15_wire\;
    DEBUG_2 <= \DEBUG_2_wire\;
    DATA13 <= \DATA13_wire\;
    FIFO_D5 <= \FIFO_D5_wire\;
    FIFO_D4 <= \FIFO_D4_wire\;
    FIFO_D18 <= \FIFO_D18_wire\;
    DATA23 <= \DATA23_wire\;
    \FIFO_D0_wire\ <= FIFO_D0;
    \ICE_SYSCLK_wire\ <= ICE_SYSCLK;
    FIFO_D30 <= \FIFO_D30_wire\;
    DATA0 <= \DATA0_wire\;
    \clock_inst.pll_config_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';

    \clock_inst.pll_config\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0001",
            DIVQ => "100",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__5214\,
            RESETB => \N__10186\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \clock_inst.pll_config_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => pll_clk_unbuf
        );

    \FIFO_CLK_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__13546\,
            GLOBALBUFFEROUTPUT => \FIFO_CLK_c\
        );

    \FIFO_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13548\,
            DIN => \N__13547\,
            DOUT => \N__13546\,
            PACKAGEPIN => \FIFO_CLK_wire\
        );

    \FIFO_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13548\,
            PADOUT => \N__13547\,
            PADIN => \N__13546\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_BE1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13537\,
            DIN => \N__13536\,
            DOUT => \N__13535\,
            PACKAGEPIN => \FIFO_BE1_wire\
        );

    \FIFO_BE1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13537\,
            PADOUT => \N__13536\,
            PADIN => \N__13535\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VALID_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13528\,
            DIN => \N__13527\,
            DOUT => \N__13526\,
            PACKAGEPIN => \VALID_wire\
        );

    \VALID_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13528\,
            PADOUT => \N__13527\,
            PADIN => \N__13526\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D14_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13519\,
            DIN => \N__13518\,
            DOUT => \N__13517\,
            PACKAGEPIN => \FIFO_D14_wire\
        );

    \FIFO_D14_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13519\,
            PADOUT => \N__13518\,
            PADIN => \N__13517\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA30_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13510\,
            DIN => \N__13509\,
            DOUT => \N__13508\,
            PACKAGEPIN => \DATA30_wire\
        );

    \DATA30_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13510\,
            PADOUT => \N__13509\,
            PADIN => \N__13508\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10030\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_9_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13501\,
            DIN => \N__13500\,
            DOUT => \N__13499\,
            PACKAGEPIN => \DEBUG_9_wire\
        );

    \DEBUG_9_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13501\,
            PADOUT => \N__13500\,
            PADIN => \N__13499\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5322\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13492\,
            DIN => \N__13491\,
            DOUT => \N__13490\,
            PACKAGEPIN => \FIFO_D8_wire\
        );

    \FIFO_D8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13492\,
            PADOUT => \N__13491\,
            PADIN => \N__13490\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13483\,
            DIN => \N__13482\,
            DOUT => \N__13481\,
            PACKAGEPIN => \DATA7_wire\
        );

    \DATA7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13483\,
            PADOUT => \N__13482\,
            PADIN => \N__13481\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10216\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13474\,
            DIN => \N__13473\,
            DOUT => \N__13472\,
            PACKAGEPIN => \DEBUG_1_wire\
        );

    \DEBUG_1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13474\,
            PADOUT => \N__13473\,
            PADIN => \N__13472\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11007\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA4_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13465\,
            DIN => \N__13464\,
            DOUT => \N__13463\,
            PACKAGEPIN => \DATA4_wire\
        );

    \DATA4_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13465\,
            PADOUT => \N__13464\,
            PADIN => \N__13463\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10189\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D26_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13456\,
            DIN => \N__13455\,
            DOUT => \N__13454\,
            PACKAGEPIN => \FIFO_D26_wire\
        );

    \FIFO_D26_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13456\,
            PADOUT => \N__13455\,
            PADIN => \N__13454\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA24_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13447\,
            DIN => \N__13446\,
            DOUT => \N__13445\,
            PACKAGEPIN => \DATA24_wire\
        );

    \DATA24_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13447\,
            PADOUT => \N__13446\,
            PADIN => \N__13445\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10187\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DTR_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13438\,
            DIN => \N__13437\,
            DOUT => \N__13436\,
            PACKAGEPIN => \DTR_wire\
        );

    \DTR_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13438\,
            PADOUT => \N__13437\,
            PADIN => \N__13436\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA29_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13429\,
            DIN => \N__13428\,
            DOUT => \N__13427\,
            PACKAGEPIN => \DATA29_wire\
        );

    \DATA29_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13429\,
            PADOUT => \N__13428\,
            PADIN => \N__13427\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10027\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D16_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13420\,
            DIN => \N__13419\,
            DOUT => \N__13418\,
            PACKAGEPIN => \FIFO_D16_wire\
        );

    \FIFO_D16_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13420\,
            PADOUT => \N__13419\,
            PADIN => \N__13418\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_SIWU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13411\,
            DIN => \N__13410\,
            DOUT => \N__13409\,
            PACKAGEPIN => \FT_SIWU_wire\
        );

    \FT_SIWU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13411\,
            PADOUT => \N__13410\,
            PADIN => \N__13409\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_6_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13402\,
            DIN => \N__13401\,
            DOUT => \N__13400\,
            PACKAGEPIN => \DEBUG_6_wire\
        );

    \DEBUG_6_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13402\,
            PADOUT => \N__13401\,
            PADIN => \N__13400\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9114\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA17_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13393\,
            DIN => \N__13392\,
            DOUT => \N__13391\,
            PACKAGEPIN => \DATA17_wire\
        );

    \DATA17_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13393\,
            PADOUT => \N__13392\,
            PADIN => \N__13391\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10230\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA21_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13384\,
            DIN => \N__13383\,
            DOUT => \N__13382\,
            PACKAGEPIN => \DATA21_wire\
        );

    \DATA21_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13384\,
            PADOUT => \N__13383\,
            PADIN => \N__13382\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10218\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13375\,
            DIN => \N__13374\,
            DOUT => \N__13373\,
            PACKAGEPIN => \SYNC_wire\
        );

    \SYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13375\,
            PADOUT => \N__13374\,
            PADIN => \N__13373\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13366\,
            DIN => \N__13365\,
            DOUT => \N__13364\,
            PACKAGEPIN => \SCK_wire\
        );

    \SCK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13366\,
            PADOUT => \N__13365\,
            PADIN => \N__13364\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9110\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UPDATE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13357\,
            DIN => \N__13356\,
            DOUT => \N__13355\,
            PACKAGEPIN => \UPDATE_wire\
        );

    \UPDATE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13357\,
            PADOUT => \N__13356\,
            PADIN => \N__13355\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13348\,
            DIN => \N__13347\,
            DOUT => \N__13346\,
            PACKAGEPIN => \DATA3_wire\
        );

    \DATA3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13348\,
            PADOUT => \N__13347\,
            PADIN => \N__13346\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10142\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA18_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13339\,
            DIN => \N__13338\,
            DOUT => \N__13337\,
            PACKAGEPIN => \DATA18_wire\
        );

    \DATA18_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13339\,
            PADOUT => \N__13338\,
            PADIN => \N__13337\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10229\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA25_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13330\,
            DIN => \N__13329\,
            DOUT => \N__13328\,
            PACKAGEPIN => \DATA25_wire\
        );

    \DATA25_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13330\,
            PADOUT => \N__13329\,
            PADIN => \N__13328\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10141\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_5_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13321\,
            DIN => \N__13320\,
            DOUT => \N__13319\,
            PACKAGEPIN => \DEBUG_5_wire\
        );

    \DEBUG_5_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13321\,
            PADOUT => \N__13320\,
            PADIN => \N__13319\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7575\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESET_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13312\,
            DIN => \N__13311\,
            DOUT => \N__13310\,
            PACKAGEPIN => \RESET_wire\
        );

    \RESET_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13312\,
            PADOUT => \N__13311\,
            PADIN => \N__13310\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5340\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA22_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13303\,
            DIN => \N__13302\,
            DOUT => \N__13301\,
            PACKAGEPIN => \DATA22_wire\
        );

    \DATA22_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13303\,
            PADOUT => \N__13302\,
            PADIN => \N__13301\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10217\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DSR_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13294\,
            DIN => \N__13293\,
            DOUT => \N__13292\,
            PACKAGEPIN => \DSR_wire\
        );

    \DSR_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13294\,
            PADOUT => \N__13293\,
            PADIN => \N__13292\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_WR_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13285\,
            DIN => \N__13284\,
            DOUT => \N__13283\,
            PACKAGEPIN => \FT_WR_wire\
        );

    \FT_WR_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13285\,
            PADOUT => \N__13284\,
            PADIN => \N__13283\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA12_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13276\,
            DIN => \N__13275\,
            DOUT => \N__13274\,
            PACKAGEPIN => \DATA12_wire\
        );

    \DATA12_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13276\,
            PADOUT => \N__13275\,
            PADIN => \N__13274\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10185\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D31_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13267\,
            DIN => \N__13266\,
            DOUT => \N__13265\,
            PACKAGEPIN => \FIFO_D31_wire\
        );

    \FIFO_D31_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13267\,
            PADOUT => \N__13266\,
            PADIN => \N__13265\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA11_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13258\,
            DIN => \N__13257\,
            DOUT => \N__13256\,
            PACKAGEPIN => \DATA11_wire\
        );

    \DATA11_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13258\,
            PADOUT => \N__13257\,
            PADIN => \N__13256\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10184\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA26_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13249\,
            DIN => \N__13248\,
            DOUT => \N__13247\,
            PACKAGEPIN => \DATA26_wire\
        );

    \DATA26_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13249\,
            PADOUT => \N__13248\,
            PADIN => \N__13247\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10140\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_RD_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13240\,
            DIN => \N__13239\,
            DOUT => \N__13238\,
            PACKAGEPIN => \FT_RD_wire\
        );

    \FT_RD_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13240\,
            PADOUT => \N__13239\,
            PADIN => \N__13238\,
            CLOCKENABLE => \VCCG0\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5276\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5255\
        );

    \DATA1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13231\,
            DIN => \N__13230\,
            DOUT => \N__13229\,
            PACKAGEPIN => \DATA1_wire\
        );

    \DATA1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13231\,
            PADOUT => \N__13230\,
            PADIN => \N__13229\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10028\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA31_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13222\,
            DIN => \N__13221\,
            DOUT => \N__13220\,
            PACKAGEPIN => \DATA31_wire\
        );

    \DATA31_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13222\,
            PADOUT => \N__13221\,
            PADIN => \N__13220\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10029\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D10_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13213\,
            DIN => \N__13212\,
            DOUT => \N__13211\,
            PACKAGEPIN => \FIFO_D10_wire\
        );

    \FIFO_D10_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13213\,
            PADOUT => \N__13212\,
            PADIN => \N__13211\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA5_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13204\,
            DIN => \N__13203\,
            DOUT => \N__13202\,
            PACKAGEPIN => \DATA5_wire\
        );

    \DATA5_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13204\,
            PADOUT => \N__13203\,
            PADIN => \N__13202\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10219\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \INVERT_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13195\,
            DIN => \N__13194\,
            DOUT => \N__13193\,
            PACKAGEPIN => \INVERT_wire\
        );

    \INVERT_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13195\,
            PADOUT => \N__13194\,
            PADIN => \N__13193\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D13_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13186\,
            DIN => \N__13185\,
            DOUT => \N__13184\,
            PACKAGEPIN => \FIFO_D13_wire\
        );

    \FIFO_D13_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13186\,
            PADOUT => \N__13185\,
            PADIN => \N__13184\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ICE_CREST_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13177\,
            DIN => \N__13176\,
            DOUT => \N__13175\,
            PACKAGEPIN => \ICE_CREST_wire\
        );

    \ICE_CREST_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13177\,
            PADOUT => \N__13176\,
            PADIN => \N__13175\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13168\,
            DIN => \N__13167\,
            DOUT => \N__13166\,
            PACKAGEPIN => \DEBUG_3_wire\
        );

    \DEBUG_3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13168\,
            PADOUT => \N__13167\,
            PADIN => \N__13166\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D17_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13159\,
            DIN => \N__13158\,
            DOUT => \N__13157\,
            PACKAGEPIN => \FIFO_D17_wire\
        );

    \FIFO_D17_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13159\,
            PADOUT => \N__13158\,
            PADIN => \N__13157\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13150\,
            DIN => \N__13149\,
            DOUT => \N__13148\,
            PACKAGEPIN => \DATA8_wire\
        );

    \DATA8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13150\,
            PADOUT => \N__13149\,
            PADIN => \N__13148\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10174\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D27_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13141\,
            DIN => \N__13140\,
            DOUT => \N__13139\,
            PACKAGEPIN => \FIFO_D27_wire\
        );

    \FIFO_D27_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13141\,
            PADOUT => \N__13140\,
            PADIN => \N__13139\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13132\,
            DIN => \N__13131\,
            DOUT => \N__13130\,
            PACKAGEPIN => \FIFO_D1_wire\
        );

    \FIFO_D1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13132\,
            PADOUT => \N__13131\,
            PADIN => \N__13130\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA15_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13123\,
            DIN => \N__13122\,
            DOUT => \N__13121\,
            PACKAGEPIN => \DATA15_wire\
        );

    \DATA15_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13123\,
            PADOUT => \N__13122\,
            PADIN => \N__13121\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10214\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA20_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13114\,
            DIN => \N__13113\,
            DOUT => \N__13112\,
            PACKAGEPIN => \DATA20_wire\
        );

    \DATA20_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13114\,
            PADOUT => \N__13113\,
            PADIN => \N__13112\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10220\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_5_c_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13105\,
            DIN => \N__13104\,
            DOUT => \N__13103\,
            PACKAGEPIN => \SOUT_wire\
        );

    \DEBUG_5_c_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13105\,
            PADOUT => \N__13104\,
            PADIN => \N__13103\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_5_c_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA16_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13096\,
            DIN => \N__13095\,
            DOUT => \N__13094\,
            PACKAGEPIN => \DATA16_wire\
        );

    \DATA16_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13096\,
            PADOUT => \N__13095\,
            PADIN => \N__13094\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10215\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA28_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13087\,
            DIN => \N__13086\,
            DOUT => \N__13085\,
            PACKAGEPIN => \DATA28_wire\
        );

    \DATA28_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13087\,
            PADOUT => \N__13086\,
            PADIN => \N__13085\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9980\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D23_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13078\,
            DIN => \N__13077\,
            DOUT => \N__13076\,
            PACKAGEPIN => \FIFO_D23_wire\
        );

    \FIFO_D23_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13078\,
            PADOUT => \N__13077\,
            PADIN => \N__13076\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ICE_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13069\,
            DIN => \N__13068\,
            DOUT => \N__13067\,
            PACKAGEPIN => \ICE_CLK_wire\
        );

    \ICE_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13069\,
            PADOUT => \N__13068\,
            PADIN => \N__13067\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CTS_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13060\,
            DIN => \N__13059\,
            DOUT => \N__13058\,
            PACKAGEPIN => \CTS_wire\
        );

    \CTS_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13060\,
            PADOUT => \N__13059\,
            PADIN => \N__13058\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_9_c_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13051\,
            DIN => \N__13050\,
            DOUT => \N__13049\,
            PACKAGEPIN => \FR_RXF_wire\
        );

    \DEBUG_9_c_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13051\,
            PADOUT => \N__13050\,
            PADIN => \N__13049\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_9_c_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SLM_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13042\,
            DIN => \N__13041\,
            DOUT => \N__13040\,
            PACKAGEPIN => \SLM_CLK_wire\
        );

    \SLM_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13042\,
            PADOUT => \N__13041\,
            PADIN => \N__13040\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12321\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D20_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13033\,
            DIN => \N__13032\,
            DOUT => \N__13031\,
            PACKAGEPIN => \FIFO_D20_wire\
        );

    \FIFO_D20_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13033\,
            PADOUT => \N__13032\,
            PADIN => \N__13031\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FT_OE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13024\,
            DIN => \N__13023\,
            DOUT => \N__13022\,
            PACKAGEPIN => \FT_OE_wire\
        );

    \FT_OE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13024\,
            PADOUT => \N__13023\,
            PADIN => \N__13022\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5280\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_BE3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13015\,
            DIN => \N__13014\,
            DOUT => \N__13013\,
            PACKAGEPIN => \FIFO_BE3_wire\
        );

    \FIFO_BE3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13015\,
            PADOUT => \N__13014\,
            PADIN => \N__13013\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D19_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13006\,
            DIN => \N__13005\,
            DOUT => \N__13004\,
            PACKAGEPIN => \FIFO_D19_wire\
        );

    \FIFO_D19_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13006\,
            PADOUT => \N__13005\,
            PADIN => \N__13004\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12997\,
            DIN => \N__12996\,
            DOUT => \N__12995\,
            PACKAGEPIN => \FIFO_D7_wire\
        );

    \FIFO_D7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12997\,
            PADOUT => \N__12996\,
            PADIN => \N__12995\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UART_RX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12988\,
            DIN => \N__12987\,
            DOUT => \N__12986\,
            PACKAGEPIN => \UART_RX_wire\
        );

    \UART_RX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12988\,
            PADOUT => \N__12987\,
            PADIN => \N__12986\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \UART_RX_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D6_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12979\,
            DIN => \N__12978\,
            DOUT => \N__12977\,
            PACKAGEPIN => \FIFO_D6_wire\
        );

    \FIFO_D6_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12979\,
            PADOUT => \N__12978\,
            PADIN => \N__12977\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SDAT_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12970\,
            DIN => \N__12969\,
            DOUT => \N__12968\,
            PACKAGEPIN => \SDAT_wire\
        );

    \SDAT_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12970\,
            PADOUT => \N__12969\,
            PADIN => \N__12968\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6195\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_BE0_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12961\,
            DIN => \N__12960\,
            DOUT => \N__12959\,
            PACKAGEPIN => \FIFO_BE0_wire\
        );

    \FIFO_BE0_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12961\,
            PADOUT => \N__12960\,
            PADIN => \N__12959\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA19_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12952\,
            DIN => \N__12951\,
            DOUT => \N__12950\,
            PACKAGEPIN => \DATA19_wire\
        );

    \DATA19_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12952\,
            PADOUT => \N__12951\,
            PADIN => \N__12950\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10221\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D28_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12943\,
            DIN => \N__12942\,
            DOUT => \N__12941\,
            PACKAGEPIN => \FIFO_D28_wire\
        );

    \FIFO_D28_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12943\,
            PADOUT => \N__12942\,
            PADIN => \N__12941\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA14_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12934\,
            DIN => \N__12933\,
            DOUT => \N__12932\,
            PACKAGEPIN => \DATA14_wire\
        );

    \DATA14_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12934\,
            PADOUT => \N__12933\,
            PADIN => \N__12932\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10173\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA10_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12925\,
            DIN => \N__12924\,
            DOUT => \N__12923\,
            PACKAGEPIN => \DATA10_wire\
        );

    \DATA10_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12925\,
            PADOUT => \N__12924\,
            PADIN => \N__12923\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10213\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA6_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12916\,
            DIN => \N__12915\,
            DOUT => \N__12914\,
            PACKAGEPIN => \DATA6_wire\
        );

    \DATA6_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12916\,
            PADOUT => \N__12915\,
            PADIN => \N__12914\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10222\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_BE2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12907\,
            DIN => \N__12906\,
            DOUT => \N__12905\,
            PACKAGEPIN => \FIFO_BE2_wire\
        );

    \FIFO_BE2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12907\,
            PADOUT => \N__12906\,
            PADIN => \N__12905\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D11_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12898\,
            DIN => \N__12897\,
            DOUT => \N__12896\,
            PACKAGEPIN => \FIFO_D11_wire\
        );

    \FIFO_D11_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12898\,
            PADOUT => \N__12897\,
            PADIN => \N__12896\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12889\,
            DIN => \N__12888\,
            DOUT => \N__12887\,
            PACKAGEPIN => \FIFO_D3_wire\
        );

    \FIFO_D3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12889\,
            PADOUT => \N__12888\,
            PADIN => \N__12887\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12880\,
            DIN => \N__12879\,
            DOUT => \N__12878\,
            PACKAGEPIN => \RST_wire\
        );

    \RST_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12880\,
            PADOUT => \N__12879\,
            PADIN => \N__12878\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D25_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12871\,
            DIN => \N__12870\,
            DOUT => \N__12869\,
            PACKAGEPIN => \FIFO_D25_wire\
        );

    \FIFO_D25_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12871\,
            PADOUT => \N__12870\,
            PADIN => \N__12869\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ICE_CDONE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12862\,
            DIN => \N__12861\,
            DOUT => \N__12860\,
            PACKAGEPIN => \ICE_CDONE_wire\
        );

    \ICE_CDONE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12862\,
            PADOUT => \N__12861\,
            PADIN => \N__12860\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SEN_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12853\,
            DIN => \N__12852\,
            DOUT => \N__12851\,
            PACKAGEPIN => \SEN_wire\
        );

    \SEN_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12853\,
            PADOUT => \N__12852\,
            PADIN => \N__12851\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9135\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DCD_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12844\,
            DIN => \N__12843\,
            DOUT => \N__12842\,
            PACKAGEPIN => \DCD_wire\
        );

    \DCD_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12844\,
            PADOUT => \N__12843\,
            PADIN => \N__12842\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D9_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12835\,
            DIN => \N__12834\,
            DOUT => \N__12833\,
            PACKAGEPIN => \FIFO_D9_wire\
        );

    \FIFO_D9_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12835\,
            PADOUT => \N__12834\,
            PADIN => \N__12833\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA9_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12826\,
            DIN => \N__12825\,
            DOUT => \N__12824\,
            PACKAGEPIN => \DATA9_wire\
        );

    \DATA9_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12826\,
            PADOUT => \N__12825\,
            PADIN => \N__12824\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10168\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D12_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12817\,
            DIN => \N__12816\,
            DOUT => \N__12815\,
            PACKAGEPIN => \FIFO_D12_wire\
        );

    \FIFO_D12_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12817\,
            PADOUT => \N__12816\,
            PADIN => \N__12815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA27_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12808\,
            DIN => \N__12807\,
            DOUT => \N__12806\,
            PACKAGEPIN => \DATA27_wire\
        );

    \DATA27_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12808\,
            PADOUT => \N__12807\,
            PADIN => \N__12806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10084\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_0_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12799\,
            DIN => \N__12798\,
            DOUT => \N__12797\,
            PACKAGEPIN => \DEBUG_0_wire\
        );

    \DEBUG_0_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12799\,
            PADOUT => \N__12798\,
            PADIN => \N__12797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12552\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12790\,
            DIN => \N__12789\,
            DOUT => \N__12788\,
            PACKAGEPIN => \DATA2_wire\
        );

    \DATA2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12790\,
            PADOUT => \N__12789\,
            PADIN => \N__12788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10085\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D24_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12781\,
            DIN => \N__12780\,
            DOUT => \N__12779\,
            PACKAGEPIN => \FIFO_D24_wire\
        );

    \FIFO_D24_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12781\,
            PADOUT => \N__12780\,
            PADIN => \N__12779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12772\,
            DIN => \N__12771\,
            DOUT => \N__12770\,
            PACKAGEPIN => \FIFO_D2_wire\
        );

    \FIFO_D2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12772\,
            PADOUT => \N__12771\,
            PADIN => \N__12770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D22_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12763\,
            DIN => \N__12762\,
            DOUT => \N__12761\,
            PACKAGEPIN => \FIFO_D22_wire\
        );

    \FIFO_D22_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12763\,
            PADOUT => \N__12762\,
            PADIN => \N__12761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UART_TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12754\,
            DIN => \N__12753\,
            DOUT => \N__12752\,
            PACKAGEPIN => \UART_TX_wire\
        );

    \UART_TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12754\,
            PADOUT => \N__12753\,
            PADIN => \N__12752\,
            CLOCKENABLE => \N__7314\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5730\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__12524\
        );

    \FIFO_D29_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12745\,
            DIN => \N__12744\,
            DOUT => \N__12743\,
            PACKAGEPIN => \FIFO_D29_wire\
        );

    \FIFO_D29_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12745\,
            PADOUT => \N__12744\,
            PADIN => \N__12743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D21_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12736\,
            DIN => \N__12735\,
            DOUT => \N__12734\,
            PACKAGEPIN => \FIFO_D21_wire\
        );

    \FIFO_D21_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12736\,
            PADOUT => \N__12735\,
            PADIN => \N__12734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12727\,
            DIN => \N__12726\,
            DOUT => \N__12725\,
            PACKAGEPIN => \DEBUG_8_wire\
        );

    \DEBUG_8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12727\,
            PADOUT => \N__12726\,
            PADIN => \N__12725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5193\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D15_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12718\,
            DIN => \N__12717\,
            DOUT => \N__12716\,
            PACKAGEPIN => \FIFO_D15_wire\
        );

    \FIFO_D15_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12718\,
            PADOUT => \N__12717\,
            PADIN => \N__12716\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12709\,
            DIN => \N__12708\,
            DOUT => \N__12707\,
            PACKAGEPIN => \DEBUG_2_wire\
        );

    \DEBUG_2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12709\,
            PADOUT => \N__12708\,
            PADIN => \N__12707\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11946\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA13_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12700\,
            DIN => \N__12699\,
            DOUT => \N__12698\,
            PACKAGEPIN => \DATA13_wire\
        );

    \DATA13_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12700\,
            PADOUT => \N__12699\,
            PADIN => \N__12698\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10172\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D5_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12691\,
            DIN => \N__12690\,
            DOUT => \N__12689\,
            PACKAGEPIN => \FIFO_D5_wire\
        );

    \FIFO_D5_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12691\,
            PADOUT => \N__12690\,
            PADIN => \N__12689\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D4_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12682\,
            DIN => \N__12681\,
            DOUT => \N__12680\,
            PACKAGEPIN => \FIFO_D4_wire\
        );

    \FIFO_D4_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12682\,
            PADOUT => \N__12681\,
            PADIN => \N__12680\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D18_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12673\,
            DIN => \N__12672\,
            DOUT => \N__12671\,
            PACKAGEPIN => \FIFO_D18_wire\
        );

    \FIFO_D18_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12673\,
            PADOUT => \N__12672\,
            PADIN => \N__12671\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA23_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12664\,
            DIN => \N__12663\,
            DOUT => \N__12662\,
            PACKAGEPIN => \DATA23_wire\
        );

    \DATA23_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12664\,
            PADOUT => \N__12663\,
            PADIN => \N__12662\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10188\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_8_c_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12655\,
            DIN => \N__12654\,
            DOUT => \N__12653\,
            PACKAGEPIN => \FIFO_D0_wire\
        );

    \DEBUG_8_c_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12655\,
            PADOUT => \N__12654\,
            PADIN => \N__12653\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_8_c_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ICE_SYSCLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12646\,
            DIN => \N__12645\,
            DOUT => \N__12644\,
            PACKAGEPIN => \ICE_SYSCLK_wire\
        );

    \ICE_SYSCLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12646\,
            PADOUT => \N__12645\,
            PADIN => \N__12644\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ICE_SYSCLK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \FIFO_D30_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12637\,
            DIN => \N__12636\,
            DOUT => \N__12635\,
            PACKAGEPIN => \FIFO_D30_wire\
        );

    \FIFO_D30_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12637\,
            PADOUT => \N__12636\,
            PADIN => \N__12635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DATA0_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12628\,
            DIN => \N__12627\,
            DOUT => \N__12626\,
            PACKAGEPIN => \DATA0_wire\
        );

    \DATA0_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__12628\,
            PADOUT => \N__12627\,
            PADIN => \N__12626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10083\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2921\ : InMux
    port map (
            O => \N__12609\,
            I => \N__12606\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__12606\,
            I => n7
        );

    \I__2919\ : InMux
    port map (
            O => \N__12603\,
            I => n2955
        );

    \I__2918\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12597\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__12597\,
            I => n6
        );

    \I__2916\ : InMux
    port map (
            O => \N__12594\,
            I => n2956
        );

    \I__2915\ : InMux
    port map (
            O => \N__12591\,
            I => \N__12588\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__12588\,
            I => n5
        );

    \I__2913\ : InMux
    port map (
            O => \N__12585\,
            I => n2957
        );

    \I__2912\ : InMux
    port map (
            O => \N__12582\,
            I => \N__12579\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__12579\,
            I => n4_adj_502
        );

    \I__2910\ : InMux
    port map (
            O => \N__12576\,
            I => n2958
        );

    \I__2909\ : InMux
    port map (
            O => \N__12573\,
            I => \N__12570\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__12570\,
            I => n3
        );

    \I__2907\ : InMux
    port map (
            O => \N__12567\,
            I => n2959
        );

    \I__2906\ : InMux
    port map (
            O => \N__12564\,
            I => \N__12561\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__12561\,
            I => n2_adj_503
        );

    \I__2904\ : InMux
    port map (
            O => \N__12558\,
            I => n2960
        );

    \I__2903\ : InMux
    port map (
            O => \N__12555\,
            I => \bfn_24_9_0_\
        );

    \I__2902\ : IoInMux
    port map (
            O => \N__12552\,
            I => \N__12549\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__12549\,
            I => \N__12546\
        );

    \I__2900\ : IoSpan4Mux
    port map (
            O => \N__12546\,
            I => \N__12543\
        );

    \I__2899\ : Span4Mux_s3_h
    port map (
            O => \N__12543\,
            I => \N__12540\
        );

    \I__2898\ : Span4Mux_v
    port map (
            O => \N__12540\,
            I => \N__12536\
        );

    \I__2897\ : InMux
    port map (
            O => \N__12539\,
            I => \N__12533\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__12536\,
            I => \DEBUG_0_c_24\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__12533\,
            I => \DEBUG_0_c_24\
        );

    \I__2894\ : InMux
    port map (
            O => \N__12528\,
            I => \N__12525\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__12525\,
            I => \N__12516\
        );

    \I__2892\ : ClkMux
    port map (
            O => \N__12524\,
            I => \N__12327\
        );

    \I__2891\ : ClkMux
    port map (
            O => \N__12523\,
            I => \N__12327\
        );

    \I__2890\ : ClkMux
    port map (
            O => \N__12522\,
            I => \N__12327\
        );

    \I__2889\ : ClkMux
    port map (
            O => \N__12521\,
            I => \N__12327\
        );

    \I__2888\ : ClkMux
    port map (
            O => \N__12520\,
            I => \N__12327\
        );

    \I__2887\ : ClkMux
    port map (
            O => \N__12519\,
            I => \N__12327\
        );

    \I__2886\ : Glb2LocalMux
    port map (
            O => \N__12516\,
            I => \N__12327\
        );

    \I__2885\ : ClkMux
    port map (
            O => \N__12515\,
            I => \N__12327\
        );

    \I__2884\ : ClkMux
    port map (
            O => \N__12514\,
            I => \N__12327\
        );

    \I__2883\ : ClkMux
    port map (
            O => \N__12513\,
            I => \N__12327\
        );

    \I__2882\ : ClkMux
    port map (
            O => \N__12512\,
            I => \N__12327\
        );

    \I__2881\ : ClkMux
    port map (
            O => \N__12511\,
            I => \N__12327\
        );

    \I__2880\ : ClkMux
    port map (
            O => \N__12510\,
            I => \N__12327\
        );

    \I__2879\ : ClkMux
    port map (
            O => \N__12509\,
            I => \N__12327\
        );

    \I__2878\ : ClkMux
    port map (
            O => \N__12508\,
            I => \N__12327\
        );

    \I__2877\ : ClkMux
    port map (
            O => \N__12507\,
            I => \N__12327\
        );

    \I__2876\ : ClkMux
    port map (
            O => \N__12506\,
            I => \N__12327\
        );

    \I__2875\ : ClkMux
    port map (
            O => \N__12505\,
            I => \N__12327\
        );

    \I__2874\ : ClkMux
    port map (
            O => \N__12504\,
            I => \N__12327\
        );

    \I__2873\ : ClkMux
    port map (
            O => \N__12503\,
            I => \N__12327\
        );

    \I__2872\ : ClkMux
    port map (
            O => \N__12502\,
            I => \N__12327\
        );

    \I__2871\ : ClkMux
    port map (
            O => \N__12501\,
            I => \N__12327\
        );

    \I__2870\ : ClkMux
    port map (
            O => \N__12500\,
            I => \N__12327\
        );

    \I__2869\ : ClkMux
    port map (
            O => \N__12499\,
            I => \N__12327\
        );

    \I__2868\ : ClkMux
    port map (
            O => \N__12498\,
            I => \N__12327\
        );

    \I__2867\ : ClkMux
    port map (
            O => \N__12497\,
            I => \N__12327\
        );

    \I__2866\ : ClkMux
    port map (
            O => \N__12496\,
            I => \N__12327\
        );

    \I__2865\ : ClkMux
    port map (
            O => \N__12495\,
            I => \N__12327\
        );

    \I__2864\ : ClkMux
    port map (
            O => \N__12494\,
            I => \N__12327\
        );

    \I__2863\ : ClkMux
    port map (
            O => \N__12493\,
            I => \N__12327\
        );

    \I__2862\ : ClkMux
    port map (
            O => \N__12492\,
            I => \N__12327\
        );

    \I__2861\ : ClkMux
    port map (
            O => \N__12491\,
            I => \N__12327\
        );

    \I__2860\ : ClkMux
    port map (
            O => \N__12490\,
            I => \N__12327\
        );

    \I__2859\ : ClkMux
    port map (
            O => \N__12489\,
            I => \N__12327\
        );

    \I__2858\ : ClkMux
    port map (
            O => \N__12488\,
            I => \N__12327\
        );

    \I__2857\ : ClkMux
    port map (
            O => \N__12487\,
            I => \N__12327\
        );

    \I__2856\ : ClkMux
    port map (
            O => \N__12486\,
            I => \N__12327\
        );

    \I__2855\ : ClkMux
    port map (
            O => \N__12485\,
            I => \N__12327\
        );

    \I__2854\ : ClkMux
    port map (
            O => \N__12484\,
            I => \N__12327\
        );

    \I__2853\ : ClkMux
    port map (
            O => \N__12483\,
            I => \N__12327\
        );

    \I__2852\ : ClkMux
    port map (
            O => \N__12482\,
            I => \N__12327\
        );

    \I__2851\ : ClkMux
    port map (
            O => \N__12481\,
            I => \N__12327\
        );

    \I__2850\ : ClkMux
    port map (
            O => \N__12480\,
            I => \N__12327\
        );

    \I__2849\ : ClkMux
    port map (
            O => \N__12479\,
            I => \N__12327\
        );

    \I__2848\ : ClkMux
    port map (
            O => \N__12478\,
            I => \N__12327\
        );

    \I__2847\ : ClkMux
    port map (
            O => \N__12477\,
            I => \N__12327\
        );

    \I__2846\ : ClkMux
    port map (
            O => \N__12476\,
            I => \N__12327\
        );

    \I__2845\ : ClkMux
    port map (
            O => \N__12475\,
            I => \N__12327\
        );

    \I__2844\ : ClkMux
    port map (
            O => \N__12474\,
            I => \N__12327\
        );

    \I__2843\ : ClkMux
    port map (
            O => \N__12473\,
            I => \N__12327\
        );

    \I__2842\ : ClkMux
    port map (
            O => \N__12472\,
            I => \N__12327\
        );

    \I__2841\ : ClkMux
    port map (
            O => \N__12471\,
            I => \N__12327\
        );

    \I__2840\ : ClkMux
    port map (
            O => \N__12470\,
            I => \N__12327\
        );

    \I__2839\ : ClkMux
    port map (
            O => \N__12469\,
            I => \N__12327\
        );

    \I__2838\ : ClkMux
    port map (
            O => \N__12468\,
            I => \N__12327\
        );

    \I__2837\ : ClkMux
    port map (
            O => \N__12467\,
            I => \N__12327\
        );

    \I__2836\ : ClkMux
    port map (
            O => \N__12466\,
            I => \N__12327\
        );

    \I__2835\ : ClkMux
    port map (
            O => \N__12465\,
            I => \N__12327\
        );

    \I__2834\ : ClkMux
    port map (
            O => \N__12464\,
            I => \N__12327\
        );

    \I__2833\ : ClkMux
    port map (
            O => \N__12463\,
            I => \N__12327\
        );

    \I__2832\ : ClkMux
    port map (
            O => \N__12462\,
            I => \N__12327\
        );

    \I__2831\ : ClkMux
    port map (
            O => \N__12461\,
            I => \N__12327\
        );

    \I__2830\ : ClkMux
    port map (
            O => \N__12460\,
            I => \N__12327\
        );

    \I__2829\ : ClkMux
    port map (
            O => \N__12459\,
            I => \N__12327\
        );

    \I__2828\ : ClkMux
    port map (
            O => \N__12458\,
            I => \N__12327\
        );

    \I__2827\ : GlobalMux
    port map (
            O => \N__12327\,
            I => \N__12324\
        );

    \I__2826\ : gio2CtrlBuf
    port map (
            O => \N__12324\,
            I => \SLM_CLK_c\
        );

    \I__2825\ : IoInMux
    port map (
            O => \N__12321\,
            I => \N__12318\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__12318\,
            I => \N__12315\
        );

    \I__2823\ : Span4Mux_s3_h
    port map (
            O => \N__12315\,
            I => \N__12312\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__12312\,
            I => \GB_BUFFER_SLM_CLK_c_THRU_CO\
        );

    \I__2821\ : InMux
    port map (
            O => \N__12309\,
            I => \N__12306\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__12306\,
            I => n16
        );

    \I__2819\ : InMux
    port map (
            O => \N__12303\,
            I => n2946
        );

    \I__2818\ : InMux
    port map (
            O => \N__12300\,
            I => \N__12297\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__12297\,
            I => n15
        );

    \I__2816\ : InMux
    port map (
            O => \N__12294\,
            I => n2947
        );

    \I__2815\ : InMux
    port map (
            O => \N__12291\,
            I => \N__12288\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__12288\,
            I => n14
        );

    \I__2813\ : InMux
    port map (
            O => \N__12285\,
            I => n2948
        );

    \I__2812\ : InMux
    port map (
            O => \N__12282\,
            I => \N__12279\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__12279\,
            I => n13
        );

    \I__2810\ : InMux
    port map (
            O => \N__12276\,
            I => n2949
        );

    \I__2809\ : InMux
    port map (
            O => \N__12273\,
            I => \N__12270\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__12270\,
            I => n12
        );

    \I__2807\ : InMux
    port map (
            O => \N__12267\,
            I => n2950
        );

    \I__2806\ : InMux
    port map (
            O => \N__12264\,
            I => \N__12261\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__12261\,
            I => n11
        );

    \I__2804\ : InMux
    port map (
            O => \N__12258\,
            I => n2951
        );

    \I__2803\ : InMux
    port map (
            O => \N__12255\,
            I => \N__12252\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__12252\,
            I => n10
        );

    \I__2801\ : InMux
    port map (
            O => \N__12249\,
            I => n2952
        );

    \I__2800\ : InMux
    port map (
            O => \N__12246\,
            I => \N__12243\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__12243\,
            I => n9
        );

    \I__2798\ : InMux
    port map (
            O => \N__12240\,
            I => \bfn_24_8_0_\
        );

    \I__2797\ : InMux
    port map (
            O => \N__12237\,
            I => \N__12234\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__12234\,
            I => n8_adj_501
        );

    \I__2795\ : InMux
    port map (
            O => \N__12231\,
            I => n2954
        );

    \I__2794\ : InMux
    port map (
            O => \N__12228\,
            I => \N__12225\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__12225\,
            I => n24
        );

    \I__2792\ : InMux
    port map (
            O => \N__12222\,
            I => n2938
        );

    \I__2791\ : InMux
    port map (
            O => \N__12219\,
            I => \N__12216\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__12216\,
            I => n23
        );

    \I__2789\ : InMux
    port map (
            O => \N__12213\,
            I => n2939
        );

    \I__2788\ : InMux
    port map (
            O => \N__12210\,
            I => \N__12207\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__12207\,
            I => n22
        );

    \I__2786\ : InMux
    port map (
            O => \N__12204\,
            I => n2940
        );

    \I__2785\ : InMux
    port map (
            O => \N__12201\,
            I => \N__12198\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__12198\,
            I => n21
        );

    \I__2783\ : InMux
    port map (
            O => \N__12195\,
            I => n2941
        );

    \I__2782\ : InMux
    port map (
            O => \N__12192\,
            I => \N__12189\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__12189\,
            I => n20
        );

    \I__2780\ : InMux
    port map (
            O => \N__12186\,
            I => n2942
        );

    \I__2779\ : InMux
    port map (
            O => \N__12183\,
            I => \N__12180\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__12180\,
            I => n19
        );

    \I__2777\ : InMux
    port map (
            O => \N__12177\,
            I => n2943
        );

    \I__2776\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12171\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__12171\,
            I => n18
        );

    \I__2774\ : InMux
    port map (
            O => \N__12168\,
            I => n2944
        );

    \I__2773\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12162\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__12162\,
            I => n17
        );

    \I__2771\ : InMux
    port map (
            O => \N__12159\,
            I => \bfn_24_7_0_\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__12156\,
            I => \N__12153\
        );

    \I__2769\ : InMux
    port map (
            O => \N__12153\,
            I => \N__12150\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__12150\,
            I => n4_adj_506
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__12147\,
            I => \n4_adj_506_cascade_\
        );

    \I__2766\ : InMux
    port map (
            O => \N__12144\,
            I => \N__12141\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__12141\,
            I => \N__12138\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__12138\,
            I => \N__12134\
        );

    \I__2763\ : InMux
    port map (
            O => \N__12137\,
            I => \N__12131\
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__12134\,
            I => pc_data_rx_5
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__12131\,
            I => pc_data_rx_5
        );

    \I__2760\ : InMux
    port map (
            O => \N__12126\,
            I => \N__12118\
        );

    \I__2759\ : InMux
    port map (
            O => \N__12125\,
            I => \N__12113\
        );

    \I__2758\ : InMux
    port map (
            O => \N__12124\,
            I => \N__12113\
        );

    \I__2757\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12110\
        );

    \I__2756\ : InMux
    port map (
            O => \N__12122\,
            I => \N__12107\
        );

    \I__2755\ : InMux
    port map (
            O => \N__12121\,
            I => \N__12104\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__12118\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__12113\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__12110\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__12107\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__12104\,
            I => \pc_rx.r_Bit_Index_2\
        );

    \I__2749\ : InMux
    port map (
            O => \N__12093\,
            I => \N__12084\
        );

    \I__2748\ : InMux
    port map (
            O => \N__12092\,
            I => \N__12079\
        );

    \I__2747\ : InMux
    port map (
            O => \N__12091\,
            I => \N__12079\
        );

    \I__2746\ : InMux
    port map (
            O => \N__12090\,
            I => \N__12076\
        );

    \I__2745\ : InMux
    port map (
            O => \N__12089\,
            I => \N__12073\
        );

    \I__2744\ : InMux
    port map (
            O => \N__12088\,
            I => \N__12068\
        );

    \I__2743\ : InMux
    port map (
            O => \N__12087\,
            I => \N__12068\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__12084\,
            I => \pc_rx.r_Bit_Index_1\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__12079\,
            I => \pc_rx.r_Bit_Index_1\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__12076\,
            I => \pc_rx.r_Bit_Index_1\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__12073\,
            I => \pc_rx.r_Bit_Index_1\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__12068\,
            I => \pc_rx.r_Bit_Index_1\
        );

    \I__2737\ : InMux
    port map (
            O => \N__12057\,
            I => \N__12054\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__12054\,
            I => n4_adj_500
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__12051\,
            I => \n4_adj_500_cascade_\
        );

    \I__2734\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12042\
        );

    \I__2733\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12042\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__12042\,
            I => n1754
        );

    \I__2731\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12036\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__12036\,
            I => \N__12033\
        );

    \I__2729\ : Span4Mux_v
    port map (
            O => \N__12033\,
            I => \N__12029\
        );

    \I__2728\ : InMux
    port map (
            O => \N__12032\,
            I => \N__12026\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__12029\,
            I => pc_data_rx_1
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__12026\,
            I => pc_data_rx_1
        );

    \I__2725\ : InMux
    port map (
            O => \N__12021\,
            I => \N__12018\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__12018\,
            I => \N__12005\
        );

    \I__2723\ : InMux
    port map (
            O => \N__12017\,
            I => \N__12000\
        );

    \I__2722\ : InMux
    port map (
            O => \N__12016\,
            I => \N__12000\
        );

    \I__2721\ : InMux
    port map (
            O => \N__12015\,
            I => \N__11993\
        );

    \I__2720\ : InMux
    port map (
            O => \N__12014\,
            I => \N__11993\
        );

    \I__2719\ : InMux
    port map (
            O => \N__12013\,
            I => \N__11993\
        );

    \I__2718\ : InMux
    port map (
            O => \N__12012\,
            I => \N__11990\
        );

    \I__2717\ : InMux
    port map (
            O => \N__12011\,
            I => \N__11987\
        );

    \I__2716\ : InMux
    port map (
            O => \N__12010\,
            I => \N__11984\
        );

    \I__2715\ : InMux
    port map (
            O => \N__12009\,
            I => \N__11981\
        );

    \I__2714\ : InMux
    port map (
            O => \N__12008\,
            I => \N__11977\
        );

    \I__2713\ : Span4Mux_h
    port map (
            O => \N__12005\,
            I => \N__11962\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__12000\,
            I => \N__11962\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__11993\,
            I => \N__11962\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__11990\,
            I => \N__11962\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__11987\,
            I => \N__11962\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__11984\,
            I => \N__11962\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11981\,
            I => \N__11962\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11980\,
            I => \N__11959\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__11977\,
            I => \N__11956\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__11962\,
            I => \N__11951\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__11959\,
            I => \N__11951\
        );

    \I__2702\ : Odrv12
    port map (
            O => \N__11956\,
            I => \r_Rx_Data\
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__11951\,
            I => \r_Rx_Data\
        );

    \I__2700\ : IoInMux
    port map (
            O => \N__11946\,
            I => \N__11942\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__11945\,
            I => \N__11939\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__11942\,
            I => \N__11935\
        );

    \I__2697\ : InMux
    port map (
            O => \N__11939\,
            I => \N__11932\
        );

    \I__2696\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11929\
        );

    \I__2695\ : Span4Mux_s2_h
    port map (
            O => \N__11935\,
            I => \N__11926\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__11932\,
            I => \N__11921\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__11929\,
            I => \N__11921\
        );

    \I__2692\ : Span4Mux_v
    port map (
            O => \N__11926\,
            I => \N__11918\
        );

    \I__2691\ : Span4Mux_v
    port map (
            O => \N__11921\,
            I => \N__11915\
        );

    \I__2690\ : Span4Mux_h
    port map (
            O => \N__11918\,
            I => \N__11912\
        );

    \I__2689\ : Span4Mux_h
    port map (
            O => \N__11915\,
            I => \N__11909\
        );

    \I__2688\ : Odrv4
    port map (
            O => \N__11912\,
            I => \DEBUG_2_c\
        );

    \I__2687\ : Odrv4
    port map (
            O => \N__11909\,
            I => \DEBUG_2_c\
        );

    \I__2686\ : InMux
    port map (
            O => \N__11904\,
            I => \N__11895\
        );

    \I__2685\ : InMux
    port map (
            O => \N__11903\,
            I => \N__11890\
        );

    \I__2684\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11890\
        );

    \I__2683\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11887\
        );

    \I__2682\ : InMux
    port map (
            O => \N__11900\,
            I => \N__11884\
        );

    \I__2681\ : InMux
    port map (
            O => \N__11899\,
            I => \N__11873\
        );

    \I__2680\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11873\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__11895\,
            I => \N__11870\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__11890\,
            I => \N__11863\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11887\,
            I => \N__11863\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__11884\,
            I => \N__11863\
        );

    \I__2675\ : InMux
    port map (
            O => \N__11883\,
            I => \N__11860\
        );

    \I__2674\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11855\
        );

    \I__2673\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11855\
        );

    \I__2672\ : InMux
    port map (
            O => \N__11880\,
            I => \N__11850\
        );

    \I__2671\ : InMux
    port map (
            O => \N__11879\,
            I => \N__11850\
        );

    \I__2670\ : InMux
    port map (
            O => \N__11878\,
            I => \N__11846\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__11873\,
            I => \N__11841\
        );

    \I__2668\ : Span4Mux_h
    port map (
            O => \N__11870\,
            I => \N__11833\
        );

    \I__2667\ : Span4Mux_v
    port map (
            O => \N__11863\,
            I => \N__11833\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__11860\,
            I => \N__11833\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__11855\,
            I => \N__11828\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__11850\,
            I => \N__11828\
        );

    \I__2663\ : InMux
    port map (
            O => \N__11849\,
            I => \N__11825\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__11846\,
            I => \N__11822\
        );

    \I__2661\ : InMux
    port map (
            O => \N__11845\,
            I => \N__11819\
        );

    \I__2660\ : InMux
    port map (
            O => \N__11844\,
            I => \N__11816\
        );

    \I__2659\ : Span4Mux_v
    port map (
            O => \N__11841\,
            I => \N__11812\
        );

    \I__2658\ : InMux
    port map (
            O => \N__11840\,
            I => \N__11809\
        );

    \I__2657\ : Span4Mux_h
    port map (
            O => \N__11833\,
            I => \N__11798\
        );

    \I__2656\ : Span4Mux_v
    port map (
            O => \N__11828\,
            I => \N__11798\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__11825\,
            I => \N__11798\
        );

    \I__2654\ : Span4Mux_v
    port map (
            O => \N__11822\,
            I => \N__11798\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__11819\,
            I => \N__11798\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__11816\,
            I => \N__11795\
        );

    \I__2651\ : InMux
    port map (
            O => \N__11815\,
            I => \N__11792\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__11812\,
            I => \N__11789\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__11809\,
            I => \N__11786\
        );

    \I__2648\ : Span4Mux_v
    port map (
            O => \N__11798\,
            I => \N__11783\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__11795\,
            I => \N__11778\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__11792\,
            I => \N__11778\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__11789\,
            I => uart_rx_complete_rising_edge
        );

    \I__2644\ : Odrv12
    port map (
            O => \N__11786\,
            I => uart_rx_complete_rising_edge
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__11783\,
            I => uart_rx_complete_rising_edge
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__11778\,
            I => uart_rx_complete_rising_edge
        );

    \I__2641\ : InMux
    port map (
            O => \N__11769\,
            I => \N__11765\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11762\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__11765\,
            I => even_byte_flag
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__11762\,
            I => even_byte_flag
        );

    \I__2637\ : InMux
    port map (
            O => \N__11757\,
            I => \N__11754\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__11754\,
            I => \N__11751\
        );

    \I__2635\ : Span4Mux_v
    port map (
            O => \N__11751\,
            I => \N__11748\
        );

    \I__2634\ : Span4Mux_h
    port map (
            O => \N__11748\,
            I => \N__11745\
        );

    \I__2633\ : Span4Mux_v
    port map (
            O => \N__11745\,
            I => \N__11742\
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__11742\,
            I => \UART_RX_c\
        );

    \I__2631\ : InMux
    port map (
            O => \N__11739\,
            I => \N__11736\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__11736\,
            I => \N__11733\
        );

    \I__2629\ : Span12Mux_v
    port map (
            O => \N__11733\,
            I => \N__11730\
        );

    \I__2628\ : Odrv12
    port map (
            O => \N__11730\,
            I => \pc_rx.r_Rx_Data_R\
        );

    \I__2627\ : InMux
    port map (
            O => \N__11727\,
            I => \N__11724\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__11724\,
            I => n25
        );

    \I__2625\ : InMux
    port map (
            O => \N__11721\,
            I => \bfn_24_6_0_\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__11718\,
            I => \n4_adj_504_cascade_\
        );

    \I__2623\ : InMux
    port map (
            O => \N__11715\,
            I => \N__11712\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__11712\,
            I => \N__11709\
        );

    \I__2621\ : Span4Mux_v
    port map (
            O => \N__11709\,
            I => \N__11706\
        );

    \I__2620\ : Span4Mux_v
    port map (
            O => \N__11706\,
            I => \N__11702\
        );

    \I__2619\ : InMux
    port map (
            O => \N__11705\,
            I => \N__11699\
        );

    \I__2618\ : Odrv4
    port map (
            O => \N__11702\,
            I => pc_data_rx_2
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__11699\,
            I => pc_data_rx_2
        );

    \I__2616\ : CascadeMux
    port map (
            O => \N__11694\,
            I => \pc_rx.n3334_cascade_\
        );

    \I__2615\ : SRMux
    port map (
            O => \N__11691\,
            I => \N__11688\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__11688\,
            I => \pc_rx.n1900\
        );

    \I__2613\ : SRMux
    port map (
            O => \N__11685\,
            I => \N__11682\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__11682\,
            I => \N__11676\
        );

    \I__2611\ : InMux
    port map (
            O => \N__11681\,
            I => \N__11671\
        );

    \I__2610\ : InMux
    port map (
            O => \N__11680\,
            I => \N__11671\
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__11679\,
            I => \N__11665\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__11676\,
            I => \N__11660\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__11671\,
            I => \N__11657\
        );

    \I__2606\ : InMux
    port map (
            O => \N__11670\,
            I => \N__11654\
        );

    \I__2605\ : InMux
    port map (
            O => \N__11669\,
            I => \N__11649\
        );

    \I__2604\ : InMux
    port map (
            O => \N__11668\,
            I => \N__11649\
        );

    \I__2603\ : InMux
    port map (
            O => \N__11665\,
            I => \N__11646\
        );

    \I__2602\ : InMux
    port map (
            O => \N__11664\,
            I => \N__11641\
        );

    \I__2601\ : InMux
    port map (
            O => \N__11663\,
            I => \N__11641\
        );

    \I__2600\ : Odrv4
    port map (
            O => \N__11660\,
            I => \r_SM_Main_2\
        );

    \I__2599\ : Odrv4
    port map (
            O => \N__11657\,
            I => \r_SM_Main_2\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__11654\,
            I => \r_SM_Main_2\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__11649\,
            I => \r_SM_Main_2\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__11646\,
            I => \r_SM_Main_2\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__11641\,
            I => \r_SM_Main_2\
        );

    \I__2594\ : InMux
    port map (
            O => \N__11628\,
            I => \N__11623\
        );

    \I__2593\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11618\
        );

    \I__2592\ : InMux
    port map (
            O => \N__11626\,
            I => \N__11618\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__11623\,
            I => \N__11611\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__11618\,
            I => \N__11608\
        );

    \I__2589\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11605\
        );

    \I__2588\ : InMux
    port map (
            O => \N__11616\,
            I => \N__11601\
        );

    \I__2587\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11598\
        );

    \I__2586\ : InMux
    port map (
            O => \N__11614\,
            I => \N__11595\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__11611\,
            I => \N__11588\
        );

    \I__2584\ : Span4Mux_v
    port map (
            O => \N__11608\,
            I => \N__11588\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__11605\,
            I => \N__11588\
        );

    \I__2582\ : InMux
    port map (
            O => \N__11604\,
            I => \N__11585\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__11601\,
            I => \r_SM_Main_2_N_108_2\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__11598\,
            I => \r_SM_Main_2_N_108_2\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__11595\,
            I => \r_SM_Main_2_N_108_2\
        );

    \I__2578\ : Odrv4
    port map (
            O => \N__11588\,
            I => \r_SM_Main_2_N_108_2\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__11585\,
            I => \r_SM_Main_2_N_108_2\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__11574\,
            I => \N__11571\
        );

    \I__2575\ : InMux
    port map (
            O => \N__11571\,
            I => \N__11559\
        );

    \I__2574\ : InMux
    port map (
            O => \N__11570\,
            I => \N__11559\
        );

    \I__2573\ : InMux
    port map (
            O => \N__11569\,
            I => \N__11559\
        );

    \I__2572\ : InMux
    port map (
            O => \N__11568\,
            I => \N__11551\
        );

    \I__2571\ : InMux
    port map (
            O => \N__11567\,
            I => \N__11551\
        );

    \I__2570\ : InMux
    port map (
            O => \N__11566\,
            I => \N__11551\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__11559\,
            I => \N__11544\
        );

    \I__2568\ : InMux
    port map (
            O => \N__11558\,
            I => \N__11541\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__11551\,
            I => \N__11538\
        );

    \I__2566\ : InMux
    port map (
            O => \N__11550\,
            I => \N__11535\
        );

    \I__2565\ : InMux
    port map (
            O => \N__11549\,
            I => \N__11532\
        );

    \I__2564\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11527\
        );

    \I__2563\ : InMux
    port map (
            O => \N__11547\,
            I => \N__11527\
        );

    \I__2562\ : Odrv4
    port map (
            O => \N__11544\,
            I => \r_SM_Main_0\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__11541\,
            I => \r_SM_Main_0\
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__11538\,
            I => \r_SM_Main_0\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__11535\,
            I => \r_SM_Main_0\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__11532\,
            I => \r_SM_Main_0\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__11527\,
            I => \r_SM_Main_0\
        );

    \I__2556\ : CEMux
    port map (
            O => \N__11514\,
            I => \N__11511\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__11511\,
            I => \N__11508\
        );

    \I__2554\ : Span4Mux_v
    port map (
            O => \N__11508\,
            I => \N__11505\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__11505\,
            I => n3293
        );

    \I__2552\ : InMux
    port map (
            O => \N__11502\,
            I => \N__11492\
        );

    \I__2551\ : InMux
    port map (
            O => \N__11501\,
            I => \N__11492\
        );

    \I__2550\ : InMux
    port map (
            O => \N__11500\,
            I => \N__11492\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__11499\,
            I => \N__11488\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__11492\,
            I => \N__11482\
        );

    \I__2547\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11475\
        );

    \I__2546\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11475\
        );

    \I__2545\ : InMux
    port map (
            O => \N__11487\,
            I => \N__11475\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__11486\,
            I => \N__11471\
        );

    \I__2543\ : InMux
    port map (
            O => \N__11485\,
            I => \N__11466\
        );

    \I__2542\ : Span4Mux_h
    port map (
            O => \N__11482\,
            I => \N__11461\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__11475\,
            I => \N__11461\
        );

    \I__2540\ : InMux
    port map (
            O => \N__11474\,
            I => \N__11458\
        );

    \I__2539\ : InMux
    port map (
            O => \N__11471\,
            I => \N__11455\
        );

    \I__2538\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11450\
        );

    \I__2537\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11450\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__11466\,
            I => \r_SM_Main_1\
        );

    \I__2535\ : Odrv4
    port map (
            O => \N__11461\,
            I => \r_SM_Main_1\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__11458\,
            I => \r_SM_Main_1\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__11455\,
            I => \r_SM_Main_1\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__11450\,
            I => \r_SM_Main_1\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__11439\,
            I => \n3293_cascade_\
        );

    \I__2530\ : InMux
    port map (
            O => \N__11436\,
            I => \N__11427\
        );

    \I__2529\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11427\
        );

    \I__2528\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11427\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__11427\,
            I => \N__11419\
        );

    \I__2526\ : InMux
    port map (
            O => \N__11426\,
            I => \N__11414\
        );

    \I__2525\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11414\
        );

    \I__2524\ : InMux
    port map (
            O => \N__11424\,
            I => \N__11411\
        );

    \I__2523\ : InMux
    port map (
            O => \N__11423\,
            I => \N__11406\
        );

    \I__2522\ : InMux
    port map (
            O => \N__11422\,
            I => \N__11406\
        );

    \I__2521\ : Odrv4
    port map (
            O => \N__11419\,
            I => \r_Bit_Index_0\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__11414\,
            I => \r_Bit_Index_0\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__11411\,
            I => \r_Bit_Index_0\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__11406\,
            I => \r_Bit_Index_0\
        );

    \I__2517\ : InMux
    port map (
            O => \N__11397\,
            I => \N__11393\
        );

    \I__2516\ : InMux
    port map (
            O => \N__11396\,
            I => \N__11389\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__11393\,
            I => \N__11386\
        );

    \I__2514\ : InMux
    port map (
            O => \N__11392\,
            I => \N__11383\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__11389\,
            I => \N__11380\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__11386\,
            I => n2540
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__11383\,
            I => n2540
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__11380\,
            I => n2540
        );

    \I__2509\ : InMux
    port map (
            O => \N__11373\,
            I => \N__11370\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__11370\,
            I => \N__11366\
        );

    \I__2507\ : InMux
    port map (
            O => \N__11369\,
            I => \N__11363\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__11366\,
            I => pc_data_rx_4
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__11363\,
            I => pc_data_rx_4
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__11358\,
            I => \N__11355\
        );

    \I__2503\ : InMux
    port map (
            O => \N__11355\,
            I => \N__11352\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__11352\,
            I => \N__11347\
        );

    \I__2501\ : InMux
    port map (
            O => \N__11351\,
            I => \N__11344\
        );

    \I__2500\ : InMux
    port map (
            O => \N__11350\,
            I => \N__11341\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__11347\,
            I => n1750
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__11344\,
            I => n1750
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__11341\,
            I => n1750
        );

    \I__2496\ : InMux
    port map (
            O => \N__11334\,
            I => \N__11331\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__11331\,
            I => \N__11328\
        );

    \I__2494\ : Span4Mux_h
    port map (
            O => \N__11328\,
            I => \N__11324\
        );

    \I__2493\ : InMux
    port map (
            O => \N__11327\,
            I => \N__11321\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__11324\,
            I => pc_data_rx_0
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__11321\,
            I => pc_data_rx_0
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__11316\,
            I => \n1754_cascade_\
        );

    \I__2489\ : InMux
    port map (
            O => \N__11313\,
            I => \N__11310\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__11310\,
            I => \N__11306\
        );

    \I__2487\ : InMux
    port map (
            O => \N__11309\,
            I => \N__11303\
        );

    \I__2486\ : Odrv12
    port map (
            O => \N__11306\,
            I => pc_data_rx_3
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__11303\,
            I => pc_data_rx_3
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__11298\,
            I => \N__11295\
        );

    \I__2483\ : InMux
    port map (
            O => \N__11295\,
            I => \N__11292\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__11292\,
            I => n1747
        );

    \I__2481\ : InMux
    port map (
            O => \N__11289\,
            I => \N__11286\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__11286\,
            I => \N__11282\
        );

    \I__2479\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11279\
        );

    \I__2478\ : Odrv4
    port map (
            O => \N__11282\,
            I => pc_data_rx_7
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__11279\,
            I => pc_data_rx_7
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__11274\,
            I => \N__11271\
        );

    \I__2475\ : InMux
    port map (
            O => \N__11271\,
            I => \N__11268\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__11268\,
            I => \N__11264\
        );

    \I__2473\ : InMux
    port map (
            O => \N__11267\,
            I => \N__11261\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__11264\,
            I => \N__11258\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__11261\,
            I => \N__11255\
        );

    \I__2470\ : Span4Mux_h
    port map (
            O => \N__11258\,
            I => \N__11251\
        );

    \I__2469\ : Span4Mux_h
    port map (
            O => \N__11255\,
            I => \N__11248\
        );

    \I__2468\ : InMux
    port map (
            O => \N__11254\,
            I => \N__11245\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__11251\,
            I => tx_data_byte_7
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__11248\,
            I => tx_data_byte_7
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__11245\,
            I => tx_data_byte_7
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__11238\,
            I => \N__11235\
        );

    \I__2463\ : InMux
    port map (
            O => \N__11235\,
            I => \N__11232\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__11232\,
            I => \pc_rx.n3271\
        );

    \I__2461\ : InMux
    port map (
            O => \N__11229\,
            I => \N__11226\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__11226\,
            I => \N__11223\
        );

    \I__2459\ : Span4Mux_v
    port map (
            O => \N__11223\,
            I => \N__11217\
        );

    \I__2458\ : InMux
    port map (
            O => \N__11222\,
            I => \N__11214\
        );

    \I__2457\ : InMux
    port map (
            O => \N__11221\,
            I => \N__11211\
        );

    \I__2456\ : InMux
    port map (
            O => \N__11220\,
            I => \N__11208\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__11217\,
            I => \pc_rx.r_SM_Main_2_N_114_0\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__11214\,
            I => \pc_rx.r_SM_Main_2_N_114_0\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__11211\,
            I => \pc_rx.r_SM_Main_2_N_114_0\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__11208\,
            I => \pc_rx.r_SM_Main_2_N_114_0\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__11199\,
            I => \pc_rx.n1_cascade_\
        );

    \I__2450\ : InMux
    port map (
            O => \N__11196\,
            I => \N__11193\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__11193\,
            I => \pc_rx.n2578\
        );

    \I__2448\ : InMux
    port map (
            O => \N__11190\,
            I => \N__11184\
        );

    \I__2447\ : InMux
    port map (
            O => \N__11189\,
            I => \N__11184\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__11184\,
            I => \N__11180\
        );

    \I__2445\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11177\
        );

    \I__2444\ : Odrv12
    port map (
            O => \N__11180\,
            I => \pc_rx.n1715\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__11177\,
            I => \pc_rx.n1715\
        );

    \I__2442\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11169\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__11169\,
            I => \N__11166\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__11166\,
            I => n4_adj_504
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__11163\,
            I => \pc_rx.n3273_cascade_\
        );

    \I__2438\ : SRMux
    port map (
            O => \N__11160\,
            I => \N__11156\
        );

    \I__2437\ : SRMux
    port map (
            O => \N__11159\,
            I => \N__11153\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__11156\,
            I => \N__11150\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__11153\,
            I => \N__11147\
        );

    \I__2434\ : Span4Mux_v
    port map (
            O => \N__11150\,
            I => \N__11144\
        );

    \I__2433\ : Sp12to4
    port map (
            O => \N__11147\,
            I => \N__11141\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__11144\,
            I => \pc_rx.n1910\
        );

    \I__2431\ : Odrv12
    port map (
            O => \N__11141\,
            I => \pc_rx.n1910\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__11136\,
            I => \pc_rx.n6_adj_492_cascade_\
        );

    \I__2429\ : CEMux
    port map (
            O => \N__11133\,
            I => \N__11130\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__11130\,
            I => \N__11126\
        );

    \I__2427\ : CEMux
    port map (
            O => \N__11129\,
            I => \N__11123\
        );

    \I__2426\ : Span4Mux_v
    port map (
            O => \N__11126\,
            I => \N__11120\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__11123\,
            I => \N__11117\
        );

    \I__2424\ : Span4Mux_h
    port map (
            O => \N__11120\,
            I => \N__11114\
        );

    \I__2423\ : Span4Mux_h
    port map (
            O => \N__11117\,
            I => \N__11111\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__11114\,
            I => \pc_rx.n1815\
        );

    \I__2421\ : Odrv4
    port map (
            O => \N__11111\,
            I => \pc_rx.n1815\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__11106\,
            I => \n1747_cascade_\
        );

    \I__2419\ : InMux
    port map (
            O => \N__11103\,
            I => \N__11100\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__11100\,
            I => \N__11096\
        );

    \I__2417\ : InMux
    port map (
            O => \N__11099\,
            I => \N__11093\
        );

    \I__2416\ : Odrv4
    port map (
            O => \N__11096\,
            I => pc_data_rx_6
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__11093\,
            I => pc_data_rx_6
        );

    \I__2414\ : InMux
    port map (
            O => \N__11088\,
            I => \N__11085\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__11085\,
            I => \N__11081\
        );

    \I__2412\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11078\
        );

    \I__2411\ : Span4Mux_v
    port map (
            O => \N__11081\,
            I => \N__11074\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__11078\,
            I => \N__11071\
        );

    \I__2409\ : InMux
    port map (
            O => \N__11077\,
            I => \N__11068\
        );

    \I__2408\ : Odrv4
    port map (
            O => \N__11074\,
            I => tx_data_byte_5
        );

    \I__2407\ : Odrv4
    port map (
            O => \N__11071\,
            I => tx_data_byte_5
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__11068\,
            I => tx_data_byte_5
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__11061\,
            I => \N__11058\
        );

    \I__2404\ : InMux
    port map (
            O => \N__11058\,
            I => \N__11055\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__11055\,
            I => \N__11052\
        );

    \I__2402\ : Span4Mux_h
    port map (
            O => \N__11052\,
            I => \N__11048\
        );

    \I__2401\ : InMux
    port map (
            O => \N__11051\,
            I => \N__11045\
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__11048\,
            I => tx_addr_byte_2
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__11045\,
            I => tx_addr_byte_2
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__11040\,
            I => \N__11037\
        );

    \I__2397\ : InMux
    port map (
            O => \N__11037\,
            I => \N__11034\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__11034\,
            I => \N__11031\
        );

    \I__2395\ : Span4Mux_h
    port map (
            O => \N__11031\,
            I => \N__11026\
        );

    \I__2394\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11021\
        );

    \I__2393\ : InMux
    port map (
            O => \N__11029\,
            I => \N__11021\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__11026\,
            I => tx_data_byte_2
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__11021\,
            I => tx_data_byte_2
        );

    \I__2390\ : InMux
    port map (
            O => \N__11016\,
            I => \N__11013\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__11013\,
            I => uart_rx_complete_prev
        );

    \I__2388\ : CascadeMux
    port map (
            O => \N__11010\,
            I => \n1764_cascade_\
        );

    \I__2387\ : IoInMux
    port map (
            O => \N__11007\,
            I => \N__11004\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__11004\,
            I => \N__11001\
        );

    \I__2385\ : Span4Mux_s0_h
    port map (
            O => \N__11001\,
            I => \N__10998\
        );

    \I__2384\ : Sp12to4
    port map (
            O => \N__10998\,
            I => \N__10995\
        );

    \I__2383\ : Span12Mux_v
    port map (
            O => \N__10995\,
            I => \N__10989\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10982\
        );

    \I__2381\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10982\
        );

    \I__2380\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10982\
        );

    \I__2379\ : Odrv12
    port map (
            O => \N__10989\,
            I => \DEBUG_1_c\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10982\,
            I => \DEBUG_1_c\
        );

    \I__2377\ : InMux
    port map (
            O => \N__10977\,
            I => \pc_rx.n2920\
        );

    \I__2376\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10967\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10967\
        );

    \I__2374\ : InMux
    port map (
            O => \N__10972\,
            I => \N__10964\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__10967\,
            I => \pc_rx.r_Clock_Count_2\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10964\,
            I => \pc_rx.r_Clock_Count_2\
        );

    \I__2371\ : InMux
    port map (
            O => \N__10959\,
            I => \pc_rx.n2921\
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__10956\,
            I => \N__10953\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10953\,
            I => \N__10946\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10952\,
            I => \N__10946\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10951\,
            I => \N__10943\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__10946\,
            I => \pc_rx.r_Clock_Count_3\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__10943\,
            I => \pc_rx.r_Clock_Count_3\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10938\,
            I => \pc_rx.n2922\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10935\,
            I => \N__10931\
        );

    \I__2362\ : InMux
    port map (
            O => \N__10934\,
            I => \N__10927\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__10931\,
            I => \N__10924\
        );

    \I__2360\ : InMux
    port map (
            O => \N__10930\,
            I => \N__10921\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10927\,
            I => \pc_rx.r_Clock_Count_4\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__10924\,
            I => \pc_rx.r_Clock_Count_4\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10921\,
            I => \pc_rx.r_Clock_Count_4\
        );

    \I__2356\ : InMux
    port map (
            O => \N__10914\,
            I => \pc_rx.n2923\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10904\
        );

    \I__2354\ : InMux
    port map (
            O => \N__10910\,
            I => \N__10904\
        );

    \I__2353\ : InMux
    port map (
            O => \N__10909\,
            I => \N__10901\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__10904\,
            I => \pc_rx.r_Clock_Count_5\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__10901\,
            I => \pc_rx.r_Clock_Count_5\
        );

    \I__2350\ : InMux
    port map (
            O => \N__10896\,
            I => \pc_rx.n2924\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10893\,
            I => \N__10886\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10892\,
            I => \N__10886\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10891\,
            I => \N__10883\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10886\,
            I => \pc_rx.r_Clock_Count_6\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10883\,
            I => \pc_rx.r_Clock_Count_6\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10878\,
            I => \pc_rx.n2925\
        );

    \I__2343\ : InMux
    port map (
            O => \N__10875\,
            I => \N__10868\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10874\,
            I => \N__10868\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10873\,
            I => \N__10865\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__10868\,
            I => \pc_rx.r_Clock_Count_7\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10865\,
            I => \pc_rx.r_Clock_Count_7\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10860\,
            I => \pc_rx.n2926\
        );

    \I__2337\ : InMux
    port map (
            O => \N__10857\,
            I => \N__10851\
        );

    \I__2336\ : InMux
    port map (
            O => \N__10856\,
            I => \N__10851\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__10851\,
            I => \N__10847\
        );

    \I__2334\ : InMux
    port map (
            O => \N__10850\,
            I => \N__10844\
        );

    \I__2333\ : Odrv4
    port map (
            O => \N__10847\,
            I => \pc_rx.r_Clock_Count_8\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__10844\,
            I => \pc_rx.r_Clock_Count_8\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10839\,
            I => \bfn_18_12_0_\
        );

    \I__2330\ : InMux
    port map (
            O => \N__10836\,
            I => \pc_rx.n2928\
        );

    \I__2329\ : InMux
    port map (
            O => \N__10833\,
            I => \N__10827\
        );

    \I__2328\ : InMux
    port map (
            O => \N__10832\,
            I => \N__10827\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__10827\,
            I => \N__10823\
        );

    \I__2326\ : InMux
    port map (
            O => \N__10826\,
            I => \N__10820\
        );

    \I__2325\ : Odrv12
    port map (
            O => \N__10823\,
            I => \pc_rx.r_Clock_Count_9\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__10820\,
            I => \pc_rx.r_Clock_Count_9\
        );

    \I__2323\ : InMux
    port map (
            O => \N__10815\,
            I => \N__10803\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10803\
        );

    \I__2321\ : InMux
    port map (
            O => \N__10813\,
            I => \N__10803\
        );

    \I__2320\ : InMux
    port map (
            O => \N__10812\,
            I => \N__10796\
        );

    \I__2319\ : InMux
    port map (
            O => \N__10811\,
            I => \N__10796\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10810\,
            I => \N__10796\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__10803\,
            I => \N__10790\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__10796\,
            I => \N__10787\
        );

    \I__2315\ : InMux
    port map (
            O => \N__10795\,
            I => \N__10780\
        );

    \I__2314\ : InMux
    port map (
            O => \N__10794\,
            I => \N__10780\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10780\
        );

    \I__2312\ : Span4Mux_h
    port map (
            O => \N__10790\,
            I => \N__10763\
        );

    \I__2311\ : Span4Mux_h
    port map (
            O => \N__10787\,
            I => \N__10758\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__10780\,
            I => \N__10758\
        );

    \I__2309\ : InMux
    port map (
            O => \N__10779\,
            I => \N__10743\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10778\,
            I => \N__10743\
        );

    \I__2307\ : InMux
    port map (
            O => \N__10777\,
            I => \N__10743\
        );

    \I__2306\ : InMux
    port map (
            O => \N__10776\,
            I => \N__10743\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10775\,
            I => \N__10743\
        );

    \I__2304\ : InMux
    port map (
            O => \N__10774\,
            I => \N__10743\
        );

    \I__2303\ : InMux
    port map (
            O => \N__10773\,
            I => \N__10743\
        );

    \I__2302\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10738\
        );

    \I__2301\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10738\
        );

    \I__2300\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10727\
        );

    \I__2299\ : InMux
    port map (
            O => \N__10769\,
            I => \N__10727\
        );

    \I__2298\ : InMux
    port map (
            O => \N__10768\,
            I => \N__10727\
        );

    \I__2297\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10727\
        );

    \I__2296\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10727\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__10763\,
            I => n3279
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__10758\,
            I => n3279
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__10743\,
            I => n3279
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__10738\,
            I => n3279
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__10727\,
            I => n3279
        );

    \I__2290\ : InMux
    port map (
            O => \N__10716\,
            I => \N__10712\
        );

    \I__2289\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10709\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__10712\,
            I => rx_shift_reg_6
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__10709\,
            I => rx_shift_reg_6
        );

    \I__2286\ : ClkMux
    port map (
            O => \N__10704\,
            I => \N__10694\
        );

    \I__2285\ : ClkMux
    port map (
            O => \N__10703\,
            I => \N__10691\
        );

    \I__2284\ : ClkMux
    port map (
            O => \N__10702\,
            I => \N__10681\
        );

    \I__2283\ : ClkMux
    port map (
            O => \N__10701\,
            I => \N__10678\
        );

    \I__2282\ : ClkMux
    port map (
            O => \N__10700\,
            I => \N__10675\
        );

    \I__2281\ : ClkMux
    port map (
            O => \N__10699\,
            I => \N__10672\
        );

    \I__2280\ : ClkMux
    port map (
            O => \N__10698\,
            I => \N__10669\
        );

    \I__2279\ : ClkMux
    port map (
            O => \N__10697\,
            I => \N__10666\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__10694\,
            I => \N__10661\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__10691\,
            I => \N__10661\
        );

    \I__2276\ : ClkMux
    port map (
            O => \N__10690\,
            I => \N__10658\
        );

    \I__2275\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10655\
        );

    \I__2274\ : ClkMux
    port map (
            O => \N__10688\,
            I => \N__10652\
        );

    \I__2273\ : ClkMux
    port map (
            O => \N__10687\,
            I => \N__10649\
        );

    \I__2272\ : ClkMux
    port map (
            O => \N__10686\,
            I => \N__10646\
        );

    \I__2271\ : ClkMux
    port map (
            O => \N__10685\,
            I => \N__10643\
        );

    \I__2270\ : ClkMux
    port map (
            O => \N__10684\,
            I => \N__10640\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__10681\,
            I => \N__10635\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__10678\,
            I => \N__10635\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__10675\,
            I => \N__10628\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__10672\,
            I => \N__10628\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__10669\,
            I => \N__10628\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__10666\,
            I => \N__10624\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__10661\,
            I => \N__10621\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__10658\,
            I => \N__10618\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__10655\,
            I => \N__10609\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__10652\,
            I => \N__10609\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__10649\,
            I => \N__10609\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__10646\,
            I => \N__10609\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__10643\,
            I => \N__10604\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__10640\,
            I => \N__10604\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__10635\,
            I => \N__10599\
        );

    \I__2254\ : Span4Mux_v
    port map (
            O => \N__10628\,
            I => \N__10599\
        );

    \I__2253\ : ClkMux
    port map (
            O => \N__10627\,
            I => \N__10596\
        );

    \I__2252\ : Span4Mux_v
    port map (
            O => \N__10624\,
            I => \N__10593\
        );

    \I__2251\ : Span4Mux_h
    port map (
            O => \N__10621\,
            I => \N__10585\
        );

    \I__2250\ : Span4Mux_v
    port map (
            O => \N__10618\,
            I => \N__10585\
        );

    \I__2249\ : Span4Mux_v
    port map (
            O => \N__10609\,
            I => \N__10585\
        );

    \I__2248\ : Span4Mux_v
    port map (
            O => \N__10604\,
            I => \N__10582\
        );

    \I__2247\ : Sp12to4
    port map (
            O => \N__10599\,
            I => \N__10577\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__10596\,
            I => \N__10577\
        );

    \I__2245\ : Span4Mux_h
    port map (
            O => \N__10593\,
            I => \N__10574\
        );

    \I__2244\ : InMux
    port map (
            O => \N__10592\,
            I => \N__10571\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__10585\,
            I => \spi0.spi_clk\
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__10582\,
            I => \spi0.spi_clk\
        );

    \I__2241\ : Odrv12
    port map (
            O => \N__10577\,
            I => \spi0.spi_clk\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__10574\,
            I => \spi0.spi_clk\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__10571\,
            I => \spi0.spi_clk\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__10560\,
            I => \pc_rx.n3291_cascade_\
        );

    \I__2237\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10554\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__10554\,
            I => \pc_rx.n6\
        );

    \I__2235\ : InMux
    port map (
            O => \N__10551\,
            I => \N__10548\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__10548\,
            I => \pc_rx.n3260\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__10545\,
            I => \pc_rx.n3261_cascade_\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__10542\,
            I => \pc_rx.n2558_cascade_\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__10539\,
            I => \N__10535\
        );

    \I__2230\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10529\
        );

    \I__2229\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10529\
        );

    \I__2228\ : InMux
    port map (
            O => \N__10534\,
            I => \N__10526\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__10529\,
            I => \pc_rx.r_Clock_Count_0\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__10526\,
            I => \pc_rx.r_Clock_Count_0\
        );

    \I__2225\ : InMux
    port map (
            O => \N__10521\,
            I => \bfn_18_11_0_\
        );

    \I__2224\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10513\
        );

    \I__2223\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10510\
        );

    \I__2222\ : InMux
    port map (
            O => \N__10516\,
            I => \N__10507\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__10513\,
            I => \pc_rx.r_Clock_Count_1\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__10510\,
            I => \pc_rx.r_Clock_Count_1\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__10507\,
            I => \pc_rx.r_Clock_Count_1\
        );

    \I__2218\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10496\
        );

    \I__2217\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10493\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__10496\,
            I => \N__10488\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__10493\,
            I => \N__10488\
        );

    \I__2214\ : Span4Mux_h
    port map (
            O => \N__10488\,
            I => \N__10485\
        );

    \I__2213\ : Odrv4
    port map (
            O => \N__10485\,
            I => rx_shift_reg_2
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__10482\,
            I => \N__10478\
        );

    \I__2211\ : InMux
    port map (
            O => \N__10481\,
            I => \N__10473\
        );

    \I__2210\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10473\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__10473\,
            I => \N__10468\
        );

    \I__2208\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10465\
        );

    \I__2207\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10462\
        );

    \I__2206\ : Span4Mux_v
    port map (
            O => \N__10468\,
            I => \N__10459\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__10465\,
            I => \N__10454\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__10462\,
            I => \N__10454\
        );

    \I__2203\ : Span4Mux_h
    port map (
            O => \N__10459\,
            I => \N__10450\
        );

    \I__2202\ : Span4Mux_v
    port map (
            O => \N__10454\,
            I => \N__10447\
        );

    \I__2201\ : InMux
    port map (
            O => \N__10453\,
            I => \N__10444\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__10450\,
            I => rx_buf_byte_7
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__10447\,
            I => rx_buf_byte_7
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__10444\,
            I => rx_buf_byte_7
        );

    \I__2197\ : InMux
    port map (
            O => \N__10437\,
            I => \N__10431\
        );

    \I__2196\ : InMux
    port map (
            O => \N__10436\,
            I => \N__10431\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__10431\,
            I => \N__10427\
        );

    \I__2194\ : InMux
    port map (
            O => \N__10430\,
            I => \N__10424\
        );

    \I__2193\ : Span4Mux_h
    port map (
            O => \N__10427\,
            I => \N__10418\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__10424\,
            I => \N__10418\
        );

    \I__2191\ : InMux
    port map (
            O => \N__10423\,
            I => \N__10415\
        );

    \I__2190\ : Span4Mux_v
    port map (
            O => \N__10418\,
            I => \N__10410\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__10415\,
            I => \N__10410\
        );

    \I__2188\ : Span4Mux_h
    port map (
            O => \N__10410\,
            I => \N__10406\
        );

    \I__2187\ : InMux
    port map (
            O => \N__10409\,
            I => \N__10403\
        );

    \I__2186\ : Odrv4
    port map (
            O => \N__10406\,
            I => rx_buf_byte_4
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__10403\,
            I => rx_buf_byte_4
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__10398\,
            I => \N__10395\
        );

    \I__2183\ : InMux
    port map (
            O => \N__10395\,
            I => \N__10386\
        );

    \I__2182\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10386\
        );

    \I__2181\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10386\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__10386\,
            I => \N__10382\
        );

    \I__2179\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10379\
        );

    \I__2178\ : Span4Mux_h
    port map (
            O => \N__10382\,
            I => \N__10374\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__10379\,
            I => \N__10374\
        );

    \I__2176\ : Span4Mux_h
    port map (
            O => \N__10374\,
            I => \N__10370\
        );

    \I__2175\ : InMux
    port map (
            O => \N__10373\,
            I => \N__10367\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__10370\,
            I => rx_buf_byte_2
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__10367\,
            I => rx_buf_byte_2
        );

    \I__2172\ : InMux
    port map (
            O => \N__10362\,
            I => \N__10347\
        );

    \I__2171\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10347\
        );

    \I__2170\ : InMux
    port map (
            O => \N__10360\,
            I => \N__10347\
        );

    \I__2169\ : InMux
    port map (
            O => \N__10359\,
            I => \N__10347\
        );

    \I__2168\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10340\
        );

    \I__2167\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10340\
        );

    \I__2166\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10340\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__10347\,
            I => \rx_shift_reg_15__N_319\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__10340\,
            I => \rx_shift_reg_15__N_319\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__10335\,
            I => \N__10331\
        );

    \I__2162\ : InMux
    port map (
            O => \N__10334\,
            I => \N__10325\
        );

    \I__2161\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10325\
        );

    \I__2160\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10322\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__10325\,
            I => \N__10318\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__10322\,
            I => \N__10315\
        );

    \I__2157\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10312\
        );

    \I__2156\ : Span4Mux_h
    port map (
            O => \N__10318\,
            I => \N__10305\
        );

    \I__2155\ : Span4Mux_v
    port map (
            O => \N__10315\,
            I => \N__10305\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__10312\,
            I => \N__10305\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__10305\,
            I => \N__10301\
        );

    \I__2152\ : InMux
    port map (
            O => \N__10304\,
            I => \N__10298\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__10301\,
            I => rx_buf_byte_5
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__10298\,
            I => rx_buf_byte_5
        );

    \I__2149\ : InMux
    port map (
            O => \N__10293\,
            I => \N__10289\
        );

    \I__2148\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10286\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__10289\,
            I => rx_shift_reg_3
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__10286\,
            I => rx_shift_reg_3
        );

    \I__2145\ : InMux
    port map (
            O => \N__10281\,
            I => \N__10277\
        );

    \I__2144\ : InMux
    port map (
            O => \N__10280\,
            I => \N__10274\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__10277\,
            I => rx_shift_reg_4
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__10274\,
            I => rx_shift_reg_4
        );

    \I__2141\ : InMux
    port map (
            O => \N__10269\,
            I => \N__10265\
        );

    \I__2140\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10262\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__10265\,
            I => rx_shift_reg_7
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__10262\,
            I => rx_shift_reg_7
        );

    \I__2137\ : InMux
    port map (
            O => \N__10257\,
            I => \N__10254\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__10254\,
            I => rx_shift_reg_8
        );

    \I__2135\ : InMux
    port map (
            O => \N__10251\,
            I => \N__10247\
        );

    \I__2134\ : InMux
    port map (
            O => \N__10250\,
            I => \N__10244\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__10247\,
            I => rx_shift_reg_5
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__10244\,
            I => rx_shift_reg_5
        );

    \I__2131\ : InMux
    port map (
            O => \N__10239\,
            I => \spi0.n2916\
        );

    \I__2130\ : InMux
    port map (
            O => \N__10236\,
            I => \spi0.n2917\
        );

    \I__2129\ : InMux
    port map (
            O => \N__10233\,
            I => \spi0.n2918\
        );

    \I__2128\ : IoInMux
    port map (
            O => \N__10230\,
            I => \N__10226\
        );

    \I__2127\ : IoInMux
    port map (
            O => \N__10229\,
            I => \N__10223\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__10226\,
            I => \N__10208\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__10223\,
            I => \N__10208\
        );

    \I__2124\ : IoInMux
    port map (
            O => \N__10222\,
            I => \N__10205\
        );

    \I__2123\ : IoInMux
    port map (
            O => \N__10221\,
            I => \N__10202\
        );

    \I__2122\ : IoInMux
    port map (
            O => \N__10220\,
            I => \N__10199\
        );

    \I__2121\ : IoInMux
    port map (
            O => \N__10219\,
            I => \N__10196\
        );

    \I__2120\ : IoInMux
    port map (
            O => \N__10218\,
            I => \N__10193\
        );

    \I__2119\ : IoInMux
    port map (
            O => \N__10217\,
            I => \N__10190\
        );

    \I__2118\ : IoInMux
    port map (
            O => \N__10216\,
            I => \N__10181\
        );

    \I__2117\ : IoInMux
    port map (
            O => \N__10215\,
            I => \N__10178\
        );

    \I__2116\ : IoInMux
    port map (
            O => \N__10214\,
            I => \N__10175\
        );

    \I__2115\ : IoInMux
    port map (
            O => \N__10213\,
            I => \N__10169\
        );

    \I__2114\ : IoSpan4Mux
    port map (
            O => \N__10208\,
            I => \N__10155\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__10205\,
            I => \N__10155\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__10202\,
            I => \N__10155\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__10199\,
            I => \N__10155\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__10196\,
            I => \N__10155\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__10193\,
            I => \N__10155\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__10190\,
            I => \N__10152\
        );

    \I__2107\ : IoInMux
    port map (
            O => \N__10189\,
            I => \N__10149\
        );

    \I__2106\ : IoInMux
    port map (
            O => \N__10188\,
            I => \N__10146\
        );

    \I__2105\ : IoInMux
    port map (
            O => \N__10187\,
            I => \N__10143\
        );

    \I__2104\ : IoInMux
    port map (
            O => \N__10186\,
            I => \N__10137\
        );

    \I__2103\ : IoInMux
    port map (
            O => \N__10185\,
            I => \N__10134\
        );

    \I__2102\ : IoInMux
    port map (
            O => \N__10184\,
            I => \N__10131\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__10181\,
            I => \N__10124\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__10178\,
            I => \N__10124\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__10175\,
            I => \N__10124\
        );

    \I__2098\ : IoInMux
    port map (
            O => \N__10174\,
            I => \N__10121\
        );

    \I__2097\ : IoInMux
    port map (
            O => \N__10173\,
            I => \N__10118\
        );

    \I__2096\ : IoInMux
    port map (
            O => \N__10172\,
            I => \N__10115\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__10169\,
            I => \N__10112\
        );

    \I__2094\ : IoInMux
    port map (
            O => \N__10168\,
            I => \N__10109\
        );

    \I__2093\ : IoSpan4Mux
    port map (
            O => \N__10155\,
            I => \N__10095\
        );

    \I__2092\ : IoSpan4Mux
    port map (
            O => \N__10152\,
            I => \N__10095\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__10149\,
            I => \N__10095\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__10146\,
            I => \N__10095\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__10143\,
            I => \N__10095\
        );

    \I__2088\ : IoInMux
    port map (
            O => \N__10142\,
            I => \N__10092\
        );

    \I__2087\ : IoInMux
    port map (
            O => \N__10141\,
            I => \N__10089\
        );

    \I__2086\ : IoInMux
    port map (
            O => \N__10140\,
            I => \N__10086\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__10137\,
            I => \N__10080\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__10134\,
            I => \N__10075\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__10131\,
            I => \N__10075\
        );

    \I__2082\ : IoSpan4Mux
    port map (
            O => \N__10124\,
            I => \N__10066\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__10121\,
            I => \N__10066\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__10118\,
            I => \N__10066\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__10115\,
            I => \N__10066\
        );

    \I__2078\ : IoSpan4Mux
    port map (
            O => \N__10112\,
            I => \N__10061\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__10109\,
            I => \N__10061\
        );

    \I__2076\ : CascadeMux
    port map (
            O => \N__10108\,
            I => \N__10058\
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__10107\,
            I => \N__10054\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__10106\,
            I => \N__10050\
        );

    \I__2073\ : IoSpan4Mux
    port map (
            O => \N__10095\,
            I => \N__10043\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__10092\,
            I => \N__10043\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__10089\,
            I => \N__10043\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__10086\,
            I => \N__10040\
        );

    \I__2069\ : IoInMux
    port map (
            O => \N__10085\,
            I => \N__10037\
        );

    \I__2068\ : IoInMux
    port map (
            O => \N__10084\,
            I => \N__10034\
        );

    \I__2067\ : IoInMux
    port map (
            O => \N__10083\,
            I => \N__10031\
        );

    \I__2066\ : IoSpan4Mux
    port map (
            O => \N__10080\,
            I => \N__10024\
        );

    \I__2065\ : Span4Mux_s3_h
    port map (
            O => \N__10075\,
            I => \N__10021\
        );

    \I__2064\ : IoSpan4Mux
    port map (
            O => \N__10066\,
            I => \N__10016\
        );

    \I__2063\ : IoSpan4Mux
    port map (
            O => \N__10061\,
            I => \N__10016\
        );

    \I__2062\ : InMux
    port map (
            O => \N__10058\,
            I => \N__10005\
        );

    \I__2061\ : InMux
    port map (
            O => \N__10057\,
            I => \N__10005\
        );

    \I__2060\ : InMux
    port map (
            O => \N__10054\,
            I => \N__10005\
        );

    \I__2059\ : InMux
    port map (
            O => \N__10053\,
            I => \N__10005\
        );

    \I__2058\ : InMux
    port map (
            O => \N__10050\,
            I => \N__10005\
        );

    \I__2057\ : IoSpan4Mux
    port map (
            O => \N__10043\,
            I => \N__9996\
        );

    \I__2056\ : IoSpan4Mux
    port map (
            O => \N__10040\,
            I => \N__9996\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__10037\,
            I => \N__9996\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__10034\,
            I => \N__9996\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__10031\,
            I => \N__9993\
        );

    \I__2052\ : IoInMux
    port map (
            O => \N__10030\,
            I => \N__9990\
        );

    \I__2051\ : IoInMux
    port map (
            O => \N__10029\,
            I => \N__9987\
        );

    \I__2050\ : IoInMux
    port map (
            O => \N__10028\,
            I => \N__9984\
        );

    \I__2049\ : IoInMux
    port map (
            O => \N__10027\,
            I => \N__9981\
        );

    \I__2048\ : Span4Mux_s2_v
    port map (
            O => \N__10024\,
            I => \N__9977\
        );

    \I__2047\ : Span4Mux_v
    port map (
            O => \N__10021\,
            I => \N__9972\
        );

    \I__2046\ : Span4Mux_s3_h
    port map (
            O => \N__10016\,
            I => \N__9972\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__10005\,
            I => \N__9969\
        );

    \I__2044\ : IoSpan4Mux
    port map (
            O => \N__9996\,
            I => \N__9966\
        );

    \I__2043\ : IoSpan4Mux
    port map (
            O => \N__9993\,
            I => \N__9955\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9990\,
            I => \N__9955\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__9987\,
            I => \N__9955\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9984\,
            I => \N__9955\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__9981\,
            I => \N__9955\
        );

    \I__2038\ : IoInMux
    port map (
            O => \N__9980\,
            I => \N__9952\
        );

    \I__2037\ : Sp12to4
    port map (
            O => \N__9977\,
            I => \N__9949\
        );

    \I__2036\ : Span4Mux_h
    port map (
            O => \N__9972\,
            I => \N__9946\
        );

    \I__2035\ : Span4Mux_v
    port map (
            O => \N__9969\,
            I => \N__9943\
        );

    \I__2034\ : IoSpan4Mux
    port map (
            O => \N__9966\,
            I => \N__9938\
        );

    \I__2033\ : IoSpan4Mux
    port map (
            O => \N__9955\,
            I => \N__9938\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9952\,
            I => \N__9935\
        );

    \I__2031\ : Span12Mux_v
    port map (
            O => \N__9949\,
            I => \N__9932\
        );

    \I__2030\ : Span4Mux_h
    port map (
            O => \N__9946\,
            I => \N__9927\
        );

    \I__2029\ : Span4Mux_v
    port map (
            O => \N__9943\,
            I => \N__9927\
        );

    \I__2028\ : Span4Mux_s0_v
    port map (
            O => \N__9938\,
            I => \N__9922\
        );

    \I__2027\ : Span4Mux_s0_v
    port map (
            O => \N__9935\,
            I => \N__9922\
        );

    \I__2026\ : Span12Mux_h
    port map (
            O => \N__9932\,
            I => \N__9919\
        );

    \I__2025\ : Sp12to4
    port map (
            O => \N__9927\,
            I => \N__9916\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__9922\,
            I => \N__9913\
        );

    \I__2023\ : Odrv12
    port map (
            O => \N__9919\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2022\ : Odrv12
    port map (
            O => \N__9916\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2021\ : Odrv4
    port map (
            O => \N__9913\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9906\,
            I => \spi0.n2919\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9903\,
            I => \N__9899\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9902\,
            I => \N__9896\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__9899\,
            I => \spi0.spi_clk_counter_1\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9896\,
            I => \spi0.spi_clk_counter_1\
        );

    \I__2015\ : InMux
    port map (
            O => \N__9891\,
            I => \N__9887\
        );

    \I__2014\ : InMux
    port map (
            O => \N__9890\,
            I => \N__9884\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__9887\,
            I => \spi0.spi_clk_counter_5\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__9884\,
            I => \spi0.spi_clk_counter_5\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__9879\,
            I => \N__9876\
        );

    \I__2010\ : InMux
    port map (
            O => \N__9876\,
            I => \N__9873\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__9873\,
            I => \N__9869\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9866\
        );

    \I__2007\ : Odrv12
    port map (
            O => \N__9869\,
            I => \spi0.spi_clk_counter_0\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__9866\,
            I => \spi0.spi_clk_counter_0\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__9861\,
            I => \N__9857\
        );

    \I__2004\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9854\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9857\,
            I => \N__9851\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9854\,
            I => \spi0.spi_clk_counter_2\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9851\,
            I => \spi0.spi_clk_counter_2\
        );

    \I__2000\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9842\
        );

    \I__1999\ : InMux
    port map (
            O => \N__9845\,
            I => \N__9839\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__9842\,
            I => \spi0.spi_clk_counter_3\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__9839\,
            I => \spi0.spi_clk_counter_3\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__9834\,
            I => \spi0.n10_cascade_\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__9831\,
            I => \N__9827\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9824\
        );

    \I__1993\ : InMux
    port map (
            O => \N__9827\,
            I => \N__9821\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__9824\,
            I => \spi0.spi_clk_counter_4\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__9821\,
            I => \spi0.spi_clk_counter_4\
        );

    \I__1990\ : InMux
    port map (
            O => \N__9816\,
            I => \N__9812\
        );

    \I__1989\ : SRMux
    port map (
            O => \N__9815\,
            I => \N__9809\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9812\,
            I => \N__9806\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__9809\,
            I => \N__9803\
        );

    \I__1986\ : Span4Mux_h
    port map (
            O => \N__9806\,
            I => \N__9800\
        );

    \I__1985\ : Span4Mux_v
    port map (
            O => \N__9803\,
            I => \N__9797\
        );

    \I__1984\ : Odrv4
    port map (
            O => \N__9800\,
            I => \spi0.n1896\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__9797\,
            I => \spi0.n1896\
        );

    \I__1982\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9789\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__9789\,
            I => \N__9784\
        );

    \I__1980\ : InMux
    port map (
            O => \N__9788\,
            I => \N__9779\
        );

    \I__1979\ : InMux
    port map (
            O => \N__9787\,
            I => \N__9779\
        );

    \I__1978\ : Odrv12
    port map (
            O => \N__9784\,
            I => tx_data_byte_1
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__9779\,
            I => tx_data_byte_1
        );

    \I__1976\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9771\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__9771\,
            I => \N__9768\
        );

    \I__1974\ : Span4Mux_v
    port map (
            O => \N__9768\,
            I => \N__9764\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9761\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__9764\,
            I => tx_addr_byte_1
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__9761\,
            I => tx_addr_byte_1
        );

    \I__1970\ : InMux
    port map (
            O => \N__9756\,
            I => \N__9751\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9748\
        );

    \I__1968\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9745\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__9751\,
            I => \spi0.state_next_2__N_310\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__9748\,
            I => \spi0.state_next_2__N_310\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__9745\,
            I => \spi0.state_next_2__N_310\
        );

    \I__1964\ : InMux
    port map (
            O => \N__9738\,
            I => \N__9719\
        );

    \I__1963\ : InMux
    port map (
            O => \N__9737\,
            I => \N__9719\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9736\,
            I => \N__9712\
        );

    \I__1961\ : InMux
    port map (
            O => \N__9735\,
            I => \N__9712\
        );

    \I__1960\ : InMux
    port map (
            O => \N__9734\,
            I => \N__9712\
        );

    \I__1959\ : InMux
    port map (
            O => \N__9733\,
            I => \N__9705\
        );

    \I__1958\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9705\
        );

    \I__1957\ : InMux
    port map (
            O => \N__9731\,
            I => \N__9705\
        );

    \I__1956\ : InMux
    port map (
            O => \N__9730\,
            I => \N__9696\
        );

    \I__1955\ : InMux
    port map (
            O => \N__9729\,
            I => \N__9696\
        );

    \I__1954\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9696\
        );

    \I__1953\ : InMux
    port map (
            O => \N__9727\,
            I => \N__9696\
        );

    \I__1952\ : InMux
    port map (
            O => \N__9726\,
            I => \N__9689\
        );

    \I__1951\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9689\
        );

    \I__1950\ : InMux
    port map (
            O => \N__9724\,
            I => \N__9689\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__9719\,
            I => \spi0.n4\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__9712\,
            I => \spi0.n4\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__9705\,
            I => \spi0.n4\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__9696\,
            I => \spi0.n4\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__9689\,
            I => \spi0.n4\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__9678\,
            I => \N__9668\
        );

    \I__1943\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9657\
        );

    \I__1942\ : InMux
    port map (
            O => \N__9676\,
            I => \N__9652\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9675\,
            I => \N__9652\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9674\,
            I => \N__9649\
        );

    \I__1939\ : InMux
    port map (
            O => \N__9673\,
            I => \N__9638\
        );

    \I__1938\ : InMux
    port map (
            O => \N__9672\,
            I => \N__9638\
        );

    \I__1937\ : InMux
    port map (
            O => \N__9671\,
            I => \N__9638\
        );

    \I__1936\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9638\
        );

    \I__1935\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9638\
        );

    \I__1934\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9623\
        );

    \I__1933\ : InMux
    port map (
            O => \N__9665\,
            I => \N__9623\
        );

    \I__1932\ : InMux
    port map (
            O => \N__9664\,
            I => \N__9623\
        );

    \I__1931\ : InMux
    port map (
            O => \N__9663\,
            I => \N__9623\
        );

    \I__1930\ : InMux
    port map (
            O => \N__9662\,
            I => \N__9623\
        );

    \I__1929\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9623\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9623\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__9657\,
            I => \spi0.state_next_1\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__9652\,
            I => \spi0.state_next_1\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__9649\,
            I => \spi0.state_next_1\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9638\,
            I => \spi0.state_next_1\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__9623\,
            I => \spi0.state_next_1\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__9612\,
            I => \N__9609\
        );

    \I__1921\ : InMux
    port map (
            O => \N__9609\,
            I => \N__9606\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__9606\,
            I => \N__9603\
        );

    \I__1919\ : Span4Mux_h
    port map (
            O => \N__9603\,
            I => \N__9600\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__9600\,
            I => \spi0.n499\
        );

    \I__1917\ : InMux
    port map (
            O => \N__9597\,
            I => \N__9584\
        );

    \I__1916\ : InMux
    port map (
            O => \N__9596\,
            I => \N__9581\
        );

    \I__1915\ : InMux
    port map (
            O => \N__9595\,
            I => \N__9578\
        );

    \I__1914\ : InMux
    port map (
            O => \N__9594\,
            I => \N__9574\
        );

    \I__1913\ : SRMux
    port map (
            O => \N__9593\,
            I => \N__9570\
        );

    \I__1912\ : SRMux
    port map (
            O => \N__9592\,
            I => \N__9564\
        );

    \I__1911\ : SRMux
    port map (
            O => \N__9591\,
            I => \N__9561\
        );

    \I__1910\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9558\
        );

    \I__1909\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9551\
        );

    \I__1908\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9551\
        );

    \I__1907\ : SRMux
    port map (
            O => \N__9587\,
            I => \N__9551\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__9584\,
            I => \N__9544\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__9581\,
            I => \N__9544\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__9578\,
            I => \N__9544\
        );

    \I__1903\ : SRMux
    port map (
            O => \N__9577\,
            I => \N__9541\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__9574\,
            I => \N__9537\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__9573\,
            I => \N__9533\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__9570\,
            I => \N__9527\
        );

    \I__1899\ : InMux
    port map (
            O => \N__9569\,
            I => \N__9520\
        );

    \I__1898\ : InMux
    port map (
            O => \N__9568\,
            I => \N__9520\
        );

    \I__1897\ : InMux
    port map (
            O => \N__9567\,
            I => \N__9520\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__9564\,
            I => \N__9515\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__9561\,
            I => \N__9515\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__9558\,
            I => \N__9510\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__9551\,
            I => \N__9510\
        );

    \I__1892\ : Span4Mux_v
    port map (
            O => \N__9544\,
            I => \N__9505\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__9541\,
            I => \N__9505\
        );

    \I__1890\ : SRMux
    port map (
            O => \N__9540\,
            I => \N__9502\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__9537\,
            I => \N__9499\
        );

    \I__1888\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9494\
        );

    \I__1887\ : InMux
    port map (
            O => \N__9533\,
            I => \N__9494\
        );

    \I__1886\ : InMux
    port map (
            O => \N__9532\,
            I => \N__9490\
        );

    \I__1885\ : InMux
    port map (
            O => \N__9531\,
            I => \N__9487\
        );

    \I__1884\ : InMux
    port map (
            O => \N__9530\,
            I => \N__9484\
        );

    \I__1883\ : Span4Mux_v
    port map (
            O => \N__9527\,
            I => \N__9478\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__9520\,
            I => \N__9475\
        );

    \I__1881\ : Span4Mux_v
    port map (
            O => \N__9515\,
            I => \N__9472\
        );

    \I__1880\ : Span4Mux_v
    port map (
            O => \N__9510\,
            I => \N__9469\
        );

    \I__1879\ : Span4Mux_v
    port map (
            O => \N__9505\,
            I => \N__9464\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__9502\,
            I => \N__9464\
        );

    \I__1877\ : Span4Mux_h
    port map (
            O => \N__9499\,
            I => \N__9459\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__9494\,
            I => \N__9459\
        );

    \I__1875\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9456\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__9490\,
            I => \N__9449\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__9487\,
            I => \N__9449\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__9484\,
            I => \N__9449\
        );

    \I__1871\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9442\
        );

    \I__1870\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9442\
        );

    \I__1869\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9442\
        );

    \I__1868\ : Span4Mux_h
    port map (
            O => \N__9478\,
            I => \N__9437\
        );

    \I__1867\ : Span4Mux_v
    port map (
            O => \N__9475\,
            I => \N__9437\
        );

    \I__1866\ : Span4Mux_h
    port map (
            O => \N__9472\,
            I => \N__9430\
        );

    \I__1865\ : Span4Mux_v
    port map (
            O => \N__9469\,
            I => \N__9430\
        );

    \I__1864\ : Span4Mux_h
    port map (
            O => \N__9464\,
            I => \N__9430\
        );

    \I__1863\ : Span4Mux_v
    port map (
            O => \N__9459\,
            I => \N__9425\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__9456\,
            I => \N__9425\
        );

    \I__1861\ : Span12Mux_h
    port map (
            O => \N__9449\,
            I => \N__9420\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__9442\,
            I => \N__9420\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__9437\,
            I => reset_all_w
        );

    \I__1858\ : Odrv4
    port map (
            O => \N__9430\,
            I => reset_all_w
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__9425\,
            I => reset_all_w
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__9420\,
            I => reset_all_w
        );

    \I__1855\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9407\
        );

    \I__1854\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9403\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__9407\,
            I => \N__9390\
        );

    \I__1852\ : InMux
    port map (
            O => \N__9406\,
            I => \N__9387\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__9403\,
            I => \N__9384\
        );

    \I__1850\ : InMux
    port map (
            O => \N__9402\,
            I => \N__9379\
        );

    \I__1849\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9379\
        );

    \I__1848\ : InMux
    port map (
            O => \N__9400\,
            I => \N__9372\
        );

    \I__1847\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9372\
        );

    \I__1846\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9372\
        );

    \I__1845\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9367\
        );

    \I__1844\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9367\
        );

    \I__1843\ : InMux
    port map (
            O => \N__9395\,
            I => \N__9364\
        );

    \I__1842\ : InMux
    port map (
            O => \N__9394\,
            I => \N__9359\
        );

    \I__1841\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9359\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__9390\,
            I => state_reg_0
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__9387\,
            I => state_reg_0
        );

    \I__1838\ : Odrv4
    port map (
            O => \N__9384\,
            I => state_reg_0
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__9379\,
            I => state_reg_0
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__9372\,
            I => state_reg_0
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__9367\,
            I => state_reg_0
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__9364\,
            I => state_reg_0
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__9359\,
            I => state_reg_0
        );

    \I__1832\ : InMux
    port map (
            O => \N__9342\,
            I => \N__9338\
        );

    \I__1831\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9335\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__9338\,
            I => \N__9318\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__9335\,
            I => \N__9315\
        );

    \I__1828\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9308\
        );

    \I__1827\ : InMux
    port map (
            O => \N__9333\,
            I => \N__9308\
        );

    \I__1826\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9308\
        );

    \I__1825\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9305\
        );

    \I__1824\ : InMux
    port map (
            O => \N__9330\,
            I => \N__9298\
        );

    \I__1823\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9298\
        );

    \I__1822\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9298\
        );

    \I__1821\ : InMux
    port map (
            O => \N__9327\,
            I => \N__9295\
        );

    \I__1820\ : InMux
    port map (
            O => \N__9326\,
            I => \N__9284\
        );

    \I__1819\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9284\
        );

    \I__1818\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9284\
        );

    \I__1817\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9284\
        );

    \I__1816\ : InMux
    port map (
            O => \N__9322\,
            I => \N__9284\
        );

    \I__1815\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9281\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__9318\,
            I => state_reg_2
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__9315\,
            I => state_reg_2
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__9308\,
            I => state_reg_2
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__9305\,
            I => state_reg_2
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__9298\,
            I => state_reg_2
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__9295\,
            I => state_reg_2
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__9284\,
            I => state_reg_2
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__9281\,
            I => state_reg_2
        );

    \I__1806\ : SRMux
    port map (
            O => \N__9264\,
            I => \N__9261\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__9261\,
            I => \N__9257\
        );

    \I__1804\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9241\
        );

    \I__1803\ : Span4Mux_v
    port map (
            O => \N__9257\,
            I => \N__9222\
        );

    \I__1802\ : InMux
    port map (
            O => \N__9256\,
            I => \N__9209\
        );

    \I__1801\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9209\
        );

    \I__1800\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9209\
        );

    \I__1799\ : InMux
    port map (
            O => \N__9253\,
            I => \N__9209\
        );

    \I__1798\ : InMux
    port map (
            O => \N__9252\,
            I => \N__9209\
        );

    \I__1797\ : InMux
    port map (
            O => \N__9251\,
            I => \N__9209\
        );

    \I__1796\ : InMux
    port map (
            O => \N__9250\,
            I => \N__9194\
        );

    \I__1795\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9194\
        );

    \I__1794\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9194\
        );

    \I__1793\ : InMux
    port map (
            O => \N__9247\,
            I => \N__9194\
        );

    \I__1792\ : InMux
    port map (
            O => \N__9246\,
            I => \N__9194\
        );

    \I__1791\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9194\
        );

    \I__1790\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9194\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__9241\,
            I => \N__9191\
        );

    \I__1788\ : InMux
    port map (
            O => \N__9240\,
            I => \N__9182\
        );

    \I__1787\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9182\
        );

    \I__1786\ : InMux
    port map (
            O => \N__9238\,
            I => \N__9182\
        );

    \I__1785\ : InMux
    port map (
            O => \N__9237\,
            I => \N__9182\
        );

    \I__1784\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9171\
        );

    \I__1783\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9171\
        );

    \I__1782\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9171\
        );

    \I__1781\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9171\
        );

    \I__1780\ : InMux
    port map (
            O => \N__9232\,
            I => \N__9171\
        );

    \I__1779\ : InMux
    port map (
            O => \N__9231\,
            I => \N__9168\
        );

    \I__1778\ : InMux
    port map (
            O => \N__9230\,
            I => \N__9157\
        );

    \I__1777\ : InMux
    port map (
            O => \N__9229\,
            I => \N__9157\
        );

    \I__1776\ : InMux
    port map (
            O => \N__9228\,
            I => \N__9157\
        );

    \I__1775\ : InMux
    port map (
            O => \N__9227\,
            I => \N__9157\
        );

    \I__1774\ : InMux
    port map (
            O => \N__9226\,
            I => \N__9157\
        );

    \I__1773\ : InMux
    port map (
            O => \N__9225\,
            I => \N__9154\
        );

    \I__1772\ : Odrv4
    port map (
            O => \N__9222\,
            I => state_reg_1
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__9209\,
            I => state_reg_1
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__9194\,
            I => state_reg_1
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__9191\,
            I => state_reg_1
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__9182\,
            I => state_reg_1
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__9171\,
            I => state_reg_1
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__9168\,
            I => state_reg_1
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__9157\,
            I => state_reg_1
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__9154\,
            I => state_reg_1
        );

    \I__1763\ : IoInMux
    port map (
            O => \N__9135\,
            I => \N__9132\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__9132\,
            I => \N__9129\
        );

    \I__1761\ : Span12Mux_s8_v
    port map (
            O => \N__9129\,
            I => \N__9126\
        );

    \I__1760\ : Span12Mux_h
    port map (
            O => \N__9126\,
            I => \N__9122\
        );

    \I__1759\ : InMux
    port map (
            O => \N__9125\,
            I => \N__9119\
        );

    \I__1758\ : Odrv12
    port map (
            O => \N__9122\,
            I => \SEN_c\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__9119\,
            I => \SEN_c\
        );

    \I__1756\ : IoInMux
    port map (
            O => \N__9114\,
            I => \N__9111\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__9111\,
            I => \N__9107\
        );

    \I__1754\ : IoInMux
    port map (
            O => \N__9110\,
            I => \N__9104\
        );

    \I__1753\ : IoSpan4Mux
    port map (
            O => \N__9107\,
            I => \N__9101\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__9104\,
            I => \N__9098\
        );

    \I__1751\ : Span4Mux_s1_h
    port map (
            O => \N__9101\,
            I => \N__9095\
        );

    \I__1750\ : Span4Mux_s2_v
    port map (
            O => \N__9098\,
            I => \N__9092\
        );

    \I__1749\ : Sp12to4
    port map (
            O => \N__9095\,
            I => \N__9089\
        );

    \I__1748\ : Span4Mux_h
    port map (
            O => \N__9092\,
            I => \N__9086\
        );

    \I__1747\ : Span12Mux_h
    port map (
            O => \N__9089\,
            I => \N__9083\
        );

    \I__1746\ : Sp12to4
    port map (
            O => \N__9086\,
            I => \N__9080\
        );

    \I__1745\ : Span12Mux_v
    port map (
            O => \N__9083\,
            I => \N__9075\
        );

    \I__1744\ : Span12Mux_h
    port map (
            O => \N__9080\,
            I => \N__9075\
        );

    \I__1743\ : Odrv12
    port map (
            O => \N__9075\,
            I => \DEBUG_6_c\
        );

    \I__1742\ : InMux
    port map (
            O => \N__9072\,
            I => \N__9069\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__9069\,
            I => \N__9065\
        );

    \I__1740\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9062\
        );

    \I__1739\ : Span4Mux_h
    port map (
            O => \N__9065\,
            I => \N__9059\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__9062\,
            I => \N__9056\
        );

    \I__1737\ : Span4Mux_v
    port map (
            O => \N__9059\,
            I => \N__9052\
        );

    \I__1736\ : Span4Mux_h
    port map (
            O => \N__9056\,
            I => \N__9049\
        );

    \I__1735\ : InMux
    port map (
            O => \N__9055\,
            I => \N__9046\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__9052\,
            I => tx_data_byte_4
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__9049\,
            I => tx_data_byte_4
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__9046\,
            I => tx_data_byte_4
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__9039\,
            I => \N__9036\
        );

    \I__1730\ : InMux
    port map (
            O => \N__9036\,
            I => \N__9033\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__9033\,
            I => \N__9029\
        );

    \I__1728\ : InMux
    port map (
            O => \N__9032\,
            I => \N__9026\
        );

    \I__1727\ : Span4Mux_v
    port map (
            O => \N__9029\,
            I => \N__9020\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__9026\,
            I => \N__9020\
        );

    \I__1725\ : InMux
    port map (
            O => \N__9025\,
            I => \N__9017\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__9020\,
            I => tx_data_byte_6
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__9017\,
            I => tx_data_byte_6
        );

    \I__1722\ : InMux
    port map (
            O => \N__9012\,
            I => \N__9009\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__9009\,
            I => \N__9006\
        );

    \I__1720\ : Odrv12
    port map (
            O => \N__9006\,
            I => start_transfer_prev
        );

    \I__1719\ : InMux
    port map (
            O => \N__9003\,
            I => \N__9000\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__9000\,
            I => \N__8997\
        );

    \I__1717\ : Span4Mux_v
    port map (
            O => \N__8997\,
            I => \N__8993\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8990\
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__8993\,
            I => n5_adj_507
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8990\,
            I => n5_adj_507
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__8985\,
            I => \N__8982\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8982\,
            I => \N__8979\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8979\,
            I => \N__8976\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__8976\,
            I => \N__8972\
        );

    \I__1709\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8969\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__8972\,
            I => start_transfer_edge
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__8969\,
            I => start_transfer_edge
        );

    \I__1706\ : InMux
    port map (
            O => \N__8964\,
            I => \bfn_17_14_0_\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8961\,
            I => \spi0.n2915\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8958\,
            I => \N__8952\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8957\,
            I => \N__8952\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8952\,
            I => \N__8949\
        );

    \I__1701\ : Odrv12
    port map (
            O => \N__8949\,
            I => spi_busy
        );

    \I__1700\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8941\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8945\,
            I => \N__8938\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8944\,
            I => \N__8935\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8941\,
            I => \N__8929\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__8938\,
            I => \N__8929\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8935\,
            I => \N__8926\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8934\,
            I => \N__8923\
        );

    \I__1693\ : Span4Mux_v
    port map (
            O => \N__8929\,
            I => \N__8920\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__8926\,
            I => \N__8917\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__8923\,
            I => \N__8914\
        );

    \I__1690\ : Span4Mux_h
    port map (
            O => \N__8920\,
            I => \N__8910\
        );

    \I__1689\ : Span4Mux_h
    port map (
            O => \N__8917\,
            I => \N__8905\
        );

    \I__1688\ : Span4Mux_v
    port map (
            O => \N__8914\,
            I => \N__8905\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8902\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__8910\,
            I => rx_buf_byte_6
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__8905\,
            I => rx_buf_byte_6
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__8902\,
            I => rx_buf_byte_6
        );

    \I__1683\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8890\
        );

    \I__1682\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8887\
        );

    \I__1681\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8883\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8890\,
            I => \N__8878\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8887\,
            I => \N__8878\
        );

    \I__1678\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8875\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8883\,
            I => \N__8872\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__8878\,
            I => \N__8867\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__8875\,
            I => \N__8867\
        );

    \I__1674\ : Span4Mux_v
    port map (
            O => \N__8872\,
            I => \N__8863\
        );

    \I__1673\ : Span4Mux_h
    port map (
            O => \N__8867\,
            I => \N__8860\
        );

    \I__1672\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8857\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__8863\,
            I => rx_buf_byte_3
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__8860\,
            I => rx_buf_byte_3
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8857\,
            I => rx_buf_byte_3
        );

    \I__1668\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8847\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__8847\,
            I => \spi0.n906\
        );

    \I__1666\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8837\
        );

    \I__1665\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8834\
        );

    \I__1664\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8827\
        );

    \I__1663\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8827\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8840\,
            I => \N__8827\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__8837\,
            I => n883
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__8834\,
            I => n883
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__8827\,
            I => n883
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__8820\,
            I => \spi0.n906_cascade_\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__8817\,
            I => \N__8814\
        );

    \I__1656\ : InMux
    port map (
            O => \N__8814\,
            I => \N__8811\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__8811\,
            I => \N__8808\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__8808\,
            I => \spi0.n492\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__8805\,
            I => \N__8802\
        );

    \I__1652\ : InMux
    port map (
            O => \N__8802\,
            I => \N__8799\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8799\,
            I => \N__8796\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__8796\,
            I => \spi0.n493\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__8793\,
            I => \N__8790\
        );

    \I__1648\ : InMux
    port map (
            O => \N__8790\,
            I => \N__8787\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__8787\,
            I => \spi0.n494\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__8784\,
            I => \N__8781\
        );

    \I__1645\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8776\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__8780\,
            I => \N__8772\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__8779\,
            I => \N__8769\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__8776\,
            I => \N__8766\
        );

    \I__1641\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8763\
        );

    \I__1640\ : InMux
    port map (
            O => \N__8772\,
            I => \N__8760\
        );

    \I__1639\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8757\
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__8766\,
            I => \state_next_2__N_312\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__8763\,
            I => \state_next_2__N_312\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__8760\,
            I => \state_next_2__N_312\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__8757\,
            I => \state_next_2__N_312\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__8748\,
            I => \N__8745\
        );

    \I__1633\ : InMux
    port map (
            O => \N__8745\,
            I => \N__8742\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__8742\,
            I => \spi0.n495\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__8739\,
            I => \N__8736\
        );

    \I__1630\ : InMux
    port map (
            O => \N__8736\,
            I => \N__8733\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__8733\,
            I => \spi0.n502\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8730\,
            I => \N__8724\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8729\,
            I => \N__8724\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__8724\,
            I => \spi0.state_next_2__N_311\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__8721\,
            I => \N__8718\
        );

    \I__1624\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8715\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8715\,
            I => \spi0.n487\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__8712\,
            I => \N__8709\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8709\,
            I => \N__8706\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__8706\,
            I => \spi0.n488\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__8703\,
            I => \N__8700\
        );

    \I__1618\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8697\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__8697\,
            I => \spi0.n489\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__8694\,
            I => \N__8691\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8691\,
            I => \N__8688\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__8688\,
            I => \spi0.n490\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__8685\,
            I => \N__8682\
        );

    \I__1612\ : InMux
    port map (
            O => \N__8682\,
            I => \N__8679\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__8679\,
            I => \spi0.n491\
        );

    \I__1610\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8673\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__8673\,
            I => \N__8670\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__8670\,
            I => \N__8666\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8663\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__8666\,
            I => rx_shift_reg_1
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__8663\,
            I => rx_shift_reg_1
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__8658\,
            I => \rx_shift_reg_15__N_319_cascade_\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__8655\,
            I => \N__8651\
        );

    \I__1602\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8646\
        );

    \I__1601\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8643\
        );

    \I__1600\ : InMux
    port map (
            O => \N__8650\,
            I => \N__8640\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8637\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__8646\,
            I => \N__8634\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__8643\,
            I => \N__8631\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__8640\,
            I => \N__8628\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__8637\,
            I => \N__8625\
        );

    \I__1594\ : Span4Mux_v
    port map (
            O => \N__8634\,
            I => \N__8622\
        );

    \I__1593\ : Span4Mux_h
    port map (
            O => \N__8631\,
            I => \N__8617\
        );

    \I__1592\ : Span4Mux_v
    port map (
            O => \N__8628\,
            I => \N__8617\
        );

    \I__1591\ : Span4Mux_v
    port map (
            O => \N__8625\,
            I => \N__8614\
        );

    \I__1590\ : Span4Mux_v
    port map (
            O => \N__8622\,
            I => \N__8610\
        );

    \I__1589\ : Span4Mux_v
    port map (
            O => \N__8617\,
            I => \N__8605\
        );

    \I__1588\ : Span4Mux_h
    port map (
            O => \N__8614\,
            I => \N__8605\
        );

    \I__1587\ : InMux
    port map (
            O => \N__8613\,
            I => \N__8602\
        );

    \I__1586\ : Odrv4
    port map (
            O => \N__8610\,
            I => rx_buf_byte_0
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__8605\,
            I => rx_buf_byte_0
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__8602\,
            I => rx_buf_byte_0
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__8595\,
            I => \N__8590\
        );

    \I__1582\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8586\
        );

    \I__1581\ : InMux
    port map (
            O => \N__8593\,
            I => \N__8579\
        );

    \I__1580\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8579\
        );

    \I__1579\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8579\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__8586\,
            I => \N__8574\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__8579\,
            I => \N__8574\
        );

    \I__1576\ : Span4Mux_h
    port map (
            O => \N__8574\,
            I => \N__8570\
        );

    \I__1575\ : InMux
    port map (
            O => \N__8573\,
            I => \N__8567\
        );

    \I__1574\ : Odrv4
    port map (
            O => \N__8570\,
            I => rx_buf_byte_1
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__8567\,
            I => rx_buf_byte_1
        );

    \I__1572\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__8559\,
            I => \spi0.state_next_2\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__8556\,
            I => \spi0.state_next_0_cascade_\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__8553\,
            I => \spi0.n4_cascade_\
        );

    \I__1568\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8547\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__8547\,
            I => \spi0.CS_w\
        );

    \I__1566\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8541\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__8541\,
            I => spi_busy_prev
        );

    \I__1564\ : InMux
    port map (
            O => \N__8538\,
            I => \N__8535\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__8535\,
            I => spi_busy_falling_edge
        );

    \I__1562\ : InMux
    port map (
            O => \N__8532\,
            I => \N__8529\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__8529\,
            I => \N__8524\
        );

    \I__1560\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8521\
        );

    \I__1559\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8518\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__8524\,
            I => tx_data_byte_0
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__8521\,
            I => tx_data_byte_0
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__8518\,
            I => tx_data_byte_0
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__8511\,
            I => \N__8508\
        );

    \I__1554\ : InMux
    port map (
            O => \N__8508\,
            I => \N__8505\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__8505\,
            I => \N__8502\
        );

    \I__1552\ : Span4Mux_h
    port map (
            O => \N__8502\,
            I => \N__8498\
        );

    \I__1551\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8495\
        );

    \I__1550\ : Odrv4
    port map (
            O => \N__8498\,
            I => tx_addr_byte_5
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__8495\,
            I => tx_addr_byte_5
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__8490\,
            I => \N__8487\
        );

    \I__1547\ : InMux
    port map (
            O => \N__8487\,
            I => \N__8484\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__8484\,
            I => \spi0.n497\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__8481\,
            I => \N__8478\
        );

    \I__1544\ : InMux
    port map (
            O => \N__8478\,
            I => \N__8475\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__8475\,
            I => \spi0.n498\
        );

    \I__1542\ : CascadeMux
    port map (
            O => \N__8472\,
            I => \n883_cascade_\
        );

    \I__1541\ : InMux
    port map (
            O => \N__8469\,
            I => \N__8466\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__8466\,
            I => \spi0.n2433\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__8463\,
            I => \spi0.n3337_cascade_\
        );

    \I__1538\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8457\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__8457\,
            I => \spi0.n13\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__8454\,
            I => \N__8450\
        );

    \I__1535\ : InMux
    port map (
            O => \N__8453\,
            I => \N__8446\
        );

    \I__1534\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8441\
        );

    \I__1533\ : InMux
    port map (
            O => \N__8449\,
            I => \N__8441\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__8446\,
            I => \spi0.n1429\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__8441\,
            I => \spi0.n1429\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__8436\,
            I => \spi0.n13_cascade_\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__8433\,
            I => \N__8429\
        );

    \I__1528\ : CascadeMux
    port map (
            O => \N__8432\,
            I => \N__8426\
        );

    \I__1527\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8421\
        );

    \I__1526\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8421\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__8421\,
            I => \N__8417\
        );

    \I__1524\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8414\
        );

    \I__1523\ : Span4Mux_v
    port map (
            O => \N__8417\,
            I => \N__8405\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__8414\,
            I => \N__8405\
        );

    \I__1521\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8402\
        );

    \I__1520\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8395\
        );

    \I__1519\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8395\
        );

    \I__1518\ : InMux
    port map (
            O => \N__8410\,
            I => \N__8395\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__8405\,
            I => is_tx_fifo_full_flag
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__8402\,
            I => is_tx_fifo_full_flag
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__8395\,
            I => is_tx_fifo_full_flag
        );

    \I__1514\ : InMux
    port map (
            O => \N__8388\,
            I => \N__8383\
        );

    \I__1513\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8378\
        );

    \I__1512\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8378\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__8383\,
            I => \N__8374\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__8378\,
            I => \N__8371\
        );

    \I__1509\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8368\
        );

    \I__1508\ : Span4Mux_v
    port map (
            O => \N__8374\,
            I => \N__8363\
        );

    \I__1507\ : Span12Mux_v
    port map (
            O => \N__8371\,
            I => \N__8358\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__8368\,
            I => \N__8358\
        );

    \I__1505\ : InMux
    port map (
            O => \N__8367\,
            I => \N__8355\
        );

    \I__1504\ : InMux
    port map (
            O => \N__8366\,
            I => \N__8352\
        );

    \I__1503\ : Odrv4
    port map (
            O => \N__8363\,
            I => fifo_write_cmd
        );

    \I__1502\ : Odrv12
    port map (
            O => \N__8358\,
            I => fifo_write_cmd
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__8355\,
            I => fifo_write_cmd
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__8352\,
            I => fifo_write_cmd
        );

    \I__1499\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8339\
        );

    \I__1498\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8336\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__8339\,
            I => wr_fifo_en_w
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__8336\,
            I => wr_fifo_en_w
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__8331\,
            I => \wr_fifo_en_w_cascade_\
        );

    \I__1494\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8319\
        );

    \I__1493\ : InMux
    port map (
            O => \N__8327\,
            I => \N__8319\
        );

    \I__1492\ : InMux
    port map (
            O => \N__8326\,
            I => \N__8314\
        );

    \I__1491\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8314\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__8324\,
            I => \N__8311\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__8319\,
            I => \N__8308\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__8314\,
            I => \N__8305\
        );

    \I__1487\ : InMux
    port map (
            O => \N__8311\,
            I => \N__8302\
        );

    \I__1486\ : Span4Mux_v
    port map (
            O => \N__8308\,
            I => \N__8290\
        );

    \I__1485\ : Span4Mux_h
    port map (
            O => \N__8305\,
            I => \N__8290\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__8302\,
            I => \N__8290\
        );

    \I__1483\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8287\
        );

    \I__1482\ : InMux
    port map (
            O => \N__8300\,
            I => \N__8282\
        );

    \I__1481\ : InMux
    port map (
            O => \N__8299\,
            I => \N__8282\
        );

    \I__1480\ : InMux
    port map (
            O => \N__8298\,
            I => \N__8277\
        );

    \I__1479\ : InMux
    port map (
            O => \N__8297\,
            I => \N__8277\
        );

    \I__1478\ : Odrv4
    port map (
            O => \N__8290\,
            I => wr_addr_r_0
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__8287\,
            I => wr_addr_r_0
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__8282\,
            I => wr_addr_r_0
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__8277\,
            I => wr_addr_r_0
        );

    \I__1474\ : InMux
    port map (
            O => \N__8268\,
            I => \N__8252\
        );

    \I__1473\ : InMux
    port map (
            O => \N__8267\,
            I => \N__8249\
        );

    \I__1472\ : InMux
    port map (
            O => \N__8266\,
            I => \N__8246\
        );

    \I__1471\ : InMux
    port map (
            O => \N__8265\,
            I => \N__8234\
        );

    \I__1470\ : InMux
    port map (
            O => \N__8264\,
            I => \N__8234\
        );

    \I__1469\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8234\
        );

    \I__1468\ : InMux
    port map (
            O => \N__8262\,
            I => \N__8234\
        );

    \I__1467\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8229\
        );

    \I__1466\ : InMux
    port map (
            O => \N__8260\,
            I => \N__8229\
        );

    \I__1465\ : InMux
    port map (
            O => \N__8259\,
            I => \N__8226\
        );

    \I__1464\ : InMux
    port map (
            O => \N__8258\,
            I => \N__8221\
        );

    \I__1463\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8221\
        );

    \I__1462\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8216\
        );

    \I__1461\ : InMux
    port map (
            O => \N__8255\,
            I => \N__8216\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__8252\,
            I => \N__8209\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__8249\,
            I => \N__8209\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__8246\,
            I => \N__8206\
        );

    \I__1457\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8199\
        );

    \I__1456\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8199\
        );

    \I__1455\ : InMux
    port map (
            O => \N__8243\,
            I => \N__8199\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__8234\,
            I => \N__8191\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__8229\,
            I => \N__8191\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__8226\,
            I => \N__8191\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__8221\,
            I => \N__8186\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__8216\,
            I => \N__8186\
        );

    \I__1449\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8181\
        );

    \I__1448\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8181\
        );

    \I__1447\ : Span4Mux_v
    port map (
            O => \N__8209\,
            I => \N__8172\
        );

    \I__1446\ : Span4Mux_v
    port map (
            O => \N__8206\,
            I => \N__8172\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__8199\,
            I => \N__8169\
        );

    \I__1444\ : InMux
    port map (
            O => \N__8198\,
            I => \N__8166\
        );

    \I__1443\ : Span4Mux_v
    port map (
            O => \N__8191\,
            I => \N__8159\
        );

    \I__1442\ : Span4Mux_v
    port map (
            O => \N__8186\,
            I => \N__8159\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__8181\,
            I => \N__8159\
        );

    \I__1440\ : InMux
    port map (
            O => \N__8180\,
            I => \N__8154\
        );

    \I__1439\ : InMux
    port map (
            O => \N__8179\,
            I => \N__8154\
        );

    \I__1438\ : InMux
    port map (
            O => \N__8178\,
            I => \N__8149\
        );

    \I__1437\ : InMux
    port map (
            O => \N__8177\,
            I => \N__8149\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__8172\,
            I => wr_addr_r_1
        );

    \I__1435\ : Odrv12
    port map (
            O => \N__8169\,
            I => wr_addr_r_1
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__8166\,
            I => wr_addr_r_1
        );

    \I__1433\ : Odrv4
    port map (
            O => \N__8159\,
            I => wr_addr_r_1
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__8154\,
            I => wr_addr_r_1
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__8149\,
            I => wr_addr_r_1
        );

    \I__1430\ : InMux
    port map (
            O => \N__8136\,
            I => \N__8133\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__8133\,
            I => \N__8130\
        );

    \I__1428\ : Span4Mux_v
    port map (
            O => \N__8130\,
            I => \N__8126\
        );

    \I__1427\ : InMux
    port map (
            O => \N__8129\,
            I => \N__8123\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__8126\,
            I => tx_addr_byte_6
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__8123\,
            I => tx_addr_byte_6
        );

    \I__1424\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8115\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__8115\,
            I => tx_shift_reg_0
        );

    \I__1422\ : SRMux
    port map (
            O => \N__8112\,
            I => \N__8109\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__8109\,
            I => \spi0.n890\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__8106\,
            I => \spi0.n3328_cascade_\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__8103\,
            I => \spi0.n1429_cascade_\
        );

    \I__1418\ : InMux
    port map (
            O => \N__8100\,
            I => \N__8097\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__8097\,
            I => \spi0.n3328\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__8094\,
            I => \tx_fifo.lscc_fifo_inst.n2_cascade_\
        );

    \I__1415\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8088\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__8088\,
            I => \N__8083\
        );

    \I__1413\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8080\
        );

    \I__1412\ : InMux
    port map (
            O => \N__8086\,
            I => \N__8077\
        );

    \I__1411\ : Odrv4
    port map (
            O => \N__8083\,
            I => rd_addr_r_2
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__8080\,
            I => rd_addr_r_2
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__8077\,
            I => rd_addr_r_2
        );

    \I__1408\ : InMux
    port map (
            O => \N__8070\,
            I => \N__8067\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__8067\,
            I => wr_addr_p1_w_2
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__8064\,
            I => \wr_addr_p1_w_2_cascade_\
        );

    \I__1405\ : InMux
    port map (
            O => \N__8061\,
            I => \N__8058\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__8058\,
            I => \N__8053\
        );

    \I__1403\ : InMux
    port map (
            O => \N__8057\,
            I => \N__8048\
        );

    \I__1402\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8048\
        );

    \I__1401\ : Odrv4
    port map (
            O => \N__8053\,
            I => wr_addr_r_2
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__8048\,
            I => wr_addr_r_2
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__8043\,
            I => \N__8034\
        );

    \I__1398\ : InMux
    port map (
            O => \N__8042\,
            I => \N__8031\
        );

    \I__1397\ : InMux
    port map (
            O => \N__8041\,
            I => \N__8020\
        );

    \I__1396\ : InMux
    port map (
            O => \N__8040\,
            I => \N__8020\
        );

    \I__1395\ : InMux
    port map (
            O => \N__8039\,
            I => \N__8020\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__8038\,
            I => \N__8017\
        );

    \I__1393\ : InMux
    port map (
            O => \N__8037\,
            I => \N__8014\
        );

    \I__1392\ : InMux
    port map (
            O => \N__8034\,
            I => \N__8011\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__8031\,
            I => \N__8008\
        );

    \I__1390\ : InMux
    port map (
            O => \N__8030\,
            I => \N__8005\
        );

    \I__1389\ : InMux
    port map (
            O => \N__8029\,
            I => \N__7998\
        );

    \I__1388\ : InMux
    port map (
            O => \N__8028\,
            I => \N__7998\
        );

    \I__1387\ : InMux
    port map (
            O => \N__8027\,
            I => \N__7998\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__8020\,
            I => \N__7991\
        );

    \I__1385\ : InMux
    port map (
            O => \N__8017\,
            I => \N__7988\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__8014\,
            I => \N__7983\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__8011\,
            I => \N__7983\
        );

    \I__1382\ : Span4Mux_v
    port map (
            O => \N__8008\,
            I => \N__7976\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__8005\,
            I => \N__7976\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7998\,
            I => \N__7976\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7997\,
            I => \N__7973\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7996\,
            I => \N__7968\
        );

    \I__1377\ : InMux
    port map (
            O => \N__7995\,
            I => \N__7968\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7994\,
            I => \N__7965\
        );

    \I__1375\ : Odrv4
    port map (
            O => \N__7991\,
            I => rd_addr_r_0
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7988\,
            I => rd_addr_r_0
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__7983\,
            I => rd_addr_r_0
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__7976\,
            I => rd_addr_r_0
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7973\,
            I => rd_addr_r_0
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__7968\,
            I => rd_addr_r_0
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__7965\,
            I => rd_addr_r_0
        );

    \I__1368\ : InMux
    port map (
            O => \N__7950\,
            I => \N__7947\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7947\,
            I => n1
        );

    \I__1366\ : InMux
    port map (
            O => \N__7944\,
            I => \N__7940\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__7943\,
            I => \N__7934\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7940\,
            I => \N__7931\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7926\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7926\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7923\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7934\,
            I => \N__7920\
        );

    \I__1359\ : Span4Mux_v
    port map (
            O => \N__7931\,
            I => \N__7915\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__7926\,
            I => \N__7912\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7923\,
            I => \N__7909\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7920\,
            I => \N__7906\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7903\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7918\,
            I => \N__7900\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__7915\,
            I => fifo_read_cmd
        );

    \I__1352\ : Odrv12
    port map (
            O => \N__7912\,
            I => fifo_read_cmd
        );

    \I__1351\ : Odrv4
    port map (
            O => \N__7909\,
            I => fifo_read_cmd
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__7906\,
            I => fifo_read_cmd
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__7903\,
            I => fifo_read_cmd
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__7900\,
            I => fifo_read_cmd
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__7887\,
            I => \n1_cascade_\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7884\,
            I => \N__7871\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7868\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7863\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7863\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7860\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7879\,
            I => \N__7857\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7852\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7852\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7845\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__7875\,
            I => \N__7841\
        );

    \I__1336\ : InMux
    port map (
            O => \N__7874\,
            I => \N__7836\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7871\,
            I => \N__7831\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7868\,
            I => \N__7831\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7863\,
            I => \N__7828\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__7860\,
            I => \N__7821\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__7857\,
            I => \N__7821\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__7852\,
            I => \N__7821\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__7851\,
            I => \N__7818\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__7850\,
            I => \N__7814\
        );

    \I__1327\ : InMux
    port map (
            O => \N__7849\,
            I => \N__7809\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7848\,
            I => \N__7809\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7845\,
            I => \N__7806\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7801\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7841\,
            I => \N__7801\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__7840\,
            I => \N__7795\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__7839\,
            I => \N__7792\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__7836\,
            I => \N__7789\
        );

    \I__1319\ : Span4Mux_v
    port map (
            O => \N__7831\,
            I => \N__7786\
        );

    \I__1318\ : Span4Mux_v
    port map (
            O => \N__7828\,
            I => \N__7781\
        );

    \I__1317\ : Span4Mux_v
    port map (
            O => \N__7821\,
            I => \N__7781\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7818\,
            I => \N__7778\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7773\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7773\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__7809\,
            I => \N__7770\
        );

    \I__1312\ : Span4Mux_v
    port map (
            O => \N__7806\,
            I => \N__7765\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7801\,
            I => \N__7765\
        );

    \I__1310\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7762\
        );

    \I__1309\ : InMux
    port map (
            O => \N__7799\,
            I => \N__7759\
        );

    \I__1308\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7756\
        );

    \I__1307\ : InMux
    port map (
            O => \N__7795\,
            I => \N__7751\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7792\,
            I => \N__7751\
        );

    \I__1305\ : Odrv4
    port map (
            O => \N__7789\,
            I => rd_addr_r_1
        );

    \I__1304\ : Odrv4
    port map (
            O => \N__7786\,
            I => rd_addr_r_1
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__7781\,
            I => rd_addr_r_1
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__7778\,
            I => rd_addr_r_1
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__7773\,
            I => rd_addr_r_1
        );

    \I__1300\ : Odrv12
    port map (
            O => \N__7770\,
            I => rd_addr_r_1
        );

    \I__1299\ : Odrv4
    port map (
            O => \N__7765\,
            I => rd_addr_r_1
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__7762\,
            I => rd_addr_r_1
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__7759\,
            I => rd_addr_r_1
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__7756\,
            I => rd_addr_r_1
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__7751\,
            I => rd_addr_r_1
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__7728\,
            I => \n3275_cascade_\
        );

    \I__1293\ : InMux
    port map (
            O => \N__7725\,
            I => \N__7722\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__7722\,
            I => n2968
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__7719\,
            I => \n15_adj_509_cascade_\
        );

    \I__1290\ : InMux
    port map (
            O => \N__7716\,
            I => \N__7713\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__7713\,
            I => tx_shift_reg_1
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__7710\,
            I => \N__7707\
        );

    \I__1287\ : InMux
    port map (
            O => \N__7707\,
            I => \N__7704\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__7704\,
            I => tx_shift_reg_2
        );

    \I__1285\ : InMux
    port map (
            O => \N__7701\,
            I => \N__7698\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__7698\,
            I => tx_shift_reg_4
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__7695\,
            I => \n1728_cascade_\
        );

    \I__1282\ : InMux
    port map (
            O => \N__7692\,
            I => \N__7689\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__7689\,
            I => tx_shift_reg_5
        );

    \I__1280\ : InMux
    port map (
            O => \N__7686\,
            I => \N__7683\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__7683\,
            I => \N__7680\
        );

    \I__1278\ : Span4Mux_v
    port map (
            O => \N__7680\,
            I => \N__7676\
        );

    \I__1277\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7673\
        );

    \I__1276\ : Odrv4
    port map (
            O => \N__7676\,
            I => tx_addr_byte_0
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__7673\,
            I => tx_addr_byte_0
        );

    \I__1274\ : InMux
    port map (
            O => \N__7668\,
            I => \N__7665\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__7665\,
            I => tx_shift_reg_6
        );

    \I__1272\ : InMux
    port map (
            O => \N__7662\,
            I => \N__7659\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__7659\,
            I => tx_shift_reg_7
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__7656\,
            I => \N__7649\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__7655\,
            I => \N__7640\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__7654\,
            I => \N__7637\
        );

    \I__1267\ : CascadeMux
    port map (
            O => \N__7653\,
            I => \N__7632\
        );

    \I__1266\ : InMux
    port map (
            O => \N__7652\,
            I => \N__7628\
        );

    \I__1265\ : InMux
    port map (
            O => \N__7649\,
            I => \N__7621\
        );

    \I__1264\ : InMux
    port map (
            O => \N__7648\,
            I => \N__7621\
        );

    \I__1263\ : InMux
    port map (
            O => \N__7647\,
            I => \N__7621\
        );

    \I__1262\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7612\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7645\,
            I => \N__7612\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7644\,
            I => \N__7612\
        );

    \I__1259\ : InMux
    port map (
            O => \N__7643\,
            I => \N__7612\
        );

    \I__1258\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7599\
        );

    \I__1257\ : InMux
    port map (
            O => \N__7637\,
            I => \N__7599\
        );

    \I__1256\ : InMux
    port map (
            O => \N__7636\,
            I => \N__7599\
        );

    \I__1255\ : InMux
    port map (
            O => \N__7635\,
            I => \N__7599\
        );

    \I__1254\ : InMux
    port map (
            O => \N__7632\,
            I => \N__7599\
        );

    \I__1253\ : InMux
    port map (
            O => \N__7631\,
            I => \N__7599\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__7628\,
            I => \N__7596\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__7621\,
            I => n1728
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__7612\,
            I => n1728
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__7599\,
            I => n1728
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__7596\,
            I => n1728
        );

    \I__1247\ : InMux
    port map (
            O => \N__7587\,
            I => \N__7584\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__7584\,
            I => tx_shift_reg_8
        );

    \I__1245\ : InMux
    port map (
            O => \N__7581\,
            I => \N__7578\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__7578\,
            I => tx_shift_reg_9
        );

    \I__1243\ : IoInMux
    port map (
            O => \N__7575\,
            I => \N__7572\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__7572\,
            I => \N__7569\
        );

    \I__1241\ : Span12Mux_s2_h
    port map (
            O => \N__7569\,
            I => \N__7566\
        );

    \I__1240\ : Span12Mux_h
    port map (
            O => \N__7566\,
            I => \N__7562\
        );

    \I__1239\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7559\
        );

    \I__1238\ : Span12Mux_h
    port map (
            O => \N__7562\,
            I => \N__7556\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__7559\,
            I => \N__7553\
        );

    \I__1236\ : Span12Mux_v
    port map (
            O => \N__7556\,
            I => \N__7550\
        );

    \I__1235\ : Span12Mux_v
    port map (
            O => \N__7553\,
            I => \N__7547\
        );

    \I__1234\ : Span12Mux_v
    port map (
            O => \N__7550\,
            I => \N__7542\
        );

    \I__1233\ : Span12Mux_h
    port map (
            O => \N__7547\,
            I => \N__7542\
        );

    \I__1232\ : Odrv12
    port map (
            O => \N__7542\,
            I => \DEBUG_5_c_c\
        );

    \I__1231\ : InMux
    port map (
            O => \N__7539\,
            I => \N__7536\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__7536\,
            I => rx_shift_reg_0
        );

    \I__1229\ : InMux
    port map (
            O => \N__7533\,
            I => \N__7521\
        );

    \I__1228\ : InMux
    port map (
            O => \N__7532\,
            I => \N__7521\
        );

    \I__1227\ : InMux
    port map (
            O => \N__7531\,
            I => \N__7518\
        );

    \I__1226\ : InMux
    port map (
            O => \N__7530\,
            I => \N__7513\
        );

    \I__1225\ : InMux
    port map (
            O => \N__7529\,
            I => \N__7513\
        );

    \I__1224\ : InMux
    port map (
            O => \N__7528\,
            I => \N__7510\
        );

    \I__1223\ : InMux
    port map (
            O => \N__7527\,
            I => \N__7507\
        );

    \I__1222\ : InMux
    port map (
            O => \N__7526\,
            I => \N__7504\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__7521\,
            I => \N__7497\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__7518\,
            I => \N__7497\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__7513\,
            I => \N__7497\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__7510\,
            I => \N__7494\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__7507\,
            I => \N__7489\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__7504\,
            I => \N__7489\
        );

    \I__1215\ : Span4Mux_v
    port map (
            O => \N__7497\,
            I => \N__7486\
        );

    \I__1214\ : Span4Mux_v
    port map (
            O => \N__7494\,
            I => \N__7481\
        );

    \I__1213\ : Span4Mux_v
    port map (
            O => \N__7489\,
            I => \N__7481\
        );

    \I__1212\ : Odrv4
    port map (
            O => \N__7486\,
            I => n4_adj_494
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__7481\,
            I => n4_adj_494
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__7476\,
            I => \N__7473\
        );

    \I__1209\ : InMux
    port map (
            O => \N__7473\,
            I => \N__7470\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__7470\,
            I => \N__7467\
        );

    \I__1207\ : Span4Mux_v
    port map (
            O => \N__7467\,
            I => \N__7463\
        );

    \I__1206\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7460\
        );

    \I__1205\ : Odrv4
    port map (
            O => \N__7463\,
            I => \mem_LUT_mem_1_7\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__7460\,
            I => \mem_LUT_mem_1_7\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__7455\,
            I => \n3279_cascade_\
        );

    \I__1202\ : InMux
    port map (
            O => \N__7452\,
            I => \N__7449\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__7449\,
            I => \spi0.tx_shift_reg_14\
        );

    \I__1200\ : InMux
    port map (
            O => \N__7446\,
            I => \N__7443\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__7443\,
            I => \N__7440\
        );

    \I__1198\ : Odrv4
    port map (
            O => \N__7440\,
            I => tx_shift_reg_12
        );

    \I__1197\ : InMux
    port map (
            O => \N__7437\,
            I => \N__7434\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__7434\,
            I => tx_shift_reg_13
        );

    \I__1195\ : InMux
    port map (
            O => \N__7431\,
            I => \N__7428\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__7428\,
            I => tx_shift_reg_3
        );

    \I__1193\ : InMux
    port map (
            O => \N__7425\,
            I => \N__7421\
        );

    \I__1192\ : InMux
    port map (
            O => \N__7424\,
            I => \N__7418\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__7421\,
            I => \pc_tx.r_Clock_Count_3\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__7418\,
            I => \pc_tx.r_Clock_Count_3\
        );

    \I__1189\ : InMux
    port map (
            O => \N__7413\,
            I => \pc_tx.n2931\
        );

    \I__1188\ : InMux
    port map (
            O => \N__7410\,
            I => \N__7406\
        );

    \I__1187\ : InMux
    port map (
            O => \N__7409\,
            I => \N__7403\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__7406\,
            I => \pc_tx.r_Clock_Count_4\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__7403\,
            I => \pc_tx.r_Clock_Count_4\
        );

    \I__1184\ : InMux
    port map (
            O => \N__7398\,
            I => \pc_tx.n2932\
        );

    \I__1183\ : InMux
    port map (
            O => \N__7395\,
            I => \N__7391\
        );

    \I__1182\ : InMux
    port map (
            O => \N__7394\,
            I => \N__7388\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__7391\,
            I => \pc_tx.r_Clock_Count_5\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__7388\,
            I => \pc_tx.r_Clock_Count_5\
        );

    \I__1179\ : InMux
    port map (
            O => \N__7383\,
            I => \pc_tx.n2933\
        );

    \I__1178\ : InMux
    port map (
            O => \N__7380\,
            I => \N__7376\
        );

    \I__1177\ : InMux
    port map (
            O => \N__7379\,
            I => \N__7373\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__7376\,
            I => \pc_tx.r_Clock_Count_6\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__7373\,
            I => \pc_tx.r_Clock_Count_6\
        );

    \I__1174\ : InMux
    port map (
            O => \N__7368\,
            I => \pc_tx.n2934\
        );

    \I__1173\ : InMux
    port map (
            O => \N__7365\,
            I => \N__7361\
        );

    \I__1172\ : InMux
    port map (
            O => \N__7364\,
            I => \N__7358\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__7361\,
            I => \pc_tx.r_Clock_Count_7\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__7358\,
            I => \pc_tx.r_Clock_Count_7\
        );

    \I__1169\ : InMux
    port map (
            O => \N__7353\,
            I => \pc_tx.n2935\
        );

    \I__1168\ : InMux
    port map (
            O => \N__7350\,
            I => \N__7347\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__7347\,
            I => \N__7343\
        );

    \I__1166\ : InMux
    port map (
            O => \N__7346\,
            I => \N__7340\
        );

    \I__1165\ : Odrv12
    port map (
            O => \N__7343\,
            I => \pc_tx.r_Clock_Count_8\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__7340\,
            I => \pc_tx.r_Clock_Count_8\
        );

    \I__1163\ : InMux
    port map (
            O => \N__7335\,
            I => \bfn_14_13_0_\
        );

    \I__1162\ : InMux
    port map (
            O => \N__7332\,
            I => \pc_tx.n2937\
        );

    \I__1161\ : InMux
    port map (
            O => \N__7329\,
            I => \N__7326\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__7326\,
            I => \N__7322\
        );

    \I__1159\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7319\
        );

    \I__1158\ : Odrv12
    port map (
            O => \N__7322\,
            I => \pc_tx.r_Clock_Count_9\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__7319\,
            I => \pc_tx.r_Clock_Count_9\
        );

    \I__1156\ : CEMux
    port map (
            O => \N__7314\,
            I => \N__7311\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__7311\,
            I => \N__7306\
        );

    \I__1154\ : CEMux
    port map (
            O => \N__7310\,
            I => \N__7303\
        );

    \I__1153\ : CEMux
    port map (
            O => \N__7309\,
            I => \N__7300\
        );

    \I__1152\ : Span12Mux_s5_h
    port map (
            O => \N__7306\,
            I => \N__7297\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__7303\,
            I => \N__7294\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__7300\,
            I => \N__7291\
        );

    \I__1149\ : Span12Mux_v
    port map (
            O => \N__7297\,
            I => \N__7288\
        );

    \I__1148\ : Span4Mux_v
    port map (
            O => \N__7294\,
            I => \N__7283\
        );

    \I__1147\ : Span4Mux_v
    port map (
            O => \N__7291\,
            I => \N__7283\
        );

    \I__1146\ : Odrv12
    port map (
            O => \N__7288\,
            I => \pc_tx.n1\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__7283\,
            I => \pc_tx.n1\
        );

    \I__1144\ : SRMux
    port map (
            O => \N__7278\,
            I => \N__7274\
        );

    \I__1143\ : SRMux
    port map (
            O => \N__7277\,
            I => \N__7271\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__7274\,
            I => \N__7268\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__7271\,
            I => \N__7265\
        );

    \I__1140\ : Span4Mux_h
    port map (
            O => \N__7268\,
            I => \N__7262\
        );

    \I__1139\ : Span12Mux_h
    port map (
            O => \N__7265\,
            I => \N__7259\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__7262\,
            I => \pc_tx.n1919\
        );

    \I__1137\ : Odrv12
    port map (
            O => \N__7259\,
            I => \pc_tx.n1919\
        );

    \I__1136\ : SRMux
    port map (
            O => \N__7254\,
            I => \N__7250\
        );

    \I__1135\ : SRMux
    port map (
            O => \N__7253\,
            I => \N__7247\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__7250\,
            I => \N__7238\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__7247\,
            I => \N__7235\
        );

    \I__1132\ : InMux
    port map (
            O => \N__7246\,
            I => \N__7230\
        );

    \I__1131\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7230\
        );

    \I__1130\ : InMux
    port map (
            O => \N__7244\,
            I => \N__7225\
        );

    \I__1129\ : InMux
    port map (
            O => \N__7243\,
            I => \N__7225\
        );

    \I__1128\ : InMux
    port map (
            O => \N__7242\,
            I => \N__7222\
        );

    \I__1127\ : InMux
    port map (
            O => \N__7241\,
            I => \N__7219\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__7238\,
            I => \r_SM_Main_2_adj_495\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__7235\,
            I => \r_SM_Main_2_adj_495\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__7230\,
            I => \r_SM_Main_2_adj_495\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__7225\,
            I => \r_SM_Main_2_adj_495\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__7222\,
            I => \r_SM_Main_2_adj_495\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__7219\,
            I => \r_SM_Main_2_adj_495\
        );

    \I__1120\ : InMux
    port map (
            O => \N__7206\,
            I => \N__7199\
        );

    \I__1119\ : InMux
    port map (
            O => \N__7205\,
            I => \N__7195\
        );

    \I__1118\ : InMux
    port map (
            O => \N__7204\,
            I => \N__7190\
        );

    \I__1117\ : InMux
    port map (
            O => \N__7203\,
            I => \N__7190\
        );

    \I__1116\ : InMux
    port map (
            O => \N__7202\,
            I => \N__7187\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__7199\,
            I => \N__7183\
        );

    \I__1114\ : InMux
    port map (
            O => \N__7198\,
            I => \N__7180\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__7195\,
            I => \N__7173\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__7190\,
            I => \N__7173\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__7187\,
            I => \N__7173\
        );

    \I__1110\ : InMux
    port map (
            O => \N__7186\,
            I => \N__7170\
        );

    \I__1109\ : Span4Mux_v
    port map (
            O => \N__7183\,
            I => \N__7165\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__7180\,
            I => \N__7165\
        );

    \I__1107\ : Span4Mux_v
    port map (
            O => \N__7173\,
            I => \N__7160\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__7170\,
            I => \N__7160\
        );

    \I__1105\ : Odrv4
    port map (
            O => \N__7165\,
            I => n2
        );

    \I__1104\ : Odrv4
    port map (
            O => \N__7160\,
            I => n2
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__7155\,
            I => \n2_cascade_\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__7152\,
            I => \pc_tx.n2981_cascade_\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__7149\,
            I => \pc_tx.n2564_cascade_\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__7146\,
            I => \N__7142\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__7145\,
            I => \N__7136\
        );

    \I__1098\ : InMux
    port map (
            O => \N__7142\,
            I => \N__7131\
        );

    \I__1097\ : InMux
    port map (
            O => \N__7141\,
            I => \N__7131\
        );

    \I__1096\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7126\
        );

    \I__1095\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7126\
        );

    \I__1094\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7122\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__7131\,
            I => \N__7117\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__7126\,
            I => \N__7117\
        );

    \I__1091\ : InMux
    port map (
            O => \N__7125\,
            I => \N__7114\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__7122\,
            I => \N__7111\
        );

    \I__1089\ : Span4Mux_h
    port map (
            O => \N__7117\,
            I => \N__7107\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__7114\,
            I => \N__7104\
        );

    \I__1087\ : Span4Mux_v
    port map (
            O => \N__7111\,
            I => \N__7101\
        );

    \I__1086\ : InMux
    port map (
            O => \N__7110\,
            I => \N__7098\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__7107\,
            I => \r_SM_Main_2_N_184_1\
        );

    \I__1084\ : Odrv12
    port map (
            O => \N__7104\,
            I => \r_SM_Main_2_N_184_1\
        );

    \I__1083\ : Odrv4
    port map (
            O => \N__7101\,
            I => \r_SM_Main_2_N_184_1\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__7098\,
            I => \r_SM_Main_2_N_184_1\
        );

    \I__1081\ : InMux
    port map (
            O => \N__7089\,
            I => \N__7085\
        );

    \I__1080\ : InMux
    port map (
            O => \N__7088\,
            I => \N__7082\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__7085\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__7082\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__7077\,
            I => \N__7074\
        );

    \I__1076\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7068\
        );

    \I__1075\ : InMux
    port map (
            O => \N__7073\,
            I => \N__7068\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__7068\,
            I => \mem_LUT_mem_3_0\
        );

    \I__1073\ : InMux
    port map (
            O => \N__7065\,
            I => \N__7062\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__7062\,
            I => \N__7059\
        );

    \I__1071\ : Span4Mux_v
    port map (
            O => \N__7059\,
            I => \N__7056\
        );

    \I__1070\ : Odrv4
    port map (
            O => \N__7056\,
            I => \tx_fifo.lscc_fifo_inst.n3421\
        );

    \I__1069\ : InMux
    port map (
            O => \N__7053\,
            I => \N__7050\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__7050\,
            I => \N__7046\
        );

    \I__1067\ : InMux
    port map (
            O => \N__7049\,
            I => \N__7043\
        );

    \I__1066\ : Odrv4
    port map (
            O => \N__7046\,
            I => \pc_tx.r_Clock_Count_0\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__7043\,
            I => \pc_tx.r_Clock_Count_0\
        );

    \I__1064\ : InMux
    port map (
            O => \N__7038\,
            I => \bfn_14_12_0_\
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__7035\,
            I => \N__7032\
        );

    \I__1062\ : InMux
    port map (
            O => \N__7032\,
            I => \N__7028\
        );

    \I__1061\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7025\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__7028\,
            I => \pc_tx.r_Clock_Count_1\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__7025\,
            I => \pc_tx.r_Clock_Count_1\
        );

    \I__1058\ : InMux
    port map (
            O => \N__7020\,
            I => \pc_tx.n2929\
        );

    \I__1057\ : InMux
    port map (
            O => \N__7017\,
            I => \N__7013\
        );

    \I__1056\ : InMux
    port map (
            O => \N__7016\,
            I => \N__7010\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__7013\,
            I => \pc_tx.r_Clock_Count_2\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__7010\,
            I => \pc_tx.r_Clock_Count_2\
        );

    \I__1053\ : InMux
    port map (
            O => \N__7005\,
            I => \pc_tx.n2930\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__7002\,
            I => \N__6999\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6995\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6998\,
            I => \N__6992\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6995\,
            I => \mem_LUT_mem_1_3\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6992\,
            I => \mem_LUT_mem_1_3\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6987\,
            I => \N__6984\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6984\,
            I => \N__6980\
        );

    \I__1045\ : InMux
    port map (
            O => \N__6983\,
            I => \N__6977\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__6980\,
            I => \mem_LUT_mem_1_4\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6977\,
            I => \mem_LUT_mem_1_4\
        );

    \I__1042\ : CascadeMux
    port map (
            O => \N__6972\,
            I => \N__6969\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6969\,
            I => \N__6966\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6966\,
            I => \N__6962\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6959\
        );

    \I__1038\ : Odrv4
    port map (
            O => \N__6962\,
            I => tx_addr_byte_4
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6959\,
            I => tx_addr_byte_4
        );

    \I__1036\ : SRMux
    port map (
            O => \N__6954\,
            I => \N__6951\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6951\,
            I => \spi0.n3176\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6948\,
            I => \N__6944\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6947\,
            I => \N__6941\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6944\,
            I => \N__6935\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6941\,
            I => \N__6935\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6932\
        );

    \I__1029\ : Odrv12
    port map (
            O => \N__6935\,
            I => tx_data_byte_3
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__6932\,
            I => tx_data_byte_3
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__6927\,
            I => \N__6924\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6920\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6917\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__6920\,
            I => tx_addr_byte_3
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6917\,
            I => tx_addr_byte_3
        );

    \I__1022\ : InMux
    port map (
            O => \N__6912\,
            I => \N__6909\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6909\,
            I => tx_shift_reg_11
        );

    \I__1020\ : InMux
    port map (
            O => \N__6906\,
            I => \N__6903\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6903\,
            I => tx_shift_reg_10
        );

    \I__1018\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6896\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6899\,
            I => \N__6893\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__6896\,
            I => \N__6888\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6893\,
            I => \N__6885\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__6892\,
            I => \N__6882\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__6891\,
            I => \N__6877\
        );

    \I__1012\ : Span4Mux_h
    port map (
            O => \N__6888\,
            I => \N__6872\
        );

    \I__1011\ : Span4Mux_v
    port map (
            O => \N__6885\,
            I => \N__6869\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6882\,
            I => \N__6862\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6862\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6862\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6877\,
            I => \N__6859\
        );

    \I__1006\ : InMux
    port map (
            O => \N__6876\,
            I => \N__6856\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6875\,
            I => \N__6853\
        );

    \I__1004\ : Odrv4
    port map (
            O => \N__6872\,
            I => \r_SM_Main_0_adj_497\
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__6869\,
            I => \r_SM_Main_0_adj_497\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6862\,
            I => \r_SM_Main_0_adj_497\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__6859\,
            I => \r_SM_Main_0_adj_497\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__6856\,
            I => \r_SM_Main_0_adj_497\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__6853\,
            I => \r_SM_Main_0_adj_497\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__6840\,
            I => \N__6830\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__6839\,
            I => \N__6827\
        );

    \I__996\ : InMux
    port map (
            O => \N__6838\,
            I => \N__6817\
        );

    \I__995\ : InMux
    port map (
            O => \N__6837\,
            I => \N__6817\
        );

    \I__994\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6817\
        );

    \I__993\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6817\
        );

    \I__992\ : InMux
    port map (
            O => \N__6834\,
            I => \N__6814\
        );

    \I__991\ : InMux
    port map (
            O => \N__6833\,
            I => \N__6807\
        );

    \I__990\ : InMux
    port map (
            O => \N__6830\,
            I => \N__6807\
        );

    \I__989\ : InMux
    port map (
            O => \N__6827\,
            I => \N__6807\
        );

    \I__988\ : InMux
    port map (
            O => \N__6826\,
            I => \N__6804\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__6817\,
            I => \N__6796\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__6814\,
            I => \N__6796\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__6807\,
            I => \N__6796\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__6804\,
            I => \N__6793\
        );

    \I__983\ : InMux
    port map (
            O => \N__6803\,
            I => \N__6790\
        );

    \I__982\ : Odrv12
    port map (
            O => \N__6796\,
            I => \r_SM_Main_1_adj_496\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__6793\,
            I => \r_SM_Main_1_adj_496\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__6790\,
            I => \r_SM_Main_1_adj_496\
        );

    \I__979\ : InMux
    port map (
            O => \N__6783\,
            I => \N__6779\
        );

    \I__978\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6776\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__6779\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__6776\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1\
        );

    \I__975\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6763\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__6770\,
            I => \N__6759\
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__6769\,
            I => \N__6755\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__6768\,
            I => \N__6751\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__6767\,
            I => \N__6748\
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__6766\,
            I => \N__6745\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6763\,
            I => \N__6742\
        );

    \I__968\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6733\
        );

    \I__967\ : InMux
    port map (
            O => \N__6759\,
            I => \N__6733\
        );

    \I__966\ : InMux
    port map (
            O => \N__6758\,
            I => \N__6733\
        );

    \I__965\ : InMux
    port map (
            O => \N__6755\,
            I => \N__6733\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__6754\,
            I => \N__6727\
        );

    \I__963\ : InMux
    port map (
            O => \N__6751\,
            I => \N__6721\
        );

    \I__962\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6718\
        );

    \I__961\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6715\
        );

    \I__960\ : Span4Mux_h
    port map (
            O => \N__6742\,
            I => \N__6710\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__6733\,
            I => \N__6710\
        );

    \I__958\ : InMux
    port map (
            O => \N__6732\,
            I => \N__6707\
        );

    \I__957\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6702\
        );

    \I__956\ : InMux
    port map (
            O => \N__6730\,
            I => \N__6702\
        );

    \I__955\ : InMux
    port map (
            O => \N__6727\,
            I => \N__6697\
        );

    \I__954\ : InMux
    port map (
            O => \N__6726\,
            I => \N__6697\
        );

    \I__953\ : InMux
    port map (
            O => \N__6725\,
            I => \N__6692\
        );

    \I__952\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6692\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__6721\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__6718\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__6715\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__948\ : Odrv4
    port map (
            O => \N__6710\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__6707\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__6702\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__6697\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__6692\,
            I => \tx_fifo.lscc_fifo_inst.n4\
        );

    \I__943\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6672\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__6672\,
            I => \N__6668\
        );

    \I__941\ : InMux
    port map (
            O => \N__6671\,
            I => \N__6665\
        );

    \I__940\ : Odrv4
    port map (
            O => \N__6668\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__6665\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7\
        );

    \I__938\ : InMux
    port map (
            O => \N__6660\,
            I => \N__6657\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__6657\,
            I => \N__6648\
        );

    \I__936\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6643\
        );

    \I__935\ : InMux
    port map (
            O => \N__6655\,
            I => \N__6643\
        );

    \I__934\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6636\
        );

    \I__933\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6636\
        );

    \I__932\ : InMux
    port map (
            O => \N__6652\,
            I => \N__6636\
        );

    \I__931\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6633\
        );

    \I__930\ : Span4Mux_v
    port map (
            O => \N__6648\,
            I => \N__6628\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__6643\,
            I => \N__6628\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__6636\,
            I => n1795
        );

    \I__927\ : LocalMux
    port map (
            O => \N__6633\,
            I => n1795
        );

    \I__926\ : Odrv4
    port map (
            O => \N__6628\,
            I => n1795
        );

    \I__925\ : InMux
    port map (
            O => \N__6621\,
            I => \N__6618\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__6618\,
            I => \N__6615\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__6615\,
            I => \mem_LUT_data_raw_r_1\
        );

    \I__922\ : InMux
    port map (
            O => \N__6612\,
            I => \N__6608\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__6611\,
            I => \N__6605\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__6608\,
            I => \N__6602\
        );

    \I__919\ : InMux
    port map (
            O => \N__6605\,
            I => \N__6599\
        );

    \I__918\ : Odrv4
    port map (
            O => \N__6602\,
            I => fifo_temp_output_1
        );

    \I__917\ : LocalMux
    port map (
            O => \N__6599\,
            I => fifo_temp_output_1
        );

    \I__916\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6591\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__6591\,
            I => \N__6587\
        );

    \I__914\ : InMux
    port map (
            O => \N__6590\,
            I => \N__6584\
        );

    \I__913\ : Odrv4
    port map (
            O => \N__6587\,
            I => \mem_LUT_mem_3_6\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__6584\,
            I => \mem_LUT_mem_3_6\
        );

    \I__911\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6575\
        );

    \I__910\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6572\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__6575\,
            I => \mem_LUT_mem_3_3\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__6572\,
            I => \mem_LUT_mem_3_3\
        );

    \I__907\ : InMux
    port map (
            O => \N__6567\,
            I => \N__6564\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__6564\,
            I => \N__6560\
        );

    \I__905\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6557\
        );

    \I__904\ : Odrv12
    port map (
            O => \N__6560\,
            I => \mem_LUT_mem_1_2\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__6557\,
            I => \mem_LUT_mem_1_2\
        );

    \I__902\ : InMux
    port map (
            O => \N__6552\,
            I => \N__6548\
        );

    \I__901\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6545\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__6548\,
            I => tx_addr_byte_7
        );

    \I__899\ : LocalMux
    port map (
            O => \N__6545\,
            I => tx_addr_byte_7
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__6540\,
            I => \rd_addr_p1_w_2_cascade_\
        );

    \I__897\ : CEMux
    port map (
            O => \N__6537\,
            I => \N__6533\
        );

    \I__896\ : CEMux
    port map (
            O => \N__6536\,
            I => \N__6530\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__6533\,
            I => \N__6524\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__6530\,
            I => \N__6521\
        );

    \I__893\ : CEMux
    port map (
            O => \N__6529\,
            I => \N__6518\
        );

    \I__892\ : CEMux
    port map (
            O => \N__6528\,
            I => \N__6515\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__6527\,
            I => \N__6512\
        );

    \I__890\ : Span4Mux_v
    port map (
            O => \N__6524\,
            I => \N__6503\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__6521\,
            I => \N__6503\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__6518\,
            I => \N__6503\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__6515\,
            I => \N__6500\
        );

    \I__886\ : InMux
    port map (
            O => \N__6512\,
            I => \N__6497\
        );

    \I__885\ : InMux
    port map (
            O => \N__6511\,
            I => \N__6494\
        );

    \I__884\ : CEMux
    port map (
            O => \N__6510\,
            I => \N__6491\
        );

    \I__883\ : Span4Mux_v
    port map (
            O => \N__6503\,
            I => \N__6488\
        );

    \I__882\ : Span4Mux_v
    port map (
            O => \N__6500\,
            I => \N__6479\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__6497\,
            I => \N__6479\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__6494\,
            I => \N__6479\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__6491\,
            I => \N__6479\
        );

    \I__878\ : Sp12to4
    port map (
            O => \N__6488\,
            I => \N__6476\
        );

    \I__877\ : Span4Mux_v
    port map (
            O => \N__6479\,
            I => \N__6473\
        );

    \I__876\ : Odrv12
    port map (
            O => \N__6476\,
            I => rd_fifo_en_w
        );

    \I__875\ : Odrv4
    port map (
            O => \N__6473\,
            I => rd_fifo_en_w
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__6468\,
            I => \n3448_cascade_\
        );

    \I__873\ : InMux
    port map (
            O => \N__6465\,
            I => \N__6462\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__6462\,
            I => rd_addr_p1_w_2
        );

    \I__871\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6456\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__6456\,
            I => n3289
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__6453\,
            I => \N__6450\
        );

    \I__868\ : InMux
    port map (
            O => \N__6450\,
            I => \N__6447\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__6447\,
            I => \N__6443\
        );

    \I__866\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6440\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__6443\,
            I => \mem_LUT_mem_3_1\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__6440\,
            I => \mem_LUT_mem_3_1\
        );

    \I__863\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6432\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__6432\,
            I => \tx_fifo.lscc_fifo_inst.n3427\
        );

    \I__861\ : CascadeMux
    port map (
            O => \N__6429\,
            I => \N__6426\
        );

    \I__860\ : InMux
    port map (
            O => \N__6426\,
            I => \N__6423\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__6423\,
            I => \N__6419\
        );

    \I__858\ : InMux
    port map (
            O => \N__6422\,
            I => \N__6416\
        );

    \I__857\ : Odrv12
    port map (
            O => \N__6419\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__6416\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1\
        );

    \I__855\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6408\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__6408\,
            I => \N__6404\
        );

    \I__853\ : InMux
    port map (
            O => \N__6407\,
            I => \N__6401\
        );

    \I__852\ : Odrv4
    port map (
            O => \N__6404\,
            I => \mem_LUT_mem_1_1\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__6401\,
            I => \mem_LUT_mem_1_1\
        );

    \I__850\ : InMux
    port map (
            O => \N__6396\,
            I => \N__6393\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__6393\,
            I => \N__6389\
        );

    \I__848\ : InMux
    port map (
            O => \N__6392\,
            I => \N__6386\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__6389\,
            I => \mem_LUT_mem_1_5\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__6386\,
            I => \mem_LUT_mem_1_5\
        );

    \I__845\ : InMux
    port map (
            O => \N__6381\,
            I => \N__6378\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__6378\,
            I => \N__6375\
        );

    \I__843\ : Span4Mux_v
    port map (
            O => \N__6375\,
            I => \N__6371\
        );

    \I__842\ : InMux
    port map (
            O => \N__6374\,
            I => \N__6368\
        );

    \I__841\ : Odrv4
    port map (
            O => \N__6371\,
            I => fifo_temp_output_6
        );

    \I__840\ : LocalMux
    port map (
            O => \N__6368\,
            I => fifo_temp_output_6
        );

    \I__839\ : InMux
    port map (
            O => \N__6363\,
            I => \N__6360\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__6360\,
            I => \N__6356\
        );

    \I__837\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6353\
        );

    \I__836\ : Span4Mux_h
    port map (
            O => \N__6356\,
            I => \N__6343\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__6353\,
            I => \N__6343\
        );

    \I__834\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6338\
        );

    \I__833\ : InMux
    port map (
            O => \N__6351\,
            I => \N__6338\
        );

    \I__832\ : InMux
    port map (
            O => \N__6350\,
            I => \N__6334\
        );

    \I__831\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6331\
        );

    \I__830\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6328\
        );

    \I__829\ : Sp12to4
    port map (
            O => \N__6343\,
            I => \N__6323\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__6338\,
            I => \N__6323\
        );

    \I__827\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6320\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__6334\,
            I => \N__6317\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__6331\,
            I => \N__6312\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__6328\,
            I => \N__6312\
        );

    \I__823\ : Span12Mux_v
    port map (
            O => \N__6323\,
            I => \N__6307\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__6320\,
            I => \N__6307\
        );

    \I__821\ : Odrv4
    port map (
            O => \N__6317\,
            I => n1636
        );

    \I__820\ : Odrv4
    port map (
            O => \N__6312\,
            I => n1636
        );

    \I__819\ : Odrv12
    port map (
            O => \N__6307\,
            I => n1636
        );

    \I__818\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6297\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__6297\,
            I => \N__6294\
        );

    \I__816\ : Span4Mux_v
    port map (
            O => \N__6294\,
            I => \N__6290\
        );

    \I__815\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6287\
        );

    \I__814\ : Odrv4
    port map (
            O => \N__6290\,
            I => \r_Tx_Data_6\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__6287\,
            I => \r_Tx_Data_6\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__6282\,
            I => \N__6278\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__6281\,
            I => \N__6275\
        );

    \I__810\ : InMux
    port map (
            O => \N__6278\,
            I => \N__6272\
        );

    \I__809\ : InMux
    port map (
            O => \N__6275\,
            I => \N__6269\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__6272\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__6269\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4\
        );

    \I__806\ : InMux
    port map (
            O => \N__6264\,
            I => \N__6260\
        );

    \I__805\ : InMux
    port map (
            O => \N__6263\,
            I => \N__6257\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__6260\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__6257\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2\
        );

    \I__802\ : InMux
    port map (
            O => \N__6252\,
            I => \N__6248\
        );

    \I__801\ : InMux
    port map (
            O => \N__6251\,
            I => \N__6245\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__6248\,
            I => \mem_LUT_mem_3_2\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__6245\,
            I => \mem_LUT_mem_3_2\
        );

    \I__798\ : InMux
    port map (
            O => \N__6240\,
            I => \N__6237\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__6237\,
            I => \N__6234\
        );

    \I__796\ : Odrv4
    port map (
            O => \N__6234\,
            I => \tx_fifo.lscc_fifo_inst.n3415\
        );

    \I__795\ : InMux
    port map (
            O => \N__6231\,
            I => \N__6228\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__6228\,
            I => \mem_LUT_data_raw_r_7\
        );

    \I__793\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6222\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__6222\,
            I => \N__6219\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__6219\,
            I => \tx_fifo.lscc_fifo_inst.n3391\
        );

    \I__790\ : InMux
    port map (
            O => \N__6216\,
            I => \N__6212\
        );

    \I__789\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6209\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__6212\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__6209\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3\
        );

    \I__786\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6201\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__6201\,
            I => \N__6198\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__6198\,
            I => \mem_LUT_data_raw_r_3\
        );

    \I__783\ : IoInMux
    port map (
            O => \N__6195\,
            I => \N__6192\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__6192\,
            I => \N__6189\
        );

    \I__781\ : Span12Mux_s2_v
    port map (
            O => \N__6189\,
            I => \N__6186\
        );

    \I__780\ : Span12Mux_h
    port map (
            O => \N__6186\,
            I => \N__6183\
        );

    \I__779\ : Odrv12
    port map (
            O => \N__6183\,
            I => \SDAT_c\
        );

    \I__778\ : InMux
    port map (
            O => \N__6180\,
            I => \N__6174\
        );

    \I__777\ : InMux
    port map (
            O => \N__6179\,
            I => \N__6174\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__6174\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5\
        );

    \I__775\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6167\
        );

    \I__774\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6164\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__6167\,
            I => \mem_LUT_mem_3_5\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__6164\,
            I => \mem_LUT_mem_3_5\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__6159\,
            I => \N__6155\
        );

    \I__770\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6152\
        );

    \I__769\ : InMux
    port map (
            O => \N__6155\,
            I => \N__6149\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__6152\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__6149\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3\
        );

    \I__766\ : InMux
    port map (
            O => \N__6144\,
            I => \N__6138\
        );

    \I__765\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6138\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__6138\,
            I => \mem_LUT_mem_3_7\
        );

    \I__763\ : InMux
    port map (
            O => \N__6135\,
            I => \N__6129\
        );

    \I__762\ : InMux
    port map (
            O => \N__6134\,
            I => \N__6129\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__6129\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__6126\,
            I => \N__6123\
        );

    \I__759\ : InMux
    port map (
            O => \N__6123\,
            I => \N__6120\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__6120\,
            I => \N__6116\
        );

    \I__757\ : InMux
    port map (
            O => \N__6119\,
            I => \N__6113\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__6116\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__6113\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__6108\,
            I => \N__6105\
        );

    \I__753\ : InMux
    port map (
            O => \N__6105\,
            I => \N__6099\
        );

    \I__752\ : InMux
    port map (
            O => \N__6104\,
            I => \N__6099\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__6099\,
            I => \N__6096\
        );

    \I__750\ : Odrv4
    port map (
            O => \N__6096\,
            I => \mem_LUT_mem_3_4\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__6093\,
            I => \N__6089\
        );

    \I__748\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6084\
        );

    \I__747\ : InMux
    port map (
            O => \N__6089\,
            I => \N__6084\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__6084\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4\
        );

    \I__745\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6071\
        );

    \I__744\ : InMux
    port map (
            O => \N__6080\,
            I => \N__6071\
        );

    \I__743\ : CascadeMux
    port map (
            O => \N__6079\,
            I => \N__6068\
        );

    \I__742\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6065\
        );

    \I__741\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6062\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__6076\,
            I => \N__6057\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__6071\,
            I => \N__6054\
        );

    \I__738\ : InMux
    port map (
            O => \N__6068\,
            I => \N__6051\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__6065\,
            I => \N__6046\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__6062\,
            I => \N__6046\
        );

    \I__735\ : InMux
    port map (
            O => \N__6061\,
            I => \N__6043\
        );

    \I__734\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6038\
        );

    \I__733\ : InMux
    port map (
            O => \N__6057\,
            I => \N__6038\
        );

    \I__732\ : Odrv4
    port map (
            O => \N__6054\,
            I => is_fifo_empty_flag
        );

    \I__731\ : LocalMux
    port map (
            O => \N__6051\,
            I => is_fifo_empty_flag
        );

    \I__730\ : Odrv4
    port map (
            O => \N__6046\,
            I => is_fifo_empty_flag
        );

    \I__729\ : LocalMux
    port map (
            O => \N__6043\,
            I => is_fifo_empty_flag
        );

    \I__728\ : LocalMux
    port map (
            O => \N__6038\,
            I => is_fifo_empty_flag
        );

    \I__727\ : InMux
    port map (
            O => \N__6027\,
            I => \N__6024\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__6024\,
            I => n4_adj_511
        );

    \I__725\ : InMux
    port map (
            O => \N__6021\,
            I => \N__6018\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__6018\,
            I => \tx_fifo.lscc_fifo_inst.n3409\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__6015\,
            I => \tx_fifo.lscc_fifo_inst.n4_cascade_\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__6012\,
            I => \N__6009\
        );

    \I__721\ : InMux
    port map (
            O => \N__6009\,
            I => \N__6005\
        );

    \I__720\ : InMux
    port map (
            O => \N__6008\,
            I => \N__6002\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__6005\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__6002\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5\
        );

    \I__717\ : InMux
    port map (
            O => \N__5997\,
            I => \N__5993\
        );

    \I__716\ : InMux
    port map (
            O => \N__5996\,
            I => \N__5990\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5993\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__5990\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0\
        );

    \I__713\ : InMux
    port map (
            O => \N__5985\,
            I => \N__5982\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5982\,
            I => \N__5978\
        );

    \I__711\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5975\
        );

    \I__710\ : Odrv12
    port map (
            O => \N__5978\,
            I => \r_Tx_Data_7\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__5975\,
            I => \r_Tx_Data_7\
        );

    \I__708\ : InMux
    port map (
            O => \N__5970\,
            I => \N__5966\
        );

    \I__707\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5961\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5966\,
            I => \N__5958\
        );

    \I__705\ : InMux
    port map (
            O => \N__5965\,
            I => \N__5955\
        );

    \I__704\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5952\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5961\,
            I => \N__5945\
        );

    \I__702\ : Span12Mux_h
    port map (
            O => \N__5958\,
            I => \N__5942\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5955\,
            I => \N__5937\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5952\,
            I => \N__5937\
        );

    \I__699\ : InMux
    port map (
            O => \N__5951\,
            I => \N__5932\
        );

    \I__698\ : InMux
    port map (
            O => \N__5950\,
            I => \N__5932\
        );

    \I__697\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5927\
        );

    \I__696\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5927\
        );

    \I__695\ : Odrv12
    port map (
            O => \N__5945\,
            I => \r_Bit_Index_0_adj_498\
        );

    \I__694\ : Odrv12
    port map (
            O => \N__5942\,
            I => \r_Bit_Index_0_adj_498\
        );

    \I__693\ : Odrv4
    port map (
            O => \N__5937\,
            I => \r_Bit_Index_0_adj_498\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5932\,
            I => \r_Bit_Index_0_adj_498\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__5927\,
            I => \r_Bit_Index_0_adj_498\
        );

    \I__690\ : CascadeMux
    port map (
            O => \N__5916\,
            I => \N__5913\
        );

    \I__689\ : InMux
    port map (
            O => \N__5913\,
            I => \N__5910\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__5910\,
            I => \N__5907\
        );

    \I__687\ : Odrv12
    port map (
            O => \N__5907\,
            I => \pc_tx.n3320\
        );

    \I__686\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5901\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__5901\,
            I => \tx_fifo.lscc_fifo_inst.n3433\
        );

    \I__684\ : InMux
    port map (
            O => \N__5898\,
            I => \N__5895\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__5895\,
            I => \mem_LUT_data_raw_r_4\
        );

    \I__682\ : InMux
    port map (
            O => \N__5892\,
            I => \N__5889\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5889\,
            I => \N__5886\
        );

    \I__680\ : Span4Mux_v
    port map (
            O => \N__5886\,
            I => \N__5882\
        );

    \I__679\ : InMux
    port map (
            O => \N__5885\,
            I => \N__5879\
        );

    \I__678\ : Odrv4
    port map (
            O => \N__5882\,
            I => fifo_temp_output_7
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5879\,
            I => fifo_temp_output_7
        );

    \I__676\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5871\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5871\,
            I => \N__5868\
        );

    \I__674\ : Span4Mux_v
    port map (
            O => \N__5868\,
            I => \N__5865\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__5865\,
            I => \tx_fifo.lscc_fifo_inst.n3403\
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__5862\,
            I => \n32_cascade_\
        );

    \I__671\ : CascadeMux
    port map (
            O => \N__5859\,
            I => \n24_adj_510_cascade_\
        );

    \I__670\ : InMux
    port map (
            O => \N__5856\,
            I => \N__5853\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5853\,
            I => \N__5850\
        );

    \I__668\ : Span4Mux_v
    port map (
            O => \N__5850\,
            I => \N__5847\
        );

    \I__667\ : Odrv4
    port map (
            O => \N__5847\,
            I => \mem_LUT_data_raw_r_5\
        );

    \I__666\ : InMux
    port map (
            O => \N__5844\,
            I => \N__5841\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5841\,
            I => \tx_fifo.lscc_fifo_inst.n3397\
        );

    \I__664\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5832\
        );

    \I__663\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5832\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__5832\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6\
        );

    \I__661\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5825\
        );

    \I__660\ : InMux
    port map (
            O => \N__5828\,
            I => \N__5822\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__5825\,
            I => \r_Tx_Data_1\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__5822\,
            I => \r_Tx_Data_1\
        );

    \I__657\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5814\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__5814\,
            I => \N__5810\
        );

    \I__655\ : InMux
    port map (
            O => \N__5813\,
            I => \N__5807\
        );

    \I__654\ : Odrv12
    port map (
            O => \N__5810\,
            I => \mem_LUT_mem_1_0\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__5807\,
            I => \mem_LUT_mem_1_0\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__5802\,
            I => \N__5798\
        );

    \I__651\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5795\
        );

    \I__650\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5792\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__5795\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__5792\,
            I => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6\
        );

    \I__647\ : CascadeMux
    port map (
            O => \N__5787\,
            I => \N__5784\
        );

    \I__646\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5781\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__5781\,
            I => rd_fifo_en_prev_r
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__5778\,
            I => \n1795_cascade_\
        );

    \I__643\ : CascadeMux
    port map (
            O => \N__5775\,
            I => \n4_cascade_\
        );

    \I__642\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5767\
        );

    \I__641\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5762\
        );

    \I__640\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5762\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__5767\,
            I => tx_uart_active_flag
        );

    \I__638\ : LocalMux
    port map (
            O => \N__5762\,
            I => tx_uart_active_flag
        );

    \I__637\ : InMux
    port map (
            O => \N__5757\,
            I => \N__5749\
        );

    \I__636\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5749\
        );

    \I__635\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5744\
        );

    \I__634\ : InMux
    port map (
            O => \N__5754\,
            I => \N__5744\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5749\,
            I => \r_SM_Main_2_N_187_0\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__5744\,
            I => \r_SM_Main_2_N_187_0\
        );

    \I__631\ : InMux
    port map (
            O => \N__5739\,
            I => \N__5736\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__5736\,
            I => \N__5733\
        );

    \I__629\ : Odrv4
    port map (
            O => \N__5733\,
            I => \pc_tx.o_Tx_Serial_N_216\
        );

    \I__628\ : IoInMux
    port map (
            O => \N__5730\,
            I => \N__5727\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__5727\,
            I => \N__5724\
        );

    \I__626\ : Span12Mux_s8_h
    port map (
            O => \N__5724\,
            I => \N__5721\
        );

    \I__625\ : Span12Mux_v
    port map (
            O => \N__5721\,
            I => \N__5718\
        );

    \I__624\ : Odrv12
    port map (
            O => \N__5718\,
            I => \pc_tx.n3\
        );

    \I__623\ : CascadeMux
    port map (
            O => \N__5715\,
            I => \N__5712\
        );

    \I__622\ : InMux
    port map (
            O => \N__5712\,
            I => \N__5709\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__5709\,
            I => \N__5706\
        );

    \I__620\ : Odrv4
    port map (
            O => \N__5706\,
            I => \mem_LUT_data_raw_r_0\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__5703\,
            I => \N__5700\
        );

    \I__618\ : InMux
    port map (
            O => \N__5700\,
            I => \N__5697\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__5697\,
            I => \mem_LUT_data_raw_r_6\
        );

    \I__616\ : InMux
    port map (
            O => \N__5694\,
            I => \N__5688\
        );

    \I__615\ : InMux
    port map (
            O => \N__5693\,
            I => \N__5688\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__5688\,
            I => \r_Tx_Data_4\
        );

    \I__613\ : InMux
    port map (
            O => \N__5685\,
            I => \N__5679\
        );

    \I__612\ : InMux
    port map (
            O => \N__5684\,
            I => \N__5679\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__5679\,
            I => \r_Tx_Data_5\
        );

    \I__610\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5673\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__5673\,
            I => \N__5670\
        );

    \I__608\ : Odrv12
    port map (
            O => \N__5670\,
            I => \pc_tx.n3319\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__5667\,
            I => \reset_all_w_N_61_cascade_\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__5664\,
            I => \n2_adj_505_cascade_\
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__5661\,
            I => \N__5658\
        );

    \I__604\ : InMux
    port map (
            O => \N__5658\,
            I => \N__5649\
        );

    \I__603\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5649\
        );

    \I__602\ : InMux
    port map (
            O => \N__5656\,
            I => \N__5649\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__5649\,
            I => \reset_all_w_N_61\
        );

    \I__600\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5638\
        );

    \I__599\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5638\
        );

    \I__598\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5633\
        );

    \I__597\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5633\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__5638\,
            I => reset_clk_counter_2
        );

    \I__595\ : LocalMux
    port map (
            O => \N__5633\,
            I => reset_clk_counter_2
        );

    \I__594\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5619\
        );

    \I__593\ : InMux
    port map (
            O => \N__5627\,
            I => \N__5619\
        );

    \I__592\ : InMux
    port map (
            O => \N__5626\,
            I => \N__5619\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__5619\,
            I => reset_clk_counter_3
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__5616\,
            I => \N__5610\
        );

    \I__589\ : InMux
    port map (
            O => \N__5615\,
            I => \N__5598\
        );

    \I__588\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5598\
        );

    \I__587\ : InMux
    port map (
            O => \N__5613\,
            I => \N__5598\
        );

    \I__586\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5598\
        );

    \I__585\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5598\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__5598\,
            I => reset_clk_counter_1
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__5595\,
            I => \N__5588\
        );

    \I__582\ : InMux
    port map (
            O => \N__5594\,
            I => \N__5574\
        );

    \I__581\ : InMux
    port map (
            O => \N__5593\,
            I => \N__5574\
        );

    \I__580\ : InMux
    port map (
            O => \N__5592\,
            I => \N__5574\
        );

    \I__579\ : InMux
    port map (
            O => \N__5591\,
            I => \N__5574\
        );

    \I__578\ : InMux
    port map (
            O => \N__5588\,
            I => \N__5574\
        );

    \I__577\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5574\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__5574\,
            I => reset_clk_counter_0
        );

    \I__575\ : InMux
    port map (
            O => \N__5571\,
            I => \N__5565\
        );

    \I__574\ : InMux
    port map (
            O => \N__5570\,
            I => \N__5565\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__5565\,
            I => fifo_temp_output_0
        );

    \I__572\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5556\
        );

    \I__571\ : InMux
    port map (
            O => \N__5561\,
            I => \N__5556\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__5556\,
            I => \r_Tx_Data_0\
        );

    \I__569\ : InMux
    port map (
            O => \N__5553\,
            I => \N__5550\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__5550\,
            I => \mem_LUT_data_raw_r_2\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__5547\,
            I => \N__5544\
        );

    \I__566\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5540\
        );

    \I__565\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5537\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__5540\,
            I => \mem_LUT_mem_1_6\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__5537\,
            I => \mem_LUT_mem_1_6\
        );

    \I__562\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5528\
        );

    \I__561\ : CascadeMux
    port map (
            O => \N__5531\,
            I => \N__5525\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__5528\,
            I => \N__5522\
        );

    \I__559\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5519\
        );

    \I__558\ : Odrv4
    port map (
            O => \N__5522\,
            I => fifo_temp_output_3
        );

    \I__557\ : LocalMux
    port map (
            O => \N__5519\,
            I => fifo_temp_output_3
        );

    \I__556\ : CascadeMux
    port map (
            O => \N__5514\,
            I => \N__5511\
        );

    \I__555\ : InMux
    port map (
            O => \N__5511\,
            I => \N__5507\
        );

    \I__554\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5504\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__5507\,
            I => fifo_temp_output_4
        );

    \I__552\ : LocalMux
    port map (
            O => \N__5504\,
            I => fifo_temp_output_4
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__5499\,
            I => \N__5495\
        );

    \I__550\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5492\
        );

    \I__549\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5489\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__5492\,
            I => fifo_temp_output_5
        );

    \I__547\ : LocalMux
    port map (
            O => \N__5489\,
            I => fifo_temp_output_5
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__5484\,
            I => \n1819_cascade_\
        );

    \I__545\ : SRMux
    port map (
            O => \N__5481\,
            I => \N__5478\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__5478\,
            I => \N__5475\
        );

    \I__543\ : Sp12to4
    port map (
            O => \N__5475\,
            I => \N__5472\
        );

    \I__542\ : Odrv12
    port map (
            O => \N__5472\,
            I => n1898
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__5469\,
            I => \n1898_cascade_\
        );

    \I__540\ : CEMux
    port map (
            O => \N__5466\,
            I => \N__5463\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__5463\,
            I => \N__5460\
        );

    \I__538\ : Span4Mux_v
    port map (
            O => \N__5460\,
            I => \N__5456\
        );

    \I__537\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5453\
        );

    \I__536\ : Odrv4
    port map (
            O => \N__5456\,
            I => n1819
        );

    \I__535\ : LocalMux
    port map (
            O => \N__5453\,
            I => n1819
        );

    \I__534\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5445\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__5445\,
            I => \pc_tx.n2550\
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__5442\,
            I => \pc_tx.n2550_cascade_\
        );

    \I__531\ : InMux
    port map (
            O => \N__5439\,
            I => \N__5436\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__5436\,
            I => \pc_tx.n1484\
        );

    \I__529\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5430\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__5430\,
            I => \N__5424\
        );

    \I__527\ : InMux
    port map (
            O => \N__5429\,
            I => \N__5421\
        );

    \I__526\ : InMux
    port map (
            O => \N__5428\,
            I => \N__5416\
        );

    \I__525\ : InMux
    port map (
            O => \N__5427\,
            I => \N__5416\
        );

    \I__524\ : Odrv4
    port map (
            O => \N__5424\,
            I => \pc_tx.r_Bit_Index_1\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__5421\,
            I => \pc_tx.r_Bit_Index_1\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__5416\,
            I => \pc_tx.r_Bit_Index_1\
        );

    \I__521\ : InMux
    port map (
            O => \N__5409\,
            I => \N__5403\
        );

    \I__520\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5403\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__5403\,
            I => \N__5398\
        );

    \I__518\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5395\
        );

    \I__517\ : InMux
    port map (
            O => \N__5401\,
            I => \N__5392\
        );

    \I__516\ : Odrv4
    port map (
            O => \N__5398\,
            I => \pc_tx.r_Bit_Index_2\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__5395\,
            I => \pc_tx.r_Bit_Index_2\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__5392\,
            I => \pc_tx.r_Bit_Index_2\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__5385\,
            I => \pc_tx.n3385_cascade_\
        );

    \I__512\ : InMux
    port map (
            O => \N__5382\,
            I => \N__5379\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__5379\,
            I => \pc_tx.n3323\
        );

    \I__510\ : InMux
    port map (
            O => \N__5376\,
            I => \N__5373\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__5373\,
            I => \pc_tx.n3322\
        );

    \I__508\ : InMux
    port map (
            O => \N__5370\,
            I => \N__5364\
        );

    \I__507\ : InMux
    port map (
            O => \N__5369\,
            I => \N__5364\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__5364\,
            I => \r_Tx_Data_3\
        );

    \I__505\ : InMux
    port map (
            O => \N__5361\,
            I => \N__5357\
        );

    \I__504\ : InMux
    port map (
            O => \N__5360\,
            I => \N__5354\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__5357\,
            I => \r_Tx_Data_2\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__5354\,
            I => \r_Tx_Data_2\
        );

    \I__501\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5343\
        );

    \I__500\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5343\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__5343\,
            I => fifo_temp_output_2
        );

    \I__498\ : IoInMux
    port map (
            O => \N__5340\,
            I => \N__5337\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__5337\,
            I => \N__5334\
        );

    \I__496\ : IoSpan4Mux
    port map (
            O => \N__5334\,
            I => \N__5331\
        );

    \I__495\ : Sp12to4
    port map (
            O => \N__5331\,
            I => \N__5328\
        );

    \I__494\ : Span12Mux_s6_v
    port map (
            O => \N__5328\,
            I => \N__5325\
        );

    \I__493\ : Odrv12
    port map (
            O => \N__5325\,
            I => \RESET_c\
        );

    \I__492\ : IoInMux
    port map (
            O => \N__5322\,
            I => \N__5319\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__5319\,
            I => \N__5316\
        );

    \I__490\ : Span4Mux_s2_v
    port map (
            O => \N__5316\,
            I => \N__5313\
        );

    \I__489\ : Sp12to4
    port map (
            O => \N__5313\,
            I => \N__5310\
        );

    \I__488\ : Span12Mux_h
    port map (
            O => \N__5310\,
            I => \N__5306\
        );

    \I__487\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5303\
        );

    \I__486\ : Span12Mux_h
    port map (
            O => \N__5306\,
            I => \N__5300\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__5303\,
            I => \N__5297\
        );

    \I__484\ : Span12Mux_v
    port map (
            O => \N__5300\,
            I => \N__5294\
        );

    \I__483\ : Span4Mux_v
    port map (
            O => \N__5297\,
            I => \N__5291\
        );

    \I__482\ : Span12Mux_v
    port map (
            O => \N__5294\,
            I => \N__5288\
        );

    \I__481\ : Span4Mux_h
    port map (
            O => \N__5291\,
            I => \N__5285\
        );

    \I__480\ : Odrv12
    port map (
            O => \N__5288\,
            I => \DEBUG_9_c_c\
        );

    \I__479\ : Odrv4
    port map (
            O => \N__5285\,
            I => \DEBUG_9_c_c\
        );

    \I__478\ : IoInMux
    port map (
            O => \N__5280\,
            I => \N__5277\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__5277\,
            I => \N__5273\
        );

    \I__476\ : IoInMux
    port map (
            O => \N__5276\,
            I => \N__5270\
        );

    \I__475\ : IoSpan4Mux
    port map (
            O => \N__5273\,
            I => \N__5265\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__5270\,
            I => \N__5265\
        );

    \I__473\ : IoSpan4Mux
    port map (
            O => \N__5265\,
            I => \N__5262\
        );

    \I__472\ : Span4Mux_s1_h
    port map (
            O => \N__5262\,
            I => \N__5259\
        );

    \I__471\ : Odrv4
    port map (
            O => \N__5259\,
            I => \FT_OE_c\
        );

    \I__470\ : ClkMux
    port map (
            O => \N__5256\,
            I => \N__5250\
        );

    \I__469\ : ClkMux
    port map (
            O => \N__5255\,
            I => \N__5250\
        );

    \I__468\ : GlobalMux
    port map (
            O => \N__5250\,
            I => \N__5247\
        );

    \I__467\ : gio2CtrlBuf
    port map (
            O => \N__5247\,
            I => \FIFO_CLK_c\
        );

    \I__466\ : InMux
    port map (
            O => \N__5244\,
            I => \N__5241\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__464\ : Glb2LocalMux
    port map (
            O => \N__5238\,
            I => \N__5235\
        );

    \I__463\ : GlobalMux
    port map (
            O => \N__5235\,
            I => pll_clk_unbuf
        );

    \I__462\ : IoInMux
    port map (
            O => \N__5232\,
            I => \N__5229\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__5229\,
            I => \N__5226\
        );

    \I__460\ : IoSpan4Mux
    port map (
            O => \N__5226\,
            I => \N__5223\
        );

    \I__459\ : Sp12to4
    port map (
            O => \N__5223\,
            I => \N__5220\
        );

    \I__458\ : Span12Mux_h
    port map (
            O => \N__5220\,
            I => \N__5217\
        );

    \I__457\ : Odrv12
    port map (
            O => \N__5217\,
            I => \GB_BUFFER_pll_clk_unbuf_THRU_CO\
        );

    \I__456\ : IoInMux
    port map (
            O => \N__5214\,
            I => \N__5211\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__5211\,
            I => \N__5208\
        );

    \I__454\ : Span4Mux_s3_v
    port map (
            O => \N__5208\,
            I => \N__5205\
        );

    \I__453\ : Sp12to4
    port map (
            O => \N__5205\,
            I => \N__5202\
        );

    \I__452\ : Span12Mux_h
    port map (
            O => \N__5202\,
            I => \N__5199\
        );

    \I__451\ : Span12Mux_v
    port map (
            O => \N__5199\,
            I => \N__5196\
        );

    \I__450\ : Odrv12
    port map (
            O => \N__5196\,
            I => \ICE_SYSCLK_c\
        );

    \I__449\ : IoInMux
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__5190\,
            I => \N__5187\
        );

    \I__447\ : Odrv4
    port map (
            O => \N__5187\,
            I => \DEBUG_8_c_c\
        );

    \INVspi0.tx_shift_reg_i0C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i0C_net\,
            I => \N__10627\
        );

    \INVspi0.tx_shift_reg_i6C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i6C_net\,
            I => \N__10684\
        );

    \INVspi0.tx_shift_reg_i14C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i14C_net\,
            I => \N__10697\
        );

    \INVspi0.tx_shift_reg_i12C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i12C_net\,
            I => \N__10685\
        );

    \INVspi0.tx_shift_reg_i15C\ : INV
    port map (
            O => \INVspi0.tx_shift_reg_i15C_net\,
            I => \N__10690\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pc_tx.n2936\,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pc_rx.n2927\,
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_24_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_6_0_\
        );

    \IN_MUX_bfv_24_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2945,
            carryinitout => \bfn_24_7_0_\
        );

    \IN_MUX_bfv_24_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2953,
            carryinitout => \bfn_24_8_0_\
        );

    \IN_MUX_bfv_24_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2961,
            carryinitout => \bfn_24_9_0_\
        );

    \clk_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5232\,
            GLOBALBUFFEROUTPUT => \SLM_CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \FT_OE_r_200_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5309\,
            lcout => \FT_OE_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_pll_clk_unbuf_THRU_LUT4_0_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5244\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_pll_clk_unbuf_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Bit_Index_i2_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__5951\,
            in1 => \N__5401\,
            in2 => \_gnd_net_\,
            in3 => \N__5428\,
            lcout => \pc_tx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12459\,
            ce => \N__5466\,
            sr => \N__5481\
        );

    \pc_tx.r_Bit_Index_i1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__5427\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5950\,
            lcout => \pc_tx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12459\,
            ce => \N__5466\,
            sr => \N__5481\
        );

    \pc_tx.i2936_3_lut_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__5965\,
            in1 => \N__5369\,
            in2 => \_gnd_net_\,
            in3 => \N__5361\,
            lcout => \pc_tx.n3323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i3_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5370\,
            in1 => \N__5532\,
            in2 => \_gnd_net_\,
            in3 => \N__6349\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i2_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5360\,
            in1 => \N__6359\,
            in2 => \_gnd_net_\,
            in3 => \N__5348\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12464\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i5_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__5856\,
            in1 => \N__9536\,
            in2 => \N__5499\,
            in3 => \N__6656\,
            lcout => fifo_temp_output_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12464\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i2_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__6655\,
            in1 => \N__5349\,
            in2 => \N__9573\,
            in3 => \N__5553\,
            lcout => fifo_temp_output_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12464\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i1722_1_lut_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9493\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESET_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i1_3_lut_4_lut_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__6837\,
            in1 => \N__6876\,
            in2 => \N__7146\,
            in3 => \N__7245\,
            lcout => n1819,
            ltout => \n1819_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i1545_3_lut_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6836\,
            in2 => \N__5484\,
            in3 => \N__5448\,
            lcout => n1898,
            ltout => \n1898_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Bit_Index_i0_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5949\,
            in2 => \N__5469\,
            in3 => \N__5459\,
            lcout => \r_Bit_Index_0_adj_498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12462\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2_3_lut_4_lut_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__6838\,
            in1 => \N__7246\,
            in2 => \N__6891\,
            in3 => \N__5757\,
            lcout => n1636,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2_2_lut_3_lut_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5402\,
            in1 => \N__5429\,
            in2 => \_gnd_net_\,
            in3 => \N__5948\,
            lcout => \pc_tx.n2550\,
            ltout => \pc_tx.n2550_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i1132_4_lut_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__5756\,
            in1 => \N__7141\,
            in2 => \N__5442\,
            in3 => \N__6835\,
            lcout => \pc_tx.n1484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_SM_Main_i0_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__5439\,
            in1 => \N__7125\,
            in2 => \_gnd_net_\,
            in3 => \N__6875\,
            lcout => \r_SM_Main_0_adj_497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12458\,
            ce => 'H',
            sr => \N__7253\
        );

    \pc_tx.r_Bit_Index_1__bdd_4_lut_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__5433\,
            in1 => \N__5409\,
            in2 => \N__5916\,
            in3 => \N__5676\,
            lcout => OPEN,
            ltout => \pc_tx.n3385_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.n3385_bdd_4_lut_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__5408\,
            in1 => \N__5376\,
            in2 => \N__5385\,
            in3 => \N__5382\,
            lcout => \pc_tx.o_Tx_Serial_N_216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2935_3_lut_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__5964\,
            in1 => \N__5829\,
            in2 => \_gnd_net_\,
            in3 => \N__5561\,
            lcout => \pc_tx.n3322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i152_153_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5543\,
            in1 => \N__7527\,
            in2 => \_gnd_net_\,
            in3 => \N__8944\,
            lcout => \mem_LUT_mem_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i0_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__5571\,
            in1 => \N__9530\,
            in2 => \N__5715\,
            in3 => \N__6651\,
            lcout => fifo_temp_output_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i0_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5562\,
            in1 => \N__6348\,
            in2 => \_gnd_net_\,
            in3 => \N__5570\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i3_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__6567\,
            in1 => \N__5904\,
            in2 => \N__6126\,
            in3 => \N__7881\,
            lcout => \mem_LUT_data_raw_r_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12469\,
            ce => \N__6536\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i7_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__5801\,
            in1 => \N__5844\,
            in2 => \N__5547\,
            in3 => \N__7882\,
            lcout => \mem_LUT_data_raw_r_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12469\,
            ce => \N__6536\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i3_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__6204\,
            in1 => \N__9481\,
            in2 => \N__5531\,
            in3 => \N__6652\,
            lcout => fifo_temp_output_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i4_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6351\,
            in1 => \N__5694\,
            in2 => \_gnd_net_\,
            in3 => \N__5510\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i4_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__5898\,
            in1 => \N__9482\,
            in2 => \N__5514\,
            in3 => \N__6653\,
            lcout => fifo_temp_output_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i5_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5498\,
            in1 => \N__5685\,
            in2 => \_gnd_net_\,
            in3 => \N__6352\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i6_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__6374\,
            in1 => \N__9483\,
            in2 => \N__5703\,
            in3 => \N__6654\,
            lcout => fifo_temp_output_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2932_3_lut_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5693\,
            in1 => \N__5684\,
            in2 => \_gnd_net_\,
            in3 => \N__5969\,
            lcout => \pc_tx.n3319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5626\,
            in1 => \N__5609\,
            in2 => \N__5595\,
            in3 => \N__5643\,
            lcout => \reset_all_w_N_61\,
            ltout => \reset_all_w_N_61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_clk_counter_i3_582__i1_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001011010"
        )
    port map (
            in0 => \N__5613\,
            in1 => \_gnd_net_\,
            in2 => \N__5667\,
            in3 => \N__5593\,
            lcout => reset_clk_counter_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_clk_counter_i3_582__i2_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010011100"
        )
    port map (
            in0 => \N__5614\,
            in1 => \N__5645\,
            in2 => \N__5661\,
            in3 => \N__5594\,
            lcout => reset_clk_counter_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2550_2_lut_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__5587\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5656\,
            lcout => OPEN,
            ltout => \n2_adj_505_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_clk_counter_i3_582__i3_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001001"
        )
    port map (
            in0 => \N__5615\,
            in1 => \N__5628\,
            in2 => \N__5664\,
            in3 => \N__5646\,
            lcout => reset_clk_counter_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_clk_counter_i3_582__i0_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__5592\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5657\,
            lcout => reset_clk_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_all_r_198_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5644\,
            in1 => \N__5627\,
            in2 => \N__5616\,
            in3 => \N__5591\,
            lcout => reset_all_w,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_read_cmd_205_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6078\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5772\,
            lcout => fifo_read_cmd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_SM_Main_i2_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7241\,
            in1 => \N__6833\,
            in2 => \N__6892\,
            in3 => \N__7140\,
            lcout => \r_SM_Main_2_adj_495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2966_4_lut_4_lut_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000001100"
        )
    port map (
            in0 => \N__7139\,
            in1 => \N__5754\,
            in2 => \N__6839\,
            in3 => \N__6880\,
            lcout => OPEN,
            ltout => \n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Active_46_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011100"
        )
    port map (
            in0 => \N__6834\,
            in1 => \N__5770\,
            in2 => \N__5775\,
            in3 => \N__7242\,
            lcout => tx_uart_active_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \start_tx_206_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__5755\,
            in1 => \N__7918\,
            in2 => \N__6079\,
            in3 => \N__5771\,
            lcout => \r_SM_Main_2_N_187_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_SM_Main_2__I_0_55_i3_3_lut_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101111"
        )
    port map (
            in0 => \N__5739\,
            in1 => \_gnd_net_\,
            in2 => \N__6840\,
            in3 => \N__6881\,
            lcout => \pc_tx.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i8_2_lut_3_lut_4_lut_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__8297\,
            in1 => \N__8266\,
            in2 => \N__8432\,
            in3 => \N__8386\,
            lcout => n4_adj_494,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_r__i0_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110100110"
        )
    port map (
            in0 => \N__8298\,
            in1 => \N__8387\,
            in2 => \N__8433\,
            in3 => \N__9589\,
            lcout => wr_addr_r_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12460\,
            ce => 'H',
            sr => \N__9587\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r__i0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000110110"
        )
    port map (
            in0 => \N__9588\,
            in1 => \N__7994\,
            in2 => \N__7943\,
            in3 => \N__6061\,
            lcout => rd_addr_r_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12460\,
            ce => 'H',
            sr => \N__9587\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100100"
        )
    port map (
            in0 => \N__7065\,
            in1 => \N__5997\,
            in2 => \N__7850\,
            in3 => \N__5817\,
            lcout => \mem_LUT_data_raw_r_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12467\,
            ce => \N__6529\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i6_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__7817\,
            in1 => \N__6021\,
            in2 => \N__6012\,
            in3 => \N__6396\,
            lcout => \mem_LUT_data_raw_r_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12467\,
            ce => \N__6529\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3014_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__5838\,
            in1 => \N__7799\,
            in2 => \N__8043\,
            in3 => \N__6594\,
            lcout => \tx_fifo.lscc_fifo_inst.n3397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i248_249_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__8946\,
            in1 => \N__8267\,
            in2 => \N__6767\,
            in3 => \N__5837\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6350\,
            in1 => \N__5828\,
            in2 => \_gnd_net_\,
            in3 => \N__6612\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i134_135_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5813\,
            in1 => \N__7526\,
            in2 => \_gnd_net_\,
            in3 => \N__8649\,
            lcout => \mem_LUT_mem_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12476\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i56_57_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__6771\,
            in1 => \N__8268\,
            in2 => \N__5802\,
            in3 => \N__8945\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12476\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_fifo_en_prev_r_86_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7939\,
            in1 => \N__9569\,
            in2 => \_gnd_net_\,
            in3 => \N__6081\,
            lcout => rd_fifo_en_prev_r,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12476\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_28_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__7938\,
            in1 => \N__9567\,
            in2 => \N__5787\,
            in3 => \N__6080\,
            lcout => n1795,
            ltout => \n1795_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i7_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__9568\,
            in1 => \N__6231\,
            in2 => \N__5778\,
            in3 => \N__5885\,
            lcout => fifo_temp_output_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12476\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__8037\,
            in1 => \N__6264\,
            in2 => \N__7851\,
            in3 => \N__6252\,
            lcout => \tx_fifo.lscc_fifo_inst.n3433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i5_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__7876\,
            in1 => \N__5874\,
            in2 => \N__6282\,
            in3 => \N__6987\,
            lcout => \mem_LUT_data_raw_r_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12481\,
            ce => \N__6537\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_en_i_I_0_2_lut_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7919\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6077\,
            lcout => rd_fifo_en_w,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2991_4_lut_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110001"
        )
    port map (
            in0 => \N__6826\,
            in1 => \N__7244\,
            in2 => \N__7145\,
            in3 => \N__6899\,
            lcout => \pc_tx.n1919\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i7_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6337\,
            in1 => \N__5981\,
            in2 => \_gnd_net_\,
            in3 => \N__5892\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i1_1_lut_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7243\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pc_tx.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3019_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__6092\,
            in1 => \N__7844\,
            in2 => \N__6108\,
            in3 => \N__7997\,
            lcout => \tx_fifo.lscc_fifo_inst.n3403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_31_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__8300\,
            in1 => \N__8257\,
            in2 => \N__7875\,
            in3 => \N__7996\,
            lcout => OPEN,
            ltout => \n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__8388\,
            in1 => \_gnd_net_\,
            in2 => \N__5862\,
            in3 => \N__6060\,
            lcout => OPEN,
            ltout => \n24_adj_510_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.empty_r_85_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__6027\,
            in1 => \N__9590\,
            in2 => \N__5859\,
            in3 => \N__6459\,
            lcout => is_fifo_empty_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i338_339_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6104\,
            in1 => \N__7186\,
            in2 => \_gnd_net_\,
            in3 => \N__10437\,
            lcout => \mem_LUT_mem_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i242_243_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__8258\,
            in1 => \N__6732\,
            in2 => \N__6093\,
            in3 => \N__10436\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000000"
        )
    port map (
            in0 => \N__8299\,
            in1 => \N__7995\,
            in2 => \N__6076\,
            in3 => \N__7937\,
            lcout => n4_adj_511,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3024_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__6180\,
            in1 => \N__7800\,
            in2 => \N__8038\,
            in3 => \N__6171\,
            lcout => \tx_fifo.lscc_fifo_inst.n3409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i4_2_lut_3_lut_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__8301\,
            in1 => \N__8420\,
            in2 => \_gnd_net_\,
            in3 => \N__8377\,
            lcout => \tx_fifo.lscc_fifo_inst.n4\,
            ltout => \tx_fifo.lscc_fifo_inst.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i53_54_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__6008\,
            in1 => \N__8245\,
            in2 => \N__6015\,
            in3 => \N__10334\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i38_39_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__8244\,
            in1 => \N__5996\,
            in2 => \N__8655\,
            in3 => \N__6725\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2933_3_lut_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6300\,
            in1 => \N__5985\,
            in2 => \_gnd_net_\,
            in3 => \N__5970\,
            lcout => \pc_tx.n3320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i329_330_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6446\,
            in1 => \N__7202\,
            in2 => \_gnd_net_\,
            in3 => \N__8594\,
            lcout => \mem_LUT_mem_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i245_246_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__8243\,
            in1 => \N__6724\,
            in2 => \N__10335\,
            in3 => \N__6179\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r__i1_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__9531\,
            in1 => \N__8041\,
            in2 => \N__6527\,
            in3 => \N__7798\,
            lcout => rd_addr_r_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i347_348_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6143\,
            in1 => \N__7204\,
            in2 => \_gnd_net_\,
            in3 => \N__10481\,
            lcout => \mem_LUT_mem_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i341_342_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7203\,
            in1 => \N__6170\,
            in2 => \_gnd_net_\,
            in3 => \N__10330\,
            lcout => \mem_LUT_mem_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3009_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__6158\,
            in1 => \N__8039\,
            in2 => \N__7839\,
            in3 => \N__6579\,
            lcout => \tx_fifo.lscc_fifo_inst.n3391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i239_240_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__8895\,
            in1 => \N__8260\,
            in2 => \N__6159\,
            in3 => \N__6730\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3029_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__6144\,
            in1 => \N__8040\,
            in2 => \N__7840\,
            in3 => \N__6135\,
            lcout => \tx_fifo.lscc_fifo_inst.n3415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i251_252_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__6134\,
            in1 => \N__8261\,
            in2 => \N__10482\,
            in3 => \N__6731\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i44_45_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__8263\,
            in1 => \N__6758\,
            in2 => \N__10398\,
            in3 => \N__6119\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Tx_Data_i6_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6381\,
            in1 => \N__6293\,
            in2 => \_gnd_net_\,
            in3 => \N__6363\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i50_51_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__8265\,
            in1 => \N__10430\,
            in2 => \N__6281\,
            in3 => \N__6762\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i236_237_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__6263\,
            in1 => \N__8262\,
            in2 => \N__6769\,
            in3 => \N__10393\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i332_333_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6251\,
            in1 => \N__7205\,
            in2 => \_gnd_net_\,
            in3 => \N__10394\,
            lcout => \mem_LUT_mem_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i47_48_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__6215\,
            in1 => \N__8264\,
            in2 => \N__6770\,
            in3 => \N__8894\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12482\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i8_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100110101000"
        )
    port map (
            in0 => \N__6240\,
            in1 => \N__7849\,
            in2 => \N__7476\,
            in3 => \N__6675\,
            lcout => \mem_LUT_data_raw_r_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12486\,
            ce => \N__6528\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i4_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__6225\,
            in1 => \N__6216\,
            in2 => \N__7002\,
            in3 => \N__7848\,
            lcout => \mem_LUT_data_raw_r_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12486\,
            ce => \N__6528\,
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i15_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6552\,
            in2 => \_gnd_net_\,
            in3 => \N__7652\,
            lcout => \SDAT_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i15C_net\,
            ce => 'H',
            sr => \N__6954\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_raw_r__i2_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__6411\,
            in1 => \N__6435\,
            in2 => \N__6429\,
            in3 => \N__7874\,
            lcout => \mem_LUT_data_raw_r_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12478\,
            ce => \N__6510\,
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i230_231_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__8256\,
            in1 => \N__7088\,
            in2 => \N__6766\,
            in3 => \N__8654\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12468\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i779_3_lut_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__8086\,
            in1 => \N__8028\,
            in2 => \_gnd_net_\,
            in3 => \N__7878\,
            lcout => rd_addr_p1_w_2,
            ltout => \rd_addr_p1_w_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r__i2_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__8087\,
            in1 => \N__9594\,
            in2 => \N__6540\,
            in3 => \N__6511\,
            lcout => rd_addr_r_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12468\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i772_rep_9_2_lut_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8027\,
            in2 => \_gnd_net_\,
            in3 => \N__7877\,
            lcout => OPEN,
            ltout => \n3448_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2902_4_lut_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__8255\,
            in1 => \N__8061\,
            in2 => \N__6468\,
            in3 => \N__6465\,
            lcout => n3289,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3039_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__7879\,
            in1 => \N__6783\,
            in2 => \N__6453\,
            in3 => \N__8029\,
            lcout => \tx_fifo.lscc_fifo_inst.n3427\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i41_42_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__6422\,
            in1 => \N__8215\,
            in2 => \N__6754\,
            in3 => \N__8593\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i137_138_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8589\,
            in1 => \N__7529\,
            in2 => \_gnd_net_\,
            in3 => \N__6407\,
            lcout => \mem_LUT_mem_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i149_150_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7530\,
            in1 => \N__6392\,
            in2 => \_gnd_net_\,
            in3 => \N__10321\,
            lcout => \mem_LUT_mem_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i233_234_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__8214\,
            in1 => \N__6726\,
            in2 => \N__8595\,
            in3 => \N__6782\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i59_60_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__10472\,
            in1 => \N__8259\,
            in2 => \N__6768\,
            in3 => \N__6671\,
            lcout => \tx_fifo.lscc_fifo_inst.mem_LUT_mem_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12483\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.mem_LUT_data_buff_r__i1_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__9532\,
            in1 => \N__6660\,
            in2 => \N__6611\,
            in3 => \N__6621\,
            lcout => fifo_temp_output_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12483\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i3_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11313\,
            in1 => \N__11904\,
            in2 => \_gnd_net_\,
            in3 => \N__6940\,
            lcout => tx_data_byte_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12483\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i344_345_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8934\,
            in1 => \N__7198\,
            in2 => \_gnd_net_\,
            in3 => \N__6590\,
            lcout => \mem_LUT_mem_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12483\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i4_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11901\,
            in1 => \N__9068\,
            in2 => \_gnd_net_\,
            in3 => \N__6965\,
            lcout => tx_addr_byte_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i335_336_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7206\,
            in1 => \N__6578\,
            in2 => \_gnd_net_\,
            in3 => \N__8893\,
            lcout => \mem_LUT_mem_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i140_141_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10385\,
            in1 => \N__7531\,
            in2 => \_gnd_net_\,
            in3 => \N__6563\,
            lcout => \mem_LUT_mem_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i7_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6551\,
            in1 => \N__11267\,
            in2 => \_gnd_net_\,
            in3 => \N__11903\,
            lcout => tx_addr_byte_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i143_144_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6998\,
            in1 => \N__7532\,
            in2 => \_gnd_net_\,
            in3 => \N__8886\,
            lcout => \mem_LUT_mem_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i3_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6947\,
            in1 => \N__11902\,
            in2 => \_gnd_net_\,
            in3 => \N__6923\,
            lcout => tx_addr_byte_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i146_147_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10423\,
            in1 => \N__7533\,
            in2 => \_gnd_net_\,
            in3 => \N__6983\,
            lcout => \mem_LUT_mem_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i12_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__10769\,
            in1 => \N__6912\,
            in2 => \N__6972\,
            in3 => \N__7645\,
            lcout => tx_shift_reg_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i12C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i1_2_lut_adj_16_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7452\,
            in2 => \_gnd_net_\,
            in3 => \N__10766\,
            lcout => \spi0.n3176\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i3_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__10770\,
            in1 => \N__6948\,
            in2 => \N__7710\,
            in3 => \N__7646\,
            lcout => tx_shift_reg_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i12C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i11_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__7644\,
            in1 => \N__6906\,
            in2 => \N__6927\,
            in3 => \N__10768\,
            lcout => tx_shift_reg_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i12C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i10_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__10767\,
            in1 => \N__7581\,
            in2 => \N__11061\,
            in3 => \N__7643\,
            lcout => tx_shift_reg_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i12C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_SM_Main_i1_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__6803\,
            in1 => \N__7110\,
            in2 => \_gnd_net_\,
            in3 => \N__6900\,
            lcout => \r_SM_Main_1_adj_496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12484\,
            ce => 'H',
            sr => \N__7254\
        );

    \tx_fifo.lscc_fifo_inst.EnabledDecoder_2_i7_2_lut_3_lut_4_lut_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__8413\,
            in1 => \N__8198\,
            in2 => \N__8324\,
            in3 => \N__8367\,
            lcout => n2,
            ltout => \n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i326_327_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__7073\,
            in1 => \_gnd_net_\,
            in2 => \N__7155\,
            in3 => \N__8650\,
            lcout => \mem_LUT_mem_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12474\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i3_4_lut_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7425\,
            in1 => \N__7017\,
            in2 => \N__7035\,
            in3 => \N__7053\,
            lcout => OPEN,
            ltout => \pc_tx.n2981_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2212_4_lut_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__7380\,
            in1 => \N__7395\,
            in2 => \N__7152\,
            in3 => \N__7410\,
            lcout => OPEN,
            ltout => \pc_tx.n2564_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.i2218_4_lut_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__7365\,
            in1 => \N__7329\,
            in2 => \N__7149\,
            in3 => \N__7350\,
            lcout => \r_SM_Main_2_N_184_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.rd_addr_r_0__bdd_4_lut_3034_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__7089\,
            in1 => \N__7880\,
            in2 => \N__7077\,
            in3 => \N__8030\,
            lcout => \tx_fifo.lscc_fifo_inst.n3421\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_tx.r_Clock_Count_586__i0_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7049\,
            in2 => \_gnd_net_\,
            in3 => \N__7038\,
            lcout => \pc_tx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \pc_tx.n2929\,
            clk => \N__12485\,
            ce => \N__7309\,
            sr => \N__7277\
        );

    \pc_tx.r_Clock_Count_586__i1_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7031\,
            in2 => \_gnd_net_\,
            in3 => \N__7020\,
            lcout => \pc_tx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \pc_tx.n2929\,
            carryout => \pc_tx.n2930\,
            clk => \N__12485\,
            ce => \N__7309\,
            sr => \N__7277\
        );

    \pc_tx.r_Clock_Count_586__i2_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7016\,
            in2 => \_gnd_net_\,
            in3 => \N__7005\,
            lcout => \pc_tx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \pc_tx.n2930\,
            carryout => \pc_tx.n2931\,
            clk => \N__12485\,
            ce => \N__7309\,
            sr => \N__7277\
        );

    \pc_tx.r_Clock_Count_586__i3_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7424\,
            in2 => \_gnd_net_\,
            in3 => \N__7413\,
            lcout => \pc_tx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \pc_tx.n2931\,
            carryout => \pc_tx.n2932\,
            clk => \N__12485\,
            ce => \N__7309\,
            sr => \N__7277\
        );

    \pc_tx.r_Clock_Count_586__i4_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7409\,
            in2 => \_gnd_net_\,
            in3 => \N__7398\,
            lcout => \pc_tx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \pc_tx.n2932\,
            carryout => \pc_tx.n2933\,
            clk => \N__12485\,
            ce => \N__7309\,
            sr => \N__7277\
        );

    \pc_tx.r_Clock_Count_586__i5_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7394\,
            in2 => \_gnd_net_\,
            in3 => \N__7383\,
            lcout => \pc_tx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \pc_tx.n2933\,
            carryout => \pc_tx.n2934\,
            clk => \N__12485\,
            ce => \N__7309\,
            sr => \N__7277\
        );

    \pc_tx.r_Clock_Count_586__i6_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7379\,
            in2 => \_gnd_net_\,
            in3 => \N__7368\,
            lcout => \pc_tx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \pc_tx.n2934\,
            carryout => \pc_tx.n2935\,
            clk => \N__12485\,
            ce => \N__7309\,
            sr => \N__7277\
        );

    \pc_tx.r_Clock_Count_586__i7_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7364\,
            in2 => \_gnd_net_\,
            in3 => \N__7353\,
            lcout => \pc_tx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \pc_tx.n2935\,
            carryout => \pc_tx.n2936\,
            clk => \N__12485\,
            ce => \N__7309\,
            sr => \N__7277\
        );

    \pc_tx.r_Clock_Count_586__i8_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7346\,
            in2 => \_gnd_net_\,
            in3 => \N__7335\,
            lcout => \pc_tx.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \pc_tx.n2937\,
            clk => \N__12488\,
            ce => \N__7310\,
            sr => \N__7278\
        );

    \pc_tx.r_Clock_Count_586__i9_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__7325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7332\,
            lcout => \pc_tx.r_Clock_Count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12488\,
            ce => \N__7310\,
            sr => \N__7278\
        );

    \tx_addr_byte_r_i0_i0_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11900\,
            in1 => \N__8532\,
            in2 => \_gnd_net_\,
            in3 => \N__7679\,
            lcout => tx_addr_byte_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.spi_clk_76_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10592\,
            in2 => \_gnd_net_\,
            in3 => \N__9816\,
            lcout => \spi0.spi_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i155_156_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7466\,
            in1 => \N__7528\,
            in2 => \_gnd_net_\,
            in3 => \N__10471\,
            lcout => \mem_LUT_mem_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i19_3_lut_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110011"
        )
    port map (
            in0 => \N__9393\,
            in1 => \N__9321\,
            in2 => \_gnd_net_\,
            in3 => \N__9225\,
            lcout => n3279,
            ltout => \n3279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i14_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__8136\,
            in1 => \N__7437\,
            in2 => \N__7455\,
            in3 => \N__7648\,
            lcout => \spi0.tx_shift_reg_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i14C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i1_1_lut_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9394\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi0.n890\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i1_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__10772\,
            in1 => \N__9792\,
            in2 => \N__7656\,
            in3 => \N__8118\,
            lcout => tx_shift_reg_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i14C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i13_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__7446\,
            in1 => \N__7647\,
            in2 => \N__8511\,
            in3 => \N__10771\,
            lcout => tx_shift_reg_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i14C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i6_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__7692\,
            in1 => \N__7635\,
            in2 => \N__9039\,
            in3 => \N__10776\,
            lcout => tx_shift_reg_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i4_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__10774\,
            in1 => \N__9072\,
            in2 => \N__7653\,
            in3 => \N__7431\,
            lcout => tx_shift_reg_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i2_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__7716\,
            in1 => \N__7631\,
            in2 => \N__11040\,
            in3 => \N__10773\,
            lcout => tx_shift_reg_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i1_2_lut_3_lut_adj_14_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__9395\,
            in1 => \N__9327\,
            in2 => \_gnd_net_\,
            in3 => \N__9231\,
            lcout => n1728,
            ltout => \n1728_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i5_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__11088\,
            in1 => \N__7701\,
            in2 => \N__7695\,
            in3 => \N__10775\,
            lcout => tx_shift_reg_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i8_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__10778\,
            in1 => \N__7686\,
            in2 => \N__7654\,
            in3 => \N__7662\,
            lcout => tx_shift_reg_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i7_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__7668\,
            in1 => \N__7636\,
            in2 => \N__11274\,
            in3 => \N__10777\,
            lcout => tx_shift_reg_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i9_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__10779\,
            in1 => \N__9774\,
            in2 => \N__7655\,
            in3 => \N__7587\,
            lcout => tx_shift_reg_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i2_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__10794\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7539\,
            lcout => rx_shift_reg_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i1_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__7565\,
            in1 => \N__10793\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rx_shift_reg_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i3_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__10795\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8669\,
            lcout => rx_shift_reg_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_p1_w_1__I_0_i2_2_lut_3_lut_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__7884\,
            in1 => \N__8326\,
            in2 => \_gnd_net_\,
            in3 => \N__8180\,
            lcout => OPEN,
            ltout => \tx_fifo.lscc_fifo_inst.n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i1_4_lut_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__8070\,
            in1 => \N__7950\,
            in2 => \N__8094\,
            in3 => \N__8091\,
            lcout => n2968,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.i757_3_lut_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__8056\,
            in1 => \N__8179\,
            in2 => \_gnd_net_\,
            in3 => \N__8325\,
            lcout => wr_addr_p1_w_2,
            ltout => \wr_addr_p1_w_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_r__i2_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__8343\,
            in1 => \N__8057\,
            in2 => \N__8064\,
            in3 => \N__9597\,
            lcout => wr_addr_r_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12480\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_write_cmd_204_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8538\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8410\,
            lcout => fifo_write_cmd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_r_1__I_0_i1_2_lut_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8042\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8327\,
            lcout => n1,
            ltout => \n1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2889_4_lut_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111110"
        )
    port map (
            in0 => \N__7944\,
            in1 => \N__8177\,
            in2 => \N__7887\,
            in3 => \N__7883\,
            lcout => OPEN,
            ltout => \n3275_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__8411\,
            in1 => \_gnd_net_\,
            in2 => \N__7728\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n15_adj_509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.full_r_84_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__7725\,
            in1 => \N__8342\,
            in2 => \N__7719\,
            in3 => \N__9595\,
            lcout => is_tx_fifo_full_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_en_i_I_0_2_lut_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8412\,
            in2 => \_gnd_net_\,
            in3 => \N__8366\,
            lcout => wr_fifo_en_w,
            ltout => \wr_fifo_en_w_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_fifo.lscc_fifo_inst.wr_addr_r__i1_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__8178\,
            in1 => \N__9596\,
            in2 => \N__8331\,
            in3 => \N__8328\,
            lcout => wr_addr_r_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i6_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9032\,
            in1 => \N__11883\,
            in2 => \_gnd_net_\,
            in3 => \N__8129\,
            lcout => tx_addr_byte_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.tx_shift_reg_i0_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__8528\,
            in1 => \N__9331\,
            in2 => \_gnd_net_\,
            in3 => \N__9260\,
            lcout => tx_shift_reg_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi0.tx_shift_reg_i0C_net\,
            ce => 'H',
            sr => \N__8112\
        );

    \spi0.i2963_2_lut_3_lut_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__9397\,
            in1 => \N__9233\,
            in2 => \_gnd_net_\,
            in3 => \N__9755\,
            lcout => \spi0.n3328\,
            ltout => \spi0.n3328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.mux_512_i3_4_lut_4_lut_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__9329\,
            in1 => \N__8840\,
            in2 => \N__8106\,
            in3 => \N__8449\,
            lcout => \spi0.state_next_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i1077_2_lut_4_lut_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__9396\,
            in1 => \N__9232\,
            in2 => \N__8780\,
            in3 => \N__9328\,
            lcout => \spi0.n1429\,
            ltout => \spi0.n1429_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.state_reg_i2_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__9330\,
            in1 => \N__8841\,
            in2 => \N__8103\,
            in3 => \N__8100\,
            lcout => state_reg_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10698\,
            ce => 'H',
            sr => \N__9591\
        );

    \spi0.state_reg_i0_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__8842\,
            in1 => \_gnd_net_\,
            in2 => \N__8454\,
            in3 => \N__8460\,
            lcout => state_reg_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10698\,
            ce => 'H',
            sr => \N__9591\
        );

    \spi0.t_FSM_i6_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__9236\,
            in1 => \N__9676\,
            in2 => \N__8490\,
            in3 => \N__9726\,
            lcout => \state_next_2__N_312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10698\,
            ce => 'H',
            sr => \N__9591\
        );

    \spi0.t_FSM_i5_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000010000"
        )
    port map (
            in0 => \N__9725\,
            in1 => \N__9235\,
            in2 => \N__8481\,
            in3 => \N__9677\,
            lcout => \spi0.n497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10698\,
            ce => 'H',
            sr => \N__9591\
        );

    \spi0.t_FSM_i4_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__9234\,
            in1 => \N__9675\,
            in2 => \N__9612\,
            in3 => \N__9724\,
            lcout => \spi0.n498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10698\,
            ce => 'H',
            sr => \N__9591\
        );

    \i529_4_lut_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__9324\,
            in1 => \N__9398\,
            in2 => \N__8779\,
            in3 => \N__9228\,
            lcout => n883,
            ltout => \n883_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.state_reg_i1_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__9229\,
            in1 => \N__8850\,
            in2 => \N__8472\,
            in3 => \N__9326\,
            lcout => state_reg_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10701\,
            ce => 'H',
            sr => \N__9593\
        );

    \spi0.i2082_2_lut_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9226\,
            lcout => \spi0.n2433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i2962_4_lut_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100111"
        )
    port map (
            in0 => \N__9227\,
            in1 => \N__8729\,
            in2 => \N__8985\,
            in3 => \N__9322\,
            lcout => OPEN,
            ltout => \spi0.n3337_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i28_4_lut_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__9754\,
            in1 => \N__8469\,
            in2 => \N__8463\,
            in3 => \N__9399\,
            lcout => \spi0.n13\,
            ltout => \spi0.n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.mux_512_i1_3_lut_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__8453\,
            in1 => \_gnd_net_\,
            in2 => \N__8436\,
            in3 => \N__8843\,
            lcout => OPEN,
            ltout => \spi0.state_next_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i1_4_lut_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__9325\,
            in1 => \N__8562\,
            in2 => \N__8556\,
            in3 => \N__9400\,
            lcout => \spi0.n4\,
            ltout => \spi0.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i2_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__9230\,
            in1 => \N__9674\,
            in2 => \N__8553\,
            in3 => \N__8730\,
            lcout => \spi0.state_next_2__N_310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10701\,
            ce => 'H',
            sr => \N__9593\
        );

    \spi0.CS_w_79_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9410\,
            in2 => \_gnd_net_\,
            in3 => \N__9341\,
            lcout => \spi0.CS_w\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10700\,
            ce => 'H',
            sr => \N__9264\
        );

    \spi0.CS_81_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8550\,
            lcout => \SEN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10702\,
            ce => 'H',
            sr => \N__9540\
        );

    \spi_busy_prev_203_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8958\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => spi_busy_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_busy_falling_edge_202_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8544\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8957\,
            lcout => spi_busy_falling_edge,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i0_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8527\,
            in1 => \N__11899\,
            in2 => \_gnd_net_\,
            in3 => \N__11334\,
            lcout => tx_data_byte_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i5_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8501\,
            in1 => \N__11898\,
            in2 => \_gnd_net_\,
            in3 => \N__11084\,
            lcout => tx_addr_byte_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i0_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111110111111110"
        )
    port map (
            in0 => \N__9660\,
            in1 => \N__9727\,
            in2 => \N__8721\,
            in3 => \N__9244\,
            lcout => \spi0.n502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10686\,
            ce => 'H',
            sr => \N__9592\
        );

    \spi0.t_FSM_i1_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000010000"
        )
    port map (
            in0 => \N__9666\,
            in1 => \N__9730\,
            in2 => \N__8739\,
            in3 => \N__9250\,
            lcout => \spi0.state_next_2__N_311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10686\,
            ce => 'H',
            sr => \N__9592\
        );

    \spi0.t_FSM_i15_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__9249\,
            in1 => \N__9665\,
            in2 => \N__8712\,
            in3 => \N__9736\,
            lcout => \spi0.n487\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10686\,
            ce => 'H',
            sr => \N__9592\
        );

    \spi0.t_FSM_i14_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000010000"
        )
    port map (
            in0 => \N__9664\,
            in1 => \N__9729\,
            in2 => \N__8703\,
            in3 => \N__9248\,
            lcout => \spi0.n488\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10686\,
            ce => 'H',
            sr => \N__9592\
        );

    \spi0.t_FSM_i13_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__9247\,
            in1 => \N__9663\,
            in2 => \N__8694\,
            in3 => \N__9735\,
            lcout => \spi0.n489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10686\,
            ce => 'H',
            sr => \N__9592\
        );

    \spi0.t_FSM_i12_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000010000"
        )
    port map (
            in0 => \N__9662\,
            in1 => \N__9728\,
            in2 => \N__8685\,
            in3 => \N__9246\,
            lcout => \spi0.n490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10686\,
            ce => 'H',
            sr => \N__9592\
        );

    \spi0.t_FSM_i11_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__9245\,
            in1 => \N__9661\,
            in2 => \N__8817\,
            in3 => \N__9734\,
            lcout => \spi0.n491\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10686\,
            ce => 'H',
            sr => \N__9592\
        );

    \spi0.state_reg_2__I_0_108_i5_3_lut_3_lut_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__9333\,
            in1 => \N__9239\,
            in2 => \_gnd_net_\,
            in3 => \N__9402\,
            lcout => \rx_shift_reg_15__N_319\,
            ltout => \rx_shift_reg_15__N_319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i0_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8676\,
            in2 => \N__8658\,
            in3 => \N__8613\,
            lcout => rx_buf_byte_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i1_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8573\,
            in1 => \N__10500\,
            in2 => \_gnd_net_\,
            in3 => \N__10356\,
            lcout => rx_buf_byte_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.busy_86_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__9240\,
            in1 => \N__9406\,
            in2 => \_gnd_net_\,
            in3 => \N__9334\,
            lcout => spi_busy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i6_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10269\,
            in1 => \N__8913\,
            in2 => \_gnd_net_\,
            in3 => \N__10358\,
            lcout => rx_buf_byte_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i3_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10357\,
            in1 => \N__8866\,
            in2 => \_gnd_net_\,
            in3 => \N__10281\,
            lcout => rx_buf_byte_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i1_2_lut_3_lut_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8775\,
            in1 => \N__9237\,
            in2 => \_gnd_net_\,
            in3 => \N__9401\,
            lcout => \spi0.n906\,
            ltout => \spi0.n906_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.mux_512_i2_4_lut_4_lut_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__9238\,
            in1 => \N__8844\,
            in2 => \N__8820\,
            in3 => \N__9332\,
            lcout => \spi0.state_next_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.t_FSM_i10_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000010000"
        )
    port map (
            in0 => \N__9667\,
            in1 => \N__9731\,
            in2 => \N__8805\,
            in3 => \N__9251\,
            lcout => \spi0.n492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10687\,
            ce => 'H',
            sr => \N__9577\
        );

    \spi0.t_FSM_i9_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__9255\,
            in1 => \N__9673\,
            in2 => \N__8793\,
            in3 => \N__9738\,
            lcout => \spi0.n493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10687\,
            ce => 'H',
            sr => \N__9577\
        );

    \spi0.t_FSM_i8_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000010000"
        )
    port map (
            in0 => \N__9672\,
            in1 => \N__9733\,
            in2 => \N__8748\,
            in3 => \N__9254\,
            lcout => \spi0.n494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10687\,
            ce => 'H',
            sr => \N__9577\
        );

    \spi0.t_FSM_i7_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__9253\,
            in1 => \N__9671\,
            in2 => \N__8784\,
            in3 => \N__9737\,
            lcout => \spi0.n495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10687\,
            ce => 'H',
            sr => \N__9577\
        );

    \spi0.t_FSM_i3_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000010"
        )
    port map (
            in0 => \N__9756\,
            in1 => \N__9732\,
            in2 => \N__9678\,
            in3 => \N__9252\,
            lcout => \spi0.n499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10687\,
            ce => 'H',
            sr => \N__9577\
        );

    \spi0.state_reg_2__I_0_101_i5_2_lut_3_lut_3_lut_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__9411\,
            in1 => \N__9342\,
            in2 => \_gnd_net_\,
            in3 => \N__9256\,
            lcout => n5_adj_507,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i2_3_lut_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__9125\,
            in1 => \N__10689\,
            in2 => \_gnd_net_\,
            in3 => \N__8996\,
            lcout => \DEBUG_6_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.start_transfer_prev_74_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11938\,
            lcout => start_transfer_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i4_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11373\,
            in1 => \N__11845\,
            in2 => \_gnd_net_\,
            in3 => \N__9055\,
            lcout => tx_data_byte_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i6_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11103\,
            in1 => \N__11849\,
            in2 => \_gnd_net_\,
            in3 => \N__9025\,
            lcout => tx_data_byte_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12500\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.start_transfer_edge_73_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__8975\,
            in1 => \N__9012\,
            in2 => \N__11945\,
            in3 => \N__9003\,
            lcout => start_transfer_edge,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12500\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.spi_clk_counter_587__i0_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9872\,
            in2 => \_gnd_net_\,
            in3 => \N__8964\,
            lcout => \spi0.spi_clk_counter_0\,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \spi0.n2915\,
            clk => \N__12503\,
            ce => 'H',
            sr => \N__9815\
        );

    \spi0.spi_clk_counter_587__i1_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9902\,
            in2 => \N__10106\,
            in3 => \N__8961\,
            lcout => \spi0.spi_clk_counter_1\,
            ltout => OPEN,
            carryin => \spi0.n2915\,
            carryout => \spi0.n2916\,
            clk => \N__12503\,
            ce => 'H',
            sr => \N__9815\
        );

    \spi0.spi_clk_counter_587__i2_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10053\,
            in2 => \N__9861\,
            in3 => \N__10239\,
            lcout => \spi0.spi_clk_counter_2\,
            ltout => OPEN,
            carryin => \spi0.n2916\,
            carryout => \spi0.n2917\,
            clk => \N__12503\,
            ce => 'H',
            sr => \N__9815\
        );

    \spi0.spi_clk_counter_587__i3_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9845\,
            in2 => \N__10107\,
            in3 => \N__10236\,
            lcout => \spi0.spi_clk_counter_3\,
            ltout => OPEN,
            carryin => \spi0.n2917\,
            carryout => \spi0.n2918\,
            clk => \N__12503\,
            ce => 'H',
            sr => \N__9815\
        );

    \spi0.spi_clk_counter_587__i4_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10057\,
            in2 => \N__9831\,
            in3 => \N__10233\,
            lcout => \spi0.spi_clk_counter_4\,
            ltout => OPEN,
            carryin => \spi0.n2918\,
            carryout => \spi0.n2919\,
            clk => \N__12503\,
            ce => 'H',
            sr => \N__9815\
        );

    \spi0.spi_clk_counter_587__i5_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__9890\,
            in1 => \_gnd_net_\,
            in2 => \N__10108\,
            in3 => \N__9906\,
            lcout => \spi0.spi_clk_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12503\,
            ce => 'H',
            sr => \N__9815\
        );

    \tx_data_byte_r_i0_i1_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11880\,
            in1 => \N__9788\,
            in2 => \_gnd_net_\,
            in3 => \N__12039\,
            lcout => tx_data_byte_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i4_4_lut_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9903\,
            in1 => \N__9891\,
            in2 => \N__9879\,
            in3 => \N__9860\,
            lcout => OPEN,
            ltout => \spi0.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.i2987_3_lut_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__9846\,
            in1 => \_gnd_net_\,
            in2 => \N__9834\,
            in3 => \N__9830\,
            lcout => \spi0.n1896\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i1_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11879\,
            in1 => \N__9787\,
            in2 => \_gnd_net_\,
            in3 => \N__9767\,
            lcout => tx_addr_byte_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i4_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10499\,
            in2 => \_gnd_net_\,
            in3 => \N__10813\,
            lcout => rx_shift_reg_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i7_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10257\,
            in1 => \N__10453\,
            in2 => \_gnd_net_\,
            in3 => \N__10362\,
            lcout => rx_buf_byte_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i4_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10360\,
            in1 => \N__10409\,
            in2 => \_gnd_net_\,
            in3 => \N__10251\,
            lcout => rx_buf_byte_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i2_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10293\,
            in1 => \N__10373\,
            in2 => \_gnd_net_\,
            in3 => \N__10359\,
            lcout => rx_buf_byte_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.Rx_Lower_Byte_i5_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10361\,
            in1 => \N__10304\,
            in2 => \_gnd_net_\,
            in3 => \N__10716\,
            lcout => rx_buf_byte_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i5_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10292\,
            in2 => \_gnd_net_\,
            in3 => \N__10814\,
            lcout => rx_shift_reg_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i6_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__10815\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10280\,
            lcout => rx_shift_reg_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i8_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__10811\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10715\,
            lcout => rx_shift_reg_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i9_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10268\,
            in2 => \_gnd_net_\,
            in3 => \N__10812\,
            lcout => rx_shift_reg_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi0.rx__5_i7_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10250\,
            in2 => \_gnd_net_\,
            in3 => \N__10810\,
            lcout => rx_shift_reg_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2904_4_lut_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10893\,
            in1 => \N__10875\,
            in2 => \N__10956\,
            in3 => \N__10934\,
            lcout => OPEN,
            ltout => \pc_rx.n3291_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i4_4_lut_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__10833\,
            in1 => \N__10557\,
            in2 => \N__10560\,
            in3 => \N__10551\,
            lcout => \pc_rx.r_SM_Main_2_N_114_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10856\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10910\,
            lcout => \pc_rx.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_3_lut_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__10974\,
            in1 => \N__10518\,
            in2 => \_gnd_net_\,
            in3 => \N__10538\,
            lcout => \pc_rx.n3260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_4_lut_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10952\,
            in1 => \N__10973\,
            in2 => \N__10539\,
            in3 => \N__10517\,
            lcout => OPEN,
            ltout => \pc_rx.n3261_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2206_4_lut_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__10911\,
            in1 => \N__10935\,
            in2 => \N__10545\,
            in3 => \N__10892\,
            lcout => OPEN,
            ltout => \pc_rx.n2558_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2220_4_lut_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__10857\,
            in1 => \N__10832\,
            in2 => \N__10542\,
            in3 => \N__10874\,
            lcout => \r_SM_Main_2_N_108_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Clock_Count_584__i0_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10534\,
            in2 => \_gnd_net_\,
            in3 => \N__10521\,
            lcout => \pc_rx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \pc_rx.n2920\,
            clk => \N__12495\,
            ce => \N__11129\,
            sr => \N__11159\
        );

    \pc_rx.r_Clock_Count_584__i1_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10516\,
            in2 => \_gnd_net_\,
            in3 => \N__10977\,
            lcout => \pc_rx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \pc_rx.n2920\,
            carryout => \pc_rx.n2921\,
            clk => \N__12495\,
            ce => \N__11129\,
            sr => \N__11159\
        );

    \pc_rx.r_Clock_Count_584__i2_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10972\,
            in2 => \_gnd_net_\,
            in3 => \N__10959\,
            lcout => \pc_rx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \pc_rx.n2921\,
            carryout => \pc_rx.n2922\,
            clk => \N__12495\,
            ce => \N__11129\,
            sr => \N__11159\
        );

    \pc_rx.r_Clock_Count_584__i3_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10951\,
            in2 => \_gnd_net_\,
            in3 => \N__10938\,
            lcout => \pc_rx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \pc_rx.n2922\,
            carryout => \pc_rx.n2923\,
            clk => \N__12495\,
            ce => \N__11129\,
            sr => \N__11159\
        );

    \pc_rx.r_Clock_Count_584__i4_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10930\,
            in2 => \_gnd_net_\,
            in3 => \N__10914\,
            lcout => \pc_rx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \pc_rx.n2923\,
            carryout => \pc_rx.n2924\,
            clk => \N__12495\,
            ce => \N__11129\,
            sr => \N__11159\
        );

    \pc_rx.r_Clock_Count_584__i5_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10909\,
            in2 => \_gnd_net_\,
            in3 => \N__10896\,
            lcout => \pc_rx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \pc_rx.n2924\,
            carryout => \pc_rx.n2925\,
            clk => \N__12495\,
            ce => \N__11129\,
            sr => \N__11159\
        );

    \pc_rx.r_Clock_Count_584__i6_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10891\,
            in2 => \_gnd_net_\,
            in3 => \N__10878\,
            lcout => \pc_rx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \pc_rx.n2925\,
            carryout => \pc_rx.n2926\,
            clk => \N__12495\,
            ce => \N__11129\,
            sr => \N__11159\
        );

    \pc_rx.r_Clock_Count_584__i7_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10873\,
            in2 => \_gnd_net_\,
            in3 => \N__10860\,
            lcout => \pc_rx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \pc_rx.n2926\,
            carryout => \pc_rx.n2927\,
            clk => \N__12495\,
            ce => \N__11129\,
            sr => \N__11159\
        );

    \pc_rx.r_Clock_Count_584__i8_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10850\,
            in2 => \_gnd_net_\,
            in3 => \N__10839\,
            lcout => \pc_rx.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \pc_rx.n2928\,
            clk => \N__12501\,
            ce => \N__11133\,
            sr => \N__11160\
        );

    \pc_rx.r_Clock_Count_584__i9_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__10826\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10836\,
            lcout => \pc_rx.r_Clock_Count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12501\,
            ce => \N__11133\,
            sr => \N__11160\
        );

    \tx_data_byte_r_i0_i5_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12144\,
            in1 => \N__11878\,
            in2 => \_gnd_net_\,
            in3 => \N__11077\,
            lcout => tx_data_byte_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_addr_byte_r_i0_i2_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11029\,
            in1 => \N__11881\,
            in2 => \_gnd_net_\,
            in3 => \N__11051\,
            lcout => tx_addr_byte_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i2_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11030\,
            in1 => \N__11882\,
            in2 => \_gnd_net_\,
            in3 => \N__11715\,
            lcout => tx_data_byte_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_complete_rising_edge_207_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__11016\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10994\,
            lcout => uart_rx_complete_rising_edge,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2885_2_lut_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12008\,
            in2 => \_gnd_net_\,
            in3 => \N__11221\,
            lcout => \pc_rx.n3271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx_complete_prev_208_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10993\,
            lcout => uart_rx_complete_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_3_lut_4_lut_LC_19_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001111"
        )
    port map (
            in0 => \N__11680\,
            in1 => \N__11614\,
            in2 => \N__11486\,
            in3 => \N__11549\,
            lcout => OPEN,
            ltout => \n1764_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_DV_52_LC_19_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__11474\,
            in1 => \N__10992\,
            in2 => \N__11010\,
            in3 => \N__11681\,
            lcout => \DEBUG_1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2887_2_lut_3_lut_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__11220\,
            in1 => \N__11558\,
            in2 => \_gnd_net_\,
            in3 => \N__12009\,
            lcout => OPEN,
            ltout => \pc_rx.n3273_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_4_lut_adj_10_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001101"
        )
    port map (
            in0 => \N__11485\,
            in1 => \N__11604\,
            in2 => \N__11163\,
            in3 => \N__11670\,
            lcout => \pc_rx.n1910\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_SM_Main_i2_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__11664\,
            in1 => \N__11616\,
            in2 => \N__11574\,
            in3 => \N__11502\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2_3_lut_4_lut_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__11501\,
            in1 => \N__11615\,
            in2 => \N__11679\,
            in3 => \N__11570\,
            lcout => \pc_rx.n1715\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2_2_lut_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12011\,
            in2 => \_gnd_net_\,
            in3 => \N__11222\,
            lcout => OPEN,
            ltout => \pc_rx.n6_adj_492_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2981_4_lut_LC_19_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__11500\,
            in1 => \N__11663\,
            in2 => \N__11136\,
            in3 => \N__11569\,
            lcout => \pc_rx.n1815\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Bit_Index_i2_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11426\,
            in1 => \N__12121\,
            in2 => \_gnd_net_\,
            in3 => \N__12088\,
            lcout => \pc_rx.r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12504\,
            ce => \N__11514\,
            sr => \N__11691\
        );

    \pc_rx.r_Bit_Index_i1_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12087\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11425\,
            lcout => \pc_rx.r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12504\,
            ce => \N__11514\,
            sr => \N__11691\
        );

    \pc_rx.i2_3_lut_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__12123\,
            in1 => \N__12090\,
            in2 => \_gnd_net_\,
            in3 => \N__11190\,
            lcout => n1747,
            ltout => \n1747_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i6_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__11435\,
            in1 => \N__11099\,
            in2 => \N__11106\,
            in3 => \N__12021\,
            lcout => pc_data_rx_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_adj_13_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11434\,
            in2 => \_gnd_net_\,
            in3 => \N__11189\,
            lcout => n1754,
            ltout => \n1754_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i3_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__12016\,
            in1 => \N__11309\,
            in2 => \N__11316\,
            in3 => \N__11172\,
            lcout => pc_data_rx_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i7_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__11285\,
            in1 => \N__12017\,
            in2 => \N__11298\,
            in3 => \N__11436\,
            lcout => pc_data_rx_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tx_data_byte_r_i0_i7_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11840\,
            in1 => \N__11254\,
            in2 => \_gnd_net_\,
            in3 => \N__11289\,
            lcout => tx_data_byte_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12513\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_SM_Main_i1_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011110101010"
        )
    port map (
            in0 => \N__11470\,
            in1 => \N__11628\,
            in2 => \N__11238\,
            in3 => \N__11548\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12510\,
            ce => 'H',
            sr => \N__11685\
        );

    \pc_rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__11229\,
            in1 => \N__11980\,
            in2 => \_gnd_net_\,
            in3 => \N__11547\,
            lcout => OPEN,
            ltout => \pc_rx.n1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_SM_Main_i0_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__11196\,
            in1 => \_gnd_net_\,
            in2 => \N__11199\,
            in3 => \N__11469\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12510\,
            ce => 'H',
            sr => \N__11685\
        );

    \pc_rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001110111"
        )
    port map (
            in0 => \N__11397\,
            in1 => \N__11617\,
            in2 => \_gnd_net_\,
            in3 => \N__11550\,
            lcout => \pc_rx.n2578\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_2_lut_adj_12_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11183\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11422\,
            lcout => n1750,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.equal_258_i4_2_lut_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__12093\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12126\,
            lcout => n4_adj_504,
            ltout => \n4_adj_504_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i2_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__11705\,
            in1 => \N__12010\,
            in2 => \N__11718\,
            in3 => \N__11350\,
            lcout => pc_data_rx_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2957_2_lut_3_lut_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11396\,
            in1 => \N__11567\,
            in2 => \_gnd_net_\,
            in3 => \N__11626\,
            lcout => OPEN,
            ltout => \pc_rx.n3334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i1_4_lut_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000010001"
        )
    port map (
            in0 => \N__11566\,
            in1 => \N__11668\,
            in2 => \N__11694\,
            in3 => \N__11487\,
            lcout => \pc_rx.n1900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2996_3_lut_4_lut_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__11669\,
            in1 => \N__11627\,
            in2 => \N__11499\,
            in3 => \N__11568\,
            lcout => n3293,
            ltout => \n3293_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Bit_Index_i0_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101000000"
        )
    port map (
            in0 => \N__11392\,
            in1 => \N__11491\,
            in2 => \N__11439\,
            in3 => \N__11423\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.i2_2_lut_3_lut_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12122\,
            in1 => \N__12089\,
            in2 => \_gnd_net_\,
            in3 => \N__11424\,
            lcout => n2540,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i4_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__12012\,
            in1 => \N__11369\,
            in2 => \N__12156\,
            in3 => \N__11351\,
            lcout => pc_data_rx_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i0_LC_20_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__12013\,
            in1 => \N__11327\,
            in2 => \N__11358\,
            in3 => \N__12057\,
            lcout => pc_data_rx_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.equal_257_i4_2_lut_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12124\,
            in2 => \_gnd_net_\,
            in3 => \N__12091\,
            lcout => n4_adj_506,
            ltout => \n4_adj_506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i5_LC_20_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__12015\,
            in1 => \N__12137\,
            in2 => \N__12147\,
            in3 => \N__12048\,
            lcout => pc_data_rx_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.equal_261_i4_2_lut_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12125\,
            in2 => \_gnd_net_\,
            in3 => \N__12092\,
            lcout => n4_adj_500,
            ltout => \n4_adj_500_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Byte_i1_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__12014\,
            in1 => \N__12032\,
            in2 => \N__12051\,
            in3 => \N__12047\,
            lcout => pc_data_rx_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Data_50_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11739\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12515\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debug_check_211_LC_22_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11769\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11815\,
            lcout => \DEBUG_2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12515\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \even_byte_flag_214_LC_22_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11844\,
            in2 => \_gnd_net_\,
            in3 => \N__11768\,
            lcout => even_byte_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc_rx.r_Rx_Data_R_49_LC_23_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11757\,
            lcout => \pc_rx.r_Rx_Data_R\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i0_LC_24_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11727\,
            in2 => \_gnd_net_\,
            in3 => \N__11721\,
            lcout => n25,
            ltout => OPEN,
            carryin => \bfn_24_6_0_\,
            carryout => n2938,
            clk => \N__12522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i1_LC_24_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12228\,
            in2 => \_gnd_net_\,
            in3 => \N__12222\,
            lcout => n24,
            ltout => OPEN,
            carryin => n2938,
            carryout => n2939,
            clk => \N__12522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i2_LC_24_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12219\,
            in2 => \_gnd_net_\,
            in3 => \N__12213\,
            lcout => n23,
            ltout => OPEN,
            carryin => n2939,
            carryout => n2940,
            clk => \N__12522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i3_LC_24_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12210\,
            in2 => \_gnd_net_\,
            in3 => \N__12204\,
            lcout => n22,
            ltout => OPEN,
            carryin => n2940,
            carryout => n2941,
            clk => \N__12522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i4_LC_24_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12201\,
            in2 => \_gnd_net_\,
            in3 => \N__12195\,
            lcout => n21,
            ltout => OPEN,
            carryin => n2941,
            carryout => n2942,
            clk => \N__12522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i5_LC_24_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12192\,
            in2 => \_gnd_net_\,
            in3 => \N__12186\,
            lcout => n20,
            ltout => OPEN,
            carryin => n2942,
            carryout => n2943,
            clk => \N__12522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i6_LC_24_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12183\,
            in2 => \_gnd_net_\,
            in3 => \N__12177\,
            lcout => n19,
            ltout => OPEN,
            carryin => n2943,
            carryout => n2944,
            clk => \N__12522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i7_LC_24_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12174\,
            in2 => \_gnd_net_\,
            in3 => \N__12168\,
            lcout => n18,
            ltout => OPEN,
            carryin => n2944,
            carryout => n2945,
            clk => \N__12522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i8_LC_24_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12165\,
            in2 => \_gnd_net_\,
            in3 => \N__12159\,
            lcout => n17,
            ltout => OPEN,
            carryin => \bfn_24_7_0_\,
            carryout => n2946,
            clk => \N__12521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i9_LC_24_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12309\,
            in2 => \_gnd_net_\,
            in3 => \N__12303\,
            lcout => n16,
            ltout => OPEN,
            carryin => n2946,
            carryout => n2947,
            clk => \N__12521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i10_LC_24_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12300\,
            in2 => \_gnd_net_\,
            in3 => \N__12294\,
            lcout => n15,
            ltout => OPEN,
            carryin => n2947,
            carryout => n2948,
            clk => \N__12521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i11_LC_24_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12291\,
            in2 => \_gnd_net_\,
            in3 => \N__12285\,
            lcout => n14,
            ltout => OPEN,
            carryin => n2948,
            carryout => n2949,
            clk => \N__12521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i12_LC_24_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12282\,
            in2 => \_gnd_net_\,
            in3 => \N__12276\,
            lcout => n13,
            ltout => OPEN,
            carryin => n2949,
            carryout => n2950,
            clk => \N__12521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i13_LC_24_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12273\,
            in2 => \_gnd_net_\,
            in3 => \N__12267\,
            lcout => n12,
            ltout => OPEN,
            carryin => n2950,
            carryout => n2951,
            clk => \N__12521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i14_LC_24_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12264\,
            in2 => \_gnd_net_\,
            in3 => \N__12258\,
            lcout => n11,
            ltout => OPEN,
            carryin => n2951,
            carryout => n2952,
            clk => \N__12521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i15_LC_24_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12255\,
            in2 => \_gnd_net_\,
            in3 => \N__12249\,
            lcout => n10,
            ltout => OPEN,
            carryin => n2952,
            carryout => n2953,
            clk => \N__12521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i16_LC_24_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12246\,
            in2 => \_gnd_net_\,
            in3 => \N__12240\,
            lcout => n9,
            ltout => OPEN,
            carryin => \bfn_24_8_0_\,
            carryout => n2954,
            clk => \N__12520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i17_LC_24_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12237\,
            in2 => \_gnd_net_\,
            in3 => \N__12231\,
            lcout => n8_adj_501,
            ltout => OPEN,
            carryin => n2954,
            carryout => n2955,
            clk => \N__12520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i18_LC_24_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12609\,
            in2 => \_gnd_net_\,
            in3 => \N__12603\,
            lcout => n7,
            ltout => OPEN,
            carryin => n2955,
            carryout => n2956,
            clk => \N__12520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i19_LC_24_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12600\,
            in2 => \_gnd_net_\,
            in3 => \N__12594\,
            lcout => n6,
            ltout => OPEN,
            carryin => n2956,
            carryout => n2957,
            clk => \N__12520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i20_LC_24_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12591\,
            in2 => \_gnd_net_\,
            in3 => \N__12585\,
            lcout => n5,
            ltout => OPEN,
            carryin => n2957,
            carryout => n2958,
            clk => \N__12520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i21_LC_24_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12582\,
            in2 => \_gnd_net_\,
            in3 => \N__12576\,
            lcout => n4_adj_502,
            ltout => OPEN,
            carryin => n2958,
            carryout => n2959,
            clk => \N__12520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i22_LC_24_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12573\,
            in2 => \_gnd_net_\,
            in3 => \N__12567\,
            lcout => n3,
            ltout => OPEN,
            carryin => n2959,
            carryout => n2960,
            clk => \N__12520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i23_LC_24_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12564\,
            in2 => \_gnd_net_\,
            in3 => \N__12558\,
            lcout => n2_adj_503,
            ltout => OPEN,
            carryin => n2960,
            carryout => n2961,
            clk => \N__12520\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_counter_581_788__i24_LC_24_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12539\,
            in2 => \_gnd_net_\,
            in3 => \N__12555\,
            lcout => \DEBUG_0_c_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12519\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_SLM_CLK_c_THRU_LUT4_0_LC_24_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_SLM_CLK_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// uart.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module uart (
		input  wire        clk_clk,                               //                        clk.clk
		input  wire        reset_reset_n,                         //                      reset.reset_n
		input  wire        rs232_0_avalon_rs232_slave_address,    // rs232_0_avalon_rs232_slave.address
		input  wire        rs232_0_avalon_rs232_slave_chipselect, //                           .chipselect
		input  wire [3:0]  rs232_0_avalon_rs232_slave_byteenable, //                           .byteenable
		input  wire        rs232_0_avalon_rs232_slave_read,       //                           .read
		input  wire        rs232_0_avalon_rs232_slave_write,      //                           .write
		input  wire [31:0] rs232_0_avalon_rs232_slave_writedata,  //                           .writedata
		output wire [31:0] rs232_0_avalon_rs232_slave_readdata,   //                           .readdata
		input  wire        rs232_0_clk_clk,                       //                rs232_0_clk.clk
		input  wire        rs232_0_external_interface_RXD,        // rs232_0_external_interface.RXD
		output wire        rs232_0_external_interface_TXD,        //                           .TXD
		output wire        rs232_0_interrupt_irq,                 //          rs232_0_interrupt.irq
		input  wire        rs232_0_reset_reset                    //              rs232_0_reset.reset
	);

	uart_rs232_0 rs232_0 (
		.clk        (rs232_0_clk_clk),                       //                clk.clk
		.reset      (rs232_0_reset_reset),                   //              reset.reset
		.address    (rs232_0_avalon_rs232_slave_address),    // avalon_rs232_slave.address
		.chipselect (rs232_0_avalon_rs232_slave_chipselect), //                   .chipselect
		.byteenable (rs232_0_avalon_rs232_slave_byteenable), //                   .byteenable
		.read       (rs232_0_avalon_rs232_slave_read),       //                   .read
		.write      (rs232_0_avalon_rs232_slave_write),      //                   .write
		.writedata  (rs232_0_avalon_rs232_slave_writedata),  //                   .writedata
		.readdata   (rs232_0_avalon_rs232_slave_readdata),   //                   .readdata
		.irq        (rs232_0_interrupt_irq),                 //          interrupt.irq
		.UART_RXD   (rs232_0_external_interface_RXD),        // external_interface.export
		.UART_TXD   (rs232_0_external_interface_TXD)         //                   .export
	);

endmodule
